
module matrix_mult_N_M_3_N16_M32 ( clk, rst, g_input, e_input, o );
  input [31:0] g_input;
  input [31:0] e_input;
  output [31:0] o;
  input clk, rst;
  wire   n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486;
  wire   [31:0] oi;

  DFF \o_reg[0]  ( .D(oi[0]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[0]) );
  DFF \o_reg[1]  ( .D(oi[1]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[1]) );
  DFF \o_reg[2]  ( .D(oi[2]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[2]) );
  DFF \o_reg[3]  ( .D(oi[3]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[3]) );
  DFF \o_reg[4]  ( .D(oi[4]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[4]) );
  DFF \o_reg[5]  ( .D(oi[5]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[5]) );
  DFF \o_reg[6]  ( .D(oi[6]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[6]) );
  DFF \o_reg[7]  ( .D(oi[7]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[7]) );
  DFF \o_reg[8]  ( .D(oi[8]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[8]) );
  DFF \o_reg[9]  ( .D(oi[9]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[9]) );
  DFF \o_reg[10]  ( .D(oi[10]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[10]) );
  DFF \o_reg[11]  ( .D(oi[11]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[11]) );
  DFF \o_reg[12]  ( .D(oi[12]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[12]) );
  DFF \o_reg[13]  ( .D(oi[13]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[13]) );
  DFF \o_reg[14]  ( .D(oi[14]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[14]) );
  DFF \o_reg[15]  ( .D(oi[15]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[15]) );
  DFF \o_reg[16]  ( .D(oi[16]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[16]) );
  DFF \o_reg[17]  ( .D(oi[17]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[17]) );
  DFF \o_reg[18]  ( .D(oi[18]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[18]) );
  DFF \o_reg[19]  ( .D(oi[19]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[19]) );
  DFF \o_reg[20]  ( .D(oi[20]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[20]) );
  DFF \o_reg[21]  ( .D(oi[21]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[21]) );
  DFF \o_reg[22]  ( .D(oi[22]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[22]) );
  DFF \o_reg[23]  ( .D(oi[23]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[23]) );
  DFF \o_reg[24]  ( .D(oi[24]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[24]) );
  DFF \o_reg[25]  ( .D(oi[25]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[25]) );
  DFF \o_reg[26]  ( .D(oi[26]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[26]) );
  DFF \o_reg[27]  ( .D(oi[27]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[27]) );
  DFF \o_reg[28]  ( .D(oi[28]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[28]) );
  DFF \o_reg[29]  ( .D(oi[29]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[29]) );
  DFF \o_reg[30]  ( .D(oi[30]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[30]) );
  DFF \o_reg[31]  ( .D(oi[31]), .CLK(clk), .RST(rst), .I(1'b0), .Q(o[31]) );
  MUX U35 ( .IN0(n1374), .IN1(n33), .SEL(n1375), .F(n1273) );
  IV U36 ( .A(n1376), .Z(n33) );
  MUX U37 ( .IN0(n1381), .IN1(n34), .SEL(n1382), .F(n1279) );
  IV U38 ( .A(n1383), .Z(n34) );
  MUX U39 ( .IN0(n1727), .IN1(n35), .SEL(n1728), .F(n1646) );
  IV U40 ( .A(n1729), .Z(n35) );
  MUX U41 ( .IN0(n1387), .IN1(n36), .SEL(n1388), .F(n1286) );
  IV U42 ( .A(n1389), .Z(n36) );
  XOR U43 ( .A(n1174), .B(n1173), .Z(n1260) );
  XOR U44 ( .A(n826), .B(n825), .Z(n930) );
  MUX U45 ( .IN0(n1294), .IN1(n37), .SEL(n1295), .F(n1183) );
  IV U46 ( .A(n1296), .Z(n37) );
  MUX U47 ( .IN0(n1301), .IN1(n38), .SEL(n1302), .F(n1193) );
  IV U48 ( .A(n1303), .Z(n38) );
  MUX U49 ( .IN0(n951), .IN1(n39), .SEL(n952), .F(n838) );
  IV U50 ( .A(n953), .Z(n39) );
  XOR U51 ( .A(n960), .B(n959), .Z(n1033) );
  MUX U52 ( .IN0(n2019), .IN1(n40), .SEL(n2020), .F(n1954) );
  IV U53 ( .A(n2021), .Z(n40) );
  MUX U54 ( .IN0(n969), .IN1(n41), .SEL(n970), .F(n856) );
  IV U55 ( .A(n971), .Z(n41) );
  MUX U56 ( .IN0(n1207), .IN1(n42), .SEL(n1208), .F(n1090) );
  IV U57 ( .A(n1209), .Z(n42) );
  XOR U58 ( .A(n978), .B(n977), .Z(n1027) );
  MUX U59 ( .IN0(n1219), .IN1(n43), .SEL(n1220), .F(n1104) );
  IV U60 ( .A(n1221), .Z(n43) );
  MUX U61 ( .IN0(n1419), .IN1(n44), .SEL(n1420), .F(n1319) );
  IV U62 ( .A(n1421), .Z(n44) );
  MUX U63 ( .IN0(n1600), .IN1(n45), .SEL(n1601), .F(n1511) );
  IV U64 ( .A(n1602), .Z(n45) );
  MUX U65 ( .IN0(n1760), .IN1(n46), .SEL(n1761), .F(n1679) );
  IV U66 ( .A(n1762), .Z(n46) );
  MUX U67 ( .IN0(n2242), .IN1(n47), .SEL(n2243), .F(n2193) );
  IV U68 ( .A(n2244), .Z(n47) );
  MUX U69 ( .IN0(n2347), .IN1(n48), .SEL(n2348), .F(n2281) );
  IV U70 ( .A(n2349), .Z(n48) );
  XOR U71 ( .A(n877), .B(n876), .Z(n913) );
  MUX U72 ( .IN0(n886), .IN1(n49), .SEL(n887), .F(n766) );
  IV U73 ( .A(n888), .Z(n49) );
  MUX U74 ( .IN0(n1561), .IN1(n50), .SEL(n1562), .F(n1468) );
  IV U75 ( .A(n1563), .Z(n50) );
  XOR U76 ( .A(n1273), .B(n1271), .Z(n1365) );
  MUX U77 ( .IN0(n1567), .IN1(n51), .SEL(n1568), .F(n1476) );
  IV U78 ( .A(n1569), .Z(n51) );
  XOR U79 ( .A(n1171), .B(n1170), .Z(n1261) );
  MUX U80 ( .IN0(n1809), .IN1(n52), .SEL(n1810), .F(n1730) );
  IV U81 ( .A(n1811), .Z(n52) );
  XOR U82 ( .A(n942), .B(n941), .Z(n1039) );
  MUX U83 ( .IN0(n1576), .IN1(n53), .SEL(n1577), .F(n1487) );
  IV U84 ( .A(n1578), .Z(n53) );
  XOR U85 ( .A(n1183), .B(n1182), .Z(n1257) );
  MUX U86 ( .IN0(n1815), .IN1(n54), .SEL(n1816), .F(n1736) );
  IV U87 ( .A(n1817), .Z(n54) );
  MUX U88 ( .IN0(n2013), .IN1(n55), .SEL(n2014), .F(n1948) );
  IV U89 ( .A(n2015), .Z(n55) );
  XOR U90 ( .A(n835), .B(n834), .Z(n927) );
  MUX U91 ( .IN0(n1196), .IN1(n56), .SEL(n1197), .F(n1078) );
  IV U92 ( .A(n1198), .Z(n56) );
  XOR U93 ( .A(n847), .B(n846), .Z(n923) );
  MUX U94 ( .IN0(n1407), .IN1(n57), .SEL(n1408), .F(n1307) );
  IV U95 ( .A(n1409), .Z(n57) );
  MUX U96 ( .IN0(n1960), .IN1(n58), .SEL(n1961), .F(n1891) );
  IV U97 ( .A(n1962), .Z(n58) );
  MUX U98 ( .IN0(n2134), .IN1(n59), .SEL(n2135), .F(n2077) );
  IV U99 ( .A(n2136), .Z(n59) );
  MUX U100 ( .IN0(n2230), .IN1(n2232), .SEL(n2231), .F(n2181) );
  XOR U101 ( .A(n1090), .B(n1088), .Z(n1142) );
  MUX U102 ( .IN0(n1897), .IN1(n60), .SEL(n1898), .F(n1824) );
  IV U103 ( .A(n1899), .Z(n60) );
  MUX U104 ( .IN0(n2083), .IN1(n61), .SEL(n2084), .F(n2022) );
  IV U105 ( .A(n2085), .Z(n61) );
  XOR U106 ( .A(n981), .B(n980), .Z(n1026) );
  MUX U107 ( .IN0(n1322), .IN1(n62), .SEL(n1323), .F(n1216) );
  IV U108 ( .A(n1324), .Z(n62) );
  MUX U109 ( .IN0(n1514), .IN1(n63), .SEL(n1515), .F(n1416) );
  IV U110 ( .A(n1516), .Z(n63) );
  MUX U111 ( .IN0(n1682), .IN1(n64), .SEL(n1683), .F(n1597) );
  IV U112 ( .A(n1684), .Z(n64) );
  MUX U113 ( .IN0(n1836), .IN1(n65), .SEL(n1837), .F(n1757) );
  IV U114 ( .A(n1838), .Z(n65) );
  MUX U115 ( .IN0(n1972), .IN1(n66), .SEL(n1973), .F(n1903) );
  IV U116 ( .A(n1974), .Z(n66) );
  MUX U117 ( .IN0(n2196), .IN1(n67), .SEL(n2197), .F(n2143) );
  IV U118 ( .A(n2198), .Z(n67) );
  MUX U119 ( .IN0(n2284), .IN1(n68), .SEL(n2285), .F(n2239) );
  IV U120 ( .A(n2286), .Z(n68) );
  MUX U121 ( .IN0(n2376), .IN1(n69), .SEL(n2377), .F(n2344) );
  IV U122 ( .A(n2378), .Z(n69) );
  MUX U123 ( .IN0(n877), .IN1(n70), .SEL(n878), .F(n757) );
  IV U124 ( .A(n879), .Z(n70) );
  MUX U125 ( .IN0(n1112), .IN1(n71), .SEL(n1113), .F(n994) );
  IV U126 ( .A(n1114), .Z(n71) );
  MUX U127 ( .IN0(n2149), .IN1(n72), .SEL(n2150), .F(n2092) );
  IV U128 ( .A(n2151), .Z(n72) );
  MUX U129 ( .IN0(n1000), .IN1(n73), .SEL(n1001), .F(n886) );
  IV U130 ( .A(n1002), .Z(n73) );
  MUX U131 ( .IN0(n1371), .IN1(n74), .SEL(n1372), .F(n1269) );
  IV U132 ( .A(n1373), .Z(n74) );
  MUX U133 ( .IN0(n1476), .IN1(n75), .SEL(n1477), .F(n1378) );
  IV U134 ( .A(n1478), .Z(n75) );
  MUX U135 ( .IN0(n1649), .IN1(n76), .SEL(n1650), .F(n1564) );
  IV U136 ( .A(n1651), .Z(n76) );
  XOR U137 ( .A(n1053), .B(n1052), .Z(n1153) );
  MUX U138 ( .IN0(n1282), .IN1(n77), .SEL(n1283), .F(n1174) );
  IV U139 ( .A(n1284), .Z(n77) );
  MUX U140 ( .IN0(n1655), .IN1(n78), .SEL(n1656), .F(n1570) );
  IV U141 ( .A(n1657), .Z(n78) );
  MUX U142 ( .IN0(n1490), .IN1(n79), .SEL(n1491), .F(n1390) );
  IV U143 ( .A(n1492), .Z(n79) );
  MUX U144 ( .IN0(n1948), .IN1(n80), .SEL(n1949), .F(n1879) );
  IV U145 ( .A(n1950), .Z(n80) );
  MUX U146 ( .IN0(n826), .IN1(n81), .SEL(n827), .F(n706) );
  IV U147 ( .A(n828), .Z(n81) );
  MUX U148 ( .IN0(n1063), .IN1(n82), .SEL(n1064), .F(n951) );
  IV U149 ( .A(n1065), .Z(n82) );
  MUX U150 ( .IN0(n1661), .IN1(n83), .SEL(n1662), .F(n1576) );
  IV U151 ( .A(n1663), .Z(n83) );
  MUX U152 ( .IN0(n1885), .IN1(n84), .SEL(n1886), .F(n1812) );
  IV U153 ( .A(n1887), .Z(n84) );
  MUX U154 ( .IN0(n832), .IN1(n85), .SEL(n833), .F(n712) );
  IV U155 ( .A(n834), .Z(n85) );
  XOR U156 ( .A(n1193), .B(n1191), .Z(n1255) );
  MUX U157 ( .IN0(n1496), .IN1(n86), .SEL(n1497), .F(n1398) );
  IV U158 ( .A(n1498), .Z(n86) );
  MUX U159 ( .IN0(n1818), .IN1(n87), .SEL(n1819), .F(n1739) );
  IV U160 ( .A(n1820), .Z(n87) );
  MUX U161 ( .IN0(n841), .IN1(n88), .SEL(n842), .F(n721) );
  IV U162 ( .A(n843), .Z(n88) );
  XOR U163 ( .A(n1082), .B(n1080), .Z(n1144) );
  MUX U164 ( .IN0(n2077), .IN1(n89), .SEL(n2078), .F(n2016) );
  IV U165 ( .A(n2079), .Z(n89) );
  MUX U166 ( .IN0(n1310), .IN1(n90), .SEL(n1311), .F(n1204) );
  IV U167 ( .A(n1312), .Z(n90) );
  MUX U168 ( .IN0(n1502), .IN1(n91), .SEL(n1503), .F(n1404) );
  IV U169 ( .A(n1504), .Z(n91) );
  XOR U170 ( .A(n850), .B(n849), .Z(n922) );
  MUX U171 ( .IN0(n1673), .IN1(n92), .SEL(n1674), .F(n1588) );
  IV U172 ( .A(n1675), .Z(n92) );
  MUX U173 ( .IN0(n1827), .IN1(n93), .SEL(n1828), .F(n1748) );
  IV U174 ( .A(n1829), .Z(n93) );
  MUX U175 ( .IN0(n1963), .IN1(n94), .SEL(n1964), .F(n1894) );
  IV U176 ( .A(n1965), .Z(n94) );
  MUX U177 ( .IN0(n2233), .IN1(n95), .SEL(n2234), .F(n2184) );
  IV U178 ( .A(n2235), .Z(n95) );
  MUX U179 ( .IN0(n1095), .IN1(n96), .SEL(n1096), .F(n978) );
  IV U180 ( .A(n1097), .Z(n96) );
  XOR U181 ( .A(n862), .B(n861), .Z(n918) );
  MUX U182 ( .IN0(n2190), .IN1(n97), .SEL(n2191), .F(n2137) );
  IV U183 ( .A(n2192), .Z(n97) );
  MUX U184 ( .IN0(n2143), .IN1(n98), .SEL(n2144), .F(n2086) );
  IV U185 ( .A(n2145), .Z(n98) );
  XOR U186 ( .A(n988), .B(n987), .Z(n1024) );
  MUX U187 ( .IN0(n1975), .IN1(n99), .SEL(n1976), .F(n1906) );
  IV U188 ( .A(n1977), .Z(n99) );
  MUX U189 ( .IN0(n2095), .IN1(n100), .SEL(n2096), .F(n2034) );
  IV U190 ( .A(n2097), .Z(n100) );
  MUX U191 ( .IN0(n2199), .IN1(n101), .SEL(n2200), .F(n2146) );
  IV U192 ( .A(n2201), .Z(n101) );
  XOR U193 ( .A(n883), .B(n882), .Z(n911) );
  MUX U194 ( .IN0(n1225), .IN1(n102), .SEL(n1226), .F(n1112) );
  IV U195 ( .A(n1227), .Z(n102) );
  MUX U196 ( .IN0(n1425), .IN1(n103), .SEL(n1426), .F(n1325) );
  IV U197 ( .A(n1427), .Z(n103) );
  MUX U198 ( .IN0(n1606), .IN1(n104), .SEL(n1607), .F(n1517) );
  IV U199 ( .A(n1608), .Z(n104) );
  MUX U200 ( .IN0(n1766), .IN1(n105), .SEL(n1767), .F(n1685) );
  IV U201 ( .A(n1768), .Z(n105) );
  MUX U202 ( .IN0(n1912), .IN1(n106), .SEL(n1913), .F(n1839) );
  IV U203 ( .A(n1914), .Z(n106) );
  MUX U204 ( .IN0(n2353), .IN1(n107), .SEL(n2354), .F(n2287) );
  IV U205 ( .A(n2355), .Z(n107) );
  MUX U206 ( .IN0(n2407), .IN1(n108), .SEL(n2408), .F(n2379) );
  IV U207 ( .A(n2409), .Z(n108) );
  MUX U208 ( .IN0(n1003), .IN1(n109), .SEL(n1004), .F(n889) );
  IV U209 ( .A(n1005), .Z(n109) );
  MUX U210 ( .IN0(n1464), .IN1(n1466), .SEL(n1465), .F(n1368) );
  MUX U211 ( .IN0(n1646), .IN1(n110), .SEL(n1647), .F(n1561) );
  IV U212 ( .A(n1648), .Z(n110) );
  MUX U213 ( .IN0(n1378), .IN1(n111), .SEL(n1379), .F(n1276) );
  IV U214 ( .A(n1380), .Z(n111) );
  MUX U215 ( .IN0(n1269), .IN1(n112), .SEL(n1270), .F(n1160) );
  IV U216 ( .A(n1271), .Z(n112) );
  MUX U217 ( .IN0(n1479), .IN1(n113), .SEL(n1480), .F(n1381) );
  IV U218 ( .A(n1481), .Z(n113) );
  MUX U219 ( .IN0(n1803), .IN1(n1805), .SEL(n1804), .F(n1724) );
  XOR U220 ( .A(n1050), .B(n1048), .Z(n1154) );
  MUX U221 ( .IN0(n1390), .IN1(n114), .SEL(n1391), .F(n1289) );
  IV U222 ( .A(n1392), .Z(n114) );
  MUX U223 ( .IN0(n1733), .IN1(n115), .SEL(n1734), .F(n1652) );
  IV U224 ( .A(n1735), .Z(n115) );
  MUX U225 ( .IN0(n1177), .IN1(n116), .SEL(n1178), .F(n1063) );
  IV U226 ( .A(n1179), .Z(n116) );
  MUX U227 ( .IN0(n1658), .IN1(n117), .SEL(n1659), .F(n1573) );
  IV U228 ( .A(n1660), .Z(n117) );
  XOR U229 ( .A(n829), .B(n828), .Z(n929) );
  MUX U230 ( .IN0(n1493), .IN1(n118), .SEL(n1494), .F(n1393) );
  IV U231 ( .A(n1495), .Z(n118) );
  MUX U232 ( .IN0(n1951), .IN1(n119), .SEL(n1952), .F(n1882) );
  IV U233 ( .A(n1953), .Z(n119) );
  XOR U234 ( .A(n712), .B(n711), .Z(n815) );
  XOR U235 ( .A(n954), .B(n953), .Z(n1035) );
  MUX U236 ( .IN0(n1401), .IN1(n120), .SEL(n1402), .F(n1301) );
  IV U237 ( .A(n1403), .Z(n120) );
  XOR U238 ( .A(n1196), .B(n1195), .Z(n1254) );
  MUX U239 ( .IN0(n1745), .IN1(n121), .SEL(n1746), .F(n1664) );
  IV U240 ( .A(n1747), .Z(n121) );
  MUX U241 ( .IN0(n1957), .IN1(n122), .SEL(n1958), .F(n1888) );
  IV U242 ( .A(n1959), .Z(n122) );
  MUX U243 ( .IN0(n2131), .IN1(n123), .SEL(n2132), .F(n2074) );
  IV U244 ( .A(n2133), .Z(n123) );
  MUX U245 ( .IN0(n1670), .IN1(n124), .SEL(n1671), .F(n1585) );
  IV U246 ( .A(n1672), .Z(n124) );
  MUX U247 ( .IN0(n1894), .IN1(n125), .SEL(n1895), .F(n1821) );
  IV U248 ( .A(n1896), .Z(n125) );
  XOR U249 ( .A(n727), .B(n726), .Z(n810) );
  MUX U250 ( .IN0(n856), .IN1(n126), .SEL(n857), .F(n736) );
  IV U251 ( .A(n858), .Z(n126) );
  MUX U252 ( .IN0(n2137), .IN1(n127), .SEL(n2138), .F(n2080) );
  IV U253 ( .A(n2139), .Z(n127) );
  MUX U254 ( .IN0(n1098), .IN1(n128), .SEL(n1099), .F(n981) );
  IV U255 ( .A(n1100), .Z(n128) );
  MUX U256 ( .IN0(n1316), .IN1(n129), .SEL(n1317), .F(n1210) );
  IV U257 ( .A(n1318), .Z(n129) );
  MUX U258 ( .IN0(n1508), .IN1(n130), .SEL(n1509), .F(n1410) );
  IV U259 ( .A(n1510), .Z(n130) );
  MUX U260 ( .IN0(n1676), .IN1(n131), .SEL(n1677), .F(n1591) );
  IV U261 ( .A(n1678), .Z(n131) );
  MUX U262 ( .IN0(n1900), .IN1(n132), .SEL(n1901), .F(n1827) );
  IV U263 ( .A(n1902), .Z(n132) );
  MUX U264 ( .IN0(n2086), .IN1(n133), .SEL(n2087), .F(n2025) );
  IV U265 ( .A(n2088), .Z(n133) );
  MUX U266 ( .IN0(n2236), .IN1(n134), .SEL(n2237), .F(n2187) );
  IV U267 ( .A(n2238), .Z(n134) );
  MUX U268 ( .IN0(n862), .IN1(n135), .SEL(n863), .F(n742) );
  IV U269 ( .A(n864), .Z(n135) );
  MUX U270 ( .IN0(n2031), .IN1(n136), .SEL(n2032), .F(n1966) );
  IV U271 ( .A(n2033), .Z(n136) );
  MUX U272 ( .IN0(n2373), .IN1(n2375), .SEL(n2374), .F(n2341) );
  MUX U273 ( .IN0(n1104), .IN1(n137), .SEL(n1105), .F(n988) );
  IV U274 ( .A(n1106), .Z(n137) );
  MUX U275 ( .IN0(n871), .IN1(n138), .SEL(n872), .F(n751) );
  IV U276 ( .A(n873), .Z(n138) );
  MUX U277 ( .IN0(n2146), .IN1(n139), .SEL(n2147), .F(n2089) );
  IV U278 ( .A(n2148), .Z(n139) );
  MUX U279 ( .IN0(n2037), .IN1(n140), .SEL(n2038), .F(n1972) );
  IV U280 ( .A(n2039), .Z(n140) );
  MUX U281 ( .IN0(n994), .IN1(n141), .SEL(n995), .F(n880) );
  IV U282 ( .A(n996), .Z(n141) );
  MUX U283 ( .IN0(n1115), .IN1(n142), .SEL(n1116), .F(n997) );
  IV U284 ( .A(n1117), .Z(n142) );
  MUX U285 ( .IN0(n1328), .IN1(n143), .SEL(n1329), .F(n1222) );
  IV U286 ( .A(n1330), .Z(n143) );
  MUX U287 ( .IN0(n1520), .IN1(n144), .SEL(n1521), .F(n1422) );
  IV U288 ( .A(n1522), .Z(n144) );
  MUX U289 ( .IN0(n1688), .IN1(n145), .SEL(n1689), .F(n1603) );
  IV U290 ( .A(n1690), .Z(n145) );
  MUX U291 ( .IN0(n1842), .IN1(n146), .SEL(n1843), .F(n1763) );
  IV U292 ( .A(n1844), .Z(n146) );
  MUX U293 ( .IN0(n1978), .IN1(n147), .SEL(n1979), .F(n1909) );
  IV U294 ( .A(n1980), .Z(n147) );
  MUX U295 ( .IN0(n2152), .IN1(n148), .SEL(n2153), .F(n2095) );
  IV U296 ( .A(n2154), .Z(n148) );
  MUX U297 ( .IN0(n2290), .IN1(n149), .SEL(n2291), .F(n2245) );
  IV U298 ( .A(n2292), .Z(n149) );
  MUX U299 ( .IN0(n2382), .IN1(n150), .SEL(n2383), .F(n2350) );
  IV U300 ( .A(n2384), .Z(n150) );
  MUX U301 ( .IN0(n2428), .IN1(n151), .SEL(n2429), .F(n2404) );
  IV U302 ( .A(n2430), .Z(n151) );
  XOR U303 ( .A(n766), .B(n765), .Z(n797) );
  MUX U304 ( .IN0(n2251), .IN1(n152), .SEL(n2252), .F(n2202) );
  IV U305 ( .A(n2253), .Z(n152) );
  MUX U306 ( .IN0(n892), .IN1(n153), .SEL(n893), .F(n772) );
  IV U307 ( .A(n894), .Z(n153) );
  MUX U308 ( .IN0(n1558), .IN1(n1560), .SEL(n1559), .F(n1464) );
  XOR U309 ( .A(n1269), .B(n1268), .Z(n1366) );
  XOR U310 ( .A(n1374), .B(n1373), .Z(n1461) );
  MUX U311 ( .IN0(n1384), .IN1(n154), .SEL(n1385), .F(n1282) );
  IV U312 ( .A(n1386), .Z(n154) );
  MUX U313 ( .IN0(n1570), .IN1(n155), .SEL(n1571), .F(n1479) );
  IV U314 ( .A(n1572), .Z(n155) );
  MUX U315 ( .IN0(n1730), .IN1(n156), .SEL(n1731), .F(n1649) );
  IV U316 ( .A(n1732), .Z(n156) );
  MUX U317 ( .IN0(n1168), .IN1(n157), .SEL(n1169), .F(n1053) );
  IV U318 ( .A(n1170), .Z(n157) );
  XOR U319 ( .A(n936), .B(n935), .Z(n1041) );
  MUX U320 ( .IN0(n1879), .IN1(n158), .SEL(n1880), .F(n1806) );
  IV U321 ( .A(n1881), .Z(n158) );
  XOR U322 ( .A(n1180), .B(n1179), .Z(n1258) );
  XOR U323 ( .A(n1063), .B(n1062), .Z(n1150) );
  MUX U324 ( .IN0(n1812), .IN1(n159), .SEL(n1813), .F(n1733) );
  IV U325 ( .A(n1814), .Z(n159) );
  MUX U326 ( .IN0(n2010), .IN1(n2012), .SEL(n2011), .F(n1945) );
  XOR U327 ( .A(n832), .B(n831), .Z(n928) );
  MUX U328 ( .IN0(n1739), .IN1(n160), .SEL(n1740), .F(n1658) );
  IV U329 ( .A(n1741), .Z(n160) );
  MUX U330 ( .IN0(n1664), .IN1(n161), .SEL(n1665), .F(n1579) );
  IV U331 ( .A(n1666), .Z(n161) );
  MUX U332 ( .IN0(n1888), .IN1(n162), .SEL(n1889), .F(n1815) );
  IV U333 ( .A(n1890), .Z(n162) );
  MUX U334 ( .IN0(n2016), .IN1(n163), .SEL(n2017), .F(n1951) );
  IV U335 ( .A(n2018), .Z(n163) );
  XOR U336 ( .A(n957), .B(n956), .Z(n1034) );
  XOR U337 ( .A(n718), .B(n717), .Z(n813) );
  XOR U338 ( .A(n1301), .B(n1300), .Z(n1357) );
  MUX U339 ( .IN0(n1585), .IN1(n164), .SEL(n1586), .F(n1496) );
  IV U340 ( .A(n1587), .Z(n164) );
  MUX U341 ( .IN0(n1821), .IN1(n165), .SEL(n1822), .F(n1742) );
  IV U342 ( .A(n1823), .Z(n165) );
  MUX U343 ( .IN0(n1204), .IN1(n166), .SEL(n1205), .F(n1086) );
  IV U344 ( .A(n1206), .Z(n166) );
  MUX U345 ( .IN0(n1748), .IN1(n167), .SEL(n1749), .F(n1667) );
  IV U346 ( .A(n1750), .Z(n167) );
  MUX U347 ( .IN0(n2080), .IN1(n168), .SEL(n2081), .F(n2019) );
  IV U348 ( .A(n2082), .Z(n168) );
  XOR U349 ( .A(n853), .B(n852), .Z(n921) );
  MUX U350 ( .IN0(n2025), .IN1(n169), .SEL(n2026), .F(n1960) );
  IV U351 ( .A(n2027), .Z(n169) );
  XOR U352 ( .A(n2131), .B(n2130), .Z(n2179) );
  XOR U353 ( .A(n736), .B(n735), .Z(n807) );
  MUX U354 ( .IN0(n1213), .IN1(n170), .SEL(n1214), .F(n1098) );
  IV U355 ( .A(n1215), .Z(n170) );
  MUX U356 ( .IN0(n1413), .IN1(n171), .SEL(n1414), .F(n1313) );
  IV U357 ( .A(n1415), .Z(n171) );
  MUX U358 ( .IN0(n1594), .IN1(n172), .SEL(n1595), .F(n1505) );
  IV U359 ( .A(n1596), .Z(n172) );
  MUX U360 ( .IN0(n1754), .IN1(n173), .SEL(n1755), .F(n1673) );
  IV U361 ( .A(n1756), .Z(n173) );
  MUX U362 ( .IN0(n1966), .IN1(n174), .SEL(n1967), .F(n1897) );
  IV U363 ( .A(n1968), .Z(n174) );
  MUX U364 ( .IN0(n2341), .IN1(n2343), .SEL(n2342), .F(n2275) );
  MUX U365 ( .IN0(n978), .IN1(n175), .SEL(n979), .F(n865) );
  IV U366 ( .A(n980), .Z(n175) );
  MUX U367 ( .IN0(n1903), .IN1(n176), .SEL(n1904), .F(n1830) );
  IV U368 ( .A(n1905), .Z(n176) );
  MUX U369 ( .IN0(n2089), .IN1(n177), .SEL(n2090), .F(n2028) );
  IV U370 ( .A(n2091), .Z(n177) );
  MUX U371 ( .IN0(n2193), .IN1(n178), .SEL(n2194), .F(n2140) );
  IV U372 ( .A(n2195), .Z(n178) );
  MUX U373 ( .IN0(n2281), .IN1(n179), .SEL(n2282), .F(n2236) );
  IV U374 ( .A(n2283), .Z(n179) );
  XOR U375 ( .A(n748), .B(n747), .Z(n803) );
  MUX U376 ( .IN0(n2034), .IN1(n180), .SEL(n2035), .F(n1969) );
  IV U377 ( .A(n2036), .Z(n180) );
  MUX U378 ( .IN0(n988), .IN1(n181), .SEL(n989), .F(n874) );
  IV U379 ( .A(n990), .Z(n181) );
  MUX U380 ( .IN0(n1222), .IN1(n182), .SEL(n1223), .F(n1107) );
  IV U381 ( .A(n1224), .Z(n182) );
  MUX U382 ( .IN0(n1422), .IN1(n183), .SEL(n1423), .F(n1322) );
  IV U383 ( .A(n1424), .Z(n183) );
  MUX U384 ( .IN0(n1603), .IN1(n184), .SEL(n1604), .F(n1514) );
  IV U385 ( .A(n1605), .Z(n184) );
  MUX U386 ( .IN0(n1763), .IN1(n185), .SEL(n1764), .F(n1682) );
  IV U387 ( .A(n1765), .Z(n185) );
  MUX U388 ( .IN0(n1909), .IN1(n186), .SEL(n1910), .F(n1836) );
  IV U389 ( .A(n1911), .Z(n186) );
  MUX U390 ( .IN0(n2245), .IN1(n187), .SEL(n2246), .F(n2196) );
  IV U391 ( .A(n2247), .Z(n187) );
  MUX U392 ( .IN0(n2350), .IN1(n188), .SEL(n2351), .F(n2284) );
  IV U393 ( .A(n2352), .Z(n188) );
  MUX U394 ( .IN0(n2404), .IN1(n189), .SEL(n2405), .F(n2376) );
  IV U395 ( .A(n2406), .Z(n189) );
  MUX U396 ( .IN0(n997), .IN1(n190), .SEL(n998), .F(n883) );
  IV U397 ( .A(n999), .Z(n190) );
  MUX U398 ( .IN0(n2040), .IN1(n191), .SEL(n2041), .F(n1975) );
  IV U399 ( .A(n2042), .Z(n191) );
  MUX U400 ( .IN0(n2202), .IN1(n192), .SEL(n2203), .F(n2149) );
  IV U401 ( .A(n2204), .Z(n192) );
  MUX U402 ( .IN0(n2445), .IN1(n2447), .SEL(n2446), .F(n2425) );
  XOR U403 ( .A(n760), .B(n759), .Z(n799) );
  MUX U404 ( .IN0(n1118), .IN1(n193), .SEL(n1119), .F(n1000) );
  IV U405 ( .A(n1120), .Z(n193) );
  MUX U406 ( .IN0(n1331), .IN1(n194), .SEL(n1332), .F(n1225) );
  IV U407 ( .A(n1333), .Z(n194) );
  MUX U408 ( .IN0(n1523), .IN1(n195), .SEL(n1524), .F(n1425) );
  IV U409 ( .A(n1525), .Z(n195) );
  MUX U410 ( .IN0(n1691), .IN1(n196), .SEL(n1692), .F(n1606) );
  IV U411 ( .A(n1693), .Z(n196) );
  MUX U412 ( .IN0(n1845), .IN1(n197), .SEL(n1846), .F(n1766) );
  IV U413 ( .A(n1847), .Z(n197) );
  MUX U414 ( .IN0(n1981), .IN1(n198), .SEL(n1982), .F(n1912) );
  IV U415 ( .A(n1983), .Z(n198) );
  MUX U416 ( .IN0(n2155), .IN1(n199), .SEL(n2156), .F(n2098) );
  IV U417 ( .A(n2157), .Z(n199) );
  MUX U418 ( .IN0(n2293), .IN1(n200), .SEL(n2294), .F(n2248) );
  IV U419 ( .A(n2295), .Z(n200) );
  MUX U420 ( .IN0(n2385), .IN1(n201), .SEL(n2386), .F(n2353) );
  IV U421 ( .A(n2387), .Z(n201) );
  MUX U422 ( .IN0(n2431), .IN1(n202), .SEL(n2432), .F(n2407) );
  IV U423 ( .A(n2433), .Z(n202) );
  XOR U424 ( .A(n772), .B(n771), .Z(n795) );
  MUX U425 ( .IN0(n2256), .IN1(n203), .SEL(n2255), .F(n2205) );
  IV U426 ( .A(n2254), .Z(n203) );
  MUX U427 ( .IN0(n791), .IN1(n789), .SEL(n790), .F(n668) );
  MUX U428 ( .IN0(n1241), .IN1(n1239), .SEL(n1240), .F(n1129) );
  MUX U429 ( .IN0(n1622), .IN1(n1620), .SEL(n1621), .F(n1534) );
  MUX U430 ( .IN0(n1928), .IN1(n1926), .SEL(n1927), .F(n1856) );
  MUX U431 ( .IN0(n2168), .IN1(n2166), .SEL(n2167), .F(n2112) );
  MUX U432 ( .IN0(n381), .IN1(n2307), .SEL(n382), .F(n2304) );
  MUX U433 ( .IN0(n389), .IN1(n2319), .SEL(n390), .F(n2316) );
  MUX U434 ( .IN0(n1643), .IN1(n1645), .SEL(n1644), .F(n1558) );
  MUX U435 ( .IN0(n1564), .IN1(n204), .SEL(n1565), .F(n1471) );
  IV U436 ( .A(n1566), .Z(n204) );
  XOR U437 ( .A(n1160), .B(n1159), .Z(n1264) );
  MUX U438 ( .IN0(n1279), .IN1(n205), .SEL(n1280), .F(n1171) );
  IV U439 ( .A(n1281), .Z(n205) );
  MUX U440 ( .IN0(n1652), .IN1(n206), .SEL(n1653), .F(n1567) );
  IV U441 ( .A(n1654), .Z(n206) );
  MUX U442 ( .IN0(n1806), .IN1(n207), .SEL(n1807), .F(n1727) );
  IV U443 ( .A(n1808), .Z(n207) );
  MUX U444 ( .IN0(n1573), .IN1(n208), .SEL(n1574), .F(n1482) );
  IV U445 ( .A(n1575), .Z(n208) );
  MUX U446 ( .IN0(n1945), .IN1(n1947), .SEL(n1946), .F(n1876) );
  MUX U447 ( .IN0(n1053), .IN1(n209), .SEL(n1054), .F(n942) );
  IV U448 ( .A(n1055), .Z(n209) );
  XOR U449 ( .A(n823), .B(n822), .Z(n931) );
  XOR U450 ( .A(n1289), .B(n1288), .Z(n1360) );
  MUX U451 ( .IN0(n1736), .IN1(n210), .SEL(n1737), .F(n1655) );
  IV U452 ( .A(n1738), .Z(n210) );
  MUX U453 ( .IN0(n1882), .IN1(n211), .SEL(n1883), .F(n1809) );
  IV U454 ( .A(n1884), .Z(n211) );
  XOR U455 ( .A(n706), .B(n705), .Z(n817) );
  MUX U456 ( .IN0(n1060), .IN1(n212), .SEL(n1061), .F(n948) );
  IV U457 ( .A(n1062), .Z(n212) );
  MUX U458 ( .IN0(n1398), .IN1(n213), .SEL(n1399), .F(n1298) );
  IV U459 ( .A(n1400), .Z(n213) );
  XOR U460 ( .A(n838), .B(n837), .Z(n926) );
  MUX U461 ( .IN0(n1582), .IN1(n214), .SEL(n1583), .F(n1493) );
  IV U462 ( .A(n1584), .Z(n214) );
  MUX U463 ( .IN0(n1742), .IN1(n215), .SEL(n1743), .F(n1661) );
  IV U464 ( .A(n1744), .Z(n215) );
  MUX U465 ( .IN0(n1954), .IN1(n216), .SEL(n1955), .F(n1885) );
  IV U466 ( .A(n1956), .Z(n216) );
  MUX U467 ( .IN0(n2074), .IN1(n217), .SEL(n2075), .F(n2013) );
  IV U468 ( .A(n2076), .Z(n217) );
  MUX U469 ( .IN0(n1069), .IN1(n218), .SEL(n1070), .F(n957) );
  IV U470 ( .A(n1071), .Z(n218) );
  MUX U471 ( .IN0(n1082), .IN1(n219), .SEL(n1083), .F(n969) );
  IV U472 ( .A(n1084), .Z(n219) );
  MUX U473 ( .IN0(n1404), .IN1(n220), .SEL(n1405), .F(n1304) );
  IV U474 ( .A(n1406), .Z(n220) );
  MUX U475 ( .IN0(n1891), .IN1(n221), .SEL(n1892), .F(n1818) );
  IV U476 ( .A(n1893), .Z(n221) );
  MUX U477 ( .IN0(n2181), .IN1(n2183), .SEL(n2182), .F(n2128) );
  XOR U478 ( .A(n721), .B(n720), .Z(n812) );
  MUX U479 ( .IN0(n1588), .IN1(n222), .SEL(n1589), .F(n1499) );
  IV U480 ( .A(n1590), .Z(n222) );
  MUX U481 ( .IN0(n1824), .IN1(n223), .SEL(n1825), .F(n1745) );
  IV U482 ( .A(n1826), .Z(n223) );
  MUX U483 ( .IN0(n2022), .IN1(n224), .SEL(n2023), .F(n1957) );
  IV U484 ( .A(n2024), .Z(n224) );
  MUX U485 ( .IN0(n963), .IN1(n225), .SEL(n964), .F(n850) );
  IV U486 ( .A(n965), .Z(n225) );
  MUX U487 ( .IN0(n1313), .IN1(n226), .SEL(n1314), .F(n1207) );
  IV U488 ( .A(n1315), .Z(n226) );
  MUX U489 ( .IN0(n1505), .IN1(n227), .SEL(n1506), .F(n1407) );
  IV U490 ( .A(n1507), .Z(n227) );
  MUX U491 ( .IN0(n2187), .IN1(n228), .SEL(n2188), .F(n2134) );
  IV U492 ( .A(n2189), .Z(n228) );
  XOR U493 ( .A(n733), .B(n732), .Z(n808) );
  MUX U494 ( .IN0(n1830), .IN1(n229), .SEL(n1831), .F(n1751) );
  IV U495 ( .A(n1832), .Z(n229) );
  MUX U496 ( .IN0(n2028), .IN1(n230), .SEL(n2029), .F(n1963) );
  IV U497 ( .A(n2030), .Z(n230) );
  MUX U498 ( .IN0(n2278), .IN1(n231), .SEL(n2279), .F(n2233) );
  IV U499 ( .A(n2280), .Z(n231) );
  MUX U500 ( .IN0(n859), .IN1(n232), .SEL(n860), .F(n739) );
  IV U501 ( .A(n861), .Z(n232) );
  XOR U502 ( .A(n868), .B(n867), .Z(n916) );
  MUX U503 ( .IN0(n1216), .IN1(n233), .SEL(n1217), .F(n1101) );
  IV U504 ( .A(n1218), .Z(n233) );
  MUX U505 ( .IN0(n1416), .IN1(n234), .SEL(n1417), .F(n1316) );
  IV U506 ( .A(n1418), .Z(n234) );
  MUX U507 ( .IN0(n1597), .IN1(n235), .SEL(n1598), .F(n1508) );
  IV U508 ( .A(n1599), .Z(n235) );
  MUX U509 ( .IN0(n1757), .IN1(n236), .SEL(n1758), .F(n1676) );
  IV U510 ( .A(n1759), .Z(n236) );
  MUX U511 ( .IN0(n1969), .IN1(n237), .SEL(n1970), .F(n1900) );
  IV U512 ( .A(n1971), .Z(n237) );
  MUX U513 ( .IN0(n2239), .IN1(n238), .SEL(n2240), .F(n2190) );
  IV U514 ( .A(n2241), .Z(n238) );
  MUX U515 ( .IN0(n1906), .IN1(n239), .SEL(n1907), .F(n1833) );
  IV U516 ( .A(n1908), .Z(n239) );
  MUX U517 ( .IN0(n2092), .IN1(n240), .SEL(n2093), .F(n2031) );
  IV U518 ( .A(n2094), .Z(n240) );
  MUX U519 ( .IN0(n2401), .IN1(n2403), .SEL(n2402), .F(n2373) );
  XOR U520 ( .A(n751), .B(n750), .Z(n802) );
  MUX U521 ( .IN0(n1325), .IN1(n241), .SEL(n1326), .F(n1219) );
  IV U522 ( .A(n1327), .Z(n241) );
  MUX U523 ( .IN0(n1517), .IN1(n242), .SEL(n1518), .F(n1419) );
  IV U524 ( .A(n1519), .Z(n242) );
  MUX U525 ( .IN0(n1685), .IN1(n243), .SEL(n1686), .F(n1600) );
  IV U526 ( .A(n1687), .Z(n243) );
  MUX U527 ( .IN0(n1839), .IN1(n244), .SEL(n1840), .F(n1760) );
  IV U528 ( .A(n1841), .Z(n244) );
  XOR U529 ( .A(n2143), .B(n2142), .Z(n2175) );
  MUX U530 ( .IN0(n2287), .IN1(n245), .SEL(n2288), .F(n2242) );
  IV U531 ( .A(n2289), .Z(n245) );
  MUX U532 ( .IN0(n2379), .IN1(n246), .SEL(n2380), .F(n2347) );
  IV U533 ( .A(n2381), .Z(n246) );
  XOR U534 ( .A(n994), .B(n993), .Z(n1022) );
  MUX U535 ( .IN0(n2098), .IN1(n247), .SEL(n2099), .F(n2037) );
  IV U536 ( .A(n2100), .Z(n247) );
  MUX U537 ( .IN0(n2248), .IN1(n248), .SEL(n2249), .F(n2199) );
  IV U538 ( .A(n2250), .Z(n248) );
  XOR U539 ( .A(n763), .B(n762), .Z(n798) );
  MUX U540 ( .IN0(n1228), .IN1(n249), .SEL(n1229), .F(n1115) );
  IV U541 ( .A(n1230), .Z(n249) );
  MUX U542 ( .IN0(n1428), .IN1(n250), .SEL(n1429), .F(n1328) );
  IV U543 ( .A(n1430), .Z(n250) );
  MUX U544 ( .IN0(n1609), .IN1(n251), .SEL(n1610), .F(n1520) );
  IV U545 ( .A(n1611), .Z(n251) );
  MUX U546 ( .IN0(n1769), .IN1(n252), .SEL(n1770), .F(n1688) );
  IV U547 ( .A(n1771), .Z(n252) );
  MUX U548 ( .IN0(n1915), .IN1(n253), .SEL(n1916), .F(n1842) );
  IV U549 ( .A(n1917), .Z(n253) );
  MUX U550 ( .IN0(n2043), .IN1(n254), .SEL(n2044), .F(n1978) );
  IV U551 ( .A(n2045), .Z(n254) );
  MUX U552 ( .IN0(n2205), .IN1(n255), .SEL(n2206), .F(n2152) );
  IV U553 ( .A(n2207), .Z(n255) );
  MUX U554 ( .IN0(n2356), .IN1(n256), .SEL(n2357), .F(n2290) );
  IV U555 ( .A(n2358), .Z(n256) );
  MUX U556 ( .IN0(n2410), .IN1(n257), .SEL(n2411), .F(n2382) );
  IV U557 ( .A(n2412), .Z(n257) );
  MUX U558 ( .IN0(n2448), .IN1(n258), .SEL(n2449), .F(n2428) );
  IV U559 ( .A(n2450), .Z(n258) );
  MUX U560 ( .IN0(n889), .IN1(n259), .SEL(n890), .F(n769) );
  IV U561 ( .A(n891), .Z(n259) );
  MUX U562 ( .IN0(n1008), .IN1(n260), .SEL(n1007), .F(n892) );
  IV U563 ( .A(n1006), .Z(n260) );
  MUX U564 ( .IN0(n2160), .IN1(n261), .SEL(n2159), .F(n2101) );
  IV U565 ( .A(n2158), .Z(n261) );
  MUX U566 ( .IN0(n2298), .IN1(n262), .SEL(n2297), .F(n2251) );
  IV U567 ( .A(n2296), .Z(n262) );
  MUX U568 ( .IN0(n905), .IN1(n903), .SEL(n904), .F(n789) );
  MUX U569 ( .IN0(n1344), .IN1(n1342), .SEL(n1343), .F(n1239) );
  MUX U570 ( .IN0(n1704), .IN1(n1702), .SEL(n1703), .F(n1620) );
  MUX U571 ( .IN0(n1994), .IN1(n1992), .SEL(n1993), .F(n1926) );
  MUX U572 ( .IN0(n2218), .IN1(n2216), .SEL(n2217), .F(n2166) );
  MUX U573 ( .IN0(n383), .IN1(n2310), .SEL(n384), .F(n2307) );
  MUX U574 ( .IN0(n391), .IN1(n2322), .SEL(n392), .F(n2319) );
  MUX U575 ( .IN0(n1368), .IN1(n1370), .SEL(n1369), .F(n1266) );
  MUX U576 ( .IN0(n1724), .IN1(n1726), .SEL(n1725), .F(n1643) );
  XOR U577 ( .A(n1046), .B(n1045), .Z(n1155) );
  XOR U578 ( .A(n1381), .B(n1380), .Z(n1459) );
  XOR U579 ( .A(n1476), .B(n1475), .Z(n1554) );
  XOR U580 ( .A(n1564), .B(n1563), .Z(n1640) );
  MUX U581 ( .IN0(n1487), .IN1(n263), .SEL(n1488), .F(n1387) );
  IV U582 ( .A(n1489), .Z(n263) );
  MUX U583 ( .IN0(n1174), .IN1(n264), .SEL(n1175), .F(n1060) );
  IV U584 ( .A(n1176), .Z(n264) );
  MUX U585 ( .IN0(n1180), .IN1(n265), .SEL(n1181), .F(n1066) );
  IV U586 ( .A(n1182), .Z(n265) );
  MUX U587 ( .IN0(n942), .IN1(n266), .SEL(n943), .F(n829) );
  IV U588 ( .A(n944), .Z(n266) );
  XOR U589 ( .A(n703), .B(n702), .Z(n818) );
  XOR U590 ( .A(n951), .B(n950), .Z(n1036) );
  XOR U591 ( .A(n1294), .B(n1293), .Z(n1359) );
  MUX U592 ( .IN0(n1579), .IN1(n267), .SEL(n1580), .F(n1490) );
  IV U593 ( .A(n1581), .Z(n267) );
  XOR U594 ( .A(n1879), .B(n1878), .Z(n1943) );
  MUX U595 ( .IN0(n2071), .IN1(n2073), .SEL(n2072), .F(n2010) );
  MUX U596 ( .IN0(n1072), .IN1(n268), .SEL(n1073), .F(n960) );
  IV U597 ( .A(n1074), .Z(n268) );
  XOR U598 ( .A(n1658), .B(n1657), .Z(n1718) );
  XOR U599 ( .A(n1736), .B(n1735), .Z(n1798) );
  XOR U600 ( .A(n715), .B(n714), .Z(n814) );
  MUX U601 ( .IN0(n1307), .IN1(n269), .SEL(n1308), .F(n1199) );
  IV U602 ( .A(n1309), .Z(n269) );
  MUX U603 ( .IN0(n1499), .IN1(n270), .SEL(n1500), .F(n1401) );
  IV U604 ( .A(n1501), .Z(n270) );
  MUX U605 ( .IN0(n1667), .IN1(n271), .SEL(n1668), .F(n1582) );
  IV U606 ( .A(n1669), .Z(n271) );
  MUX U607 ( .IN0(n1078), .IN1(n272), .SEL(n1079), .F(n966) );
  IV U608 ( .A(n1080), .Z(n272) );
  XOR U609 ( .A(n844), .B(n843), .Z(n924) );
  MUX U610 ( .IN0(n1210), .IN1(n273), .SEL(n1211), .F(n1095) );
  IV U611 ( .A(n1212), .Z(n273) );
  MUX U612 ( .IN0(n1410), .IN1(n274), .SEL(n1411), .F(n1310) );
  IV U613 ( .A(n1412), .Z(n274) );
  MUX U614 ( .IN0(n1591), .IN1(n275), .SEL(n1592), .F(n1502) );
  IV U615 ( .A(n1593), .Z(n275) );
  MUX U616 ( .IN0(n1751), .IN1(n276), .SEL(n1752), .F(n1670) );
  IV U617 ( .A(n1753), .Z(n276) );
  XOR U618 ( .A(n2019), .B(n2018), .Z(n2067) );
  MUX U619 ( .IN0(n2275), .IN1(n2277), .SEL(n2276), .F(n2230) );
  XOR U620 ( .A(n730), .B(n729), .Z(n809) );
  MUX U621 ( .IN0(n463), .IN1(n277), .SEL(n464), .F(n462) );
  IV U622 ( .A(n465), .Z(n277) );
  MUX U623 ( .IN0(n972), .IN1(n278), .SEL(n973), .F(n859) );
  IV U624 ( .A(n974), .Z(n278) );
  MUX U625 ( .IN0(n1101), .IN1(n279), .SEL(n1102), .F(n985) );
  IV U626 ( .A(n1103), .Z(n279) );
  XOR U627 ( .A(n1824), .B(n1823), .Z(n1868) );
  XOR U628 ( .A(n1894), .B(n1893), .Z(n1938) );
  MUX U629 ( .IN0(n2140), .IN1(n280), .SEL(n2141), .F(n2083) );
  IV U630 ( .A(n2142), .Z(n280) );
  MUX U631 ( .IN0(n1319), .IN1(n281), .SEL(n1320), .F(n1213) );
  IV U632 ( .A(n1321), .Z(n281) );
  MUX U633 ( .IN0(n1511), .IN1(n282), .SEL(n1512), .F(n1413) );
  IV U634 ( .A(n1513), .Z(n282) );
  MUX U635 ( .IN0(n1679), .IN1(n283), .SEL(n1680), .F(n1594) );
  IV U636 ( .A(n1681), .Z(n283) );
  MUX U637 ( .IN0(n1833), .IN1(n284), .SEL(n1834), .F(n1754) );
  IV U638 ( .A(n1835), .Z(n284) );
  XOR U639 ( .A(n2187), .B(n2186), .Z(n2227) );
  MUX U640 ( .IN0(n2344), .IN1(n285), .SEL(n2345), .F(n2278) );
  IV U641 ( .A(n2346), .Z(n285) );
  XOR U642 ( .A(n745), .B(n744), .Z(n804) );
  XOR U643 ( .A(n874), .B(n873), .Z(n914) );
  MUX U644 ( .IN0(n2425), .IN1(n2427), .SEL(n2426), .F(n2401) );
  XOR U645 ( .A(n757), .B(n756), .Z(n800) );
  XOR U646 ( .A(n1972), .B(n1971), .Z(n2000) );
  XOR U647 ( .A(n2034), .B(n2033), .Z(n2062) );
  XOR U648 ( .A(n997), .B(n996), .Z(n1021) );
  XOR U649 ( .A(n1222), .B(n1221), .Z(n1246) );
  XOR U650 ( .A(n1422), .B(n1421), .Z(n1446) );
  XOR U651 ( .A(n1603), .B(n1602), .Z(n1627) );
  XOR U652 ( .A(n1763), .B(n1762), .Z(n1789) );
  XOR U653 ( .A(n1909), .B(n1908), .Z(n1933) );
  MUX U654 ( .IN0(n2101), .IN1(n286), .SEL(n2102), .F(n2040) );
  IV U655 ( .A(n2103), .Z(n286) );
  XOR U656 ( .A(n2149), .B(n2148), .Z(n2173) );
  XOR U657 ( .A(n2199), .B(n2198), .Z(n2223) );
  XOR U658 ( .A(n2287), .B(n2286), .Z(n2336) );
  XOR U659 ( .A(n2379), .B(n2378), .Z(n2398) );
  XOR U660 ( .A(n769), .B(n768), .Z(n796) );
  MUX U661 ( .IN0(n1233), .IN1(n287), .SEL(n1232), .F(n1118) );
  IV U662 ( .A(n1231), .Z(n287) );
  MUX U663 ( .IN0(n1433), .IN1(n288), .SEL(n1432), .F(n1331) );
  IV U664 ( .A(n1431), .Z(n288) );
  MUX U665 ( .IN0(n1614), .IN1(n289), .SEL(n1613), .F(n1523) );
  IV U666 ( .A(n1612), .Z(n289) );
  MUX U667 ( .IN0(n1774), .IN1(n290), .SEL(n1773), .F(n1691) );
  IV U668 ( .A(n1772), .Z(n290) );
  MUX U669 ( .IN0(n1920), .IN1(n291), .SEL(n1919), .F(n1845) );
  IV U670 ( .A(n1918), .Z(n291) );
  MUX U671 ( .IN0(n2048), .IN1(n292), .SEL(n2047), .F(n1981) );
  IV U672 ( .A(n2046), .Z(n292) );
  MUX U673 ( .IN0(n2210), .IN1(n293), .SEL(n2209), .F(n2155) );
  IV U674 ( .A(n2208), .Z(n293) );
  MUX U675 ( .IN0(n2390), .IN1(n294), .SEL(n2389), .F(n2356) );
  IV U676 ( .A(n2388), .Z(n294) );
  MUX U677 ( .IN0(n2436), .IN1(n295), .SEL(n2435), .F(n2410) );
  IV U678 ( .A(n2434), .Z(n295) );
  MUX U679 ( .IN0(n2466), .IN1(n296), .SEL(n2465), .F(n2448) );
  IV U680 ( .A(n2464), .Z(n296) );
  MUX U681 ( .IN0(n897), .IN1(n297), .SEL(n896), .F(n775) );
  IV U682 ( .A(n895), .Z(n297) );
  MUX U683 ( .IN0(n2301), .IN1(n2299), .SEL(n2300), .F(n2254) );
  MUX U684 ( .IN0(n1016), .IN1(n1014), .SEL(n1015), .F(n903) );
  MUX U685 ( .IN0(n1441), .IN1(n1439), .SEL(n1440), .F(n1342) );
  MUX U686 ( .IN0(n1784), .IN1(n1782), .SEL(n1783), .F(n1702) );
  MUX U687 ( .IN0(n2056), .IN1(n2054), .SEL(n2055), .F(n1992) );
  MUX U688 ( .IN0(n2264), .IN1(n2262), .SEL(n2263), .F(n2216) );
  MUX U689 ( .IN0(n385), .IN1(n2313), .SEL(n386), .F(n2310) );
  MUX U690 ( .IN0(n788), .IN1(n2325), .SEL(n787), .F(n2322) );
  MUX U691 ( .IN0(n1468), .IN1(n298), .SEL(n1469), .F(n1371) );
  IV U692 ( .A(n1470), .Z(n298) );
  MUX U693 ( .IN0(n1266), .IN1(n1268), .SEL(n1267), .F(n1157) );
  MUX U694 ( .IN0(n1276), .IN1(n299), .SEL(n1277), .F(n1168) );
  IV U695 ( .A(n1278), .Z(n299) );
  MUX U696 ( .IN0(n1046), .IN1(n300), .SEL(n1047), .F(n936) );
  IV U697 ( .A(n1048), .Z(n300) );
  MUX U698 ( .IN0(n1286), .IN1(n301), .SEL(n1287), .F(n1177) );
  IV U699 ( .A(n1288), .Z(n301) );
  XOR U700 ( .A(n1384), .B(n1383), .Z(n1458) );
  XOR U701 ( .A(n1479), .B(n1478), .Z(n1553) );
  XOR U702 ( .A(n1567), .B(n1566), .Z(n1639) );
  XOR U703 ( .A(n1649), .B(n1648), .Z(n1721) );
  XOR U704 ( .A(n1727), .B(n1726), .Z(n1801) );
  MUX U705 ( .IN0(n1057), .IN1(n302), .SEL(n1058), .F(n945) );
  IV U706 ( .A(n1059), .Z(n302) );
  MUX U707 ( .IN0(n820), .IN1(n822), .SEL(n821), .F(n700) );
  XOR U708 ( .A(n1066), .B(n1065), .Z(n1149) );
  MUX U709 ( .IN0(n829), .IN1(n303), .SEL(n830), .F(n709) );
  IV U710 ( .A(n831), .Z(n303) );
  MUX U711 ( .IN0(n706), .IN1(n304), .SEL(n707), .F(n491) );
  IV U712 ( .A(n708), .Z(n304) );
  MUX U713 ( .IN0(n1304), .IN1(n305), .SEL(n1305), .F(n1196) );
  IV U714 ( .A(n1306), .Z(n305) );
  XOR U715 ( .A(n1948), .B(n1947), .Z(n2008) );
  MUX U716 ( .IN0(n835), .IN1(n306), .SEL(n836), .F(n715) );
  IV U717 ( .A(n837), .Z(n306) );
  MUX U718 ( .IN0(n721), .IN1(n307), .SEL(n722), .F(n477) );
  IV U719 ( .A(n723), .Z(n307) );
  XOR U720 ( .A(n1398), .B(n1397), .Z(n1454) );
  XOR U721 ( .A(n1493), .B(n1492), .Z(n1549) );
  XOR U722 ( .A(n1579), .B(n1578), .Z(n1635) );
  XOR U723 ( .A(n1661), .B(n1660), .Z(n1717) );
  XOR U724 ( .A(n1739), .B(n1738), .Z(n1797) );
  XOR U725 ( .A(n1815), .B(n1814), .Z(n1871) );
  XOR U726 ( .A(n1885), .B(n1884), .Z(n1941) );
  MUX U727 ( .IN0(n1075), .IN1(n308), .SEL(n1076), .F(n963) );
  IV U728 ( .A(n1077), .Z(n308) );
  MUX U729 ( .IN0(n957), .IN1(n309), .SEL(n958), .F(n844) );
  IV U730 ( .A(n959), .Z(n309) );
  XOR U731 ( .A(n2016), .B(n2015), .Z(n2068) );
  MUX U732 ( .IN0(n727), .IN1(n310), .SEL(n728), .F(n524) );
  IV U733 ( .A(n729), .Z(n310) );
  MUX U734 ( .IN0(n1086), .IN1(n311), .SEL(n1087), .F(n972) );
  IV U735 ( .A(n1088), .Z(n311) );
  MUX U736 ( .IN0(n853), .IN1(n312), .SEL(n854), .F(n733) );
  IV U737 ( .A(n855), .Z(n312) );
  XOR U738 ( .A(n1960), .B(n1959), .Z(n2004) );
  XOR U739 ( .A(n865), .B(n864), .Z(n917) );
  XOR U740 ( .A(n742), .B(n741), .Z(n805) );
  MUX U741 ( .IN0(n985), .IN1(n313), .SEL(n986), .F(n871) );
  IV U742 ( .A(n987), .Z(n313) );
  XOR U743 ( .A(n1098), .B(n1097), .Z(n1140) );
  XOR U744 ( .A(n1210), .B(n1209), .Z(n1250) );
  XOR U745 ( .A(n1313), .B(n1312), .Z(n1353) );
  XOR U746 ( .A(n1410), .B(n1409), .Z(n1450) );
  XOR U747 ( .A(n1505), .B(n1504), .Z(n1545) );
  XOR U748 ( .A(n1591), .B(n1590), .Z(n1631) );
  XOR U749 ( .A(n1673), .B(n1672), .Z(n1713) );
  XOR U750 ( .A(n1751), .B(n1750), .Z(n1793) );
  XOR U751 ( .A(n1827), .B(n1826), .Z(n1867) );
  XOR U752 ( .A(n1897), .B(n1896), .Z(n1937) );
  XOR U753 ( .A(n2083), .B(n2082), .Z(n2123) );
  XOR U754 ( .A(n2233), .B(n2232), .Z(n2273) );
  MUX U755 ( .IN0(n991), .IN1(n314), .SEL(n992), .F(n877) );
  IV U756 ( .A(n993), .Z(n314) );
  XOR U757 ( .A(n2028), .B(n2027), .Z(n2064) );
  XOR U758 ( .A(n2190), .B(n2189), .Z(n2226) );
  XOR U759 ( .A(n754), .B(n753), .Z(n801) );
  XOR U760 ( .A(n886), .B(n885), .Z(n910) );
  XOR U761 ( .A(n1112), .B(n1111), .Z(n1136) );
  XOR U762 ( .A(n1325), .B(n1324), .Z(n1349) );
  XOR U763 ( .A(n1517), .B(n1516), .Z(n1541) );
  XOR U764 ( .A(n1685), .B(n1684), .Z(n1709) );
  XOR U765 ( .A(n1839), .B(n1838), .Z(n1863) );
  XOR U766 ( .A(n1975), .B(n1974), .Z(n1999) );
  XOR U767 ( .A(n2095), .B(n2094), .Z(n2119) );
  XOR U768 ( .A(n2245), .B(n2244), .Z(n2269) );
  XOR U769 ( .A(n2350), .B(n2349), .Z(n2369) );
  XOR U770 ( .A(n2404), .B(n2403), .Z(n2423) );
  MUX U771 ( .IN0(n1123), .IN1(n315), .SEL(n1122), .F(n1003) );
  IV U772 ( .A(n1121), .Z(n315) );
  MUX U773 ( .IN0(n1336), .IN1(n316), .SEL(n1335), .F(n1228) );
  IV U774 ( .A(n1334), .Z(n316) );
  MUX U775 ( .IN0(n1528), .IN1(n317), .SEL(n1527), .F(n1428) );
  IV U776 ( .A(n1526), .Z(n317) );
  MUX U777 ( .IN0(n1696), .IN1(n318), .SEL(n1695), .F(n1609) );
  IV U778 ( .A(n1694), .Z(n318) );
  MUX U779 ( .IN0(n1850), .IN1(n319), .SEL(n1849), .F(n1769) );
  IV U780 ( .A(n1848), .Z(n319) );
  MUX U781 ( .IN0(n1986), .IN1(n320), .SEL(n1985), .F(n1915) );
  IV U782 ( .A(n1984), .Z(n320) );
  MUX U783 ( .IN0(n2106), .IN1(n321), .SEL(n2105), .F(n2043) );
  IV U784 ( .A(n2104), .Z(n321) );
  XOR U785 ( .A(n2202), .B(n2201), .Z(n2222) );
  MUX U786 ( .IN0(n2361), .IN1(n322), .SEL(n2360), .F(n2293) );
  IV U787 ( .A(n2359), .Z(n322) );
  MUX U788 ( .IN0(n2415), .IN1(n323), .SEL(n2414), .F(n2385) );
  IV U789 ( .A(n2413), .Z(n323) );
  MUX U790 ( .IN0(n2453), .IN1(n324), .SEL(n2452), .F(n2431) );
  IV U791 ( .A(n2451), .Z(n324) );
  MUX U792 ( .IN0(n325), .IN1(n2473), .SEL(n2474), .F(n2461) );
  IV U793 ( .A(n2475), .Z(n325) );
  MUX U794 ( .IN0(n783), .IN1(n781), .SEL(n782), .F(n414) );
  MUX U795 ( .IN0(n772), .IN1(n326), .SEL(n773), .F(n608) );
  IV U796 ( .A(n774), .Z(n326) );
  MUX U797 ( .IN0(n1011), .IN1(n1009), .SEL(n1010), .F(n895) );
  MUX U798 ( .IN0(n2213), .IN1(n2211), .SEL(n2212), .F(n2158) );
  MUX U799 ( .IN0(n670), .IN1(n668), .SEL(n669), .F(n399) );
  MUX U800 ( .IN0(n1131), .IN1(n1129), .SEL(n1130), .F(n1014) );
  MUX U801 ( .IN0(n1536), .IN1(n1534), .SEL(n1535), .F(n1439) );
  MUX U802 ( .IN0(n1858), .IN1(n1856), .SEL(n1857), .F(n1782) );
  MUX U803 ( .IN0(n2114), .IN1(n2112), .SEL(n2113), .F(n2054) );
  MUX U804 ( .IN0(n327), .IN1(n2304), .SEL(n380), .F(n2262) );
  IV U805 ( .A(n379), .Z(n327) );
  MUX U806 ( .IN0(n387), .IN1(n2316), .SEL(n388), .F(n2313) );
  MUX U807 ( .IN0(n1781), .IN1(n2328), .SEL(n1780), .F(n2325) );
  XOR U808 ( .A(n1378), .B(n1376), .Z(n1460) );
  MUX U809 ( .IN0(n1157), .IN1(n1159), .SEL(n1158), .F(n1043) );
  XOR U810 ( .A(n1646), .B(n1645), .Z(n1722) );
  MUX U811 ( .IN0(n1876), .IN1(n1878), .SEL(n1877), .F(n1803) );
  MUX U812 ( .IN0(n1050), .IN1(n328), .SEL(n1051), .F(n939) );
  IV U813 ( .A(n1052), .Z(n328) );
  MUX U814 ( .IN0(n1171), .IN1(n329), .SEL(n1172), .F(n1057) );
  IV U815 ( .A(n1173), .Z(n329) );
  XOR U816 ( .A(n1286), .B(n1284), .Z(n1361) );
  MUX U817 ( .IN0(n936), .IN1(n330), .SEL(n937), .F(n823) );
  IV U818 ( .A(n938), .Z(n330) );
  XOR U819 ( .A(n1482), .B(n1481), .Z(n1552) );
  XOR U820 ( .A(n1730), .B(n1729), .Z(n1800) );
  MUX U821 ( .IN0(n1066), .IN1(n331), .SEL(n1067), .F(n954) );
  IV U822 ( .A(n1068), .Z(n331) );
  XOR U823 ( .A(n709), .B(n708), .Z(n816) );
  MUX U824 ( .IN0(n700), .IN1(n702), .SEL(n701), .F(n490) );
  MUX U825 ( .IN0(n948), .IN1(n332), .SEL(n949), .F(n835) );
  IV U826 ( .A(n950), .Z(n332) );
  XOR U827 ( .A(n1393), .B(n1392), .Z(n1455) );
  XOR U828 ( .A(n1576), .B(n1575), .Z(n1636) );
  XOR U829 ( .A(n1812), .B(n1811), .Z(n1872) );
  MUX U830 ( .IN0(n2128), .IN1(n2130), .SEL(n2129), .F(n2071) );
  MUX U831 ( .IN0(n1193), .IN1(n333), .SEL(n1194), .F(n1075) );
  IV U832 ( .A(n1195), .Z(n333) );
  MUX U833 ( .IN0(n960), .IN1(n334), .SEL(n961), .F(n847) );
  IV U834 ( .A(n962), .Z(n334) );
  XOR U835 ( .A(n1951), .B(n1950), .Z(n2007) );
  MUX U836 ( .IN0(n718), .IN1(n335), .SEL(n719), .F(n525) );
  IV U837 ( .A(n720), .Z(n335) );
  XOR U838 ( .A(n1086), .B(n1084), .Z(n1143) );
  XOR U839 ( .A(n1304), .B(n1303), .Z(n1356) );
  XOR U840 ( .A(n1496), .B(n1495), .Z(n1548) );
  XOR U841 ( .A(n1664), .B(n1663), .Z(n1716) );
  XOR U842 ( .A(n1888), .B(n1887), .Z(n1940) );
  MUX U843 ( .IN0(n2184), .IN1(n336), .SEL(n2185), .F(n2131) );
  IV U844 ( .A(n2186), .Z(n336) );
  MUX U845 ( .IN0(n966), .IN1(n337), .SEL(n967), .F(n853) );
  IV U846 ( .A(n968), .Z(n337) );
  MUX U847 ( .IN0(n844), .IN1(n338), .SEL(n845), .F(n724) );
  IV U848 ( .A(n846), .Z(n338) );
  XOR U849 ( .A(n1207), .B(n1206), .Z(n1251) );
  XOR U850 ( .A(n1407), .B(n1406), .Z(n1451) );
  XOR U851 ( .A(n1588), .B(n1587), .Z(n1632) );
  XOR U852 ( .A(n1748), .B(n1747), .Z(n1794) );
  XOR U853 ( .A(n2080), .B(n2079), .Z(n2124) );
  MUX U854 ( .IN0(n730), .IN1(n339), .SEL(n731), .F(n455) );
  IV U855 ( .A(n732), .Z(n339) );
  XOR U856 ( .A(n739), .B(n738), .Z(n806) );
  MUX U857 ( .IN0(n981), .IN1(n340), .SEL(n982), .F(n868) );
  IV U858 ( .A(n983), .Z(n340) );
  XOR U859 ( .A(n1963), .B(n1962), .Z(n2003) );
  XOR U860 ( .A(n2025), .B(n2024), .Z(n2065) );
  MUX U861 ( .IN0(n865), .IN1(n341), .SEL(n866), .F(n745) );
  IV U862 ( .A(n867), .Z(n341) );
  MUX U863 ( .IN0(n751), .IN1(n342), .SEL(n752), .F(n447) );
  IV U864 ( .A(n753), .Z(n342) );
  XOR U865 ( .A(n1101), .B(n1100), .Z(n1139) );
  XOR U866 ( .A(n1316), .B(n1315), .Z(n1352) );
  XOR U867 ( .A(n1508), .B(n1507), .Z(n1544) );
  XOR U868 ( .A(n1676), .B(n1675), .Z(n1712) );
  XOR U869 ( .A(n1830), .B(n1829), .Z(n1866) );
  XOR U870 ( .A(n2140), .B(n2139), .Z(n2176) );
  XOR U871 ( .A(n2236), .B(n2235), .Z(n2272) );
  MUX U872 ( .IN0(n757), .IN1(n343), .SEL(n758), .F(n580) );
  IV U873 ( .A(n759), .Z(n343) );
  XOR U874 ( .A(n1219), .B(n1218), .Z(n1247) );
  XOR U875 ( .A(n1419), .B(n1418), .Z(n1447) );
  XOR U876 ( .A(n1600), .B(n1599), .Z(n1628) );
  XOR U877 ( .A(n1760), .B(n1759), .Z(n1790) );
  XOR U878 ( .A(n1906), .B(n1905), .Z(n1934) );
  XOR U879 ( .A(n2092), .B(n2091), .Z(n2120) );
  XOR U880 ( .A(n2284), .B(n2283), .Z(n2337) );
  XOR U881 ( .A(n2376), .B(n2375), .Z(n2399) );
  MUX U882 ( .IN0(n880), .IN1(n344), .SEL(n881), .F(n760) );
  IV U883 ( .A(n882), .Z(n344) );
  MUX U884 ( .IN0(n766), .IN1(n345), .SEL(n767), .F(n431) );
  IV U885 ( .A(n768), .Z(n345) );
  XOR U886 ( .A(n2037), .B(n2036), .Z(n2061) );
  MUX U887 ( .IN0(n2461), .IN1(n2463), .SEL(n2462), .F(n2445) );
  XOR U888 ( .A(n889), .B(n888), .Z(n909) );
  XOR U889 ( .A(n1115), .B(n1114), .Z(n1135) );
  XOR U890 ( .A(n1328), .B(n1327), .Z(n1348) );
  XOR U891 ( .A(n1520), .B(n1519), .Z(n1540) );
  XOR U892 ( .A(n1688), .B(n1687), .Z(n1708) );
  XOR U893 ( .A(n1842), .B(n1841), .Z(n1862) );
  XOR U894 ( .A(n1978), .B(n1977), .Z(n1998) );
  XOR U895 ( .A(n2152), .B(n2151), .Z(n2172) );
  XOR U896 ( .A(n2248), .B(n2247), .Z(n2268) );
  XOR U897 ( .A(n2353), .B(n2352), .Z(n2368) );
  XOR U898 ( .A(n2407), .B(n2406), .Z(n2422) );
  XOR U899 ( .A(n775), .B(n774), .Z(n794) );
  MUX U900 ( .IN0(n1126), .IN1(n1124), .SEL(n1125), .F(n1006) );
  MUX U901 ( .IN0(n1339), .IN1(n1337), .SEL(n1338), .F(n1231) );
  MUX U902 ( .IN0(n1531), .IN1(n1529), .SEL(n1530), .F(n1431) );
  MUX U903 ( .IN0(n1699), .IN1(n1697), .SEL(n1698), .F(n1612) );
  MUX U904 ( .IN0(n1853), .IN1(n1851), .SEL(n1852), .F(n1772) );
  MUX U905 ( .IN0(n1989), .IN1(n1987), .SEL(n1988), .F(n1918) );
  MUX U906 ( .IN0(n2109), .IN1(n2107), .SEL(n2108), .F(n2046) );
  MUX U907 ( .IN0(n2259), .IN1(n2257), .SEL(n2258), .F(n2208) );
  MUX U908 ( .IN0(n2364), .IN1(n2362), .SEL(n2363), .F(n2296) );
  MUX U909 ( .IN0(n2418), .IN1(n2416), .SEL(n2417), .F(n2388) );
  MUX U910 ( .IN0(n2456), .IN1(n2454), .SEL(n2455), .F(n2434) );
  MUX U911 ( .IN0(n2478), .IN1(n2479), .SEL(n2477), .F(n2464) );
  XNOR U912 ( .A(n789), .B(o[28]), .Z(n790) );
  XNOR U913 ( .A(n1129), .B(o[25]), .Z(n1130) );
  XNOR U914 ( .A(n1439), .B(o[22]), .Z(n1440) );
  XNOR U915 ( .A(n1702), .B(o[19]), .Z(n1703) );
  XNOR U916 ( .A(n1926), .B(o[16]), .Z(n1927) );
  XNOR U917 ( .A(n2112), .B(o[13]), .Z(n2113) );
  XNOR U918 ( .A(n2262), .B(o[10]), .Z(n2263) );
  XNOR U919 ( .A(n2310), .B(o[7]), .Z(n384) );
  XNOR U920 ( .A(n2319), .B(o[4]), .Z(n390) );
  XOR U921 ( .A(n1468), .B(n1466), .Z(n1556) );
  MUX U922 ( .IN0(n1273), .IN1(n346), .SEL(n1274), .F(n1163) );
  IV U923 ( .A(n1275), .Z(n346) );
  MUX U924 ( .IN0(n1160), .IN1(n347), .SEL(n1161), .F(n1046) );
  IV U925 ( .A(n1162), .Z(n347) );
  XOR U926 ( .A(n1282), .B(n1281), .Z(n1362) );
  XOR U927 ( .A(n1057), .B(n1055), .Z(n1152) );
  MUX U928 ( .IN0(n933), .IN1(n935), .SEL(n934), .F(n820) );
  XOR U929 ( .A(n1387), .B(n1386), .Z(n1457) );
  XOR U930 ( .A(n1570), .B(n1569), .Z(n1638) );
  XOR U931 ( .A(n1652), .B(n1651), .Z(n1720) );
  XOR U932 ( .A(n1806), .B(n1805), .Z(n1874) );
  XOR U933 ( .A(n948), .B(n947), .Z(n1037) );
  MUX U934 ( .IN0(n703), .IN1(n348), .SEL(n704), .F(n489) );
  IV U935 ( .A(n705), .Z(n348) );
  XOR U936 ( .A(n1069), .B(n1068), .Z(n1148) );
  XOR U937 ( .A(n1298), .B(n1296), .Z(n1358) );
  XOR U938 ( .A(n1490), .B(n1489), .Z(n1550) );
  XOR U939 ( .A(n1882), .B(n1881), .Z(n1942) );
  MUX U940 ( .IN0(n712), .IN1(n349), .SEL(n713), .F(n499) );
  IV U941 ( .A(n714), .Z(n349) );
  XOR U942 ( .A(n841), .B(n840), .Z(n925) );
  XOR U943 ( .A(n966), .B(n965), .Z(n1031) );
  XOR U944 ( .A(n1199), .B(n1198), .Z(n1253) );
  XOR U945 ( .A(n1401), .B(n1400), .Z(n1453) );
  XOR U946 ( .A(n1582), .B(n1581), .Z(n1634) );
  XOR U947 ( .A(n1742), .B(n1741), .Z(n1796) );
  XOR U948 ( .A(n1818), .B(n1817), .Z(n1870) );
  XOR U949 ( .A(n1954), .B(n1953), .Z(n2006) );
  XOR U950 ( .A(n2074), .B(n2073), .Z(n2126) );
  XOR U951 ( .A(n724), .B(n723), .Z(n811) );
  MUX U952 ( .IN0(n850), .IN1(n350), .SEL(n851), .F(n730) );
  IV U953 ( .A(n852), .Z(n350) );
  MUX U954 ( .IN0(n736), .IN1(n351), .SEL(n737), .F(n463) );
  IV U955 ( .A(n738), .Z(n351) );
  XOR U956 ( .A(n859), .B(n858), .Z(n919) );
  XOR U957 ( .A(n1095), .B(n1094), .Z(n1141) );
  XOR U958 ( .A(n1310), .B(n1309), .Z(n1354) );
  XOR U959 ( .A(n1502), .B(n1501), .Z(n1546) );
  XOR U960 ( .A(n1670), .B(n1669), .Z(n1714) );
  XOR U961 ( .A(n2022), .B(n2021), .Z(n2066) );
  XOR U962 ( .A(n2134), .B(n2133), .Z(n2178) );
  XOR U963 ( .A(n985), .B(n983), .Z(n1025) );
  MUX U964 ( .IN0(n742), .IN1(n352), .SEL(n743), .F(n552) );
  IV U965 ( .A(n744), .Z(n352) );
  XOR U966 ( .A(n1213), .B(n1212), .Z(n1249) );
  XOR U967 ( .A(n1413), .B(n1412), .Z(n1449) );
  XOR U968 ( .A(n1594), .B(n1593), .Z(n1630) );
  XOR U969 ( .A(n1754), .B(n1753), .Z(n1792) );
  XOR U970 ( .A(n1900), .B(n1899), .Z(n1936) );
  XOR U971 ( .A(n1966), .B(n1965), .Z(n2002) );
  XOR U972 ( .A(n2086), .B(n2085), .Z(n2122) );
  XOR U973 ( .A(n2278), .B(n2277), .Z(n2339) );
  MUX U974 ( .IN0(n748), .IN1(n353), .SEL(n749), .F(n581) );
  IV U975 ( .A(n750), .Z(n353) );
  XOR U976 ( .A(n2193), .B(n2192), .Z(n2225) );
  XOR U977 ( .A(n2239), .B(n2238), .Z(n2271) );
  MUX U978 ( .IN0(n874), .IN1(n354), .SEL(n875), .F(n754) );
  IV U979 ( .A(n876), .Z(n354) );
  XOR U980 ( .A(n1107), .B(n1106), .Z(n1137) );
  XOR U981 ( .A(n1322), .B(n1321), .Z(n1350) );
  XOR U982 ( .A(n1514), .B(n1513), .Z(n1542) );
  XOR U983 ( .A(n1682), .B(n1681), .Z(n1710) );
  XOR U984 ( .A(n1836), .B(n1835), .Z(n1864) );
  XOR U985 ( .A(n2146), .B(n2145), .Z(n2174) );
  XOR U986 ( .A(n2347), .B(n2346), .Z(n2370) );
  MUX U987 ( .IN0(n883), .IN1(n355), .SEL(n884), .F(n763) );
  IV U988 ( .A(n885), .Z(n355) );
  MUX U989 ( .IN0(n431), .IN1(n356), .SEL(n432), .F(n430) );
  IV U990 ( .A(n433), .Z(n356) );
  MUX U991 ( .IN0(n760), .IN1(n357), .SEL(n761), .F(n423) );
  IV U992 ( .A(n762), .Z(n357) );
  XOR U993 ( .A(n1000), .B(n999), .Z(n1020) );
  XOR U994 ( .A(n1225), .B(n1224), .Z(n1245) );
  XOR U995 ( .A(n1425), .B(n1424), .Z(n1445) );
  XOR U996 ( .A(n1606), .B(n1605), .Z(n1626) );
  XOR U997 ( .A(n1766), .B(n1765), .Z(n1788) );
  XOR U998 ( .A(n1912), .B(n1911), .Z(n1932) );
  XOR U999 ( .A(n2040), .B(n2039), .Z(n2060) );
  XOR U1000 ( .A(n2098), .B(n2097), .Z(n2118) );
  XOR U1001 ( .A(n2290), .B(n2289), .Z(n2335) );
  XOR U1002 ( .A(n2382), .B(n2381), .Z(n2397) );
  XOR U1003 ( .A(n2428), .B(n2427), .Z(n2443) );
  MUX U1004 ( .IN0(n769), .IN1(n358), .SEL(n770), .F(n623) );
  IV U1005 ( .A(n771), .Z(n358) );
  MUX U1006 ( .IN0(n900), .IN1(n898), .SEL(n899), .F(n778) );
  MUX U1007 ( .IN0(n1236), .IN1(n1234), .SEL(n1235), .F(n1121) );
  MUX U1008 ( .IN0(n1436), .IN1(n1434), .SEL(n1435), .F(n1334) );
  MUX U1009 ( .IN0(n1617), .IN1(n1615), .SEL(n1616), .F(n1526) );
  MUX U1010 ( .IN0(n1777), .IN1(n1775), .SEL(n1776), .F(n1694) );
  MUX U1011 ( .IN0(n1923), .IN1(n1921), .SEL(n1922), .F(n1848) );
  MUX U1012 ( .IN0(n2051), .IN1(n2049), .SEL(n2050), .F(n1984) );
  MUX U1013 ( .IN0(n2163), .IN1(n2161), .SEL(n2162), .F(n2104) );
  XOR U1014 ( .A(n2205), .B(n2204), .Z(n2221) );
  XOR U1015 ( .A(n2251), .B(n2250), .Z(n2267) );
  MUX U1016 ( .IN0(n2393), .IN1(n2391), .SEL(n2392), .F(n2359) );
  MUX U1017 ( .IN0(n2439), .IN1(n2437), .SEL(n2438), .F(n2413) );
  MUX U1018 ( .IN0(n2469), .IN1(n2467), .SEL(n2468), .F(n2451) );
  MUX U1019 ( .IN0(n775), .IN1(n359), .SEL(n776), .F(n405) );
  IV U1020 ( .A(n777), .Z(n359) );
  XNOR U1021 ( .A(n2486), .B(n2483), .Z(n2485) );
  XNOR U1022 ( .A(n903), .B(o[27]), .Z(n904) );
  XNOR U1023 ( .A(n1239), .B(o[24]), .Z(n1240) );
  XNOR U1024 ( .A(n1534), .B(o[21]), .Z(n1535) );
  XNOR U1025 ( .A(n1782), .B(o[18]), .Z(n1783) );
  XNOR U1026 ( .A(n1992), .B(o[15]), .Z(n1993) );
  XNOR U1027 ( .A(n2166), .B(o[12]), .Z(n2167) );
  XNOR U1028 ( .A(n2304), .B(o[9]), .Z(n380) );
  XNOR U1029 ( .A(n2313), .B(o[6]), .Z(n386) );
  XNOR U1030 ( .A(n2322), .B(o[3]), .Z(n392) );
  XOR U1031 ( .A(n1279), .B(n1278), .Z(n1363) );
  XOR U1032 ( .A(n1471), .B(n1470), .Z(n1555) );
  XOR U1033 ( .A(n1561), .B(n1560), .Z(n1641) );
  XOR U1034 ( .A(n1168), .B(n1167), .Z(n1262) );
  MUX U1035 ( .IN0(n1043), .IN1(n1045), .SEL(n1044), .F(n933) );
  MUX U1036 ( .IN0(n939), .IN1(n360), .SEL(n940), .F(n826) );
  IV U1037 ( .A(n941), .Z(n360) );
  XOR U1038 ( .A(n1060), .B(n1059), .Z(n1151) );
  MUX U1039 ( .IN0(n1298), .IN1(n361), .SEL(n1299), .F(n1187) );
  IV U1040 ( .A(n1300), .Z(n361) );
  MUX U1041 ( .IN0(n823), .IN1(n362), .SEL(n824), .F(n703) );
  IV U1042 ( .A(n825), .Z(n362) );
  MUX U1043 ( .IN0(n945), .IN1(n363), .SEL(n946), .F(n832) );
  IV U1044 ( .A(n947), .Z(n363) );
  XOR U1045 ( .A(n1390), .B(n1389), .Z(n1456) );
  XOR U1046 ( .A(n1487), .B(n1486), .Z(n1551) );
  XOR U1047 ( .A(n1573), .B(n1572), .Z(n1637) );
  XOR U1048 ( .A(n1655), .B(n1654), .Z(n1719) );
  XOR U1049 ( .A(n1733), .B(n1732), .Z(n1799) );
  XOR U1050 ( .A(n1809), .B(n1808), .Z(n1873) );
  MUX U1051 ( .IN0(n1183), .IN1(n364), .SEL(n1184), .F(n1069) );
  IV U1052 ( .A(n1185), .Z(n364) );
  MUX U1053 ( .IN0(n954), .IN1(n365), .SEL(n955), .F(n841) );
  IV U1054 ( .A(n956), .Z(n365) );
  XOR U1055 ( .A(n1078), .B(n1077), .Z(n1145) );
  MUX U1056 ( .IN0(n709), .IN1(n366), .SEL(n710), .F(n481) );
  IV U1057 ( .A(n711), .Z(n366) );
  MUX U1058 ( .IN0(n838), .IN1(n367), .SEL(n839), .F(n718) );
  IV U1059 ( .A(n840), .Z(n367) );
  XOR U1060 ( .A(n2013), .B(n2012), .Z(n2069) );
  XOR U1061 ( .A(n963), .B(n962), .Z(n1032) );
  MUX U1062 ( .IN0(n715), .IN1(n368), .SEL(n716), .F(n470) );
  IV U1063 ( .A(n717), .Z(n368) );
  MUX U1064 ( .IN0(n847), .IN1(n369), .SEL(n848), .F(n727) );
  IV U1065 ( .A(n849), .Z(n369) );
  XOR U1066 ( .A(n856), .B(n855), .Z(n920) );
  XOR U1067 ( .A(n1204), .B(n1203), .Z(n1252) );
  XOR U1068 ( .A(n1307), .B(n1306), .Z(n1355) );
  XOR U1069 ( .A(n1404), .B(n1403), .Z(n1452) );
  XOR U1070 ( .A(n1499), .B(n1498), .Z(n1547) );
  XOR U1071 ( .A(n1585), .B(n1584), .Z(n1633) );
  XOR U1072 ( .A(n1667), .B(n1666), .Z(n1715) );
  XOR U1073 ( .A(n1745), .B(n1744), .Z(n1795) );
  XOR U1074 ( .A(n1821), .B(n1820), .Z(n1869) );
  XOR U1075 ( .A(n1891), .B(n1890), .Z(n1939) );
  XOR U1076 ( .A(n1957), .B(n1956), .Z(n2005) );
  XOR U1077 ( .A(n2077), .B(n2076), .Z(n2125) );
  MUX U1078 ( .IN0(n724), .IN1(n370), .SEL(n725), .F(n539) );
  IV U1079 ( .A(n726), .Z(n370) );
  MUX U1080 ( .IN0(n975), .IN1(n371), .SEL(n976), .F(n862) );
  IV U1081 ( .A(n977), .Z(n371) );
  XOR U1082 ( .A(n2184), .B(n2183), .Z(n2228) );
  MUX U1083 ( .IN0(n733), .IN1(n372), .SEL(n734), .F(n553) );
  IV U1084 ( .A(n735), .Z(n372) );
  XOR U1085 ( .A(n2137), .B(n2136), .Z(n2177) );
  MUX U1086 ( .IN0(n739), .IN1(n373), .SEL(n740), .F(n567) );
  IV U1087 ( .A(n741), .Z(n373) );
  MUX U1088 ( .IN0(n868), .IN1(n374), .SEL(n869), .F(n748) );
  IV U1089 ( .A(n870), .Z(n374) );
  MUX U1090 ( .IN0(n745), .IN1(n375), .SEL(n746), .F(n438) );
  IV U1091 ( .A(n747), .Z(n375) );
  XOR U1092 ( .A(n991), .B(n990), .Z(n1023) );
  XOR U1093 ( .A(n1104), .B(n1103), .Z(n1138) );
  XOR U1094 ( .A(n1216), .B(n1215), .Z(n1248) );
  XOR U1095 ( .A(n1319), .B(n1318), .Z(n1351) );
  XOR U1096 ( .A(n1416), .B(n1415), .Z(n1448) );
  XOR U1097 ( .A(n1511), .B(n1510), .Z(n1543) );
  XOR U1098 ( .A(n1597), .B(n1596), .Z(n1629) );
  XOR U1099 ( .A(n1679), .B(n1678), .Z(n1711) );
  XOR U1100 ( .A(n1757), .B(n1756), .Z(n1791) );
  XOR U1101 ( .A(n1833), .B(n1832), .Z(n1865) );
  XOR U1102 ( .A(n1903), .B(n1902), .Z(n1935) );
  XOR U1103 ( .A(n1969), .B(n1968), .Z(n2001) );
  XOR U1104 ( .A(n2031), .B(n2030), .Z(n2063) );
  XOR U1105 ( .A(n2089), .B(n2088), .Z(n2121) );
  XOR U1106 ( .A(n2281), .B(n2280), .Z(n2338) );
  XOR U1107 ( .A(n2344), .B(n2343), .Z(n2371) );
  XOR U1108 ( .A(n880), .B(n879), .Z(n912) );
  XOR U1109 ( .A(n2196), .B(n2195), .Z(n2224) );
  XOR U1110 ( .A(n2242), .B(n2241), .Z(n2270) );
  MUX U1111 ( .IN0(n754), .IN1(n376), .SEL(n755), .F(n595) );
  IV U1112 ( .A(n756), .Z(n376) );
  MUX U1113 ( .IN0(n763), .IN1(n377), .SEL(n764), .F(n609) );
  IV U1114 ( .A(n765), .Z(n377) );
  XOR U1115 ( .A(n892), .B(n891), .Z(n908) );
  XOR U1116 ( .A(n1003), .B(n1002), .Z(n1019) );
  XOR U1117 ( .A(n1118), .B(n1117), .Z(n1134) );
  XOR U1118 ( .A(n1228), .B(n1227), .Z(n1244) );
  XOR U1119 ( .A(n1331), .B(n1330), .Z(n1347) );
  XOR U1120 ( .A(n1428), .B(n1427), .Z(n1444) );
  XOR U1121 ( .A(n1523), .B(n1522), .Z(n1539) );
  XOR U1122 ( .A(n1609), .B(n1608), .Z(n1625) );
  XOR U1123 ( .A(n1691), .B(n1690), .Z(n1707) );
  XOR U1124 ( .A(n1769), .B(n1768), .Z(n1787) );
  XOR U1125 ( .A(n1845), .B(n1844), .Z(n1861) );
  XOR U1126 ( .A(n1915), .B(n1914), .Z(n1931) );
  XOR U1127 ( .A(n1981), .B(n1980), .Z(n1997) );
  XOR U1128 ( .A(n2043), .B(n2042), .Z(n2059) );
  XOR U1129 ( .A(n2101), .B(n2100), .Z(n2117) );
  XOR U1130 ( .A(n2155), .B(n2154), .Z(n2171) );
  XOR U1131 ( .A(n2293), .B(n2292), .Z(n2334) );
  XOR U1132 ( .A(n2356), .B(n2355), .Z(n2367) );
  XOR U1133 ( .A(n2385), .B(n2384), .Z(n2396) );
  XOR U1134 ( .A(n2410), .B(n2409), .Z(n2421) );
  XOR U1135 ( .A(n2431), .B(n2430), .Z(n2442) );
  XOR U1136 ( .A(n2448), .B(n2447), .Z(n2459) );
  MUX U1137 ( .IN0(n378), .IN1(n778), .SEL(n779), .F(n637) );
  IV U1138 ( .A(n780), .Z(n378) );
  AND U1139 ( .A(e_input[2]), .B(g_input[9]), .Z(n2256) );
  AND U1140 ( .A(e_input[2]), .B(g_input[8]), .Z(n2298) );
  XNOR U1141 ( .A(n2485), .B(n2484), .Z(n2326) );
  XNOR U1142 ( .A(n668), .B(o[29]), .Z(n669) );
  XNOR U1143 ( .A(n1014), .B(o[26]), .Z(n1015) );
  XNOR U1144 ( .A(n1342), .B(o[23]), .Z(n1343) );
  XNOR U1145 ( .A(n1620), .B(o[20]), .Z(n1621) );
  XNOR U1146 ( .A(n1856), .B(o[17]), .Z(n1857) );
  XNOR U1147 ( .A(n2054), .B(o[14]), .Z(n2055) );
  XNOR U1148 ( .A(n2216), .B(o[11]), .Z(n2217) );
  XNOR U1149 ( .A(n2307), .B(o[8]), .Z(n382) );
  XNOR U1150 ( .A(n2316), .B(o[5]), .Z(n388) );
  XNOR U1151 ( .A(n2325), .B(o[2]), .Z(n787) );
  XOR U1152 ( .A(n379), .B(n380), .Z(oi[9]) );
  XNOR U1153 ( .A(n381), .B(n382), .Z(oi[8]) );
  XNOR U1154 ( .A(n383), .B(n384), .Z(oi[7]) );
  XNOR U1155 ( .A(n385), .B(n386), .Z(oi[6]) );
  XNOR U1156 ( .A(n387), .B(n388), .Z(oi[5]) );
  XNOR U1157 ( .A(n389), .B(n390), .Z(oi[4]) );
  XNOR U1158 ( .A(n391), .B(n392), .Z(oi[3]) );
  XOR U1159 ( .A(n393), .B(n394), .Z(oi[31]) );
  XOR U1160 ( .A(n395), .B(n396), .Z(n394) );
  XOR U1161 ( .A(n397), .B(n398), .Z(n396) );
  XOR U1162 ( .A(n399), .B(n400), .Z(n398) );
  XOR U1163 ( .A(n401), .B(n402), .Z(n400) );
  XOR U1164 ( .A(n403), .B(n404), .Z(n402) );
  XOR U1165 ( .A(n405), .B(n406), .Z(n404) );
  XOR U1166 ( .A(n407), .B(n408), .Z(n406) );
  XOR U1167 ( .A(n409), .B(n410), .Z(n408) );
  XOR U1168 ( .A(n411), .B(n412), .Z(n410) );
  XNOR U1169 ( .A(n413), .B(n414), .Z(n412) );
  ANDN U1170 ( .A(n415), .B(n416), .Z(n413) );
  XOR U1171 ( .A(n417), .B(n418), .Z(n415) );
  XOR U1172 ( .A(n419), .B(n420), .Z(n411) );
  XOR U1173 ( .A(n421), .B(n422), .Z(n420) );
  XOR U1174 ( .A(n423), .B(n424), .Z(n422) );
  XOR U1175 ( .A(n425), .B(n426), .Z(n424) );
  XOR U1176 ( .A(n427), .B(n428), .Z(n426) );
  XOR U1177 ( .A(n429), .B(n430), .Z(n428) );
  XOR U1178 ( .A(n434), .B(n435), .Z(n429) );
  XOR U1179 ( .A(n436), .B(n437), .Z(n435) );
  XOR U1180 ( .A(n438), .B(n439), .Z(n437) );
  XOR U1181 ( .A(n440), .B(n441), .Z(n439) );
  XOR U1182 ( .A(n442), .B(n443), .Z(n441) );
  XOR U1183 ( .A(n444), .B(n445), .Z(n443) );
  XOR U1184 ( .A(n446), .B(n447), .Z(n445) );
  AND U1185 ( .A(n448), .B(n449), .Z(n446) );
  XNOR U1186 ( .A(n450), .B(n447), .Z(n449) );
  XOR U1187 ( .A(n451), .B(n452), .Z(n444) );
  XOR U1188 ( .A(n453), .B(n454), .Z(n452) );
  XOR U1189 ( .A(n455), .B(n456), .Z(n454) );
  XOR U1190 ( .A(n457), .B(n458), .Z(n456) );
  XOR U1191 ( .A(n459), .B(n460), .Z(n458) );
  XOR U1192 ( .A(n461), .B(n462), .Z(n460) );
  XOR U1193 ( .A(n466), .B(n467), .Z(n461) );
  XOR U1194 ( .A(n468), .B(n469), .Z(n467) );
  XOR U1195 ( .A(n470), .B(n471), .Z(n469) );
  XOR U1196 ( .A(n472), .B(n473), .Z(n471) );
  XOR U1197 ( .A(n474), .B(n475), .Z(n473) );
  XOR U1198 ( .A(n476), .B(n477), .Z(n475) );
  AND U1199 ( .A(n478), .B(n479), .Z(n476) );
  XNOR U1200 ( .A(n480), .B(n481), .Z(n479) );
  XOR U1201 ( .A(n482), .B(n483), .Z(n474) );
  XOR U1202 ( .A(n484), .B(n485), .Z(n483) );
  XOR U1203 ( .A(n481), .B(n486), .Z(n485) );
  XOR U1204 ( .A(n487), .B(n488), .Z(n486) );
  XOR U1205 ( .A(n489), .B(n490), .Z(n488) );
  XOR U1206 ( .A(n491), .B(n492), .Z(n487) );
  XOR U1207 ( .A(n493), .B(n494), .Z(n492) );
  AND U1208 ( .A(e_input[31]), .B(g_input[0]), .Z(n494) );
  AND U1209 ( .A(n495), .B(n496), .Z(n493) );
  XNOR U1210 ( .A(n497), .B(n491), .Z(n496) );
  XOR U1211 ( .A(n498), .B(n499), .Z(n484) );
  AND U1212 ( .A(n500), .B(n501), .Z(n498) );
  XOR U1213 ( .A(n490), .B(n502), .Z(n501) );
  XOR U1214 ( .A(n503), .B(n504), .Z(n482) );
  XOR U1215 ( .A(n505), .B(n506), .Z(n504) );
  AND U1216 ( .A(e_input[30]), .B(g_input[1]), .Z(n506) );
  AND U1217 ( .A(n507), .B(n508), .Z(n505) );
  XNOR U1218 ( .A(n509), .B(n489), .Z(n508) );
  XOR U1219 ( .A(n510), .B(n511), .Z(n503) );
  AND U1220 ( .A(g_input[2]), .B(e_input[29]), .Z(n511) );
  AND U1221 ( .A(g_input[3]), .B(e_input[28]), .Z(n510) );
  XOR U1222 ( .A(n512), .B(n513), .Z(n472) );
  XOR U1223 ( .A(n514), .B(n515), .Z(n513) );
  AND U1224 ( .A(g_input[4]), .B(e_input[27]), .Z(n515) );
  AND U1225 ( .A(n516), .B(n517), .Z(n514) );
  XNOR U1226 ( .A(n518), .B(n499), .Z(n517) );
  XOR U1227 ( .A(n519), .B(n520), .Z(n512) );
  AND U1228 ( .A(g_input[5]), .B(e_input[26]), .Z(n520) );
  AND U1229 ( .A(n521), .B(n522), .Z(n519) );
  XNOR U1230 ( .A(n523), .B(n477), .Z(n522) );
  XOR U1231 ( .A(n524), .B(n525), .Z(n468) );
  XOR U1232 ( .A(n526), .B(n527), .Z(n466) );
  XOR U1233 ( .A(n528), .B(n529), .Z(n527) );
  AND U1234 ( .A(n530), .B(n531), .Z(n529) );
  XNOR U1235 ( .A(n532), .B(n470), .Z(n531) );
  AND U1236 ( .A(g_input[6]), .B(e_input[25]), .Z(n528) );
  XOR U1237 ( .A(n533), .B(n534), .Z(n526) );
  AND U1238 ( .A(n535), .B(n536), .Z(n534) );
  XNOR U1239 ( .A(n537), .B(n525), .Z(n536) );
  AND U1240 ( .A(g_input[7]), .B(e_input[24]), .Z(n533) );
  XOR U1241 ( .A(n538), .B(n539), .Z(n459) );
  AND U1242 ( .A(e_input[23]), .B(g_input[8]), .Z(n538) );
  XOR U1243 ( .A(n540), .B(n541), .Z(n457) );
  XOR U1244 ( .A(n542), .B(n543), .Z(n541) );
  AND U1245 ( .A(n544), .B(n545), .Z(n543) );
  XNOR U1246 ( .A(n546), .B(n539), .Z(n545) );
  AND U1247 ( .A(e_input[22]), .B(g_input[9]), .Z(n542) );
  XOR U1248 ( .A(n547), .B(n548), .Z(n540) );
  AND U1249 ( .A(n549), .B(n550), .Z(n548) );
  XNOR U1250 ( .A(n551), .B(n524), .Z(n550) );
  AND U1251 ( .A(g_input[10]), .B(e_input[21]), .Z(n547) );
  XOR U1252 ( .A(n552), .B(n553), .Z(n453) );
  XOR U1253 ( .A(n554), .B(n555), .Z(n451) );
  XOR U1254 ( .A(n556), .B(n557), .Z(n555) );
  AND U1255 ( .A(n558), .B(n559), .Z(n557) );
  XNOR U1256 ( .A(n560), .B(n455), .Z(n559) );
  AND U1257 ( .A(g_input[11]), .B(e_input[20]), .Z(n556) );
  XOR U1258 ( .A(n561), .B(n562), .Z(n554) );
  AND U1259 ( .A(n563), .B(n564), .Z(n562) );
  XNOR U1260 ( .A(n565), .B(n553), .Z(n564) );
  AND U1261 ( .A(g_input[12]), .B(e_input[19]), .Z(n561) );
  XOR U1262 ( .A(n566), .B(n567), .Z(n442) );
  AND U1263 ( .A(g_input[13]), .B(e_input[18]), .Z(n566) );
  XOR U1264 ( .A(n568), .B(n569), .Z(n440) );
  XOR U1265 ( .A(n570), .B(n571), .Z(n569) );
  AND U1266 ( .A(n572), .B(n573), .Z(n571) );
  XNOR U1267 ( .A(n574), .B(n567), .Z(n573) );
  AND U1268 ( .A(g_input[14]), .B(e_input[17]), .Z(n570) );
  XOR U1269 ( .A(n575), .B(n576), .Z(n568) );
  AND U1270 ( .A(n577), .B(n578), .Z(n576) );
  XNOR U1271 ( .A(n579), .B(n552), .Z(n578) );
  AND U1272 ( .A(g_input[15]), .B(e_input[16]), .Z(n575) );
  XOR U1273 ( .A(n580), .B(n581), .Z(n436) );
  XOR U1274 ( .A(n582), .B(n583), .Z(n434) );
  XOR U1275 ( .A(n584), .B(n585), .Z(n583) );
  AND U1276 ( .A(n586), .B(n587), .Z(n585) );
  XNOR U1277 ( .A(n588), .B(n438), .Z(n587) );
  AND U1278 ( .A(e_input[15]), .B(g_input[16]), .Z(n584) );
  XOR U1279 ( .A(n589), .B(n590), .Z(n582) );
  AND U1280 ( .A(n591), .B(n592), .Z(n590) );
  XNOR U1281 ( .A(n593), .B(n581), .Z(n592) );
  AND U1282 ( .A(e_input[14]), .B(g_input[17]), .Z(n589) );
  XOR U1283 ( .A(n594), .B(n595), .Z(n427) );
  AND U1284 ( .A(e_input[13]), .B(g_input[18]), .Z(n594) );
  XOR U1285 ( .A(n596), .B(n597), .Z(n425) );
  XOR U1286 ( .A(n598), .B(n599), .Z(n597) );
  AND U1287 ( .A(n600), .B(n601), .Z(n599) );
  XNOR U1288 ( .A(n602), .B(n595), .Z(n601) );
  AND U1289 ( .A(e_input[12]), .B(g_input[19]), .Z(n598) );
  XOR U1290 ( .A(n603), .B(n604), .Z(n596) );
  AND U1291 ( .A(n605), .B(n606), .Z(n604) );
  XNOR U1292 ( .A(n607), .B(n580), .Z(n606) );
  AND U1293 ( .A(e_input[11]), .B(g_input[20]), .Z(n603) );
  XOR U1294 ( .A(n608), .B(n609), .Z(n421) );
  XOR U1295 ( .A(n610), .B(n611), .Z(n419) );
  XOR U1296 ( .A(n612), .B(n613), .Z(n611) );
  AND U1297 ( .A(n614), .B(n615), .Z(n613) );
  XNOR U1298 ( .A(n616), .B(n423), .Z(n615) );
  AND U1299 ( .A(e_input[10]), .B(g_input[21]), .Z(n612) );
  XOR U1300 ( .A(n617), .B(n618), .Z(n610) );
  AND U1301 ( .A(n619), .B(n620), .Z(n618) );
  XNOR U1302 ( .A(n621), .B(n609), .Z(n620) );
  AND U1303 ( .A(e_input[9]), .B(g_input[22]), .Z(n617) );
  XOR U1304 ( .A(n622), .B(n623), .Z(n409) );
  AND U1305 ( .A(e_input[8]), .B(g_input[23]), .Z(n622) );
  XOR U1306 ( .A(n624), .B(n625), .Z(n407) );
  XOR U1307 ( .A(n626), .B(n627), .Z(n625) );
  AND U1308 ( .A(n628), .B(n629), .Z(n627) );
  XNOR U1309 ( .A(n630), .B(n623), .Z(n629) );
  AND U1310 ( .A(e_input[7]), .B(g_input[24]), .Z(n626) );
  XOR U1311 ( .A(n631), .B(n632), .Z(n624) );
  AND U1312 ( .A(n633), .B(n634), .Z(n632) );
  XNOR U1313 ( .A(n635), .B(n608), .Z(n634) );
  AND U1314 ( .A(e_input[6]), .B(g_input[25]), .Z(n631) );
  XNOR U1315 ( .A(n636), .B(n637), .Z(n403) );
  AND U1316 ( .A(n638), .B(n639), .Z(n636) );
  XNOR U1317 ( .A(n640), .B(n405), .Z(n639) );
  XOR U1318 ( .A(n641), .B(n642), .Z(n401) );
  XOR U1319 ( .A(n643), .B(n644), .Z(n642) );
  AND U1320 ( .A(e_input[5]), .B(g_input[26]), .Z(n644) );
  AND U1321 ( .A(n645), .B(n646), .Z(n643) );
  XNOR U1322 ( .A(n647), .B(n648), .Z(n646) );
  XOR U1323 ( .A(n649), .B(n650), .Z(n641) );
  AND U1324 ( .A(e_input[4]), .B(g_input[27]), .Z(n650) );
  AND U1325 ( .A(e_input[3]), .B(g_input[28]), .Z(n649) );
  XOR U1326 ( .A(n651), .B(n652), .Z(n397) );
  ANDN U1327 ( .A(n653), .B(n654), .Z(n652) );
  XOR U1328 ( .A(n655), .B(n656), .Z(n653) );
  AND U1329 ( .A(g_input[29]), .B(e_input[2]), .Z(n651) );
  XOR U1330 ( .A(n657), .B(n658), .Z(n395) );
  XOR U1331 ( .A(n659), .B(n660), .Z(n658) );
  NOR U1332 ( .A(n661), .B(n662), .Z(n660) );
  AND U1333 ( .A(e_input[1]), .B(g_input[30]), .Z(n659) );
  XNOR U1334 ( .A(n656), .B(n663), .Z(n657) );
  AND U1335 ( .A(g_input[31]), .B(e_input[0]), .Z(n663) );
  XOR U1336 ( .A(n664), .B(o[31]), .Z(n393) );
  NANDN U1337 ( .B(n665), .A(n666), .Z(n664) );
  XNOR U1338 ( .A(n667), .B(n399), .Z(n666) );
  XOR U1339 ( .A(n667), .B(n665), .Z(oi[30]) );
  XNOR U1340 ( .A(n399), .B(o[30]), .Z(n665) );
  XNOR U1341 ( .A(n662), .B(n661), .Z(n667) );
  NAND U1342 ( .A(g_input[30]), .B(e_input[0]), .Z(n661) );
  XNOR U1343 ( .A(n654), .B(n655), .Z(n662) );
  NAND U1344 ( .A(g_input[29]), .B(e_input[1]), .Z(n655) );
  XNOR U1345 ( .A(n671), .B(n416), .Z(n654) );
  XOR U1346 ( .A(n672), .B(n645), .Z(n416) );
  XNOR U1347 ( .A(n673), .B(n638), .Z(n645) );
  XNOR U1348 ( .A(n674), .B(n633), .Z(n638) );
  XNOR U1349 ( .A(n675), .B(n628), .Z(n633) );
  XNOR U1350 ( .A(n676), .B(n432), .Z(n628) );
  XNOR U1351 ( .A(n677), .B(n619), .Z(n432) );
  XNOR U1352 ( .A(n678), .B(n614), .Z(n619) );
  XNOR U1353 ( .A(n679), .B(n605), .Z(n614) );
  XNOR U1354 ( .A(n680), .B(n600), .Z(n605) );
  XNOR U1355 ( .A(n681), .B(n448), .Z(n600) );
  XNOR U1356 ( .A(n682), .B(n591), .Z(n448) );
  XNOR U1357 ( .A(n683), .B(n586), .Z(n591) );
  XNOR U1358 ( .A(n684), .B(n577), .Z(n586) );
  XNOR U1359 ( .A(n685), .B(n572), .Z(n577) );
  XNOR U1360 ( .A(n686), .B(n464), .Z(n572) );
  XNOR U1361 ( .A(n687), .B(n563), .Z(n464) );
  XNOR U1362 ( .A(n688), .B(n558), .Z(n563) );
  XNOR U1363 ( .A(n689), .B(n549), .Z(n558) );
  XNOR U1364 ( .A(n690), .B(n544), .Z(n549) );
  XNOR U1365 ( .A(n691), .B(n521), .Z(n544) );
  XNOR U1366 ( .A(n692), .B(n535), .Z(n521) );
  XNOR U1367 ( .A(n693), .B(n530), .Z(n535) );
  XNOR U1368 ( .A(n694), .B(n516), .Z(n530) );
  XNOR U1369 ( .A(n695), .B(n478), .Z(n516) );
  XNOR U1370 ( .A(n696), .B(n495), .Z(n478) );
  XNOR U1371 ( .A(n697), .B(n507), .Z(n495) );
  XNOR U1372 ( .A(n698), .B(n500), .Z(n507) );
  XNOR U1373 ( .A(n490), .B(n699), .Z(n500) );
  AND U1374 ( .A(g_input[0]), .B(e_input[30]), .Z(n699) );
  XOR U1375 ( .A(n489), .B(n502), .Z(n698) );
  NAND U1376 ( .A(e_input[29]), .B(g_input[1]), .Z(n502) );
  XOR U1377 ( .A(n491), .B(n509), .Z(n697) );
  NAND U1378 ( .A(e_input[28]), .B(g_input[2]), .Z(n509) );
  XOR U1379 ( .A(n481), .B(n497), .Z(n696) );
  NAND U1380 ( .A(e_input[27]), .B(g_input[3]), .Z(n497) );
  XOR U1381 ( .A(n499), .B(n480), .Z(n695) );
  NAND U1382 ( .A(e_input[26]), .B(g_input[4]), .Z(n480) );
  XOR U1383 ( .A(n470), .B(n518), .Z(n694) );
  NAND U1384 ( .A(e_input[25]), .B(g_input[5]), .Z(n518) );
  XOR U1385 ( .A(n525), .B(n532), .Z(n693) );
  NAND U1386 ( .A(e_input[24]), .B(g_input[6]), .Z(n532) );
  XOR U1387 ( .A(n477), .B(n537), .Z(n692) );
  NAND U1388 ( .A(e_input[23]), .B(g_input[7]), .Z(n537) );
  XOR U1389 ( .A(n539), .B(n523), .Z(n691) );
  NAND U1390 ( .A(g_input[8]), .B(e_input[22]), .Z(n523) );
  XOR U1391 ( .A(n524), .B(n546), .Z(n690) );
  NAND U1392 ( .A(g_input[9]), .B(e_input[21]), .Z(n546) );
  XOR U1393 ( .A(n455), .B(n551), .Z(n689) );
  NAND U1394 ( .A(e_input[20]), .B(g_input[10]), .Z(n551) );
  XOR U1395 ( .A(n553), .B(n560), .Z(n688) );
  NAND U1396 ( .A(e_input[19]), .B(g_input[11]), .Z(n560) );
  XOR U1397 ( .A(n463), .B(n565), .Z(n687) );
  NAND U1398 ( .A(e_input[18]), .B(g_input[12]), .Z(n565) );
  XOR U1399 ( .A(n567), .B(n465), .Z(n686) );
  NAND U1400 ( .A(e_input[17]), .B(g_input[13]), .Z(n465) );
  XOR U1401 ( .A(n552), .B(n574), .Z(n685) );
  NAND U1402 ( .A(e_input[16]), .B(g_input[14]), .Z(n574) );
  XOR U1403 ( .A(n438), .B(n579), .Z(n684) );
  NAND U1404 ( .A(e_input[15]), .B(g_input[15]), .Z(n579) );
  XOR U1405 ( .A(n581), .B(n588), .Z(n683) );
  NAND U1406 ( .A(g_input[16]), .B(e_input[14]), .Z(n588) );
  XOR U1407 ( .A(n447), .B(n593), .Z(n682) );
  NAND U1408 ( .A(g_input[17]), .B(e_input[13]), .Z(n593) );
  XOR U1409 ( .A(n595), .B(n450), .Z(n681) );
  NAND U1410 ( .A(g_input[18]), .B(e_input[12]), .Z(n450) );
  XOR U1411 ( .A(n580), .B(n602), .Z(n680) );
  NAND U1412 ( .A(g_input[19]), .B(e_input[11]), .Z(n602) );
  XOR U1413 ( .A(n423), .B(n607), .Z(n679) );
  NAND U1414 ( .A(g_input[20]), .B(e_input[10]), .Z(n607) );
  XOR U1415 ( .A(n609), .B(n616), .Z(n678) );
  NAND U1416 ( .A(g_input[21]), .B(e_input[9]), .Z(n616) );
  XOR U1417 ( .A(n431), .B(n621), .Z(n677) );
  NAND U1418 ( .A(g_input[22]), .B(e_input[8]), .Z(n621) );
  XOR U1419 ( .A(n623), .B(n433), .Z(n676) );
  NAND U1420 ( .A(g_input[23]), .B(e_input[7]), .Z(n433) );
  XOR U1421 ( .A(n608), .B(n630), .Z(n675) );
  NAND U1422 ( .A(g_input[24]), .B(e_input[6]), .Z(n630) );
  XOR U1423 ( .A(n405), .B(n635), .Z(n674) );
  NAND U1424 ( .A(g_input[25]), .B(e_input[5]), .Z(n635) );
  XOR U1425 ( .A(n648), .B(n640), .Z(n673) );
  NAND U1426 ( .A(g_input[26]), .B(e_input[4]), .Z(n640) );
  IV U1427 ( .A(n637), .Z(n648) );
  XOR U1428 ( .A(n418), .B(n647), .Z(n672) );
  NAND U1429 ( .A(g_input[27]), .B(e_input[3]), .Z(n647) );
  IV U1430 ( .A(n414), .Z(n418) );
  XOR U1431 ( .A(n417), .B(n656), .Z(n671) );
  OR U1432 ( .A(n784), .B(n785), .Z(n656) );
  ANDN U1433 ( .A(g_input[28]), .B(n786), .Z(n417) );
  XNOR U1434 ( .A(n787), .B(n788), .Z(oi[2]) );
  XNOR U1435 ( .A(n670), .B(n669), .Z(oi[29]) );
  XOR U1436 ( .A(n785), .B(n784), .Z(n670) );
  NAND U1437 ( .A(g_input[29]), .B(e_input[0]), .Z(n784) );
  XNOR U1438 ( .A(n782), .B(n783), .Z(n785) );
  NAND U1439 ( .A(g_input[28]), .B(e_input[1]), .Z(n783) );
  XNOR U1440 ( .A(n792), .B(n779), .Z(n782) );
  XOR U1441 ( .A(n793), .B(n776), .Z(n779) );
  XNOR U1442 ( .A(n794), .B(n773), .Z(n776) );
  XNOR U1443 ( .A(n795), .B(n770), .Z(n773) );
  XNOR U1444 ( .A(n796), .B(n767), .Z(n770) );
  XNOR U1445 ( .A(n797), .B(n764), .Z(n767) );
  XNOR U1446 ( .A(n798), .B(n761), .Z(n764) );
  XNOR U1447 ( .A(n799), .B(n758), .Z(n761) );
  XNOR U1448 ( .A(n800), .B(n755), .Z(n758) );
  XNOR U1449 ( .A(n801), .B(n752), .Z(n755) );
  XNOR U1450 ( .A(n802), .B(n749), .Z(n752) );
  XNOR U1451 ( .A(n803), .B(n746), .Z(n749) );
  XNOR U1452 ( .A(n804), .B(n743), .Z(n746) );
  XNOR U1453 ( .A(n805), .B(n740), .Z(n743) );
  XNOR U1454 ( .A(n806), .B(n737), .Z(n740) );
  XNOR U1455 ( .A(n807), .B(n734), .Z(n737) );
  XNOR U1456 ( .A(n808), .B(n731), .Z(n734) );
  XNOR U1457 ( .A(n809), .B(n728), .Z(n731) );
  XNOR U1458 ( .A(n810), .B(n725), .Z(n728) );
  XNOR U1459 ( .A(n811), .B(n722), .Z(n725) );
  XNOR U1460 ( .A(n812), .B(n719), .Z(n722) );
  XNOR U1461 ( .A(n813), .B(n716), .Z(n719) );
  XNOR U1462 ( .A(n814), .B(n713), .Z(n716) );
  XNOR U1463 ( .A(n815), .B(n710), .Z(n713) );
  XNOR U1464 ( .A(n816), .B(n707), .Z(n710) );
  XNOR U1465 ( .A(n817), .B(n704), .Z(n707) );
  XNOR U1466 ( .A(n818), .B(n701), .Z(n704) );
  XNOR U1467 ( .A(n700), .B(n819), .Z(n701) );
  AND U1468 ( .A(g_input[0]), .B(e_input[29]), .Z(n819) );
  NAND U1469 ( .A(e_input[28]), .B(g_input[1]), .Z(n702) );
  NAND U1470 ( .A(e_input[27]), .B(g_input[2]), .Z(n705) );
  NAND U1471 ( .A(e_input[26]), .B(g_input[3]), .Z(n708) );
  NAND U1472 ( .A(e_input[25]), .B(g_input[4]), .Z(n711) );
  NAND U1473 ( .A(e_input[24]), .B(g_input[5]), .Z(n714) );
  NAND U1474 ( .A(e_input[23]), .B(g_input[6]), .Z(n717) );
  NAND U1475 ( .A(e_input[22]), .B(g_input[7]), .Z(n720) );
  NAND U1476 ( .A(g_input[8]), .B(e_input[21]), .Z(n723) );
  NAND U1477 ( .A(g_input[9]), .B(e_input[20]), .Z(n726) );
  NAND U1478 ( .A(e_input[19]), .B(g_input[10]), .Z(n729) );
  NAND U1479 ( .A(e_input[18]), .B(g_input[11]), .Z(n732) );
  NAND U1480 ( .A(e_input[17]), .B(g_input[12]), .Z(n735) );
  NAND U1481 ( .A(e_input[16]), .B(g_input[13]), .Z(n738) );
  NAND U1482 ( .A(e_input[15]), .B(g_input[14]), .Z(n741) );
  NAND U1483 ( .A(g_input[15]), .B(e_input[14]), .Z(n744) );
  NAND U1484 ( .A(g_input[16]), .B(e_input[13]), .Z(n747) );
  NAND U1485 ( .A(g_input[17]), .B(e_input[12]), .Z(n750) );
  NAND U1486 ( .A(g_input[18]), .B(e_input[11]), .Z(n753) );
  NAND U1487 ( .A(g_input[19]), .B(e_input[10]), .Z(n756) );
  NAND U1488 ( .A(g_input[20]), .B(e_input[9]), .Z(n759) );
  NAND U1489 ( .A(g_input[21]), .B(e_input[8]), .Z(n762) );
  NAND U1490 ( .A(g_input[22]), .B(e_input[7]), .Z(n765) );
  NAND U1491 ( .A(g_input[23]), .B(e_input[6]), .Z(n768) );
  NAND U1492 ( .A(g_input[24]), .B(e_input[5]), .Z(n771) );
  NAND U1493 ( .A(g_input[25]), .B(e_input[4]), .Z(n774) );
  XNOR U1494 ( .A(n778), .B(n777), .Z(n793) );
  NAND U1495 ( .A(g_input[26]), .B(e_input[3]), .Z(n777) );
  XOR U1496 ( .A(n780), .B(n781), .Z(n792) );
  OR U1497 ( .A(n901), .B(n902), .Z(n781) );
  ANDN U1498 ( .A(g_input[27]), .B(n786), .Z(n780) );
  XNOR U1499 ( .A(n791), .B(n790), .Z(oi[28]) );
  XOR U1500 ( .A(n902), .B(n901), .Z(n791) );
  NAND U1501 ( .A(g_input[28]), .B(e_input[0]), .Z(n901) );
  XNOR U1502 ( .A(n899), .B(n900), .Z(n902) );
  NAND U1503 ( .A(g_input[27]), .B(e_input[1]), .Z(n900) );
  XNOR U1504 ( .A(n906), .B(n896), .Z(n899) );
  XOR U1505 ( .A(n907), .B(n893), .Z(n896) );
  XNOR U1506 ( .A(n908), .B(n890), .Z(n893) );
  XNOR U1507 ( .A(n909), .B(n887), .Z(n890) );
  XNOR U1508 ( .A(n910), .B(n884), .Z(n887) );
  XNOR U1509 ( .A(n911), .B(n881), .Z(n884) );
  XNOR U1510 ( .A(n912), .B(n878), .Z(n881) );
  XNOR U1511 ( .A(n913), .B(n875), .Z(n878) );
  XNOR U1512 ( .A(n914), .B(n872), .Z(n875) );
  XNOR U1513 ( .A(n915), .B(n869), .Z(n872) );
  XNOR U1514 ( .A(n916), .B(n866), .Z(n869) );
  XNOR U1515 ( .A(n917), .B(n863), .Z(n866) );
  XNOR U1516 ( .A(n918), .B(n860), .Z(n863) );
  XNOR U1517 ( .A(n919), .B(n857), .Z(n860) );
  XNOR U1518 ( .A(n920), .B(n854), .Z(n857) );
  XNOR U1519 ( .A(n921), .B(n851), .Z(n854) );
  XNOR U1520 ( .A(n922), .B(n848), .Z(n851) );
  XNOR U1521 ( .A(n923), .B(n845), .Z(n848) );
  XNOR U1522 ( .A(n924), .B(n842), .Z(n845) );
  XNOR U1523 ( .A(n925), .B(n839), .Z(n842) );
  XNOR U1524 ( .A(n926), .B(n836), .Z(n839) );
  XNOR U1525 ( .A(n927), .B(n833), .Z(n836) );
  XNOR U1526 ( .A(n928), .B(n830), .Z(n833) );
  XNOR U1527 ( .A(n929), .B(n827), .Z(n830) );
  XNOR U1528 ( .A(n930), .B(n824), .Z(n827) );
  XNOR U1529 ( .A(n931), .B(n821), .Z(n824) );
  XNOR U1530 ( .A(n820), .B(n932), .Z(n821) );
  AND U1531 ( .A(g_input[0]), .B(e_input[28]), .Z(n932) );
  NAND U1532 ( .A(e_input[27]), .B(g_input[1]), .Z(n822) );
  NAND U1533 ( .A(e_input[26]), .B(g_input[2]), .Z(n825) );
  NAND U1534 ( .A(e_input[25]), .B(g_input[3]), .Z(n828) );
  NAND U1535 ( .A(e_input[24]), .B(g_input[4]), .Z(n831) );
  NAND U1536 ( .A(e_input[23]), .B(g_input[5]), .Z(n834) );
  NAND U1537 ( .A(e_input[22]), .B(g_input[6]), .Z(n837) );
  NAND U1538 ( .A(e_input[21]), .B(g_input[7]), .Z(n840) );
  NAND U1539 ( .A(g_input[8]), .B(e_input[20]), .Z(n843) );
  NAND U1540 ( .A(g_input[9]), .B(e_input[19]), .Z(n846) );
  NAND U1541 ( .A(e_input[18]), .B(g_input[10]), .Z(n849) );
  NAND U1542 ( .A(e_input[17]), .B(g_input[11]), .Z(n852) );
  NAND U1543 ( .A(e_input[16]), .B(g_input[12]), .Z(n855) );
  NAND U1544 ( .A(e_input[15]), .B(g_input[13]), .Z(n858) );
  NAND U1545 ( .A(e_input[14]), .B(g_input[14]), .Z(n861) );
  NAND U1546 ( .A(g_input[15]), .B(e_input[13]), .Z(n864) );
  NAND U1547 ( .A(g_input[16]), .B(e_input[12]), .Z(n867) );
  XNOR U1548 ( .A(n984), .B(n870), .Z(n915) );
  NAND U1549 ( .A(g_input[17]), .B(e_input[11]), .Z(n870) );
  IV U1550 ( .A(n871), .Z(n984) );
  NAND U1551 ( .A(g_input[18]), .B(e_input[10]), .Z(n873) );
  NAND U1552 ( .A(g_input[19]), .B(e_input[9]), .Z(n876) );
  NAND U1553 ( .A(g_input[20]), .B(e_input[8]), .Z(n879) );
  NAND U1554 ( .A(g_input[21]), .B(e_input[7]), .Z(n882) );
  NAND U1555 ( .A(g_input[22]), .B(e_input[6]), .Z(n885) );
  NAND U1556 ( .A(g_input[23]), .B(e_input[5]), .Z(n888) );
  NAND U1557 ( .A(g_input[24]), .B(e_input[4]), .Z(n891) );
  XNOR U1558 ( .A(n895), .B(n894), .Z(n907) );
  NAND U1559 ( .A(g_input[25]), .B(e_input[3]), .Z(n894) );
  XOR U1560 ( .A(n897), .B(n898), .Z(n906) );
  OR U1561 ( .A(n1012), .B(n1013), .Z(n898) );
  ANDN U1562 ( .A(g_input[26]), .B(n786), .Z(n897) );
  XNOR U1563 ( .A(n905), .B(n904), .Z(oi[27]) );
  XOR U1564 ( .A(n1013), .B(n1012), .Z(n905) );
  NAND U1565 ( .A(g_input[27]), .B(e_input[0]), .Z(n1012) );
  XNOR U1566 ( .A(n1010), .B(n1011), .Z(n1013) );
  NAND U1567 ( .A(g_input[26]), .B(e_input[1]), .Z(n1011) );
  XNOR U1568 ( .A(n1017), .B(n1007), .Z(n1010) );
  XOR U1569 ( .A(n1018), .B(n1004), .Z(n1007) );
  XNOR U1570 ( .A(n1019), .B(n1001), .Z(n1004) );
  XNOR U1571 ( .A(n1020), .B(n998), .Z(n1001) );
  XNOR U1572 ( .A(n1021), .B(n995), .Z(n998) );
  XNOR U1573 ( .A(n1022), .B(n992), .Z(n995) );
  XNOR U1574 ( .A(n1023), .B(n989), .Z(n992) );
  XNOR U1575 ( .A(n1024), .B(n986), .Z(n989) );
  XNOR U1576 ( .A(n1025), .B(n982), .Z(n986) );
  XNOR U1577 ( .A(n1026), .B(n979), .Z(n982) );
  XNOR U1578 ( .A(n1027), .B(n976), .Z(n979) );
  XNOR U1579 ( .A(n1028), .B(n973), .Z(n976) );
  XNOR U1580 ( .A(n1029), .B(n970), .Z(n973) );
  XNOR U1581 ( .A(n1030), .B(n967), .Z(n970) );
  XNOR U1582 ( .A(n1031), .B(n964), .Z(n967) );
  XNOR U1583 ( .A(n1032), .B(n961), .Z(n964) );
  XNOR U1584 ( .A(n1033), .B(n958), .Z(n961) );
  XNOR U1585 ( .A(n1034), .B(n955), .Z(n958) );
  XNOR U1586 ( .A(n1035), .B(n952), .Z(n955) );
  XNOR U1587 ( .A(n1036), .B(n949), .Z(n952) );
  XNOR U1588 ( .A(n1037), .B(n946), .Z(n949) );
  XNOR U1589 ( .A(n1038), .B(n943), .Z(n946) );
  XNOR U1590 ( .A(n1039), .B(n940), .Z(n943) );
  XNOR U1591 ( .A(n1040), .B(n937), .Z(n940) );
  XNOR U1592 ( .A(n1041), .B(n934), .Z(n937) );
  XNOR U1593 ( .A(n933), .B(n1042), .Z(n934) );
  AND U1594 ( .A(g_input[0]), .B(e_input[27]), .Z(n1042) );
  NAND U1595 ( .A(e_input[26]), .B(g_input[1]), .Z(n935) );
  XNOR U1596 ( .A(n1049), .B(n938), .Z(n1040) );
  NAND U1597 ( .A(e_input[25]), .B(g_input[2]), .Z(n938) );
  IV U1598 ( .A(n939), .Z(n1049) );
  NAND U1599 ( .A(e_input[24]), .B(g_input[3]), .Z(n941) );
  XNOR U1600 ( .A(n1056), .B(n944), .Z(n1038) );
  NAND U1601 ( .A(e_input[23]), .B(g_input[4]), .Z(n944) );
  IV U1602 ( .A(n945), .Z(n1056) );
  NAND U1603 ( .A(e_input[22]), .B(g_input[5]), .Z(n947) );
  NAND U1604 ( .A(e_input[21]), .B(g_input[6]), .Z(n950) );
  NAND U1605 ( .A(e_input[20]), .B(g_input[7]), .Z(n953) );
  NAND U1606 ( .A(g_input[8]), .B(e_input[19]), .Z(n956) );
  NAND U1607 ( .A(g_input[9]), .B(e_input[18]), .Z(n959) );
  NAND U1608 ( .A(e_input[17]), .B(g_input[10]), .Z(n962) );
  NAND U1609 ( .A(e_input[16]), .B(g_input[11]), .Z(n965) );
  XNOR U1610 ( .A(n1081), .B(n968), .Z(n1030) );
  NAND U1611 ( .A(e_input[15]), .B(g_input[12]), .Z(n968) );
  IV U1612 ( .A(n969), .Z(n1081) );
  XNOR U1613 ( .A(n1085), .B(n971), .Z(n1029) );
  NAND U1614 ( .A(e_input[14]), .B(g_input[13]), .Z(n971) );
  IV U1615 ( .A(n972), .Z(n1085) );
  XNOR U1616 ( .A(n1089), .B(n974), .Z(n1028) );
  NAND U1617 ( .A(g_input[14]), .B(e_input[13]), .Z(n974) );
  IV U1618 ( .A(n975), .Z(n1089) );
  XOR U1619 ( .A(n1090), .B(n1091), .Z(n975) );
  AND U1620 ( .A(n1092), .B(n1093), .Z(n1091) );
  XNOR U1621 ( .A(n1094), .B(n1090), .Z(n1093) );
  NAND U1622 ( .A(g_input[15]), .B(e_input[12]), .Z(n977) );
  NAND U1623 ( .A(g_input[16]), .B(e_input[11]), .Z(n980) );
  NAND U1624 ( .A(g_input[17]), .B(e_input[10]), .Z(n983) );
  NAND U1625 ( .A(g_input[18]), .B(e_input[9]), .Z(n987) );
  NAND U1626 ( .A(g_input[19]), .B(e_input[8]), .Z(n990) );
  XOR U1627 ( .A(n1107), .B(n1108), .Z(n991) );
  AND U1628 ( .A(n1109), .B(n1110), .Z(n1108) );
  XNOR U1629 ( .A(n1111), .B(n1107), .Z(n1110) );
  NAND U1630 ( .A(g_input[20]), .B(e_input[7]), .Z(n993) );
  NAND U1631 ( .A(g_input[21]), .B(e_input[6]), .Z(n996) );
  NAND U1632 ( .A(g_input[22]), .B(e_input[5]), .Z(n999) );
  NAND U1633 ( .A(g_input[23]), .B(e_input[4]), .Z(n1002) );
  XNOR U1634 ( .A(n1006), .B(n1005), .Z(n1018) );
  NAND U1635 ( .A(g_input[24]), .B(e_input[3]), .Z(n1005) );
  XOR U1636 ( .A(n1008), .B(n1009), .Z(n1017) );
  OR U1637 ( .A(n1127), .B(n1128), .Z(n1009) );
  ANDN U1638 ( .A(g_input[25]), .B(n786), .Z(n1008) );
  XNOR U1639 ( .A(n1016), .B(n1015), .Z(oi[26]) );
  XOR U1640 ( .A(n1128), .B(n1127), .Z(n1016) );
  NAND U1641 ( .A(g_input[26]), .B(e_input[0]), .Z(n1127) );
  XNOR U1642 ( .A(n1125), .B(n1126), .Z(n1128) );
  NAND U1643 ( .A(g_input[25]), .B(e_input[1]), .Z(n1126) );
  XNOR U1644 ( .A(n1132), .B(n1122), .Z(n1125) );
  XOR U1645 ( .A(n1133), .B(n1119), .Z(n1122) );
  XNOR U1646 ( .A(n1134), .B(n1116), .Z(n1119) );
  XNOR U1647 ( .A(n1135), .B(n1113), .Z(n1116) );
  XNOR U1648 ( .A(n1136), .B(n1109), .Z(n1113) );
  XNOR U1649 ( .A(n1137), .B(n1105), .Z(n1109) );
  XNOR U1650 ( .A(n1138), .B(n1102), .Z(n1105) );
  XNOR U1651 ( .A(n1139), .B(n1099), .Z(n1102) );
  XNOR U1652 ( .A(n1140), .B(n1096), .Z(n1099) );
  XNOR U1653 ( .A(n1141), .B(n1092), .Z(n1096) );
  XNOR U1654 ( .A(n1142), .B(n1087), .Z(n1092) );
  XNOR U1655 ( .A(n1143), .B(n1083), .Z(n1087) );
  XNOR U1656 ( .A(n1144), .B(n1079), .Z(n1083) );
  XNOR U1657 ( .A(n1145), .B(n1076), .Z(n1079) );
  XNOR U1658 ( .A(n1146), .B(n1073), .Z(n1076) );
  XNOR U1659 ( .A(n1147), .B(n1070), .Z(n1073) );
  XNOR U1660 ( .A(n1148), .B(n1067), .Z(n1070) );
  XNOR U1661 ( .A(n1149), .B(n1064), .Z(n1067) );
  XNOR U1662 ( .A(n1150), .B(n1061), .Z(n1064) );
  XNOR U1663 ( .A(n1151), .B(n1058), .Z(n1061) );
  XNOR U1664 ( .A(n1152), .B(n1054), .Z(n1058) );
  XNOR U1665 ( .A(n1153), .B(n1051), .Z(n1054) );
  XNOR U1666 ( .A(n1154), .B(n1047), .Z(n1051) );
  XNOR U1667 ( .A(n1155), .B(n1044), .Z(n1047) );
  XNOR U1668 ( .A(n1043), .B(n1156), .Z(n1044) );
  AND U1669 ( .A(g_input[0]), .B(e_input[26]), .Z(n1156) );
  NAND U1670 ( .A(e_input[25]), .B(g_input[1]), .Z(n1045) );
  NAND U1671 ( .A(e_input[24]), .B(g_input[2]), .Z(n1048) );
  XOR U1672 ( .A(n1163), .B(n1164), .Z(n1050) );
  AND U1673 ( .A(n1165), .B(n1166), .Z(n1164) );
  XNOR U1674 ( .A(n1167), .B(n1163), .Z(n1166) );
  NAND U1675 ( .A(e_input[23]), .B(g_input[3]), .Z(n1052) );
  NAND U1676 ( .A(e_input[22]), .B(g_input[4]), .Z(n1055) );
  NAND U1677 ( .A(e_input[21]), .B(g_input[5]), .Z(n1059) );
  NAND U1678 ( .A(e_input[20]), .B(g_input[6]), .Z(n1062) );
  NAND U1679 ( .A(e_input[19]), .B(g_input[7]), .Z(n1065) );
  NAND U1680 ( .A(g_input[8]), .B(e_input[18]), .Z(n1068) );
  XNOR U1681 ( .A(n1186), .B(n1071), .Z(n1147) );
  NAND U1682 ( .A(g_input[9]), .B(e_input[17]), .Z(n1071) );
  IV U1683 ( .A(n1072), .Z(n1186) );
  XOR U1684 ( .A(n1187), .B(n1188), .Z(n1072) );
  AND U1685 ( .A(n1189), .B(n1190), .Z(n1188) );
  XNOR U1686 ( .A(n1191), .B(n1187), .Z(n1190) );
  XNOR U1687 ( .A(n1192), .B(n1074), .Z(n1146) );
  NAND U1688 ( .A(e_input[16]), .B(g_input[10]), .Z(n1074) );
  IV U1689 ( .A(n1075), .Z(n1192) );
  NAND U1690 ( .A(e_input[15]), .B(g_input[11]), .Z(n1077) );
  NAND U1691 ( .A(e_input[14]), .B(g_input[12]), .Z(n1080) );
  XOR U1692 ( .A(n1199), .B(n1200), .Z(n1082) );
  AND U1693 ( .A(n1201), .B(n1202), .Z(n1200) );
  XNOR U1694 ( .A(n1203), .B(n1199), .Z(n1202) );
  NAND U1695 ( .A(e_input[13]), .B(g_input[13]), .Z(n1084) );
  NAND U1696 ( .A(g_input[14]), .B(e_input[12]), .Z(n1088) );
  NAND U1697 ( .A(g_input[15]), .B(e_input[11]), .Z(n1094) );
  NAND U1698 ( .A(g_input[16]), .B(e_input[10]), .Z(n1097) );
  NAND U1699 ( .A(g_input[17]), .B(e_input[9]), .Z(n1100) );
  NAND U1700 ( .A(g_input[18]), .B(e_input[8]), .Z(n1103) );
  NAND U1701 ( .A(g_input[19]), .B(e_input[7]), .Z(n1106) );
  NAND U1702 ( .A(g_input[20]), .B(e_input[6]), .Z(n1111) );
  NAND U1703 ( .A(g_input[21]), .B(e_input[5]), .Z(n1114) );
  NAND U1704 ( .A(g_input[22]), .B(e_input[4]), .Z(n1117) );
  XNOR U1705 ( .A(n1121), .B(n1120), .Z(n1133) );
  NAND U1706 ( .A(g_input[23]), .B(e_input[3]), .Z(n1120) );
  XOR U1707 ( .A(n1123), .B(n1124), .Z(n1132) );
  OR U1708 ( .A(n1237), .B(n1238), .Z(n1124) );
  ANDN U1709 ( .A(g_input[24]), .B(n786), .Z(n1123) );
  XNOR U1710 ( .A(n1131), .B(n1130), .Z(oi[25]) );
  XOR U1711 ( .A(n1238), .B(n1237), .Z(n1131) );
  NAND U1712 ( .A(g_input[25]), .B(e_input[0]), .Z(n1237) );
  XNOR U1713 ( .A(n1235), .B(n1236), .Z(n1238) );
  NAND U1714 ( .A(g_input[24]), .B(e_input[1]), .Z(n1236) );
  XNOR U1715 ( .A(n1242), .B(n1232), .Z(n1235) );
  XOR U1716 ( .A(n1243), .B(n1229), .Z(n1232) );
  XNOR U1717 ( .A(n1244), .B(n1226), .Z(n1229) );
  XNOR U1718 ( .A(n1245), .B(n1223), .Z(n1226) );
  XNOR U1719 ( .A(n1246), .B(n1220), .Z(n1223) );
  XNOR U1720 ( .A(n1247), .B(n1217), .Z(n1220) );
  XNOR U1721 ( .A(n1248), .B(n1214), .Z(n1217) );
  XNOR U1722 ( .A(n1249), .B(n1211), .Z(n1214) );
  XNOR U1723 ( .A(n1250), .B(n1208), .Z(n1211) );
  XNOR U1724 ( .A(n1251), .B(n1205), .Z(n1208) );
  XNOR U1725 ( .A(n1252), .B(n1201), .Z(n1205) );
  XNOR U1726 ( .A(n1253), .B(n1197), .Z(n1201) );
  XNOR U1727 ( .A(n1254), .B(n1194), .Z(n1197) );
  XNOR U1728 ( .A(n1255), .B(n1189), .Z(n1194) );
  XNOR U1729 ( .A(n1256), .B(n1184), .Z(n1189) );
  XNOR U1730 ( .A(n1257), .B(n1181), .Z(n1184) );
  XNOR U1731 ( .A(n1258), .B(n1178), .Z(n1181) );
  XNOR U1732 ( .A(n1259), .B(n1175), .Z(n1178) );
  XNOR U1733 ( .A(n1260), .B(n1172), .Z(n1175) );
  XNOR U1734 ( .A(n1261), .B(n1169), .Z(n1172) );
  XNOR U1735 ( .A(n1262), .B(n1165), .Z(n1169) );
  XNOR U1736 ( .A(n1263), .B(n1161), .Z(n1165) );
  XNOR U1737 ( .A(n1264), .B(n1158), .Z(n1161) );
  XNOR U1738 ( .A(n1157), .B(n1265), .Z(n1158) );
  AND U1739 ( .A(g_input[0]), .B(e_input[25]), .Z(n1265) );
  NAND U1740 ( .A(e_input[24]), .B(g_input[1]), .Z(n1159) );
  XNOR U1741 ( .A(n1272), .B(n1162), .Z(n1263) );
  NAND U1742 ( .A(e_input[23]), .B(g_input[2]), .Z(n1162) );
  IV U1743 ( .A(n1163), .Z(n1272) );
  NAND U1744 ( .A(e_input[22]), .B(g_input[3]), .Z(n1167) );
  NAND U1745 ( .A(e_input[21]), .B(g_input[4]), .Z(n1170) );
  NAND U1746 ( .A(e_input[20]), .B(g_input[5]), .Z(n1173) );
  XNOR U1747 ( .A(n1285), .B(n1176), .Z(n1259) );
  NAND U1748 ( .A(e_input[19]), .B(g_input[6]), .Z(n1176) );
  IV U1749 ( .A(n1177), .Z(n1285) );
  NAND U1750 ( .A(e_input[18]), .B(g_input[7]), .Z(n1179) );
  XOR U1751 ( .A(n1289), .B(n1290), .Z(n1180) );
  AND U1752 ( .A(n1291), .B(n1292), .Z(n1290) );
  XNOR U1753 ( .A(n1293), .B(n1289), .Z(n1292) );
  NAND U1754 ( .A(g_input[8]), .B(e_input[17]), .Z(n1182) );
  XNOR U1755 ( .A(n1297), .B(n1185), .Z(n1256) );
  NAND U1756 ( .A(g_input[9]), .B(e_input[16]), .Z(n1185) );
  IV U1757 ( .A(n1187), .Z(n1297) );
  NAND U1758 ( .A(e_input[15]), .B(g_input[10]), .Z(n1191) );
  NAND U1759 ( .A(e_input[14]), .B(g_input[11]), .Z(n1195) );
  NAND U1760 ( .A(e_input[13]), .B(g_input[12]), .Z(n1198) );
  NAND U1761 ( .A(g_input[13]), .B(e_input[12]), .Z(n1203) );
  NAND U1762 ( .A(g_input[14]), .B(e_input[11]), .Z(n1206) );
  NAND U1763 ( .A(g_input[15]), .B(e_input[10]), .Z(n1209) );
  NAND U1764 ( .A(g_input[16]), .B(e_input[9]), .Z(n1212) );
  NAND U1765 ( .A(g_input[17]), .B(e_input[8]), .Z(n1215) );
  NAND U1766 ( .A(g_input[18]), .B(e_input[7]), .Z(n1218) );
  NAND U1767 ( .A(g_input[19]), .B(e_input[6]), .Z(n1221) );
  NAND U1768 ( .A(g_input[20]), .B(e_input[5]), .Z(n1224) );
  NAND U1769 ( .A(g_input[21]), .B(e_input[4]), .Z(n1227) );
  XNOR U1770 ( .A(n1231), .B(n1230), .Z(n1243) );
  NAND U1771 ( .A(g_input[22]), .B(e_input[3]), .Z(n1230) );
  XOR U1772 ( .A(n1233), .B(n1234), .Z(n1242) );
  OR U1773 ( .A(n1340), .B(n1341), .Z(n1234) );
  ANDN U1774 ( .A(g_input[23]), .B(n786), .Z(n1233) );
  XNOR U1775 ( .A(n1241), .B(n1240), .Z(oi[24]) );
  XOR U1776 ( .A(n1341), .B(n1340), .Z(n1241) );
  NAND U1777 ( .A(g_input[24]), .B(e_input[0]), .Z(n1340) );
  XNOR U1778 ( .A(n1338), .B(n1339), .Z(n1341) );
  NAND U1779 ( .A(g_input[23]), .B(e_input[1]), .Z(n1339) );
  XNOR U1780 ( .A(n1345), .B(n1335), .Z(n1338) );
  XOR U1781 ( .A(n1346), .B(n1332), .Z(n1335) );
  XNOR U1782 ( .A(n1347), .B(n1329), .Z(n1332) );
  XNOR U1783 ( .A(n1348), .B(n1326), .Z(n1329) );
  XNOR U1784 ( .A(n1349), .B(n1323), .Z(n1326) );
  XNOR U1785 ( .A(n1350), .B(n1320), .Z(n1323) );
  XNOR U1786 ( .A(n1351), .B(n1317), .Z(n1320) );
  XNOR U1787 ( .A(n1352), .B(n1314), .Z(n1317) );
  XNOR U1788 ( .A(n1353), .B(n1311), .Z(n1314) );
  XNOR U1789 ( .A(n1354), .B(n1308), .Z(n1311) );
  XNOR U1790 ( .A(n1355), .B(n1305), .Z(n1308) );
  XNOR U1791 ( .A(n1356), .B(n1302), .Z(n1305) );
  XNOR U1792 ( .A(n1357), .B(n1299), .Z(n1302) );
  XNOR U1793 ( .A(n1358), .B(n1295), .Z(n1299) );
  XNOR U1794 ( .A(n1359), .B(n1291), .Z(n1295) );
  XNOR U1795 ( .A(n1360), .B(n1287), .Z(n1291) );
  XNOR U1796 ( .A(n1361), .B(n1283), .Z(n1287) );
  XNOR U1797 ( .A(n1362), .B(n1280), .Z(n1283) );
  XNOR U1798 ( .A(n1363), .B(n1277), .Z(n1280) );
  XNOR U1799 ( .A(n1364), .B(n1274), .Z(n1277) );
  XNOR U1800 ( .A(n1365), .B(n1270), .Z(n1274) );
  XNOR U1801 ( .A(n1366), .B(n1267), .Z(n1270) );
  XNOR U1802 ( .A(n1266), .B(n1367), .Z(n1267) );
  AND U1803 ( .A(g_input[0]), .B(e_input[24]), .Z(n1367) );
  NAND U1804 ( .A(e_input[23]), .B(g_input[1]), .Z(n1268) );
  NAND U1805 ( .A(e_input[22]), .B(g_input[2]), .Z(n1271) );
  XNOR U1806 ( .A(n1377), .B(n1275), .Z(n1364) );
  NAND U1807 ( .A(e_input[21]), .B(g_input[3]), .Z(n1275) );
  IV U1808 ( .A(n1276), .Z(n1377) );
  NAND U1809 ( .A(e_input[20]), .B(g_input[4]), .Z(n1278) );
  NAND U1810 ( .A(e_input[19]), .B(g_input[5]), .Z(n1281) );
  NAND U1811 ( .A(e_input[18]), .B(g_input[6]), .Z(n1284) );
  NAND U1812 ( .A(e_input[17]), .B(g_input[7]), .Z(n1288) );
  NAND U1813 ( .A(g_input[8]), .B(e_input[16]), .Z(n1293) );
  XOR U1814 ( .A(n1393), .B(n1394), .Z(n1294) );
  AND U1815 ( .A(n1395), .B(n1396), .Z(n1394) );
  XNOR U1816 ( .A(n1397), .B(n1393), .Z(n1396) );
  NAND U1817 ( .A(g_input[9]), .B(e_input[15]), .Z(n1296) );
  NAND U1818 ( .A(e_input[14]), .B(g_input[10]), .Z(n1300) );
  NAND U1819 ( .A(e_input[13]), .B(g_input[11]), .Z(n1303) );
  NAND U1820 ( .A(e_input[12]), .B(g_input[12]), .Z(n1306) );
  NAND U1821 ( .A(g_input[13]), .B(e_input[11]), .Z(n1309) );
  NAND U1822 ( .A(g_input[14]), .B(e_input[10]), .Z(n1312) );
  NAND U1823 ( .A(g_input[15]), .B(e_input[9]), .Z(n1315) );
  NAND U1824 ( .A(g_input[16]), .B(e_input[8]), .Z(n1318) );
  NAND U1825 ( .A(g_input[17]), .B(e_input[7]), .Z(n1321) );
  NAND U1826 ( .A(g_input[18]), .B(e_input[6]), .Z(n1324) );
  NAND U1827 ( .A(g_input[19]), .B(e_input[5]), .Z(n1327) );
  NAND U1828 ( .A(g_input[20]), .B(e_input[4]), .Z(n1330) );
  XNOR U1829 ( .A(n1334), .B(n1333), .Z(n1346) );
  NAND U1830 ( .A(g_input[21]), .B(e_input[3]), .Z(n1333) );
  XOR U1831 ( .A(n1336), .B(n1337), .Z(n1345) );
  OR U1832 ( .A(n1437), .B(n1438), .Z(n1337) );
  ANDN U1833 ( .A(g_input[22]), .B(n786), .Z(n1336) );
  XNOR U1834 ( .A(n1344), .B(n1343), .Z(oi[23]) );
  XOR U1835 ( .A(n1438), .B(n1437), .Z(n1344) );
  NAND U1836 ( .A(g_input[23]), .B(e_input[0]), .Z(n1437) );
  XNOR U1837 ( .A(n1435), .B(n1436), .Z(n1438) );
  NAND U1838 ( .A(g_input[22]), .B(e_input[1]), .Z(n1436) );
  XNOR U1839 ( .A(n1442), .B(n1432), .Z(n1435) );
  XOR U1840 ( .A(n1443), .B(n1429), .Z(n1432) );
  XNOR U1841 ( .A(n1444), .B(n1426), .Z(n1429) );
  XNOR U1842 ( .A(n1445), .B(n1423), .Z(n1426) );
  XNOR U1843 ( .A(n1446), .B(n1420), .Z(n1423) );
  XNOR U1844 ( .A(n1447), .B(n1417), .Z(n1420) );
  XNOR U1845 ( .A(n1448), .B(n1414), .Z(n1417) );
  XNOR U1846 ( .A(n1449), .B(n1411), .Z(n1414) );
  XNOR U1847 ( .A(n1450), .B(n1408), .Z(n1411) );
  XNOR U1848 ( .A(n1451), .B(n1405), .Z(n1408) );
  XNOR U1849 ( .A(n1452), .B(n1402), .Z(n1405) );
  XNOR U1850 ( .A(n1453), .B(n1399), .Z(n1402) );
  XNOR U1851 ( .A(n1454), .B(n1395), .Z(n1399) );
  XNOR U1852 ( .A(n1455), .B(n1391), .Z(n1395) );
  XNOR U1853 ( .A(n1456), .B(n1388), .Z(n1391) );
  XNOR U1854 ( .A(n1457), .B(n1385), .Z(n1388) );
  XNOR U1855 ( .A(n1458), .B(n1382), .Z(n1385) );
  XNOR U1856 ( .A(n1459), .B(n1379), .Z(n1382) );
  XNOR U1857 ( .A(n1460), .B(n1375), .Z(n1379) );
  XNOR U1858 ( .A(n1461), .B(n1372), .Z(n1375) );
  XNOR U1859 ( .A(n1462), .B(n1369), .Z(n1372) );
  XNOR U1860 ( .A(n1368), .B(n1463), .Z(n1369) );
  AND U1861 ( .A(g_input[0]), .B(e_input[23]), .Z(n1463) );
  XNOR U1862 ( .A(n1467), .B(n1370), .Z(n1462) );
  NAND U1863 ( .A(e_input[22]), .B(g_input[1]), .Z(n1370) );
  IV U1864 ( .A(n1371), .Z(n1467) );
  NAND U1865 ( .A(e_input[21]), .B(g_input[2]), .Z(n1373) );
  XOR U1866 ( .A(n1471), .B(n1472), .Z(n1374) );
  AND U1867 ( .A(n1473), .B(n1474), .Z(n1472) );
  XNOR U1868 ( .A(n1475), .B(n1471), .Z(n1474) );
  NAND U1869 ( .A(e_input[20]), .B(g_input[3]), .Z(n1376) );
  NAND U1870 ( .A(e_input[19]), .B(g_input[4]), .Z(n1380) );
  NAND U1871 ( .A(e_input[18]), .B(g_input[5]), .Z(n1383) );
  XOR U1872 ( .A(n1482), .B(n1483), .Z(n1384) );
  AND U1873 ( .A(n1484), .B(n1485), .Z(n1483) );
  XNOR U1874 ( .A(n1486), .B(n1482), .Z(n1485) );
  NAND U1875 ( .A(e_input[17]), .B(g_input[6]), .Z(n1386) );
  NAND U1876 ( .A(e_input[16]), .B(g_input[7]), .Z(n1389) );
  NAND U1877 ( .A(g_input[8]), .B(e_input[15]), .Z(n1392) );
  NAND U1878 ( .A(g_input[9]), .B(e_input[14]), .Z(n1397) );
  NAND U1879 ( .A(e_input[13]), .B(g_input[10]), .Z(n1400) );
  NAND U1880 ( .A(e_input[12]), .B(g_input[11]), .Z(n1403) );
  NAND U1881 ( .A(g_input[12]), .B(e_input[11]), .Z(n1406) );
  NAND U1882 ( .A(g_input[13]), .B(e_input[10]), .Z(n1409) );
  NAND U1883 ( .A(g_input[14]), .B(e_input[9]), .Z(n1412) );
  NAND U1884 ( .A(g_input[15]), .B(e_input[8]), .Z(n1415) );
  NAND U1885 ( .A(g_input[16]), .B(e_input[7]), .Z(n1418) );
  NAND U1886 ( .A(g_input[17]), .B(e_input[6]), .Z(n1421) );
  NAND U1887 ( .A(g_input[18]), .B(e_input[5]), .Z(n1424) );
  NAND U1888 ( .A(g_input[19]), .B(e_input[4]), .Z(n1427) );
  XNOR U1889 ( .A(n1431), .B(n1430), .Z(n1443) );
  NAND U1890 ( .A(g_input[20]), .B(e_input[3]), .Z(n1430) );
  XOR U1891 ( .A(n1433), .B(n1434), .Z(n1442) );
  OR U1892 ( .A(n1532), .B(n1533), .Z(n1434) );
  ANDN U1893 ( .A(g_input[21]), .B(n786), .Z(n1433) );
  XNOR U1894 ( .A(n1441), .B(n1440), .Z(oi[22]) );
  XOR U1895 ( .A(n1533), .B(n1532), .Z(n1441) );
  NAND U1896 ( .A(g_input[22]), .B(e_input[0]), .Z(n1532) );
  XNOR U1897 ( .A(n1530), .B(n1531), .Z(n1533) );
  NAND U1898 ( .A(g_input[21]), .B(e_input[1]), .Z(n1531) );
  XNOR U1899 ( .A(n1537), .B(n1527), .Z(n1530) );
  XOR U1900 ( .A(n1538), .B(n1524), .Z(n1527) );
  XNOR U1901 ( .A(n1539), .B(n1521), .Z(n1524) );
  XNOR U1902 ( .A(n1540), .B(n1518), .Z(n1521) );
  XNOR U1903 ( .A(n1541), .B(n1515), .Z(n1518) );
  XNOR U1904 ( .A(n1542), .B(n1512), .Z(n1515) );
  XNOR U1905 ( .A(n1543), .B(n1509), .Z(n1512) );
  XNOR U1906 ( .A(n1544), .B(n1506), .Z(n1509) );
  XNOR U1907 ( .A(n1545), .B(n1503), .Z(n1506) );
  XNOR U1908 ( .A(n1546), .B(n1500), .Z(n1503) );
  XNOR U1909 ( .A(n1547), .B(n1497), .Z(n1500) );
  XNOR U1910 ( .A(n1548), .B(n1494), .Z(n1497) );
  XNOR U1911 ( .A(n1549), .B(n1491), .Z(n1494) );
  XNOR U1912 ( .A(n1550), .B(n1488), .Z(n1491) );
  XNOR U1913 ( .A(n1551), .B(n1484), .Z(n1488) );
  XNOR U1914 ( .A(n1552), .B(n1480), .Z(n1484) );
  XNOR U1915 ( .A(n1553), .B(n1477), .Z(n1480) );
  XNOR U1916 ( .A(n1554), .B(n1473), .Z(n1477) );
  XNOR U1917 ( .A(n1555), .B(n1469), .Z(n1473) );
  XNOR U1918 ( .A(n1556), .B(n1465), .Z(n1469) );
  XNOR U1919 ( .A(n1464), .B(n1557), .Z(n1465) );
  AND U1920 ( .A(g_input[0]), .B(e_input[22]), .Z(n1557) );
  NAND U1921 ( .A(e_input[21]), .B(g_input[1]), .Z(n1466) );
  NAND U1922 ( .A(e_input[20]), .B(g_input[2]), .Z(n1470) );
  NAND U1923 ( .A(e_input[19]), .B(g_input[3]), .Z(n1475) );
  NAND U1924 ( .A(e_input[18]), .B(g_input[4]), .Z(n1478) );
  NAND U1925 ( .A(e_input[17]), .B(g_input[5]), .Z(n1481) );
  NAND U1926 ( .A(e_input[16]), .B(g_input[6]), .Z(n1486) );
  NAND U1927 ( .A(e_input[15]), .B(g_input[7]), .Z(n1489) );
  NAND U1928 ( .A(g_input[8]), .B(e_input[14]), .Z(n1492) );
  NAND U1929 ( .A(g_input[9]), .B(e_input[13]), .Z(n1495) );
  NAND U1930 ( .A(e_input[12]), .B(g_input[10]), .Z(n1498) );
  NAND U1931 ( .A(e_input[11]), .B(g_input[11]), .Z(n1501) );
  NAND U1932 ( .A(g_input[12]), .B(e_input[10]), .Z(n1504) );
  NAND U1933 ( .A(g_input[13]), .B(e_input[9]), .Z(n1507) );
  NAND U1934 ( .A(g_input[14]), .B(e_input[8]), .Z(n1510) );
  NAND U1935 ( .A(g_input[15]), .B(e_input[7]), .Z(n1513) );
  NAND U1936 ( .A(g_input[16]), .B(e_input[6]), .Z(n1516) );
  NAND U1937 ( .A(g_input[17]), .B(e_input[5]), .Z(n1519) );
  NAND U1938 ( .A(g_input[18]), .B(e_input[4]), .Z(n1522) );
  XNOR U1939 ( .A(n1526), .B(n1525), .Z(n1538) );
  NAND U1940 ( .A(g_input[19]), .B(e_input[3]), .Z(n1525) );
  XOR U1941 ( .A(n1528), .B(n1529), .Z(n1537) );
  OR U1942 ( .A(n1618), .B(n1619), .Z(n1529) );
  ANDN U1943 ( .A(g_input[20]), .B(n786), .Z(n1528) );
  XNOR U1944 ( .A(n1536), .B(n1535), .Z(oi[21]) );
  XOR U1945 ( .A(n1619), .B(n1618), .Z(n1536) );
  NAND U1946 ( .A(g_input[21]), .B(e_input[0]), .Z(n1618) );
  XNOR U1947 ( .A(n1616), .B(n1617), .Z(n1619) );
  NAND U1948 ( .A(g_input[20]), .B(e_input[1]), .Z(n1617) );
  XNOR U1949 ( .A(n1623), .B(n1613), .Z(n1616) );
  XOR U1950 ( .A(n1624), .B(n1610), .Z(n1613) );
  XNOR U1951 ( .A(n1625), .B(n1607), .Z(n1610) );
  XNOR U1952 ( .A(n1626), .B(n1604), .Z(n1607) );
  XNOR U1953 ( .A(n1627), .B(n1601), .Z(n1604) );
  XNOR U1954 ( .A(n1628), .B(n1598), .Z(n1601) );
  XNOR U1955 ( .A(n1629), .B(n1595), .Z(n1598) );
  XNOR U1956 ( .A(n1630), .B(n1592), .Z(n1595) );
  XNOR U1957 ( .A(n1631), .B(n1589), .Z(n1592) );
  XNOR U1958 ( .A(n1632), .B(n1586), .Z(n1589) );
  XNOR U1959 ( .A(n1633), .B(n1583), .Z(n1586) );
  XNOR U1960 ( .A(n1634), .B(n1580), .Z(n1583) );
  XNOR U1961 ( .A(n1635), .B(n1577), .Z(n1580) );
  XNOR U1962 ( .A(n1636), .B(n1574), .Z(n1577) );
  XNOR U1963 ( .A(n1637), .B(n1571), .Z(n1574) );
  XNOR U1964 ( .A(n1638), .B(n1568), .Z(n1571) );
  XNOR U1965 ( .A(n1639), .B(n1565), .Z(n1568) );
  XNOR U1966 ( .A(n1640), .B(n1562), .Z(n1565) );
  XNOR U1967 ( .A(n1641), .B(n1559), .Z(n1562) );
  XNOR U1968 ( .A(n1558), .B(n1642), .Z(n1559) );
  AND U1969 ( .A(g_input[0]), .B(e_input[21]), .Z(n1642) );
  NAND U1970 ( .A(e_input[20]), .B(g_input[1]), .Z(n1560) );
  NAND U1971 ( .A(e_input[19]), .B(g_input[2]), .Z(n1563) );
  NAND U1972 ( .A(e_input[18]), .B(g_input[3]), .Z(n1566) );
  NAND U1973 ( .A(e_input[17]), .B(g_input[4]), .Z(n1569) );
  NAND U1974 ( .A(e_input[16]), .B(g_input[5]), .Z(n1572) );
  NAND U1975 ( .A(e_input[15]), .B(g_input[6]), .Z(n1575) );
  NAND U1976 ( .A(e_input[14]), .B(g_input[7]), .Z(n1578) );
  NAND U1977 ( .A(g_input[8]), .B(e_input[13]), .Z(n1581) );
  NAND U1978 ( .A(g_input[9]), .B(e_input[12]), .Z(n1584) );
  NAND U1979 ( .A(e_input[11]), .B(g_input[10]), .Z(n1587) );
  NAND U1980 ( .A(g_input[11]), .B(e_input[10]), .Z(n1590) );
  NAND U1981 ( .A(g_input[12]), .B(e_input[9]), .Z(n1593) );
  NAND U1982 ( .A(g_input[13]), .B(e_input[8]), .Z(n1596) );
  NAND U1983 ( .A(g_input[14]), .B(e_input[7]), .Z(n1599) );
  NAND U1984 ( .A(g_input[15]), .B(e_input[6]), .Z(n1602) );
  NAND U1985 ( .A(g_input[16]), .B(e_input[5]), .Z(n1605) );
  NAND U1986 ( .A(g_input[17]), .B(e_input[4]), .Z(n1608) );
  XNOR U1987 ( .A(n1612), .B(n1611), .Z(n1624) );
  NAND U1988 ( .A(g_input[18]), .B(e_input[3]), .Z(n1611) );
  XOR U1989 ( .A(n1614), .B(n1615), .Z(n1623) );
  OR U1990 ( .A(n1700), .B(n1701), .Z(n1615) );
  ANDN U1991 ( .A(g_input[19]), .B(n786), .Z(n1614) );
  XNOR U1992 ( .A(n1622), .B(n1621), .Z(oi[20]) );
  XOR U1993 ( .A(n1701), .B(n1700), .Z(n1622) );
  NAND U1994 ( .A(g_input[20]), .B(e_input[0]), .Z(n1700) );
  XNOR U1995 ( .A(n1698), .B(n1699), .Z(n1701) );
  NAND U1996 ( .A(g_input[19]), .B(e_input[1]), .Z(n1699) );
  XNOR U1997 ( .A(n1705), .B(n1695), .Z(n1698) );
  XOR U1998 ( .A(n1706), .B(n1692), .Z(n1695) );
  XNOR U1999 ( .A(n1707), .B(n1689), .Z(n1692) );
  XNOR U2000 ( .A(n1708), .B(n1686), .Z(n1689) );
  XNOR U2001 ( .A(n1709), .B(n1683), .Z(n1686) );
  XNOR U2002 ( .A(n1710), .B(n1680), .Z(n1683) );
  XNOR U2003 ( .A(n1711), .B(n1677), .Z(n1680) );
  XNOR U2004 ( .A(n1712), .B(n1674), .Z(n1677) );
  XNOR U2005 ( .A(n1713), .B(n1671), .Z(n1674) );
  XNOR U2006 ( .A(n1714), .B(n1668), .Z(n1671) );
  XNOR U2007 ( .A(n1715), .B(n1665), .Z(n1668) );
  XNOR U2008 ( .A(n1716), .B(n1662), .Z(n1665) );
  XNOR U2009 ( .A(n1717), .B(n1659), .Z(n1662) );
  XNOR U2010 ( .A(n1718), .B(n1656), .Z(n1659) );
  XNOR U2011 ( .A(n1719), .B(n1653), .Z(n1656) );
  XNOR U2012 ( .A(n1720), .B(n1650), .Z(n1653) );
  XNOR U2013 ( .A(n1721), .B(n1647), .Z(n1650) );
  XNOR U2014 ( .A(n1722), .B(n1644), .Z(n1647) );
  XNOR U2015 ( .A(n1643), .B(n1723), .Z(n1644) );
  AND U2016 ( .A(g_input[0]), .B(e_input[20]), .Z(n1723) );
  NAND U2017 ( .A(e_input[19]), .B(g_input[1]), .Z(n1645) );
  NAND U2018 ( .A(e_input[18]), .B(g_input[2]), .Z(n1648) );
  NAND U2019 ( .A(e_input[17]), .B(g_input[3]), .Z(n1651) );
  NAND U2020 ( .A(e_input[16]), .B(g_input[4]), .Z(n1654) );
  NAND U2021 ( .A(e_input[15]), .B(g_input[5]), .Z(n1657) );
  NAND U2022 ( .A(e_input[14]), .B(g_input[6]), .Z(n1660) );
  NAND U2023 ( .A(e_input[13]), .B(g_input[7]), .Z(n1663) );
  NAND U2024 ( .A(g_input[8]), .B(e_input[12]), .Z(n1666) );
  NAND U2025 ( .A(g_input[9]), .B(e_input[11]), .Z(n1669) );
  NAND U2026 ( .A(e_input[10]), .B(g_input[10]), .Z(n1672) );
  NAND U2027 ( .A(g_input[11]), .B(e_input[9]), .Z(n1675) );
  NAND U2028 ( .A(g_input[12]), .B(e_input[8]), .Z(n1678) );
  NAND U2029 ( .A(g_input[13]), .B(e_input[7]), .Z(n1681) );
  NAND U2030 ( .A(g_input[14]), .B(e_input[6]), .Z(n1684) );
  NAND U2031 ( .A(g_input[15]), .B(e_input[5]), .Z(n1687) );
  NAND U2032 ( .A(g_input[16]), .B(e_input[4]), .Z(n1690) );
  XNOR U2033 ( .A(n1694), .B(n1693), .Z(n1706) );
  NAND U2034 ( .A(g_input[17]), .B(e_input[3]), .Z(n1693) );
  XOR U2035 ( .A(n1696), .B(n1697), .Z(n1705) );
  OR U2036 ( .A(n1778), .B(n1779), .Z(n1697) );
  ANDN U2037 ( .A(g_input[18]), .B(n786), .Z(n1696) );
  XNOR U2038 ( .A(n1780), .B(n1781), .Z(oi[1]) );
  XNOR U2039 ( .A(n1704), .B(n1703), .Z(oi[19]) );
  XOR U2040 ( .A(n1779), .B(n1778), .Z(n1704) );
  NAND U2041 ( .A(g_input[19]), .B(e_input[0]), .Z(n1778) );
  XNOR U2042 ( .A(n1776), .B(n1777), .Z(n1779) );
  NAND U2043 ( .A(g_input[18]), .B(e_input[1]), .Z(n1777) );
  XNOR U2044 ( .A(n1785), .B(n1773), .Z(n1776) );
  XOR U2045 ( .A(n1786), .B(n1770), .Z(n1773) );
  XNOR U2046 ( .A(n1787), .B(n1767), .Z(n1770) );
  XNOR U2047 ( .A(n1788), .B(n1764), .Z(n1767) );
  XNOR U2048 ( .A(n1789), .B(n1761), .Z(n1764) );
  XNOR U2049 ( .A(n1790), .B(n1758), .Z(n1761) );
  XNOR U2050 ( .A(n1791), .B(n1755), .Z(n1758) );
  XNOR U2051 ( .A(n1792), .B(n1752), .Z(n1755) );
  XNOR U2052 ( .A(n1793), .B(n1749), .Z(n1752) );
  XNOR U2053 ( .A(n1794), .B(n1746), .Z(n1749) );
  XNOR U2054 ( .A(n1795), .B(n1743), .Z(n1746) );
  XNOR U2055 ( .A(n1796), .B(n1740), .Z(n1743) );
  XNOR U2056 ( .A(n1797), .B(n1737), .Z(n1740) );
  XNOR U2057 ( .A(n1798), .B(n1734), .Z(n1737) );
  XNOR U2058 ( .A(n1799), .B(n1731), .Z(n1734) );
  XNOR U2059 ( .A(n1800), .B(n1728), .Z(n1731) );
  XNOR U2060 ( .A(n1801), .B(n1725), .Z(n1728) );
  XNOR U2061 ( .A(n1724), .B(n1802), .Z(n1725) );
  AND U2062 ( .A(g_input[0]), .B(e_input[19]), .Z(n1802) );
  NAND U2063 ( .A(e_input[18]), .B(g_input[1]), .Z(n1726) );
  NAND U2064 ( .A(e_input[17]), .B(g_input[2]), .Z(n1729) );
  NAND U2065 ( .A(e_input[16]), .B(g_input[3]), .Z(n1732) );
  NAND U2066 ( .A(e_input[15]), .B(g_input[4]), .Z(n1735) );
  NAND U2067 ( .A(e_input[14]), .B(g_input[5]), .Z(n1738) );
  NAND U2068 ( .A(e_input[13]), .B(g_input[6]), .Z(n1741) );
  NAND U2069 ( .A(e_input[12]), .B(g_input[7]), .Z(n1744) );
  NAND U2070 ( .A(g_input[8]), .B(e_input[11]), .Z(n1747) );
  NAND U2071 ( .A(g_input[9]), .B(e_input[10]), .Z(n1750) );
  NAND U2072 ( .A(g_input[10]), .B(e_input[9]), .Z(n1753) );
  NAND U2073 ( .A(g_input[11]), .B(e_input[8]), .Z(n1756) );
  NAND U2074 ( .A(g_input[12]), .B(e_input[7]), .Z(n1759) );
  NAND U2075 ( .A(g_input[13]), .B(e_input[6]), .Z(n1762) );
  NAND U2076 ( .A(g_input[14]), .B(e_input[5]), .Z(n1765) );
  NAND U2077 ( .A(g_input[15]), .B(e_input[4]), .Z(n1768) );
  XNOR U2078 ( .A(n1772), .B(n1771), .Z(n1786) );
  NAND U2079 ( .A(g_input[16]), .B(e_input[3]), .Z(n1771) );
  XOR U2080 ( .A(n1774), .B(n1775), .Z(n1785) );
  OR U2081 ( .A(n1854), .B(n1855), .Z(n1775) );
  ANDN U2082 ( .A(g_input[17]), .B(n786), .Z(n1774) );
  XNOR U2083 ( .A(n1784), .B(n1783), .Z(oi[18]) );
  XOR U2084 ( .A(n1855), .B(n1854), .Z(n1784) );
  NAND U2085 ( .A(g_input[18]), .B(e_input[0]), .Z(n1854) );
  XNOR U2086 ( .A(n1852), .B(n1853), .Z(n1855) );
  NAND U2087 ( .A(g_input[17]), .B(e_input[1]), .Z(n1853) );
  XNOR U2088 ( .A(n1859), .B(n1849), .Z(n1852) );
  XOR U2089 ( .A(n1860), .B(n1846), .Z(n1849) );
  XNOR U2090 ( .A(n1861), .B(n1843), .Z(n1846) );
  XNOR U2091 ( .A(n1862), .B(n1840), .Z(n1843) );
  XNOR U2092 ( .A(n1863), .B(n1837), .Z(n1840) );
  XNOR U2093 ( .A(n1864), .B(n1834), .Z(n1837) );
  XNOR U2094 ( .A(n1865), .B(n1831), .Z(n1834) );
  XNOR U2095 ( .A(n1866), .B(n1828), .Z(n1831) );
  XNOR U2096 ( .A(n1867), .B(n1825), .Z(n1828) );
  XNOR U2097 ( .A(n1868), .B(n1822), .Z(n1825) );
  XNOR U2098 ( .A(n1869), .B(n1819), .Z(n1822) );
  XNOR U2099 ( .A(n1870), .B(n1816), .Z(n1819) );
  XNOR U2100 ( .A(n1871), .B(n1813), .Z(n1816) );
  XNOR U2101 ( .A(n1872), .B(n1810), .Z(n1813) );
  XNOR U2102 ( .A(n1873), .B(n1807), .Z(n1810) );
  XNOR U2103 ( .A(n1874), .B(n1804), .Z(n1807) );
  XNOR U2104 ( .A(n1803), .B(n1875), .Z(n1804) );
  AND U2105 ( .A(g_input[0]), .B(e_input[18]), .Z(n1875) );
  NAND U2106 ( .A(e_input[17]), .B(g_input[1]), .Z(n1805) );
  NAND U2107 ( .A(e_input[16]), .B(g_input[2]), .Z(n1808) );
  NAND U2108 ( .A(e_input[15]), .B(g_input[3]), .Z(n1811) );
  NAND U2109 ( .A(e_input[14]), .B(g_input[4]), .Z(n1814) );
  NAND U2110 ( .A(e_input[13]), .B(g_input[5]), .Z(n1817) );
  NAND U2111 ( .A(e_input[12]), .B(g_input[6]), .Z(n1820) );
  NAND U2112 ( .A(e_input[11]), .B(g_input[7]), .Z(n1823) );
  NAND U2113 ( .A(g_input[8]), .B(e_input[10]), .Z(n1826) );
  NAND U2114 ( .A(g_input[9]), .B(e_input[9]), .Z(n1829) );
  NAND U2115 ( .A(g_input[10]), .B(e_input[8]), .Z(n1832) );
  NAND U2116 ( .A(g_input[11]), .B(e_input[7]), .Z(n1835) );
  NAND U2117 ( .A(g_input[12]), .B(e_input[6]), .Z(n1838) );
  NAND U2118 ( .A(g_input[13]), .B(e_input[5]), .Z(n1841) );
  NAND U2119 ( .A(g_input[14]), .B(e_input[4]), .Z(n1844) );
  XNOR U2120 ( .A(n1848), .B(n1847), .Z(n1860) );
  NAND U2121 ( .A(g_input[15]), .B(e_input[3]), .Z(n1847) );
  XOR U2122 ( .A(n1850), .B(n1851), .Z(n1859) );
  OR U2123 ( .A(n1924), .B(n1925), .Z(n1851) );
  ANDN U2124 ( .A(g_input[16]), .B(n786), .Z(n1850) );
  XNOR U2125 ( .A(n1858), .B(n1857), .Z(oi[17]) );
  XOR U2126 ( .A(n1925), .B(n1924), .Z(n1858) );
  NAND U2127 ( .A(g_input[17]), .B(e_input[0]), .Z(n1924) );
  XNOR U2128 ( .A(n1922), .B(n1923), .Z(n1925) );
  NAND U2129 ( .A(g_input[16]), .B(e_input[1]), .Z(n1923) );
  XNOR U2130 ( .A(n1929), .B(n1919), .Z(n1922) );
  XOR U2131 ( .A(n1930), .B(n1916), .Z(n1919) );
  XNOR U2132 ( .A(n1931), .B(n1913), .Z(n1916) );
  XNOR U2133 ( .A(n1932), .B(n1910), .Z(n1913) );
  XNOR U2134 ( .A(n1933), .B(n1907), .Z(n1910) );
  XNOR U2135 ( .A(n1934), .B(n1904), .Z(n1907) );
  XNOR U2136 ( .A(n1935), .B(n1901), .Z(n1904) );
  XNOR U2137 ( .A(n1936), .B(n1898), .Z(n1901) );
  XNOR U2138 ( .A(n1937), .B(n1895), .Z(n1898) );
  XNOR U2139 ( .A(n1938), .B(n1892), .Z(n1895) );
  XNOR U2140 ( .A(n1939), .B(n1889), .Z(n1892) );
  XNOR U2141 ( .A(n1940), .B(n1886), .Z(n1889) );
  XNOR U2142 ( .A(n1941), .B(n1883), .Z(n1886) );
  XNOR U2143 ( .A(n1942), .B(n1880), .Z(n1883) );
  XNOR U2144 ( .A(n1943), .B(n1877), .Z(n1880) );
  XNOR U2145 ( .A(n1876), .B(n1944), .Z(n1877) );
  AND U2146 ( .A(g_input[0]), .B(e_input[17]), .Z(n1944) );
  NAND U2147 ( .A(e_input[16]), .B(g_input[1]), .Z(n1878) );
  NAND U2148 ( .A(e_input[15]), .B(g_input[2]), .Z(n1881) );
  NAND U2149 ( .A(e_input[14]), .B(g_input[3]), .Z(n1884) );
  NAND U2150 ( .A(e_input[13]), .B(g_input[4]), .Z(n1887) );
  NAND U2151 ( .A(e_input[12]), .B(g_input[5]), .Z(n1890) );
  NAND U2152 ( .A(e_input[11]), .B(g_input[6]), .Z(n1893) );
  NAND U2153 ( .A(e_input[10]), .B(g_input[7]), .Z(n1896) );
  NAND U2154 ( .A(g_input[8]), .B(e_input[9]), .Z(n1899) );
  NAND U2155 ( .A(g_input[9]), .B(e_input[8]), .Z(n1902) );
  NAND U2156 ( .A(g_input[10]), .B(e_input[7]), .Z(n1905) );
  NAND U2157 ( .A(g_input[11]), .B(e_input[6]), .Z(n1908) );
  NAND U2158 ( .A(g_input[12]), .B(e_input[5]), .Z(n1911) );
  NAND U2159 ( .A(g_input[13]), .B(e_input[4]), .Z(n1914) );
  XNOR U2160 ( .A(n1918), .B(n1917), .Z(n1930) );
  NAND U2161 ( .A(g_input[14]), .B(e_input[3]), .Z(n1917) );
  XOR U2162 ( .A(n1920), .B(n1921), .Z(n1929) );
  OR U2163 ( .A(n1990), .B(n1991), .Z(n1921) );
  ANDN U2164 ( .A(g_input[15]), .B(n786), .Z(n1920) );
  XNOR U2165 ( .A(n1928), .B(n1927), .Z(oi[16]) );
  XOR U2166 ( .A(n1991), .B(n1990), .Z(n1928) );
  NAND U2167 ( .A(g_input[16]), .B(e_input[0]), .Z(n1990) );
  XNOR U2168 ( .A(n1988), .B(n1989), .Z(n1991) );
  NAND U2169 ( .A(g_input[15]), .B(e_input[1]), .Z(n1989) );
  XNOR U2170 ( .A(n1995), .B(n1985), .Z(n1988) );
  XOR U2171 ( .A(n1996), .B(n1982), .Z(n1985) );
  XNOR U2172 ( .A(n1997), .B(n1979), .Z(n1982) );
  XNOR U2173 ( .A(n1998), .B(n1976), .Z(n1979) );
  XNOR U2174 ( .A(n1999), .B(n1973), .Z(n1976) );
  XNOR U2175 ( .A(n2000), .B(n1970), .Z(n1973) );
  XNOR U2176 ( .A(n2001), .B(n1967), .Z(n1970) );
  XNOR U2177 ( .A(n2002), .B(n1964), .Z(n1967) );
  XNOR U2178 ( .A(n2003), .B(n1961), .Z(n1964) );
  XNOR U2179 ( .A(n2004), .B(n1958), .Z(n1961) );
  XNOR U2180 ( .A(n2005), .B(n1955), .Z(n1958) );
  XNOR U2181 ( .A(n2006), .B(n1952), .Z(n1955) );
  XNOR U2182 ( .A(n2007), .B(n1949), .Z(n1952) );
  XNOR U2183 ( .A(n2008), .B(n1946), .Z(n1949) );
  XNOR U2184 ( .A(n1945), .B(n2009), .Z(n1946) );
  AND U2185 ( .A(g_input[0]), .B(e_input[16]), .Z(n2009) );
  NAND U2186 ( .A(e_input[15]), .B(g_input[1]), .Z(n1947) );
  NAND U2187 ( .A(e_input[14]), .B(g_input[2]), .Z(n1950) );
  NAND U2188 ( .A(e_input[13]), .B(g_input[3]), .Z(n1953) );
  NAND U2189 ( .A(e_input[12]), .B(g_input[4]), .Z(n1956) );
  NAND U2190 ( .A(e_input[11]), .B(g_input[5]), .Z(n1959) );
  NAND U2191 ( .A(e_input[10]), .B(g_input[6]), .Z(n1962) );
  NAND U2192 ( .A(e_input[9]), .B(g_input[7]), .Z(n1965) );
  NAND U2193 ( .A(g_input[8]), .B(e_input[8]), .Z(n1968) );
  NAND U2194 ( .A(g_input[9]), .B(e_input[7]), .Z(n1971) );
  NAND U2195 ( .A(g_input[10]), .B(e_input[6]), .Z(n1974) );
  NAND U2196 ( .A(g_input[11]), .B(e_input[5]), .Z(n1977) );
  NAND U2197 ( .A(g_input[12]), .B(e_input[4]), .Z(n1980) );
  XNOR U2198 ( .A(n1984), .B(n1983), .Z(n1996) );
  NAND U2199 ( .A(g_input[13]), .B(e_input[3]), .Z(n1983) );
  XOR U2200 ( .A(n1986), .B(n1987), .Z(n1995) );
  OR U2201 ( .A(n2052), .B(n2053), .Z(n1987) );
  ANDN U2202 ( .A(g_input[14]), .B(n786), .Z(n1986) );
  XNOR U2203 ( .A(n1994), .B(n1993), .Z(oi[15]) );
  XOR U2204 ( .A(n2053), .B(n2052), .Z(n1994) );
  NAND U2205 ( .A(g_input[15]), .B(e_input[0]), .Z(n2052) );
  XNOR U2206 ( .A(n2050), .B(n2051), .Z(n2053) );
  NAND U2207 ( .A(g_input[14]), .B(e_input[1]), .Z(n2051) );
  XNOR U2208 ( .A(n2057), .B(n2047), .Z(n2050) );
  XOR U2209 ( .A(n2058), .B(n2044), .Z(n2047) );
  XNOR U2210 ( .A(n2059), .B(n2041), .Z(n2044) );
  XNOR U2211 ( .A(n2060), .B(n2038), .Z(n2041) );
  XNOR U2212 ( .A(n2061), .B(n2035), .Z(n2038) );
  XNOR U2213 ( .A(n2062), .B(n2032), .Z(n2035) );
  XNOR U2214 ( .A(n2063), .B(n2029), .Z(n2032) );
  XNOR U2215 ( .A(n2064), .B(n2026), .Z(n2029) );
  XNOR U2216 ( .A(n2065), .B(n2023), .Z(n2026) );
  XNOR U2217 ( .A(n2066), .B(n2020), .Z(n2023) );
  XNOR U2218 ( .A(n2067), .B(n2017), .Z(n2020) );
  XNOR U2219 ( .A(n2068), .B(n2014), .Z(n2017) );
  XNOR U2220 ( .A(n2069), .B(n2011), .Z(n2014) );
  XNOR U2221 ( .A(n2010), .B(n2070), .Z(n2011) );
  AND U2222 ( .A(g_input[0]), .B(e_input[15]), .Z(n2070) );
  NAND U2223 ( .A(e_input[14]), .B(g_input[1]), .Z(n2012) );
  NAND U2224 ( .A(e_input[13]), .B(g_input[2]), .Z(n2015) );
  NAND U2225 ( .A(e_input[12]), .B(g_input[3]), .Z(n2018) );
  NAND U2226 ( .A(e_input[11]), .B(g_input[4]), .Z(n2021) );
  NAND U2227 ( .A(e_input[10]), .B(g_input[5]), .Z(n2024) );
  NAND U2228 ( .A(e_input[9]), .B(g_input[6]), .Z(n2027) );
  NAND U2229 ( .A(e_input[8]), .B(g_input[7]), .Z(n2030) );
  NAND U2230 ( .A(g_input[8]), .B(e_input[7]), .Z(n2033) );
  NAND U2231 ( .A(g_input[9]), .B(e_input[6]), .Z(n2036) );
  NAND U2232 ( .A(g_input[10]), .B(e_input[5]), .Z(n2039) );
  NAND U2233 ( .A(g_input[11]), .B(e_input[4]), .Z(n2042) );
  XNOR U2234 ( .A(n2046), .B(n2045), .Z(n2058) );
  NAND U2235 ( .A(g_input[12]), .B(e_input[3]), .Z(n2045) );
  XOR U2236 ( .A(n2048), .B(n2049), .Z(n2057) );
  OR U2237 ( .A(n2110), .B(n2111), .Z(n2049) );
  ANDN U2238 ( .A(g_input[13]), .B(n786), .Z(n2048) );
  XNOR U2239 ( .A(n2056), .B(n2055), .Z(oi[14]) );
  XOR U2240 ( .A(n2111), .B(n2110), .Z(n2056) );
  NAND U2241 ( .A(g_input[14]), .B(e_input[0]), .Z(n2110) );
  XNOR U2242 ( .A(n2108), .B(n2109), .Z(n2111) );
  NAND U2243 ( .A(g_input[13]), .B(e_input[1]), .Z(n2109) );
  XNOR U2244 ( .A(n2115), .B(n2105), .Z(n2108) );
  XOR U2245 ( .A(n2116), .B(n2102), .Z(n2105) );
  XNOR U2246 ( .A(n2117), .B(n2099), .Z(n2102) );
  XNOR U2247 ( .A(n2118), .B(n2096), .Z(n2099) );
  XNOR U2248 ( .A(n2119), .B(n2093), .Z(n2096) );
  XNOR U2249 ( .A(n2120), .B(n2090), .Z(n2093) );
  XNOR U2250 ( .A(n2121), .B(n2087), .Z(n2090) );
  XNOR U2251 ( .A(n2122), .B(n2084), .Z(n2087) );
  XNOR U2252 ( .A(n2123), .B(n2081), .Z(n2084) );
  XNOR U2253 ( .A(n2124), .B(n2078), .Z(n2081) );
  XNOR U2254 ( .A(n2125), .B(n2075), .Z(n2078) );
  XNOR U2255 ( .A(n2126), .B(n2072), .Z(n2075) );
  XNOR U2256 ( .A(n2071), .B(n2127), .Z(n2072) );
  AND U2257 ( .A(g_input[0]), .B(e_input[14]), .Z(n2127) );
  NAND U2258 ( .A(e_input[13]), .B(g_input[1]), .Z(n2073) );
  NAND U2259 ( .A(e_input[12]), .B(g_input[2]), .Z(n2076) );
  NAND U2260 ( .A(e_input[11]), .B(g_input[3]), .Z(n2079) );
  NAND U2261 ( .A(e_input[10]), .B(g_input[4]), .Z(n2082) );
  NAND U2262 ( .A(e_input[9]), .B(g_input[5]), .Z(n2085) );
  NAND U2263 ( .A(e_input[8]), .B(g_input[6]), .Z(n2088) );
  NAND U2264 ( .A(e_input[7]), .B(g_input[7]), .Z(n2091) );
  NAND U2265 ( .A(g_input[8]), .B(e_input[6]), .Z(n2094) );
  NAND U2266 ( .A(g_input[9]), .B(e_input[5]), .Z(n2097) );
  NAND U2267 ( .A(g_input[10]), .B(e_input[4]), .Z(n2100) );
  XNOR U2268 ( .A(n2104), .B(n2103), .Z(n2116) );
  NAND U2269 ( .A(g_input[11]), .B(e_input[3]), .Z(n2103) );
  XOR U2270 ( .A(n2106), .B(n2107), .Z(n2115) );
  OR U2271 ( .A(n2164), .B(n2165), .Z(n2107) );
  ANDN U2272 ( .A(g_input[12]), .B(n786), .Z(n2106) );
  XNOR U2273 ( .A(n2114), .B(n2113), .Z(oi[13]) );
  XOR U2274 ( .A(n2165), .B(n2164), .Z(n2114) );
  NAND U2275 ( .A(g_input[13]), .B(e_input[0]), .Z(n2164) );
  XNOR U2276 ( .A(n2162), .B(n2163), .Z(n2165) );
  NAND U2277 ( .A(g_input[12]), .B(e_input[1]), .Z(n2163) );
  XNOR U2278 ( .A(n2169), .B(n2159), .Z(n2162) );
  XOR U2279 ( .A(n2170), .B(n2156), .Z(n2159) );
  XNOR U2280 ( .A(n2171), .B(n2153), .Z(n2156) );
  XNOR U2281 ( .A(n2172), .B(n2150), .Z(n2153) );
  XNOR U2282 ( .A(n2173), .B(n2147), .Z(n2150) );
  XNOR U2283 ( .A(n2174), .B(n2144), .Z(n2147) );
  XNOR U2284 ( .A(n2175), .B(n2141), .Z(n2144) );
  XNOR U2285 ( .A(n2176), .B(n2138), .Z(n2141) );
  XNOR U2286 ( .A(n2177), .B(n2135), .Z(n2138) );
  XNOR U2287 ( .A(n2178), .B(n2132), .Z(n2135) );
  XNOR U2288 ( .A(n2179), .B(n2129), .Z(n2132) );
  XNOR U2289 ( .A(n2128), .B(n2180), .Z(n2129) );
  AND U2290 ( .A(g_input[0]), .B(e_input[13]), .Z(n2180) );
  NAND U2291 ( .A(e_input[12]), .B(g_input[1]), .Z(n2130) );
  NAND U2292 ( .A(e_input[11]), .B(g_input[2]), .Z(n2133) );
  NAND U2293 ( .A(e_input[10]), .B(g_input[3]), .Z(n2136) );
  NAND U2294 ( .A(e_input[9]), .B(g_input[4]), .Z(n2139) );
  NAND U2295 ( .A(e_input[8]), .B(g_input[5]), .Z(n2142) );
  NAND U2296 ( .A(e_input[7]), .B(g_input[6]), .Z(n2145) );
  NAND U2297 ( .A(g_input[7]), .B(e_input[6]), .Z(n2148) );
  NAND U2298 ( .A(g_input[8]), .B(e_input[5]), .Z(n2151) );
  NAND U2299 ( .A(g_input[9]), .B(e_input[4]), .Z(n2154) );
  XNOR U2300 ( .A(n2158), .B(n2157), .Z(n2170) );
  NAND U2301 ( .A(g_input[10]), .B(e_input[3]), .Z(n2157) );
  XOR U2302 ( .A(n2160), .B(n2161), .Z(n2169) );
  OR U2303 ( .A(n2214), .B(n2215), .Z(n2161) );
  ANDN U2304 ( .A(g_input[11]), .B(n786), .Z(n2160) );
  XNOR U2305 ( .A(n2168), .B(n2167), .Z(oi[12]) );
  XOR U2306 ( .A(n2215), .B(n2214), .Z(n2168) );
  NAND U2307 ( .A(g_input[12]), .B(e_input[0]), .Z(n2214) );
  XNOR U2308 ( .A(n2212), .B(n2213), .Z(n2215) );
  NAND U2309 ( .A(g_input[11]), .B(e_input[1]), .Z(n2213) );
  XNOR U2310 ( .A(n2219), .B(n2209), .Z(n2212) );
  XOR U2311 ( .A(n2220), .B(n2206), .Z(n2209) );
  XNOR U2312 ( .A(n2221), .B(n2203), .Z(n2206) );
  XNOR U2313 ( .A(n2222), .B(n2200), .Z(n2203) );
  XNOR U2314 ( .A(n2223), .B(n2197), .Z(n2200) );
  XNOR U2315 ( .A(n2224), .B(n2194), .Z(n2197) );
  XNOR U2316 ( .A(n2225), .B(n2191), .Z(n2194) );
  XNOR U2317 ( .A(n2226), .B(n2188), .Z(n2191) );
  XNOR U2318 ( .A(n2227), .B(n2185), .Z(n2188) );
  XNOR U2319 ( .A(n2228), .B(n2182), .Z(n2185) );
  XNOR U2320 ( .A(n2181), .B(n2229), .Z(n2182) );
  AND U2321 ( .A(g_input[0]), .B(e_input[12]), .Z(n2229) );
  NAND U2322 ( .A(e_input[11]), .B(g_input[1]), .Z(n2183) );
  NAND U2323 ( .A(e_input[10]), .B(g_input[2]), .Z(n2186) );
  NAND U2324 ( .A(e_input[9]), .B(g_input[3]), .Z(n2189) );
  NAND U2325 ( .A(e_input[8]), .B(g_input[4]), .Z(n2192) );
  NAND U2326 ( .A(e_input[7]), .B(g_input[5]), .Z(n2195) );
  NAND U2327 ( .A(e_input[6]), .B(g_input[6]), .Z(n2198) );
  NAND U2328 ( .A(g_input[7]), .B(e_input[5]), .Z(n2201) );
  NAND U2329 ( .A(g_input[8]), .B(e_input[4]), .Z(n2204) );
  XNOR U2330 ( .A(n2208), .B(n2207), .Z(n2220) );
  NAND U2331 ( .A(g_input[9]), .B(e_input[3]), .Z(n2207) );
  XOR U2332 ( .A(n2210), .B(n2211), .Z(n2219) );
  OR U2333 ( .A(n2260), .B(n2261), .Z(n2211) );
  ANDN U2334 ( .A(g_input[10]), .B(n786), .Z(n2210) );
  XNOR U2335 ( .A(n2218), .B(n2217), .Z(oi[11]) );
  XOR U2336 ( .A(n2261), .B(n2260), .Z(n2218) );
  NAND U2337 ( .A(g_input[11]), .B(e_input[0]), .Z(n2260) );
  XNOR U2338 ( .A(n2258), .B(n2259), .Z(n2261) );
  NAND U2339 ( .A(g_input[10]), .B(e_input[1]), .Z(n2259) );
  XNOR U2340 ( .A(n2265), .B(n2255), .Z(n2258) );
  XOR U2341 ( .A(n2266), .B(n2252), .Z(n2255) );
  XNOR U2342 ( .A(n2267), .B(n2249), .Z(n2252) );
  XNOR U2343 ( .A(n2268), .B(n2246), .Z(n2249) );
  XNOR U2344 ( .A(n2269), .B(n2243), .Z(n2246) );
  XNOR U2345 ( .A(n2270), .B(n2240), .Z(n2243) );
  XNOR U2346 ( .A(n2271), .B(n2237), .Z(n2240) );
  XNOR U2347 ( .A(n2272), .B(n2234), .Z(n2237) );
  XNOR U2348 ( .A(n2273), .B(n2231), .Z(n2234) );
  XNOR U2349 ( .A(n2230), .B(n2274), .Z(n2231) );
  AND U2350 ( .A(g_input[0]), .B(e_input[11]), .Z(n2274) );
  NAND U2351 ( .A(e_input[10]), .B(g_input[1]), .Z(n2232) );
  NAND U2352 ( .A(e_input[9]), .B(g_input[2]), .Z(n2235) );
  NAND U2353 ( .A(e_input[8]), .B(g_input[3]), .Z(n2238) );
  NAND U2354 ( .A(e_input[7]), .B(g_input[4]), .Z(n2241) );
  NAND U2355 ( .A(e_input[6]), .B(g_input[5]), .Z(n2244) );
  NAND U2356 ( .A(g_input[6]), .B(e_input[5]), .Z(n2247) );
  NAND U2357 ( .A(g_input[7]), .B(e_input[4]), .Z(n2250) );
  XNOR U2358 ( .A(n2254), .B(n2253), .Z(n2266) );
  NAND U2359 ( .A(g_input[8]), .B(e_input[3]), .Z(n2253) );
  XOR U2360 ( .A(n2256), .B(n2257), .Z(n2265) );
  OR U2361 ( .A(n2302), .B(n2303), .Z(n2257) );
  XNOR U2362 ( .A(n2264), .B(n2263), .Z(oi[10]) );
  XNOR U2363 ( .A(n2305), .B(n2306), .Z(n379) );
  XOR U2364 ( .A(n2308), .B(n2309), .Z(n381) );
  XOR U2365 ( .A(n2311), .B(n2312), .Z(n383) );
  XOR U2366 ( .A(n2314), .B(n2315), .Z(n385) );
  XOR U2367 ( .A(n2317), .B(n2318), .Z(n387) );
  XOR U2368 ( .A(n2320), .B(n2321), .Z(n389) );
  XOR U2369 ( .A(n2323), .B(n2324), .Z(n391) );
  XNOR U2370 ( .A(n2326), .B(n2327), .Z(n788) );
  XOR U2371 ( .A(n2329), .B(n2330), .Z(n1781) );
  XNOR U2372 ( .A(n2328), .B(o[1]), .Z(n1780) );
  ANDN U2373 ( .A(o[0]), .B(n2331), .Z(n2328) );
  XOR U2374 ( .A(n2303), .B(n2302), .Z(n2264) );
  NAND U2375 ( .A(g_input[10]), .B(e_input[0]), .Z(n2302) );
  XNOR U2376 ( .A(n2300), .B(n2301), .Z(n2303) );
  NAND U2377 ( .A(g_input[9]), .B(e_input[1]), .Z(n2301) );
  XNOR U2378 ( .A(n2332), .B(n2297), .Z(n2300) );
  XOR U2379 ( .A(n2333), .B(n2294), .Z(n2297) );
  XNOR U2380 ( .A(n2334), .B(n2291), .Z(n2294) );
  XNOR U2381 ( .A(n2335), .B(n2288), .Z(n2291) );
  XNOR U2382 ( .A(n2336), .B(n2285), .Z(n2288) );
  XNOR U2383 ( .A(n2337), .B(n2282), .Z(n2285) );
  XNOR U2384 ( .A(n2338), .B(n2279), .Z(n2282) );
  XNOR U2385 ( .A(n2339), .B(n2276), .Z(n2279) );
  XNOR U2386 ( .A(n2275), .B(n2340), .Z(n2276) );
  AND U2387 ( .A(g_input[0]), .B(e_input[10]), .Z(n2340) );
  NAND U2388 ( .A(e_input[9]), .B(g_input[1]), .Z(n2277) );
  NAND U2389 ( .A(e_input[8]), .B(g_input[2]), .Z(n2280) );
  NAND U2390 ( .A(e_input[7]), .B(g_input[3]), .Z(n2283) );
  NAND U2391 ( .A(e_input[6]), .B(g_input[4]), .Z(n2286) );
  NAND U2392 ( .A(e_input[5]), .B(g_input[5]), .Z(n2289) );
  NAND U2393 ( .A(g_input[6]), .B(e_input[4]), .Z(n2292) );
  XNOR U2394 ( .A(n2296), .B(n2295), .Z(n2333) );
  NAND U2395 ( .A(g_input[7]), .B(e_input[3]), .Z(n2295) );
  XOR U2396 ( .A(n2298), .B(n2299), .Z(n2332) );
  OR U2397 ( .A(n2306), .B(n2305), .Z(n2299) );
  XNOR U2398 ( .A(n2363), .B(n2364), .Z(n2305) );
  NAND U2399 ( .A(g_input[8]), .B(e_input[1]), .Z(n2364) );
  XNOR U2400 ( .A(n2365), .B(n2360), .Z(n2363) );
  XOR U2401 ( .A(n2366), .B(n2357), .Z(n2360) );
  XNOR U2402 ( .A(n2367), .B(n2354), .Z(n2357) );
  XNOR U2403 ( .A(n2368), .B(n2351), .Z(n2354) );
  XNOR U2404 ( .A(n2369), .B(n2348), .Z(n2351) );
  XNOR U2405 ( .A(n2370), .B(n2345), .Z(n2348) );
  XNOR U2406 ( .A(n2371), .B(n2342), .Z(n2345) );
  XNOR U2407 ( .A(n2341), .B(n2372), .Z(n2342) );
  AND U2408 ( .A(g_input[0]), .B(e_input[9]), .Z(n2372) );
  NAND U2409 ( .A(e_input[8]), .B(g_input[1]), .Z(n2343) );
  NAND U2410 ( .A(e_input[7]), .B(g_input[2]), .Z(n2346) );
  NAND U2411 ( .A(e_input[6]), .B(g_input[3]), .Z(n2349) );
  NAND U2412 ( .A(e_input[5]), .B(g_input[4]), .Z(n2352) );
  NAND U2413 ( .A(g_input[5]), .B(e_input[4]), .Z(n2355) );
  XNOR U2414 ( .A(n2359), .B(n2358), .Z(n2366) );
  NAND U2415 ( .A(g_input[6]), .B(e_input[3]), .Z(n2358) );
  XOR U2416 ( .A(n2361), .B(n2362), .Z(n2365) );
  OR U2417 ( .A(n2309), .B(n2308), .Z(n2362) );
  XNOR U2418 ( .A(n2392), .B(n2393), .Z(n2308) );
  NAND U2419 ( .A(g_input[7]), .B(e_input[1]), .Z(n2393) );
  XNOR U2420 ( .A(n2394), .B(n2389), .Z(n2392) );
  XOR U2421 ( .A(n2395), .B(n2386), .Z(n2389) );
  XNOR U2422 ( .A(n2396), .B(n2383), .Z(n2386) );
  XNOR U2423 ( .A(n2397), .B(n2380), .Z(n2383) );
  XNOR U2424 ( .A(n2398), .B(n2377), .Z(n2380) );
  XNOR U2425 ( .A(n2399), .B(n2374), .Z(n2377) );
  XNOR U2426 ( .A(n2373), .B(n2400), .Z(n2374) );
  AND U2427 ( .A(g_input[0]), .B(e_input[8]), .Z(n2400) );
  NAND U2428 ( .A(e_input[7]), .B(g_input[1]), .Z(n2375) );
  NAND U2429 ( .A(e_input[6]), .B(g_input[2]), .Z(n2378) );
  NAND U2430 ( .A(e_input[5]), .B(g_input[3]), .Z(n2381) );
  NAND U2431 ( .A(e_input[4]), .B(g_input[4]), .Z(n2384) );
  XNOR U2432 ( .A(n2388), .B(n2387), .Z(n2395) );
  NAND U2433 ( .A(g_input[5]), .B(e_input[3]), .Z(n2387) );
  XOR U2434 ( .A(n2390), .B(n2391), .Z(n2394) );
  OR U2435 ( .A(n2312), .B(n2311), .Z(n2391) );
  XNOR U2436 ( .A(n2417), .B(n2418), .Z(n2311) );
  NAND U2437 ( .A(g_input[6]), .B(e_input[1]), .Z(n2418) );
  XNOR U2438 ( .A(n2419), .B(n2414), .Z(n2417) );
  XOR U2439 ( .A(n2420), .B(n2411), .Z(n2414) );
  XNOR U2440 ( .A(n2421), .B(n2408), .Z(n2411) );
  XNOR U2441 ( .A(n2422), .B(n2405), .Z(n2408) );
  XNOR U2442 ( .A(n2423), .B(n2402), .Z(n2405) );
  XNOR U2443 ( .A(n2401), .B(n2424), .Z(n2402) );
  AND U2444 ( .A(g_input[0]), .B(e_input[7]), .Z(n2424) );
  NAND U2445 ( .A(e_input[6]), .B(g_input[1]), .Z(n2403) );
  NAND U2446 ( .A(e_input[5]), .B(g_input[2]), .Z(n2406) );
  NAND U2447 ( .A(e_input[4]), .B(g_input[3]), .Z(n2409) );
  XNOR U2448 ( .A(n2413), .B(n2412), .Z(n2420) );
  NAND U2449 ( .A(g_input[4]), .B(e_input[3]), .Z(n2412) );
  XOR U2450 ( .A(n2415), .B(n2416), .Z(n2419) );
  OR U2451 ( .A(n2315), .B(n2314), .Z(n2416) );
  XNOR U2452 ( .A(n2438), .B(n2439), .Z(n2314) );
  NAND U2453 ( .A(g_input[5]), .B(e_input[1]), .Z(n2439) );
  XNOR U2454 ( .A(n2440), .B(n2435), .Z(n2438) );
  XOR U2455 ( .A(n2441), .B(n2432), .Z(n2435) );
  XNOR U2456 ( .A(n2442), .B(n2429), .Z(n2432) );
  XNOR U2457 ( .A(n2443), .B(n2426), .Z(n2429) );
  XNOR U2458 ( .A(n2425), .B(n2444), .Z(n2426) );
  AND U2459 ( .A(g_input[0]), .B(e_input[6]), .Z(n2444) );
  NAND U2460 ( .A(e_input[5]), .B(g_input[1]), .Z(n2427) );
  NAND U2461 ( .A(e_input[4]), .B(g_input[2]), .Z(n2430) );
  XNOR U2462 ( .A(n2434), .B(n2433), .Z(n2441) );
  NAND U2463 ( .A(e_input[3]), .B(g_input[3]), .Z(n2433) );
  XOR U2464 ( .A(n2436), .B(n2437), .Z(n2440) );
  OR U2465 ( .A(n2318), .B(n2317), .Z(n2437) );
  XNOR U2466 ( .A(n2455), .B(n2456), .Z(n2317) );
  NAND U2467 ( .A(g_input[4]), .B(e_input[1]), .Z(n2456) );
  XNOR U2468 ( .A(n2457), .B(n2452), .Z(n2455) );
  XOR U2469 ( .A(n2458), .B(n2449), .Z(n2452) );
  XNOR U2470 ( .A(n2459), .B(n2446), .Z(n2449) );
  XNOR U2471 ( .A(n2445), .B(n2460), .Z(n2446) );
  AND U2472 ( .A(g_input[0]), .B(e_input[5]), .Z(n2460) );
  NAND U2473 ( .A(e_input[4]), .B(g_input[1]), .Z(n2447) );
  XNOR U2474 ( .A(n2451), .B(n2450), .Z(n2458) );
  NAND U2475 ( .A(e_input[3]), .B(g_input[2]), .Z(n2450) );
  XOR U2476 ( .A(n2453), .B(n2454), .Z(n2457) );
  OR U2477 ( .A(n2321), .B(n2320), .Z(n2454) );
  XNOR U2478 ( .A(n2468), .B(n2469), .Z(n2320) );
  NAND U2479 ( .A(g_input[3]), .B(e_input[1]), .Z(n2469) );
  XNOR U2480 ( .A(n2470), .B(n2465), .Z(n2468) );
  XOR U2481 ( .A(n2471), .B(n2462), .Z(n2465) );
  XNOR U2482 ( .A(n2461), .B(n2472), .Z(n2462) );
  AND U2483 ( .A(g_input[0]), .B(e_input[4]), .Z(n2472) );
  XNOR U2484 ( .A(n2464), .B(n2463), .Z(n2471) );
  NAND U2485 ( .A(e_input[3]), .B(g_input[1]), .Z(n2463) );
  IV U2486 ( .A(n2476), .Z(n2479) );
  XOR U2487 ( .A(n2466), .B(n2467), .Z(n2470) );
  OR U2488 ( .A(n2324), .B(n2323), .Z(n2467) );
  XNOR U2489 ( .A(n2477), .B(n2478), .Z(n2323) );
  NAND U2490 ( .A(g_input[2]), .B(e_input[1]), .Z(n2478) );
  XNOR U2491 ( .A(n2480), .B(n2474), .Z(n2477) );
  XOR U2492 ( .A(n2473), .B(n2481), .Z(n2474) );
  AND U2493 ( .A(g_input[0]), .B(e_input[3]), .Z(n2481) );
  ANDN U2494 ( .A(n2482), .B(n2483), .Z(n2473) );
  NANDN U2495 ( .B(n2484), .A(n2485), .Z(n2482) );
  XNOR U2496 ( .A(n2475), .B(n2476), .Z(n2480) );
  ANDN U2497 ( .A(n2326), .B(n2327), .Z(n2476) );
  NAND U2498 ( .A(g_input[2]), .B(e_input[0]), .Z(n2327) );
  NAND U2499 ( .A(g_input[1]), .B(e_input[1]), .Z(n2484) );
  NOR U2500 ( .A(n2329), .B(n2330), .Z(n2483) );
  NAND U2501 ( .A(e_input[1]), .B(g_input[0]), .Z(n2330) );
  NAND U2502 ( .A(e_input[0]), .B(g_input[1]), .Z(n2329) );
  NAND U2503 ( .A(e_input[2]), .B(g_input[0]), .Z(n2486) );
  ANDN U2504 ( .A(g_input[1]), .B(n786), .Z(n2475) );
  NAND U2505 ( .A(g_input[3]), .B(e_input[0]), .Z(n2324) );
  ANDN U2506 ( .A(g_input[2]), .B(n786), .Z(n2466) );
  NAND U2507 ( .A(g_input[4]), .B(e_input[0]), .Z(n2321) );
  ANDN U2508 ( .A(g_input[3]), .B(n786), .Z(n2453) );
  NAND U2509 ( .A(g_input[5]), .B(e_input[0]), .Z(n2318) );
  ANDN U2510 ( .A(g_input[4]), .B(n786), .Z(n2436) );
  NAND U2511 ( .A(g_input[6]), .B(e_input[0]), .Z(n2315) );
  ANDN U2512 ( .A(g_input[5]), .B(n786), .Z(n2415) );
  NAND U2513 ( .A(g_input[7]), .B(e_input[0]), .Z(n2312) );
  ANDN U2514 ( .A(g_input[6]), .B(n786), .Z(n2390) );
  NAND U2515 ( .A(g_input[8]), .B(e_input[0]), .Z(n2309) );
  ANDN U2516 ( .A(g_input[7]), .B(n786), .Z(n2361) );
  IV U2517 ( .A(e_input[2]), .Z(n786) );
  NAND U2518 ( .A(g_input[9]), .B(e_input[0]), .Z(n2306) );
  XNOR U2519 ( .A(o[0]), .B(n2331), .Z(oi[0]) );
  NAND U2520 ( .A(g_input[0]), .B(e_input[0]), .Z(n2331) );
endmodule

