
module stackMachine_N64 ( clk, rst, x, opcode, o );
  input [63:0] x;
  input [2:0] opcode;
  output [63:0] o;
  input clk, rst;
  wire   \stack[7][63] , \stack[7][62] , \stack[7][61] , \stack[7][60] ,
         \stack[7][59] , \stack[7][58] , \stack[7][57] , \stack[7][56] ,
         \stack[7][55] , \stack[7][54] , \stack[7][53] , \stack[7][52] ,
         \stack[7][51] , \stack[7][50] , \stack[7][49] , \stack[7][48] ,
         \stack[7][47] , \stack[7][46] , \stack[7][45] , \stack[7][44] ,
         \stack[7][43] , \stack[7][42] , \stack[7][41] , \stack[7][40] ,
         \stack[7][39] , \stack[7][38] , \stack[7][37] , \stack[7][36] ,
         \stack[7][35] , \stack[7][34] , \stack[7][33] , \stack[7][32] ,
         \stack[7][31] , \stack[7][30] , \stack[7][29] , \stack[7][28] ,
         \stack[7][27] , \stack[7][26] , \stack[7][25] , \stack[7][24] ,
         \stack[7][23] , \stack[7][22] , \stack[7][21] , \stack[7][20] ,
         \stack[7][19] , \stack[7][18] , \stack[7][17] , \stack[7][16] ,
         \stack[7][15] , \stack[7][14] , \stack[7][13] , \stack[7][12] ,
         \stack[7][11] , \stack[7][10] , \stack[7][9] , \stack[7][8] ,
         \stack[7][7] , \stack[7][6] , \stack[7][5] , \stack[7][4] ,
         \stack[7][3] , \stack[7][2] , \stack[7][1] , \stack[7][0] ,
         \stack[6][63] , \stack[6][62] , \stack[6][61] , \stack[6][60] ,
         \stack[6][59] , \stack[6][58] , \stack[6][57] , \stack[6][56] ,
         \stack[6][55] , \stack[6][54] , \stack[6][53] , \stack[6][52] ,
         \stack[6][51] , \stack[6][50] , \stack[6][49] , \stack[6][48] ,
         \stack[6][47] , \stack[6][46] , \stack[6][45] , \stack[6][44] ,
         \stack[6][43] , \stack[6][42] , \stack[6][41] , \stack[6][40] ,
         \stack[6][39] , \stack[6][38] , \stack[6][37] , \stack[6][36] ,
         \stack[6][35] , \stack[6][34] , \stack[6][33] , \stack[6][32] ,
         \stack[6][31] , \stack[6][30] , \stack[6][29] , \stack[6][28] ,
         \stack[6][27] , \stack[6][26] , \stack[6][25] , \stack[6][24] ,
         \stack[6][23] , \stack[6][22] , \stack[6][21] , \stack[6][20] ,
         \stack[6][19] , \stack[6][18] , \stack[6][17] , \stack[6][16] ,
         \stack[6][15] , \stack[6][14] , \stack[6][13] , \stack[6][12] ,
         \stack[6][11] , \stack[6][10] , \stack[6][9] , \stack[6][8] ,
         \stack[6][7] , \stack[6][6] , \stack[6][5] , \stack[6][4] ,
         \stack[6][3] , \stack[6][2] , \stack[6][1] , \stack[6][0] ,
         \stack[5][63] , \stack[5][62] , \stack[5][61] , \stack[5][60] ,
         \stack[5][59] , \stack[5][58] , \stack[5][57] , \stack[5][56] ,
         \stack[5][55] , \stack[5][54] , \stack[5][53] , \stack[5][52] ,
         \stack[5][51] , \stack[5][50] , \stack[5][49] , \stack[5][48] ,
         \stack[5][47] , \stack[5][46] , \stack[5][45] , \stack[5][44] ,
         \stack[5][43] , \stack[5][42] , \stack[5][41] , \stack[5][40] ,
         \stack[5][39] , \stack[5][38] , \stack[5][37] , \stack[5][36] ,
         \stack[5][35] , \stack[5][34] , \stack[5][33] , \stack[5][32] ,
         \stack[5][31] , \stack[5][30] , \stack[5][29] , \stack[5][28] ,
         \stack[5][27] , \stack[5][26] , \stack[5][25] , \stack[5][24] ,
         \stack[5][23] , \stack[5][22] , \stack[5][21] , \stack[5][20] ,
         \stack[5][19] , \stack[5][18] , \stack[5][17] , \stack[5][16] ,
         \stack[5][15] , \stack[5][14] , \stack[5][13] , \stack[5][12] ,
         \stack[5][11] , \stack[5][10] , \stack[5][9] , \stack[5][8] ,
         \stack[5][7] , \stack[5][6] , \stack[5][5] , \stack[5][4] ,
         \stack[5][3] , \stack[5][2] , \stack[5][1] , \stack[5][0] ,
         \stack[4][63] , \stack[4][62] , \stack[4][61] , \stack[4][60] ,
         \stack[4][59] , \stack[4][58] , \stack[4][57] , \stack[4][56] ,
         \stack[4][55] , \stack[4][54] , \stack[4][53] , \stack[4][52] ,
         \stack[4][51] , \stack[4][50] , \stack[4][49] , \stack[4][48] ,
         \stack[4][47] , \stack[4][46] , \stack[4][45] , \stack[4][44] ,
         \stack[4][43] , \stack[4][42] , \stack[4][41] , \stack[4][40] ,
         \stack[4][39] , \stack[4][38] , \stack[4][37] , \stack[4][36] ,
         \stack[4][35] , \stack[4][34] , \stack[4][33] , \stack[4][32] ,
         \stack[4][31] , \stack[4][30] , \stack[4][29] , \stack[4][28] ,
         \stack[4][27] , \stack[4][26] , \stack[4][25] , \stack[4][24] ,
         \stack[4][23] , \stack[4][22] , \stack[4][21] , \stack[4][20] ,
         \stack[4][19] , \stack[4][18] , \stack[4][17] , \stack[4][16] ,
         \stack[4][15] , \stack[4][14] , \stack[4][13] , \stack[4][12] ,
         \stack[4][11] , \stack[4][10] , \stack[4][9] , \stack[4][8] ,
         \stack[4][7] , \stack[4][6] , \stack[4][5] , \stack[4][4] ,
         \stack[4][3] , \stack[4][2] , \stack[4][1] , \stack[4][0] ,
         \stack[3][63] , \stack[3][62] , \stack[3][61] , \stack[3][60] ,
         \stack[3][59] , \stack[3][58] , \stack[3][57] , \stack[3][56] ,
         \stack[3][55] , \stack[3][54] , \stack[3][53] , \stack[3][52] ,
         \stack[3][51] , \stack[3][50] , \stack[3][49] , \stack[3][48] ,
         \stack[3][47] , \stack[3][46] , \stack[3][45] , \stack[3][44] ,
         \stack[3][43] , \stack[3][42] , \stack[3][41] , \stack[3][40] ,
         \stack[3][39] , \stack[3][38] , \stack[3][37] , \stack[3][36] ,
         \stack[3][35] , \stack[3][34] , \stack[3][33] , \stack[3][32] ,
         \stack[3][31] , \stack[3][30] , \stack[3][29] , \stack[3][28] ,
         \stack[3][27] , \stack[3][26] , \stack[3][25] , \stack[3][24] ,
         \stack[3][23] , \stack[3][22] , \stack[3][21] , \stack[3][20] ,
         \stack[3][19] , \stack[3][18] , \stack[3][17] , \stack[3][16] ,
         \stack[3][15] , \stack[3][14] , \stack[3][13] , \stack[3][12] ,
         \stack[3][11] , \stack[3][10] , \stack[3][9] , \stack[3][8] ,
         \stack[3][7] , \stack[3][6] , \stack[3][5] , \stack[3][4] ,
         \stack[3][3] , \stack[3][2] , \stack[3][1] , \stack[3][0] ,
         \stack[2][63] , \stack[2][62] , \stack[2][61] , \stack[2][60] ,
         \stack[2][59] , \stack[2][58] , \stack[2][57] , \stack[2][56] ,
         \stack[2][55] , \stack[2][54] , \stack[2][53] , \stack[2][52] ,
         \stack[2][51] , \stack[2][50] , \stack[2][49] , \stack[2][48] ,
         \stack[2][47] , \stack[2][46] , \stack[2][45] , \stack[2][44] ,
         \stack[2][43] , \stack[2][42] , \stack[2][41] , \stack[2][40] ,
         \stack[2][39] , \stack[2][38] , \stack[2][37] , \stack[2][36] ,
         \stack[2][35] , \stack[2][34] , \stack[2][33] , \stack[2][32] ,
         \stack[2][31] , \stack[2][30] , \stack[2][29] , \stack[2][28] ,
         \stack[2][27] , \stack[2][26] , \stack[2][25] , \stack[2][24] ,
         \stack[2][23] , \stack[2][22] , \stack[2][21] , \stack[2][20] ,
         \stack[2][19] , \stack[2][18] , \stack[2][17] , \stack[2][16] ,
         \stack[2][15] , \stack[2][14] , \stack[2][13] , \stack[2][12] ,
         \stack[2][11] , \stack[2][10] , \stack[2][9] , \stack[2][8] ,
         \stack[2][7] , \stack[2][6] , \stack[2][5] , \stack[2][4] ,
         \stack[2][3] , \stack[2][2] , \stack[2][1] , \stack[2][0] ,
         \stack[1][63] , \stack[1][62] , \stack[1][61] , \stack[1][60] ,
         \stack[1][59] , \stack[1][58] , \stack[1][57] , \stack[1][56] ,
         \stack[1][55] , \stack[1][54] , \stack[1][53] , \stack[1][52] ,
         \stack[1][51] , \stack[1][50] , \stack[1][49] , \stack[1][48] ,
         \stack[1][47] , \stack[1][46] , \stack[1][45] , \stack[1][44] ,
         \stack[1][43] , \stack[1][42] , \stack[1][41] , \stack[1][40] ,
         \stack[1][39] , \stack[1][38] , \stack[1][37] , \stack[1][36] ,
         \stack[1][35] , \stack[1][34] , \stack[1][33] , \stack[1][32] ,
         \stack[1][31] , \stack[1][30] , \stack[1][29] , \stack[1][28] ,
         \stack[1][27] , \stack[1][26] , \stack[1][25] , \stack[1][24] ,
         \stack[1][23] , \stack[1][22] , \stack[1][21] , \stack[1][20] ,
         \stack[1][19] , \stack[1][18] , \stack[1][17] , \stack[1][16] ,
         \stack[1][15] , \stack[1][14] , \stack[1][13] , \stack[1][12] ,
         \stack[1][11] , \stack[1][10] , \stack[1][9] , \stack[1][8] ,
         \stack[1][7] , \stack[1][6] , \stack[1][5] , \stack[1][4] ,
         \stack[1][3] , \stack[1][2] , \stack[1][1] , \stack[1][0] ,
         \C3/DATA5_0 , \C3/DATA5_1 , \C3/DATA5_2 , \C3/DATA5_3 , \C3/DATA5_4 ,
         \C3/DATA5_5 , \C3/DATA5_6 , \C3/DATA5_7 , \C3/DATA5_8 , \C3/DATA5_9 ,
         \C3/DATA5_10 , \C3/DATA5_11 , \C3/DATA5_12 , \C3/DATA5_13 ,
         \C3/DATA5_14 , \C3/DATA5_15 , \C3/DATA5_16 , \C3/DATA5_17 ,
         \C3/DATA5_18 , \C3/DATA5_19 , \C3/DATA5_20 , \C3/DATA5_21 ,
         \C3/DATA5_22 , \C3/DATA5_23 , \C3/DATA5_24 , \C3/DATA5_25 ,
         \C3/DATA5_26 , \C3/DATA5_27 , \C3/DATA5_28 , \C3/DATA5_29 ,
         \C3/DATA5_30 , \C3/DATA5_31 , \C3/DATA5_32 , \C3/DATA5_33 ,
         \C3/DATA5_34 , \C3/DATA5_35 , \C3/DATA5_36 , \C3/DATA5_37 ,
         \C3/DATA5_38 , \C3/DATA5_39 , \C3/DATA5_40 , \C3/DATA5_41 ,
         \C3/DATA5_42 , \C3/DATA5_43 , \C3/DATA5_44 , \C3/DATA5_45 ,
         \C3/DATA5_46 , \C3/DATA5_47 , \C3/DATA5_48 , \C3/DATA5_49 ,
         \C3/DATA5_50 , \C3/DATA5_51 , \C3/DATA5_52 , \C3/DATA5_53 ,
         \C3/DATA5_54 , \C3/DATA5_55 , \C3/DATA5_56 , \C3/DATA5_57 ,
         \C3/DATA5_58 , \C3/DATA5_59 , \C3/DATA5_60 , \C3/DATA5_61 ,
         \C3/DATA5_62 , \C3/DATA5_63 , n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, \C1/Z_0 ,
         \U1/RSOP_16/C3/Z_63 , \U1/RSOP_16/C3/Z_62 , \U1/RSOP_16/C3/Z_61 ,
         \U1/RSOP_16/C3/Z_60 , \U1/RSOP_16/C3/Z_59 , \U1/RSOP_16/C3/Z_58 ,
         \U1/RSOP_16/C3/Z_57 , \U1/RSOP_16/C3/Z_56 , \U1/RSOP_16/C3/Z_55 ,
         \U1/RSOP_16/C3/Z_54 , \U1/RSOP_16/C3/Z_53 , \U1/RSOP_16/C3/Z_52 ,
         \U1/RSOP_16/C3/Z_51 , \U1/RSOP_16/C3/Z_50 , \U1/RSOP_16/C3/Z_49 ,
         \U1/RSOP_16/C3/Z_48 , \U1/RSOP_16/C3/Z_47 , \U1/RSOP_16/C3/Z_46 ,
         \U1/RSOP_16/C3/Z_45 , \U1/RSOP_16/C3/Z_44 , \U1/RSOP_16/C3/Z_43 ,
         \U1/RSOP_16/C3/Z_42 , \U1/RSOP_16/C3/Z_41 , \U1/RSOP_16/C3/Z_40 ,
         \U1/RSOP_16/C3/Z_39 , \U1/RSOP_16/C3/Z_38 , \U1/RSOP_16/C3/Z_37 ,
         \U1/RSOP_16/C3/Z_36 , \U1/RSOP_16/C3/Z_35 , \U1/RSOP_16/C3/Z_34 ,
         \U1/RSOP_16/C3/Z_33 , \U1/RSOP_16/C3/Z_32 , \U1/RSOP_16/C3/Z_31 ,
         \U1/RSOP_16/C3/Z_30 , \U1/RSOP_16/C3/Z_29 , \U1/RSOP_16/C3/Z_28 ,
         \U1/RSOP_16/C3/Z_27 , \U1/RSOP_16/C3/Z_26 , \U1/RSOP_16/C3/Z_25 ,
         \U1/RSOP_16/C3/Z_24 , \U1/RSOP_16/C3/Z_23 , \U1/RSOP_16/C3/Z_22 ,
         \U1/RSOP_16/C3/Z_21 , \U1/RSOP_16/C3/Z_20 , \U1/RSOP_16/C3/Z_19 ,
         \U1/RSOP_16/C3/Z_18 , \U1/RSOP_16/C3/Z_17 , \U1/RSOP_16/C3/Z_16 ,
         \U1/RSOP_16/C3/Z_15 , \U1/RSOP_16/C3/Z_14 , \U1/RSOP_16/C3/Z_13 ,
         \U1/RSOP_16/C3/Z_12 , \U1/RSOP_16/C3/Z_11 , \U1/RSOP_16/C3/Z_10 ,
         \U1/RSOP_16/C3/Z_9 , \U1/RSOP_16/C3/Z_8 , \U1/RSOP_16/C3/Z_7 ,
         \U1/RSOP_16/C3/Z_6 , \U1/RSOP_16/C3/Z_5 , \U1/RSOP_16/C3/Z_4 ,
         \U1/RSOP_16/C3/Z_3 , \U1/RSOP_16/C3/Z_2 , \U1/RSOP_16/C3/Z_1 ,
         \U1/RSOP_16/C3/Z_0 , \U1/RSOP_16/C2/Z_63 , \U1/RSOP_16/C2/Z_62 ,
         \U1/RSOP_16/C2/Z_61 , \U1/RSOP_16/C2/Z_60 , \U1/RSOP_16/C2/Z_59 ,
         \U1/RSOP_16/C2/Z_58 , \U1/RSOP_16/C2/Z_57 , \U1/RSOP_16/C2/Z_56 ,
         \U1/RSOP_16/C2/Z_55 , \U1/RSOP_16/C2/Z_54 , \U1/RSOP_16/C2/Z_53 ,
         \U1/RSOP_16/C2/Z_52 , \U1/RSOP_16/C2/Z_51 , \U1/RSOP_16/C2/Z_50 ,
         \U1/RSOP_16/C2/Z_49 , \U1/RSOP_16/C2/Z_48 , \U1/RSOP_16/C2/Z_47 ,
         \U1/RSOP_16/C2/Z_46 , \U1/RSOP_16/C2/Z_45 , \U1/RSOP_16/C2/Z_44 ,
         \U1/RSOP_16/C2/Z_43 , \U1/RSOP_16/C2/Z_42 , \U1/RSOP_16/C2/Z_41 ,
         \U1/RSOP_16/C2/Z_40 , \U1/RSOP_16/C2/Z_39 , \U1/RSOP_16/C2/Z_38 ,
         \U1/RSOP_16/C2/Z_37 , \U1/RSOP_16/C2/Z_36 , \U1/RSOP_16/C2/Z_35 ,
         \U1/RSOP_16/C2/Z_34 , \U1/RSOP_16/C2/Z_33 , \U1/RSOP_16/C2/Z_32 ,
         \U1/RSOP_16/C2/Z_31 , \U1/RSOP_16/C2/Z_30 , \U1/RSOP_16/C2/Z_29 ,
         \U1/RSOP_16/C2/Z_28 , \U1/RSOP_16/C2/Z_27 , \U1/RSOP_16/C2/Z_26 ,
         \U1/RSOP_16/C2/Z_25 , \U1/RSOP_16/C2/Z_24 , \U1/RSOP_16/C2/Z_23 ,
         \U1/RSOP_16/C2/Z_22 , \U1/RSOP_16/C2/Z_21 , \U1/RSOP_16/C2/Z_20 ,
         \U1/RSOP_16/C2/Z_19 , \U1/RSOP_16/C2/Z_18 , \U1/RSOP_16/C2/Z_17 ,
         \U1/RSOP_16/C2/Z_16 , \U1/RSOP_16/C2/Z_15 , \U1/RSOP_16/C2/Z_14 ,
         \U1/RSOP_16/C2/Z_13 , \U1/RSOP_16/C2/Z_12 , \U1/RSOP_16/C2/Z_11 ,
         \U1/RSOP_16/C2/Z_10 , \U1/RSOP_16/C2/Z_9 , \U1/RSOP_16/C2/Z_8 ,
         \U1/RSOP_16/C2/Z_7 , \U1/RSOP_16/C2/Z_6 , \U1/RSOP_16/C2/Z_5 ,
         \U1/RSOP_16/C2/Z_4 , \U1/RSOP_16/C2/Z_3 , \U1/RSOP_16/C2/Z_2 ,
         \U1/RSOP_16/C2/Z_1 , \U1/RSOP_16/C2/Z_0 , \DP_OP_25_64_8855/n656 ,
         \DP_OP_25_64_8855/n655 , \DP_OP_25_64_8855/n654 ,
         \DP_OP_25_64_8855/n653 , \DP_OP_25_64_8855/n652 ,
         \DP_OP_25_64_8855/n651 , \DP_OP_25_64_8855/n650 ,
         \DP_OP_25_64_8855/n649 , \DP_OP_25_64_8855/n648 ,
         \DP_OP_25_64_8855/n647 , \DP_OP_25_64_8855/n646 ,
         \DP_OP_25_64_8855/n645 , \DP_OP_25_64_8855/n644 ,
         \DP_OP_25_64_8855/n643 , \DP_OP_25_64_8855/n642 ,
         \DP_OP_25_64_8855/n641 , \DP_OP_25_64_8855/n640 ,
         \DP_OP_25_64_8855/n639 , \DP_OP_25_64_8855/n638 ,
         \DP_OP_25_64_8855/n637 , \DP_OP_25_64_8855/n636 ,
         \DP_OP_25_64_8855/n635 , \DP_OP_25_64_8855/n634 ,
         \DP_OP_25_64_8855/n633 , \DP_OP_25_64_8855/n632 ,
         \DP_OP_25_64_8855/n631 , \DP_OP_25_64_8855/n630 ,
         \DP_OP_25_64_8855/n629 , \DP_OP_25_64_8855/n628 ,
         \DP_OP_25_64_8855/n627 , \DP_OP_25_64_8855/n626 ,
         \DP_OP_25_64_8855/n625 , \DP_OP_25_64_8855/n624 ,
         \DP_OP_25_64_8855/n623 , \DP_OP_25_64_8855/n622 ,
         \DP_OP_25_64_8855/n621 , \DP_OP_25_64_8855/n620 ,
         \DP_OP_25_64_8855/n619 , \DP_OP_25_64_8855/n618 ,
         \DP_OP_25_64_8855/n617 , \DP_OP_25_64_8855/n616 ,
         \DP_OP_25_64_8855/n615 , \DP_OP_25_64_8855/n614 ,
         \DP_OP_25_64_8855/n613 , \DP_OP_25_64_8855/n612 ,
         \DP_OP_25_64_8855/n611 , \DP_OP_25_64_8855/n610 ,
         \DP_OP_25_64_8855/n609 , \DP_OP_25_64_8855/n608 ,
         \DP_OP_25_64_8855/n607 , \DP_OP_25_64_8855/n606 ,
         \DP_OP_25_64_8855/n605 , \DP_OP_25_64_8855/n604 ,
         \DP_OP_25_64_8855/n603 , \DP_OP_25_64_8855/n602 ,
         \DP_OP_25_64_8855/n601 , \DP_OP_25_64_8855/n600 ,
         \DP_OP_25_64_8855/n599 , \DP_OP_25_64_8855/n598 ,
         \DP_OP_25_64_8855/n597 , \DP_OP_25_64_8855/n596 ,
         \DP_OP_25_64_8855/n595 , \DP_OP_25_64_8855/n594 ,
         \DP_OP_25_64_8855/n593 , \DP_OP_25_64_8855/n588 ,
         \DP_OP_25_64_8855/n587 , \DP_OP_25_64_8855/n586 ,
         \DP_OP_25_64_8855/n585 , \DP_OP_25_64_8855/n584 ,
         \DP_OP_25_64_8855/n583 , \DP_OP_25_64_8855/n582 ,
         \DP_OP_25_64_8855/n581 , \DP_OP_25_64_8855/n580 ,
         \DP_OP_25_64_8855/n579 , \DP_OP_25_64_8855/n578 ,
         \DP_OP_25_64_8855/n577 , \DP_OP_25_64_8855/n576 ,
         \DP_OP_25_64_8855/n575 , \DP_OP_25_64_8855/n574 ,
         \DP_OP_25_64_8855/n573 , \DP_OP_25_64_8855/n572 ,
         \DP_OP_25_64_8855/n571 , \DP_OP_25_64_8855/n570 ,
         \DP_OP_25_64_8855/n569 , \DP_OP_25_64_8855/n568 ,
         \DP_OP_25_64_8855/n567 , \DP_OP_25_64_8855/n566 ,
         \DP_OP_25_64_8855/n565 , \DP_OP_25_64_8855/n564 ,
         \DP_OP_25_64_8855/n563 , \DP_OP_25_64_8855/n562 ,
         \DP_OP_25_64_8855/n561 , \DP_OP_25_64_8855/n560 ,
         \DP_OP_25_64_8855/n559 , \DP_OP_25_64_8855/n558 ,
         \DP_OP_25_64_8855/n557 , \DP_OP_25_64_8855/n556 ,
         \DP_OP_25_64_8855/n555 , \DP_OP_25_64_8855/n554 ,
         \DP_OP_25_64_8855/n553 , \DP_OP_25_64_8855/n552 ,
         \DP_OP_25_64_8855/n551 , \DP_OP_25_64_8855/n550 ,
         \DP_OP_25_64_8855/n549 , \DP_OP_25_64_8855/n548 ,
         \DP_OP_25_64_8855/n547 , \DP_OP_25_64_8855/n546 ,
         \DP_OP_25_64_8855/n545 , \DP_OP_25_64_8855/n544 ,
         \DP_OP_25_64_8855/n543 , \DP_OP_25_64_8855/n542 ,
         \DP_OP_25_64_8855/n541 , \DP_OP_25_64_8855/n540 ,
         \DP_OP_25_64_8855/n539 , \DP_OP_25_64_8855/n538 ,
         \DP_OP_25_64_8855/n537 , \DP_OP_25_64_8855/n536 ,
         \DP_OP_25_64_8855/n535 , \DP_OP_25_64_8855/n534 ,
         \DP_OP_25_64_8855/n533 , \DP_OP_25_64_8855/n532 ,
         \DP_OP_25_64_8855/n531 , \DP_OP_25_64_8855/n530 ,
         \DP_OP_25_64_8855/n529 , \DP_OP_25_64_8855/n528 ,
         \DP_OP_25_64_8855/n527 , \DP_OP_25_64_8855/n526 ,
         \DP_OP_25_64_8855/n525 , \DP_OP_25_64_8855/n524 ,
         \DP_OP_25_64_8855/n523 , \DP_OP_25_64_8855/n522 ,
         \DP_OP_25_64_8855/n521 , \DP_OP_25_64_8855/n520 ,
         \DP_OP_25_64_8855/n519 , \DP_OP_25_64_8855/n518 ,
         \DP_OP_25_64_8855/n517 , \DP_OP_25_64_8855/n516 ,
         \DP_OP_25_64_8855/n515 , \DP_OP_25_64_8855/n514 ,
         \DP_OP_25_64_8855/n513 , \DP_OP_25_64_8855/n512 ,
         \DP_OP_25_64_8855/n511 , \DP_OP_25_64_8855/n510 ,
         \DP_OP_25_64_8855/n509 , \DP_OP_25_64_8855/n508 ,
         \DP_OP_25_64_8855/n507 , \DP_OP_25_64_8855/n506 ,
         \DP_OP_25_64_8855/n505 , \DP_OP_25_64_8855/n504 ,
         \DP_OP_25_64_8855/n503 , \DP_OP_25_64_8855/n502 ,
         \DP_OP_25_64_8855/n501 , \DP_OP_25_64_8855/n500 ,
         \DP_OP_25_64_8855/n499 , \DP_OP_25_64_8855/n498 ,
         \DP_OP_25_64_8855/n497 , \DP_OP_25_64_8855/n496 ,
         \DP_OP_25_64_8855/n495 , \DP_OP_25_64_8855/n494 ,
         \DP_OP_25_64_8855/n493 , \DP_OP_25_64_8855/n492 ,
         \DP_OP_25_64_8855/n491 , \DP_OP_25_64_8855/n490 ,
         \DP_OP_25_64_8855/n489 , \DP_OP_25_64_8855/n488 ,
         \DP_OP_25_64_8855/n487 , \DP_OP_25_64_8855/n486 ,
         \DP_OP_25_64_8855/n485 , \DP_OP_25_64_8855/n484 ,
         \DP_OP_25_64_8855/n483 , \DP_OP_25_64_8855/n482 ,
         \DP_OP_25_64_8855/n481 , \DP_OP_25_64_8855/n480 ,
         \DP_OP_25_64_8855/n479 , \DP_OP_25_64_8855/n478 ,
         \DP_OP_25_64_8855/n477 , \DP_OP_25_64_8855/n476 ,
         \DP_OP_25_64_8855/n475 , \DP_OP_25_64_8855/n474 ,
         \DP_OP_25_64_8855/n473 , \DP_OP_25_64_8855/n472 ,
         \DP_OP_25_64_8855/n471 , \DP_OP_25_64_8855/n470 ,
         \DP_OP_25_64_8855/n469 , \DP_OP_25_64_8855/n468 ,
         \DP_OP_25_64_8855/n467 , \DP_OP_25_64_8855/n466 ,
         \DP_OP_25_64_8855/n465 , \DP_OP_25_64_8855/n464 ,
         \DP_OP_25_64_8855/n463 , \DP_OP_25_64_8855/n462 ,
         \DP_OP_25_64_8855/n460 , \DP_OP_25_64_8855/n459 ,
         \DP_OP_25_64_8855/n453 , \DP_OP_25_64_8855/n452 ,
         \DP_OP_25_64_8855/n446 , \DP_OP_25_64_8855/n445 ,
         \DP_OP_25_64_8855/n439 , \DP_OP_25_64_8855/n438 ,
         \DP_OP_25_64_8855/n432 , \DP_OP_25_64_8855/n431 ,
         \DP_OP_25_64_8855/n425 , \DP_OP_25_64_8855/n424 ,
         \DP_OP_25_64_8855/n418 , \DP_OP_25_64_8855/n417 ,
         \DP_OP_25_64_8855/n411 , \DP_OP_25_64_8855/n410 ,
         \DP_OP_25_64_8855/n404 , \DP_OP_25_64_8855/n403 ,
         \DP_OP_25_64_8855/n397 , \DP_OP_25_64_8855/n396 ,
         \DP_OP_25_64_8855/n390 , \DP_OP_25_64_8855/n389 ,
         \DP_OP_25_64_8855/n383 , \DP_OP_25_64_8855/n382 ,
         \DP_OP_25_64_8855/n376 , \DP_OP_25_64_8855/n375 ,
         \DP_OP_25_64_8855/n369 , \DP_OP_25_64_8855/n368 ,
         \DP_OP_25_64_8855/n362 , \DP_OP_25_64_8855/n361 ,
         \DP_OP_25_64_8855/n355 , \DP_OP_25_64_8855/n354 ,
         \DP_OP_25_64_8855/n348 , \DP_OP_25_64_8855/n347 ,
         \DP_OP_25_64_8855/n341 , \DP_OP_25_64_8855/n340 ,
         \DP_OP_25_64_8855/n334 , \DP_OP_25_64_8855/n333 ,
         \DP_OP_25_64_8855/n327 , \DP_OP_25_64_8855/n326 ,
         \DP_OP_25_64_8855/n320 , \DP_OP_25_64_8855/n319 ,
         \DP_OP_25_64_8855/n313 , \DP_OP_25_64_8855/n312 ,
         \DP_OP_25_64_8855/n306 , \DP_OP_25_64_8855/n305 ,
         \DP_OP_25_64_8855/n299 , \DP_OP_25_64_8855/n298 ,
         \DP_OP_25_64_8855/n292 , \DP_OP_25_64_8855/n291 ,
         \DP_OP_25_64_8855/n285 , \DP_OP_25_64_8855/n284 ,
         \DP_OP_25_64_8855/n278 , \DP_OP_25_64_8855/n277 ,
         \DP_OP_25_64_8855/n271 , \DP_OP_25_64_8855/n270 ,
         \DP_OP_25_64_8855/n264 , \DP_OP_25_64_8855/n263 ,
         \DP_OP_25_64_8855/n257 , \DP_OP_25_64_8855/n256 ,
         \DP_OP_25_64_8855/n250 , \DP_OP_25_64_8855/n249 ,
         \DP_OP_25_64_8855/n243 , \DP_OP_25_64_8855/n242 ,
         \DP_OP_25_64_8855/n236 , \DP_OP_25_64_8855/n235 ,
         \DP_OP_25_64_8855/n229 , \DP_OP_25_64_8855/n228 ,
         \DP_OP_25_64_8855/n222 , \DP_OP_25_64_8855/n221 ,
         \DP_OP_25_64_8855/n215 , \DP_OP_25_64_8855/n214 ,
         \DP_OP_25_64_8855/n208 , \DP_OP_25_64_8855/n207 ,
         \DP_OP_25_64_8855/n201 , \DP_OP_25_64_8855/n200 ,
         \DP_OP_25_64_8855/n194 , \DP_OP_25_64_8855/n193 ,
         \DP_OP_25_64_8855/n187 , \DP_OP_25_64_8855/n186 ,
         \DP_OP_25_64_8855/n180 , \DP_OP_25_64_8855/n179 ,
         \DP_OP_25_64_8855/n173 , \DP_OP_25_64_8855/n172 ,
         \DP_OP_25_64_8855/n166 , \DP_OP_25_64_8855/n165 ,
         \DP_OP_25_64_8855/n159 , \DP_OP_25_64_8855/n158 ,
         \DP_OP_25_64_8855/n152 , \DP_OP_25_64_8855/n151 ,
         \DP_OP_25_64_8855/n145 , \DP_OP_25_64_8855/n144 ,
         \DP_OP_25_64_8855/n138 , \DP_OP_25_64_8855/n137 ,
         \DP_OP_25_64_8855/n131 , \DP_OP_25_64_8855/n130 ,
         \DP_OP_25_64_8855/n124 , \DP_OP_25_64_8855/n123 ,
         \DP_OP_25_64_8855/n117 , \DP_OP_25_64_8855/n116 ,
         \DP_OP_25_64_8855/n110 , \DP_OP_25_64_8855/n109 ,
         \DP_OP_25_64_8855/n103 , \DP_OP_25_64_8855/n102 ,
         \DP_OP_25_64_8855/n96 , \DP_OP_25_64_8855/n95 ,
         \DP_OP_25_64_8855/n89 , \DP_OP_25_64_8855/n88 ,
         \DP_OP_25_64_8855/n82 , \DP_OP_25_64_8855/n81 ,
         \DP_OP_25_64_8855/n57 , \DP_OP_25_64_8855/n56 ,
         \DP_OP_25_64_8855/n50 , \DP_OP_25_64_8855/n49 ,
         \DP_OP_25_64_8855/n43 , \DP_OP_25_64_8855/n42 ,
         \DP_OP_25_64_8855/n36 , \DP_OP_25_64_8855/n35 ,
         \DP_OP_25_64_8855/n29 , \DP_OP_25_64_8855/n28 ,
         \DP_OP_25_64_8855/n22 , \DP_OP_25_64_8855/n21 ,
         \DP_OP_25_64_8855/n15 , \DP_OP_25_64_8855/n14 , \DP_OP_25_64_8855/n8 ,
         \DP_OP_25_64_8855/n5 , n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
         n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
         n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
         n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
         n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
         n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
         n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
         n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
         n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
         n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
         n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
         n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
         n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
         n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
         n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
         n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
         n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
         n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
         n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
         n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
         n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
         n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
         n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
         n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
         n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
         n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
         n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
         n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
         n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
         n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
         n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
         n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
         n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
         n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
         n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
         n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
         n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
         n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
         n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
         n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
         n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
         n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
         n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
         n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
         n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
         n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
         n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
         n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
         n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
         n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
         n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
         n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
         n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
         n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
         n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
         n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
         n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
         n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
         n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
         n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
         n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
         n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
         n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
         n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
         n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
         n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
         n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
         n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
         n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
         n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
         n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
         n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
         n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
         n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
         n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
         n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
         n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
         n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
         n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
         n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
         n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
         n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
         n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
         n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
         n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
         n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
         n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
         n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
         n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
         n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
         n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
         n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
         n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
         n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
         n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
         n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
         n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
         n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
         n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
         n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
         n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
         n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
         n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
         n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
         n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
         n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
         n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
         n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
         n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
         n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
         n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
         n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
         n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
         n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
         n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
         n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
         n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
         n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
         n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479,
         n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489,
         n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499,
         n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509,
         n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519,
         n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529,
         n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539,
         n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549,
         n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559,
         n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569,
         n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579,
         n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589,
         n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599,
         n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609,
         n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619,
         n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649,
         n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659,
         n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669,
         n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679,
         n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689,
         n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699,
         n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709,
         n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719,
         n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729,
         n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739,
         n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749,
         n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759,
         n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769,
         n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779,
         n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789,
         n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799,
         n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809,
         n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819,
         n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829,
         n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839,
         n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849,
         n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859,
         n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869,
         n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879,
         n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889,
         n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899,
         n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909,
         n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919,
         n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929,
         n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939,
         n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949,
         n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959,
         n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969,
         n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979,
         n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989,
         n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999,
         n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009,
         n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019,
         n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029,
         n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059,
         n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069,
         n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079,
         n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089,
         n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099,
         n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109,
         n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119,
         n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129,
         n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139,
         n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149,
         n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159,
         n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169,
         n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179,
         n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189,
         n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199,
         n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209,
         n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219,
         n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229,
         n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239,
         n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249,
         n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259,
         n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269,
         n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279,
         n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289,
         n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299,
         n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309,
         n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319,
         n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329,
         n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339,
         n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349,
         n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359,
         n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369,
         n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379,
         n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389,
         n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399,
         n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409,
         n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419,
         n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429,
         n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439,
         n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449,
         n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459,
         n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469,
         n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479,
         n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489,
         n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499,
         n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509,
         n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519,
         n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529,
         n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539,
         n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549,
         n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323;

  DFF \stack_reg[0][0]  ( .D(n2630), .CLK(clk), .RST(rst), .Q(o[0]) );
  DFF \stack_reg[1][0]  ( .D(n2629), .CLK(clk), .RST(rst), .Q(\stack[1][0] )
         );
  DFF \stack_reg[0][1]  ( .D(n2628), .CLK(clk), .RST(rst), .Q(o[1]) );
  DFF \stack_reg[1][1]  ( .D(n2627), .CLK(clk), .RST(rst), .Q(\stack[1][1] )
         );
  DFF \stack_reg[2][1]  ( .D(n2626), .CLK(clk), .RST(rst), .Q(\stack[2][1] )
         );
  DFF \stack_reg[3][1]  ( .D(n2625), .CLK(clk), .RST(rst), .Q(\stack[3][1] )
         );
  DFF \stack_reg[4][1]  ( .D(n2624), .CLK(clk), .RST(rst), .Q(\stack[4][1] )
         );
  DFF \stack_reg[5][1]  ( .D(n2623), .CLK(clk), .RST(rst), .Q(\stack[5][1] )
         );
  DFF \stack_reg[6][1]  ( .D(n2622), .CLK(clk), .RST(rst), .Q(\stack[6][1] )
         );
  DFF \stack_reg[7][1]  ( .D(n2621), .CLK(clk), .RST(rst), .Q(\stack[7][1] )
         );
  DFF \stack_reg[0][2]  ( .D(n2620), .CLK(clk), .RST(rst), .Q(o[2]) );
  DFF \stack_reg[1][2]  ( .D(n2619), .CLK(clk), .RST(rst), .Q(\stack[1][2] )
         );
  DFF \stack_reg[2][2]  ( .D(n2618), .CLK(clk), .RST(rst), .Q(\stack[2][2] )
         );
  DFF \stack_reg[3][2]  ( .D(n2617), .CLK(clk), .RST(rst), .Q(\stack[3][2] )
         );
  DFF \stack_reg[4][2]  ( .D(n2616), .CLK(clk), .RST(rst), .Q(\stack[4][2] )
         );
  DFF \stack_reg[5][2]  ( .D(n2615), .CLK(clk), .RST(rst), .Q(\stack[5][2] )
         );
  DFF \stack_reg[6][2]  ( .D(n2614), .CLK(clk), .RST(rst), .Q(\stack[6][2] )
         );
  DFF \stack_reg[7][2]  ( .D(n2613), .CLK(clk), .RST(rst), .Q(\stack[7][2] )
         );
  DFF \stack_reg[0][3]  ( .D(n2612), .CLK(clk), .RST(rst), .Q(o[3]) );
  DFF \stack_reg[1][3]  ( .D(n2611), .CLK(clk), .RST(rst), .Q(\stack[1][3] )
         );
  DFF \stack_reg[2][3]  ( .D(n2610), .CLK(clk), .RST(rst), .Q(\stack[2][3] )
         );
  DFF \stack_reg[3][3]  ( .D(n2609), .CLK(clk), .RST(rst), .Q(\stack[3][3] )
         );
  DFF \stack_reg[4][3]  ( .D(n2608), .CLK(clk), .RST(rst), .Q(\stack[4][3] )
         );
  DFF \stack_reg[5][3]  ( .D(n2607), .CLK(clk), .RST(rst), .Q(\stack[5][3] )
         );
  DFF \stack_reg[6][3]  ( .D(n2606), .CLK(clk), .RST(rst), .Q(\stack[6][3] )
         );
  DFF \stack_reg[7][3]  ( .D(n2605), .CLK(clk), .RST(rst), .Q(\stack[7][3] )
         );
  DFF \stack_reg[0][4]  ( .D(n2604), .CLK(clk), .RST(rst), .Q(o[4]) );
  DFF \stack_reg[1][4]  ( .D(n2603), .CLK(clk), .RST(rst), .Q(\stack[1][4] )
         );
  DFF \stack_reg[2][4]  ( .D(n2602), .CLK(clk), .RST(rst), .Q(\stack[2][4] )
         );
  DFF \stack_reg[3][4]  ( .D(n2601), .CLK(clk), .RST(rst), .Q(\stack[3][4] )
         );
  DFF \stack_reg[4][4]  ( .D(n2600), .CLK(clk), .RST(rst), .Q(\stack[4][4] )
         );
  DFF \stack_reg[5][4]  ( .D(n2599), .CLK(clk), .RST(rst), .Q(\stack[5][4] )
         );
  DFF \stack_reg[6][4]  ( .D(n2598), .CLK(clk), .RST(rst), .Q(\stack[6][4] )
         );
  DFF \stack_reg[7][4]  ( .D(n2597), .CLK(clk), .RST(rst), .Q(\stack[7][4] )
         );
  DFF \stack_reg[0][5]  ( .D(n2596), .CLK(clk), .RST(rst), .Q(o[5]) );
  DFF \stack_reg[1][5]  ( .D(n2595), .CLK(clk), .RST(rst), .Q(\stack[1][5] )
         );
  DFF \stack_reg[2][5]  ( .D(n2594), .CLK(clk), .RST(rst), .Q(\stack[2][5] )
         );
  DFF \stack_reg[3][5]  ( .D(n2593), .CLK(clk), .RST(rst), .Q(\stack[3][5] )
         );
  DFF \stack_reg[4][5]  ( .D(n2592), .CLK(clk), .RST(rst), .Q(\stack[4][5] )
         );
  DFF \stack_reg[5][5]  ( .D(n2591), .CLK(clk), .RST(rst), .Q(\stack[5][5] )
         );
  DFF \stack_reg[6][5]  ( .D(n2590), .CLK(clk), .RST(rst), .Q(\stack[6][5] )
         );
  DFF \stack_reg[7][5]  ( .D(n2589), .CLK(clk), .RST(rst), .Q(\stack[7][5] )
         );
  DFF \stack_reg[0][6]  ( .D(n2588), .CLK(clk), .RST(rst), .Q(o[6]) );
  DFF \stack_reg[1][6]  ( .D(n2587), .CLK(clk), .RST(rst), .Q(\stack[1][6] )
         );
  DFF \stack_reg[2][6]  ( .D(n2586), .CLK(clk), .RST(rst), .Q(\stack[2][6] )
         );
  DFF \stack_reg[3][6]  ( .D(n2585), .CLK(clk), .RST(rst), .Q(\stack[3][6] )
         );
  DFF \stack_reg[4][6]  ( .D(n2584), .CLK(clk), .RST(rst), .Q(\stack[4][6] )
         );
  DFF \stack_reg[5][6]  ( .D(n2583), .CLK(clk), .RST(rst), .Q(\stack[5][6] )
         );
  DFF \stack_reg[6][6]  ( .D(n2582), .CLK(clk), .RST(rst), .Q(\stack[6][6] )
         );
  DFF \stack_reg[7][6]  ( .D(n2581), .CLK(clk), .RST(rst), .Q(\stack[7][6] )
         );
  DFF \stack_reg[0][7]  ( .D(n2580), .CLK(clk), .RST(rst), .Q(o[7]) );
  DFF \stack_reg[1][7]  ( .D(n2579), .CLK(clk), .RST(rst), .Q(\stack[1][7] )
         );
  DFF \stack_reg[2][7]  ( .D(n2578), .CLK(clk), .RST(rst), .Q(\stack[2][7] )
         );
  DFF \stack_reg[3][7]  ( .D(n2577), .CLK(clk), .RST(rst), .Q(\stack[3][7] )
         );
  DFF \stack_reg[4][7]  ( .D(n2576), .CLK(clk), .RST(rst), .Q(\stack[4][7] )
         );
  DFF \stack_reg[5][7]  ( .D(n2575), .CLK(clk), .RST(rst), .Q(\stack[5][7] )
         );
  DFF \stack_reg[6][7]  ( .D(n2574), .CLK(clk), .RST(rst), .Q(\stack[6][7] )
         );
  DFF \stack_reg[7][7]  ( .D(n2573), .CLK(clk), .RST(rst), .Q(\stack[7][7] )
         );
  DFF \stack_reg[0][8]  ( .D(n2572), .CLK(clk), .RST(rst), .Q(o[8]) );
  DFF \stack_reg[1][8]  ( .D(n2571), .CLK(clk), .RST(rst), .Q(\stack[1][8] )
         );
  DFF \stack_reg[2][8]  ( .D(n2570), .CLK(clk), .RST(rst), .Q(\stack[2][8] )
         );
  DFF \stack_reg[3][8]  ( .D(n2569), .CLK(clk), .RST(rst), .Q(\stack[3][8] )
         );
  DFF \stack_reg[4][8]  ( .D(n2568), .CLK(clk), .RST(rst), .Q(\stack[4][8] )
         );
  DFF \stack_reg[5][8]  ( .D(n2567), .CLK(clk), .RST(rst), .Q(\stack[5][8] )
         );
  DFF \stack_reg[6][8]  ( .D(n2566), .CLK(clk), .RST(rst), .Q(\stack[6][8] )
         );
  DFF \stack_reg[7][8]  ( .D(n2565), .CLK(clk), .RST(rst), .Q(\stack[7][8] )
         );
  DFF \stack_reg[0][9]  ( .D(n2564), .CLK(clk), .RST(rst), .Q(o[9]) );
  DFF \stack_reg[1][9]  ( .D(n2563), .CLK(clk), .RST(rst), .Q(\stack[1][9] )
         );
  DFF \stack_reg[2][9]  ( .D(n2562), .CLK(clk), .RST(rst), .Q(\stack[2][9] )
         );
  DFF \stack_reg[3][9]  ( .D(n2561), .CLK(clk), .RST(rst), .Q(\stack[3][9] )
         );
  DFF \stack_reg[4][9]  ( .D(n2560), .CLK(clk), .RST(rst), .Q(\stack[4][9] )
         );
  DFF \stack_reg[5][9]  ( .D(n2559), .CLK(clk), .RST(rst), .Q(\stack[5][9] )
         );
  DFF \stack_reg[6][9]  ( .D(n2558), .CLK(clk), .RST(rst), .Q(\stack[6][9] )
         );
  DFF \stack_reg[7][9]  ( .D(n2557), .CLK(clk), .RST(rst), .Q(\stack[7][9] )
         );
  DFF \stack_reg[0][10]  ( .D(n2556), .CLK(clk), .RST(rst), .Q(o[10]) );
  DFF \stack_reg[1][10]  ( .D(n2555), .CLK(clk), .RST(rst), .Q(\stack[1][10] )
         );
  DFF \stack_reg[2][10]  ( .D(n2554), .CLK(clk), .RST(rst), .Q(\stack[2][10] )
         );
  DFF \stack_reg[3][10]  ( .D(n2553), .CLK(clk), .RST(rst), .Q(\stack[3][10] )
         );
  DFF \stack_reg[4][10]  ( .D(n2552), .CLK(clk), .RST(rst), .Q(\stack[4][10] )
         );
  DFF \stack_reg[5][10]  ( .D(n2551), .CLK(clk), .RST(rst), .Q(\stack[5][10] )
         );
  DFF \stack_reg[6][10]  ( .D(n2550), .CLK(clk), .RST(rst), .Q(\stack[6][10] )
         );
  DFF \stack_reg[7][10]  ( .D(n2549), .CLK(clk), .RST(rst), .Q(\stack[7][10] )
         );
  DFF \stack_reg[0][11]  ( .D(n2548), .CLK(clk), .RST(rst), .Q(o[11]) );
  DFF \stack_reg[1][11]  ( .D(n2547), .CLK(clk), .RST(rst), .Q(\stack[1][11] )
         );
  DFF \stack_reg[2][11]  ( .D(n2546), .CLK(clk), .RST(rst), .Q(\stack[2][11] )
         );
  DFF \stack_reg[3][11]  ( .D(n2545), .CLK(clk), .RST(rst), .Q(\stack[3][11] )
         );
  DFF \stack_reg[4][11]  ( .D(n2544), .CLK(clk), .RST(rst), .Q(\stack[4][11] )
         );
  DFF \stack_reg[5][11]  ( .D(n2543), .CLK(clk), .RST(rst), .Q(\stack[5][11] )
         );
  DFF \stack_reg[6][11]  ( .D(n2542), .CLK(clk), .RST(rst), .Q(\stack[6][11] )
         );
  DFF \stack_reg[7][11]  ( .D(n2541), .CLK(clk), .RST(rst), .Q(\stack[7][11] )
         );
  DFF \stack_reg[0][12]  ( .D(n2540), .CLK(clk), .RST(rst), .Q(o[12]) );
  DFF \stack_reg[1][12]  ( .D(n2539), .CLK(clk), .RST(rst), .Q(\stack[1][12] )
         );
  DFF \stack_reg[2][12]  ( .D(n2538), .CLK(clk), .RST(rst), .Q(\stack[2][12] )
         );
  DFF \stack_reg[3][12]  ( .D(n2537), .CLK(clk), .RST(rst), .Q(\stack[3][12] )
         );
  DFF \stack_reg[4][12]  ( .D(n2536), .CLK(clk), .RST(rst), .Q(\stack[4][12] )
         );
  DFF \stack_reg[5][12]  ( .D(n2535), .CLK(clk), .RST(rst), .Q(\stack[5][12] )
         );
  DFF \stack_reg[6][12]  ( .D(n2534), .CLK(clk), .RST(rst), .Q(\stack[6][12] )
         );
  DFF \stack_reg[7][12]  ( .D(n2533), .CLK(clk), .RST(rst), .Q(\stack[7][12] )
         );
  DFF \stack_reg[0][13]  ( .D(n2532), .CLK(clk), .RST(rst), .Q(o[13]) );
  DFF \stack_reg[1][13]  ( .D(n2531), .CLK(clk), .RST(rst), .Q(\stack[1][13] )
         );
  DFF \stack_reg[2][13]  ( .D(n2530), .CLK(clk), .RST(rst), .Q(\stack[2][13] )
         );
  DFF \stack_reg[3][13]  ( .D(n2529), .CLK(clk), .RST(rst), .Q(\stack[3][13] )
         );
  DFF \stack_reg[4][13]  ( .D(n2528), .CLK(clk), .RST(rst), .Q(\stack[4][13] )
         );
  DFF \stack_reg[5][13]  ( .D(n2527), .CLK(clk), .RST(rst), .Q(\stack[5][13] )
         );
  DFF \stack_reg[6][13]  ( .D(n2526), .CLK(clk), .RST(rst), .Q(\stack[6][13] )
         );
  DFF \stack_reg[7][13]  ( .D(n2525), .CLK(clk), .RST(rst), .Q(\stack[7][13] )
         );
  DFF \stack_reg[0][14]  ( .D(n2524), .CLK(clk), .RST(rst), .Q(o[14]) );
  DFF \stack_reg[1][14]  ( .D(n2523), .CLK(clk), .RST(rst), .Q(\stack[1][14] )
         );
  DFF \stack_reg[2][14]  ( .D(n2522), .CLK(clk), .RST(rst), .Q(\stack[2][14] )
         );
  DFF \stack_reg[3][14]  ( .D(n2521), .CLK(clk), .RST(rst), .Q(\stack[3][14] )
         );
  DFF \stack_reg[4][14]  ( .D(n2520), .CLK(clk), .RST(rst), .Q(\stack[4][14] )
         );
  DFF \stack_reg[5][14]  ( .D(n2519), .CLK(clk), .RST(rst), .Q(\stack[5][14] )
         );
  DFF \stack_reg[6][14]  ( .D(n2518), .CLK(clk), .RST(rst), .Q(\stack[6][14] )
         );
  DFF \stack_reg[7][14]  ( .D(n2517), .CLK(clk), .RST(rst), .Q(\stack[7][14] )
         );
  DFF \stack_reg[0][15]  ( .D(n2516), .CLK(clk), .RST(rst), .Q(o[15]) );
  DFF \stack_reg[1][15]  ( .D(n2515), .CLK(clk), .RST(rst), .Q(\stack[1][15] )
         );
  DFF \stack_reg[2][15]  ( .D(n2514), .CLK(clk), .RST(rst), .Q(\stack[2][15] )
         );
  DFF \stack_reg[3][15]  ( .D(n2513), .CLK(clk), .RST(rst), .Q(\stack[3][15] )
         );
  DFF \stack_reg[4][15]  ( .D(n2512), .CLK(clk), .RST(rst), .Q(\stack[4][15] )
         );
  DFF \stack_reg[5][15]  ( .D(n2511), .CLK(clk), .RST(rst), .Q(\stack[5][15] )
         );
  DFF \stack_reg[6][15]  ( .D(n2510), .CLK(clk), .RST(rst), .Q(\stack[6][15] )
         );
  DFF \stack_reg[7][15]  ( .D(n2509), .CLK(clk), .RST(rst), .Q(\stack[7][15] )
         );
  DFF \stack_reg[0][16]  ( .D(n2508), .CLK(clk), .RST(rst), .Q(o[16]) );
  DFF \stack_reg[1][16]  ( .D(n2507), .CLK(clk), .RST(rst), .Q(\stack[1][16] )
         );
  DFF \stack_reg[2][16]  ( .D(n2506), .CLK(clk), .RST(rst), .Q(\stack[2][16] )
         );
  DFF \stack_reg[3][16]  ( .D(n2505), .CLK(clk), .RST(rst), .Q(\stack[3][16] )
         );
  DFF \stack_reg[4][16]  ( .D(n2504), .CLK(clk), .RST(rst), .Q(\stack[4][16] )
         );
  DFF \stack_reg[5][16]  ( .D(n2503), .CLK(clk), .RST(rst), .Q(\stack[5][16] )
         );
  DFF \stack_reg[6][16]  ( .D(n2502), .CLK(clk), .RST(rst), .Q(\stack[6][16] )
         );
  DFF \stack_reg[7][16]  ( .D(n2501), .CLK(clk), .RST(rst), .Q(\stack[7][16] )
         );
  DFF \stack_reg[0][17]  ( .D(n2500), .CLK(clk), .RST(rst), .Q(o[17]) );
  DFF \stack_reg[1][17]  ( .D(n2499), .CLK(clk), .RST(rst), .Q(\stack[1][17] )
         );
  DFF \stack_reg[2][17]  ( .D(n2498), .CLK(clk), .RST(rst), .Q(\stack[2][17] )
         );
  DFF \stack_reg[3][17]  ( .D(n2497), .CLK(clk), .RST(rst), .Q(\stack[3][17] )
         );
  DFF \stack_reg[4][17]  ( .D(n2496), .CLK(clk), .RST(rst), .Q(\stack[4][17] )
         );
  DFF \stack_reg[5][17]  ( .D(n2495), .CLK(clk), .RST(rst), .Q(\stack[5][17] )
         );
  DFF \stack_reg[6][17]  ( .D(n2494), .CLK(clk), .RST(rst), .Q(\stack[6][17] )
         );
  DFF \stack_reg[7][17]  ( .D(n2493), .CLK(clk), .RST(rst), .Q(\stack[7][17] )
         );
  DFF \stack_reg[0][18]  ( .D(n2492), .CLK(clk), .RST(rst), .Q(o[18]) );
  DFF \stack_reg[1][18]  ( .D(n2491), .CLK(clk), .RST(rst), .Q(\stack[1][18] )
         );
  DFF \stack_reg[2][18]  ( .D(n2490), .CLK(clk), .RST(rst), .Q(\stack[2][18] )
         );
  DFF \stack_reg[3][18]  ( .D(n2489), .CLK(clk), .RST(rst), .Q(\stack[3][18] )
         );
  DFF \stack_reg[4][18]  ( .D(n2488), .CLK(clk), .RST(rst), .Q(\stack[4][18] )
         );
  DFF \stack_reg[5][18]  ( .D(n2487), .CLK(clk), .RST(rst), .Q(\stack[5][18] )
         );
  DFF \stack_reg[6][18]  ( .D(n2486), .CLK(clk), .RST(rst), .Q(\stack[6][18] )
         );
  DFF \stack_reg[7][18]  ( .D(n2485), .CLK(clk), .RST(rst), .Q(\stack[7][18] )
         );
  DFF \stack_reg[0][19]  ( .D(n2484), .CLK(clk), .RST(rst), .Q(o[19]) );
  DFF \stack_reg[1][19]  ( .D(n2483), .CLK(clk), .RST(rst), .Q(\stack[1][19] )
         );
  DFF \stack_reg[2][19]  ( .D(n2482), .CLK(clk), .RST(rst), .Q(\stack[2][19] )
         );
  DFF \stack_reg[3][19]  ( .D(n2481), .CLK(clk), .RST(rst), .Q(\stack[3][19] )
         );
  DFF \stack_reg[4][19]  ( .D(n2480), .CLK(clk), .RST(rst), .Q(\stack[4][19] )
         );
  DFF \stack_reg[5][19]  ( .D(n2479), .CLK(clk), .RST(rst), .Q(\stack[5][19] )
         );
  DFF \stack_reg[6][19]  ( .D(n2478), .CLK(clk), .RST(rst), .Q(\stack[6][19] )
         );
  DFF \stack_reg[7][19]  ( .D(n2477), .CLK(clk), .RST(rst), .Q(\stack[7][19] )
         );
  DFF \stack_reg[0][20]  ( .D(n2476), .CLK(clk), .RST(rst), .Q(o[20]) );
  DFF \stack_reg[1][20]  ( .D(n2475), .CLK(clk), .RST(rst), .Q(\stack[1][20] )
         );
  DFF \stack_reg[2][20]  ( .D(n2474), .CLK(clk), .RST(rst), .Q(\stack[2][20] )
         );
  DFF \stack_reg[3][20]  ( .D(n2473), .CLK(clk), .RST(rst), .Q(\stack[3][20] )
         );
  DFF \stack_reg[4][20]  ( .D(n2472), .CLK(clk), .RST(rst), .Q(\stack[4][20] )
         );
  DFF \stack_reg[5][20]  ( .D(n2471), .CLK(clk), .RST(rst), .Q(\stack[5][20] )
         );
  DFF \stack_reg[6][20]  ( .D(n2470), .CLK(clk), .RST(rst), .Q(\stack[6][20] )
         );
  DFF \stack_reg[7][20]  ( .D(n2469), .CLK(clk), .RST(rst), .Q(\stack[7][20] )
         );
  DFF \stack_reg[0][21]  ( .D(n2468), .CLK(clk), .RST(rst), .Q(o[21]) );
  DFF \stack_reg[1][21]  ( .D(n2467), .CLK(clk), .RST(rst), .Q(\stack[1][21] )
         );
  DFF \stack_reg[2][21]  ( .D(n2466), .CLK(clk), .RST(rst), .Q(\stack[2][21] )
         );
  DFF \stack_reg[3][21]  ( .D(n2465), .CLK(clk), .RST(rst), .Q(\stack[3][21] )
         );
  DFF \stack_reg[4][21]  ( .D(n2464), .CLK(clk), .RST(rst), .Q(\stack[4][21] )
         );
  DFF \stack_reg[5][21]  ( .D(n2463), .CLK(clk), .RST(rst), .Q(\stack[5][21] )
         );
  DFF \stack_reg[6][21]  ( .D(n2462), .CLK(clk), .RST(rst), .Q(\stack[6][21] )
         );
  DFF \stack_reg[7][21]  ( .D(n2461), .CLK(clk), .RST(rst), .Q(\stack[7][21] )
         );
  DFF \stack_reg[0][22]  ( .D(n2460), .CLK(clk), .RST(rst), .Q(o[22]) );
  DFF \stack_reg[1][22]  ( .D(n2459), .CLK(clk), .RST(rst), .Q(\stack[1][22] )
         );
  DFF \stack_reg[2][22]  ( .D(n2458), .CLK(clk), .RST(rst), .Q(\stack[2][22] )
         );
  DFF \stack_reg[3][22]  ( .D(n2457), .CLK(clk), .RST(rst), .Q(\stack[3][22] )
         );
  DFF \stack_reg[4][22]  ( .D(n2456), .CLK(clk), .RST(rst), .Q(\stack[4][22] )
         );
  DFF \stack_reg[5][22]  ( .D(n2455), .CLK(clk), .RST(rst), .Q(\stack[5][22] )
         );
  DFF \stack_reg[6][22]  ( .D(n2454), .CLK(clk), .RST(rst), .Q(\stack[6][22] )
         );
  DFF \stack_reg[7][22]  ( .D(n2453), .CLK(clk), .RST(rst), .Q(\stack[7][22] )
         );
  DFF \stack_reg[0][23]  ( .D(n2452), .CLK(clk), .RST(rst), .Q(o[23]) );
  DFF \stack_reg[1][23]  ( .D(n2451), .CLK(clk), .RST(rst), .Q(\stack[1][23] )
         );
  DFF \stack_reg[2][23]  ( .D(n2450), .CLK(clk), .RST(rst), .Q(\stack[2][23] )
         );
  DFF \stack_reg[3][23]  ( .D(n2449), .CLK(clk), .RST(rst), .Q(\stack[3][23] )
         );
  DFF \stack_reg[4][23]  ( .D(n2448), .CLK(clk), .RST(rst), .Q(\stack[4][23] )
         );
  DFF \stack_reg[5][23]  ( .D(n2447), .CLK(clk), .RST(rst), .Q(\stack[5][23] )
         );
  DFF \stack_reg[6][23]  ( .D(n2446), .CLK(clk), .RST(rst), .Q(\stack[6][23] )
         );
  DFF \stack_reg[7][23]  ( .D(n2445), .CLK(clk), .RST(rst), .Q(\stack[7][23] )
         );
  DFF \stack_reg[0][24]  ( .D(n2444), .CLK(clk), .RST(rst), .Q(o[24]) );
  DFF \stack_reg[1][24]  ( .D(n2443), .CLK(clk), .RST(rst), .Q(\stack[1][24] )
         );
  DFF \stack_reg[2][24]  ( .D(n2442), .CLK(clk), .RST(rst), .Q(\stack[2][24] )
         );
  DFF \stack_reg[3][24]  ( .D(n2441), .CLK(clk), .RST(rst), .Q(\stack[3][24] )
         );
  DFF \stack_reg[4][24]  ( .D(n2440), .CLK(clk), .RST(rst), .Q(\stack[4][24] )
         );
  DFF \stack_reg[5][24]  ( .D(n2439), .CLK(clk), .RST(rst), .Q(\stack[5][24] )
         );
  DFF \stack_reg[6][24]  ( .D(n2438), .CLK(clk), .RST(rst), .Q(\stack[6][24] )
         );
  DFF \stack_reg[7][24]  ( .D(n2437), .CLK(clk), .RST(rst), .Q(\stack[7][24] )
         );
  DFF \stack_reg[0][25]  ( .D(n2436), .CLK(clk), .RST(rst), .Q(o[25]) );
  DFF \stack_reg[1][25]  ( .D(n2435), .CLK(clk), .RST(rst), .Q(\stack[1][25] )
         );
  DFF \stack_reg[2][25]  ( .D(n2434), .CLK(clk), .RST(rst), .Q(\stack[2][25] )
         );
  DFF \stack_reg[3][25]  ( .D(n2433), .CLK(clk), .RST(rst), .Q(\stack[3][25] )
         );
  DFF \stack_reg[4][25]  ( .D(n2432), .CLK(clk), .RST(rst), .Q(\stack[4][25] )
         );
  DFF \stack_reg[5][25]  ( .D(n2431), .CLK(clk), .RST(rst), .Q(\stack[5][25] )
         );
  DFF \stack_reg[6][25]  ( .D(n2430), .CLK(clk), .RST(rst), .Q(\stack[6][25] )
         );
  DFF \stack_reg[7][25]  ( .D(n2429), .CLK(clk), .RST(rst), .Q(\stack[7][25] )
         );
  DFF \stack_reg[0][26]  ( .D(n2428), .CLK(clk), .RST(rst), .Q(o[26]) );
  DFF \stack_reg[1][26]  ( .D(n2427), .CLK(clk), .RST(rst), .Q(\stack[1][26] )
         );
  DFF \stack_reg[2][26]  ( .D(n2426), .CLK(clk), .RST(rst), .Q(\stack[2][26] )
         );
  DFF \stack_reg[3][26]  ( .D(n2425), .CLK(clk), .RST(rst), .Q(\stack[3][26] )
         );
  DFF \stack_reg[4][26]  ( .D(n2424), .CLK(clk), .RST(rst), .Q(\stack[4][26] )
         );
  DFF \stack_reg[5][26]  ( .D(n2423), .CLK(clk), .RST(rst), .Q(\stack[5][26] )
         );
  DFF \stack_reg[6][26]  ( .D(n2422), .CLK(clk), .RST(rst), .Q(\stack[6][26] )
         );
  DFF \stack_reg[7][26]  ( .D(n2421), .CLK(clk), .RST(rst), .Q(\stack[7][26] )
         );
  DFF \stack_reg[0][27]  ( .D(n2420), .CLK(clk), .RST(rst), .Q(o[27]) );
  DFF \stack_reg[1][27]  ( .D(n2419), .CLK(clk), .RST(rst), .Q(\stack[1][27] )
         );
  DFF \stack_reg[2][27]  ( .D(n2418), .CLK(clk), .RST(rst), .Q(\stack[2][27] )
         );
  DFF \stack_reg[3][27]  ( .D(n2417), .CLK(clk), .RST(rst), .Q(\stack[3][27] )
         );
  DFF \stack_reg[4][27]  ( .D(n2416), .CLK(clk), .RST(rst), .Q(\stack[4][27] )
         );
  DFF \stack_reg[5][27]  ( .D(n2415), .CLK(clk), .RST(rst), .Q(\stack[5][27] )
         );
  DFF \stack_reg[6][27]  ( .D(n2414), .CLK(clk), .RST(rst), .Q(\stack[6][27] )
         );
  DFF \stack_reg[7][27]  ( .D(n2413), .CLK(clk), .RST(rst), .Q(\stack[7][27] )
         );
  DFF \stack_reg[0][28]  ( .D(n2412), .CLK(clk), .RST(rst), .Q(o[28]) );
  DFF \stack_reg[1][28]  ( .D(n2411), .CLK(clk), .RST(rst), .Q(\stack[1][28] )
         );
  DFF \stack_reg[2][28]  ( .D(n2410), .CLK(clk), .RST(rst), .Q(\stack[2][28] )
         );
  DFF \stack_reg[3][28]  ( .D(n2409), .CLK(clk), .RST(rst), .Q(\stack[3][28] )
         );
  DFF \stack_reg[4][28]  ( .D(n2408), .CLK(clk), .RST(rst), .Q(\stack[4][28] )
         );
  DFF \stack_reg[5][28]  ( .D(n2407), .CLK(clk), .RST(rst), .Q(\stack[5][28] )
         );
  DFF \stack_reg[6][28]  ( .D(n2406), .CLK(clk), .RST(rst), .Q(\stack[6][28] )
         );
  DFF \stack_reg[7][28]  ( .D(n2405), .CLK(clk), .RST(rst), .Q(\stack[7][28] )
         );
  DFF \stack_reg[0][29]  ( .D(n2404), .CLK(clk), .RST(rst), .Q(o[29]) );
  DFF \stack_reg[1][29]  ( .D(n2403), .CLK(clk), .RST(rst), .Q(\stack[1][29] )
         );
  DFF \stack_reg[2][29]  ( .D(n2402), .CLK(clk), .RST(rst), .Q(\stack[2][29] )
         );
  DFF \stack_reg[3][29]  ( .D(n2401), .CLK(clk), .RST(rst), .Q(\stack[3][29] )
         );
  DFF \stack_reg[4][29]  ( .D(n2400), .CLK(clk), .RST(rst), .Q(\stack[4][29] )
         );
  DFF \stack_reg[5][29]  ( .D(n2399), .CLK(clk), .RST(rst), .Q(\stack[5][29] )
         );
  DFF \stack_reg[6][29]  ( .D(n2398), .CLK(clk), .RST(rst), .Q(\stack[6][29] )
         );
  DFF \stack_reg[7][29]  ( .D(n2397), .CLK(clk), .RST(rst), .Q(\stack[7][29] )
         );
  DFF \stack_reg[0][30]  ( .D(n2396), .CLK(clk), .RST(rst), .Q(o[30]) );
  DFF \stack_reg[1][30]  ( .D(n2395), .CLK(clk), .RST(rst), .Q(\stack[1][30] )
         );
  DFF \stack_reg[2][30]  ( .D(n2394), .CLK(clk), .RST(rst), .Q(\stack[2][30] )
         );
  DFF \stack_reg[3][30]  ( .D(n2393), .CLK(clk), .RST(rst), .Q(\stack[3][30] )
         );
  DFF \stack_reg[4][30]  ( .D(n2392), .CLK(clk), .RST(rst), .Q(\stack[4][30] )
         );
  DFF \stack_reg[5][30]  ( .D(n2391), .CLK(clk), .RST(rst), .Q(\stack[5][30] )
         );
  DFF \stack_reg[6][30]  ( .D(n2390), .CLK(clk), .RST(rst), .Q(\stack[6][30] )
         );
  DFF \stack_reg[7][30]  ( .D(n2389), .CLK(clk), .RST(rst), .Q(\stack[7][30] )
         );
  DFF \stack_reg[0][31]  ( .D(n2388), .CLK(clk), .RST(rst), .Q(o[31]) );
  DFF \stack_reg[1][31]  ( .D(n2387), .CLK(clk), .RST(rst), .Q(\stack[1][31] )
         );
  DFF \stack_reg[2][31]  ( .D(n2386), .CLK(clk), .RST(rst), .Q(\stack[2][31] )
         );
  DFF \stack_reg[3][31]  ( .D(n2385), .CLK(clk), .RST(rst), .Q(\stack[3][31] )
         );
  DFF \stack_reg[4][31]  ( .D(n2384), .CLK(clk), .RST(rst), .Q(\stack[4][31] )
         );
  DFF \stack_reg[5][31]  ( .D(n2383), .CLK(clk), .RST(rst), .Q(\stack[5][31] )
         );
  DFF \stack_reg[6][31]  ( .D(n2382), .CLK(clk), .RST(rst), .Q(\stack[6][31] )
         );
  DFF \stack_reg[7][31]  ( .D(n2381), .CLK(clk), .RST(rst), .Q(\stack[7][31] )
         );
  DFF \stack_reg[0][32]  ( .D(n2380), .CLK(clk), .RST(rst), .Q(o[32]) );
  DFF \stack_reg[1][32]  ( .D(n2379), .CLK(clk), .RST(rst), .Q(\stack[1][32] )
         );
  DFF \stack_reg[2][32]  ( .D(n2378), .CLK(clk), .RST(rst), .Q(\stack[2][32] )
         );
  DFF \stack_reg[3][32]  ( .D(n2377), .CLK(clk), .RST(rst), .Q(\stack[3][32] )
         );
  DFF \stack_reg[4][32]  ( .D(n2376), .CLK(clk), .RST(rst), .Q(\stack[4][32] )
         );
  DFF \stack_reg[5][32]  ( .D(n2375), .CLK(clk), .RST(rst), .Q(\stack[5][32] )
         );
  DFF \stack_reg[6][32]  ( .D(n2374), .CLK(clk), .RST(rst), .Q(\stack[6][32] )
         );
  DFF \stack_reg[7][32]  ( .D(n2373), .CLK(clk), .RST(rst), .Q(\stack[7][32] )
         );
  DFF \stack_reg[0][33]  ( .D(n2372), .CLK(clk), .RST(rst), .Q(o[33]) );
  DFF \stack_reg[1][33]  ( .D(n2371), .CLK(clk), .RST(rst), .Q(\stack[1][33] )
         );
  DFF \stack_reg[2][33]  ( .D(n2370), .CLK(clk), .RST(rst), .Q(\stack[2][33] )
         );
  DFF \stack_reg[3][33]  ( .D(n2369), .CLK(clk), .RST(rst), .Q(\stack[3][33] )
         );
  DFF \stack_reg[4][33]  ( .D(n2368), .CLK(clk), .RST(rst), .Q(\stack[4][33] )
         );
  DFF \stack_reg[5][33]  ( .D(n2367), .CLK(clk), .RST(rst), .Q(\stack[5][33] )
         );
  DFF \stack_reg[6][33]  ( .D(n2366), .CLK(clk), .RST(rst), .Q(\stack[6][33] )
         );
  DFF \stack_reg[7][33]  ( .D(n2365), .CLK(clk), .RST(rst), .Q(\stack[7][33] )
         );
  DFF \stack_reg[0][34]  ( .D(n2364), .CLK(clk), .RST(rst), .Q(o[34]) );
  DFF \stack_reg[1][34]  ( .D(n2363), .CLK(clk), .RST(rst), .Q(\stack[1][34] )
         );
  DFF \stack_reg[2][34]  ( .D(n2362), .CLK(clk), .RST(rst), .Q(\stack[2][34] )
         );
  DFF \stack_reg[3][34]  ( .D(n2361), .CLK(clk), .RST(rst), .Q(\stack[3][34] )
         );
  DFF \stack_reg[4][34]  ( .D(n2360), .CLK(clk), .RST(rst), .Q(\stack[4][34] )
         );
  DFF \stack_reg[5][34]  ( .D(n2359), .CLK(clk), .RST(rst), .Q(\stack[5][34] )
         );
  DFF \stack_reg[6][34]  ( .D(n2358), .CLK(clk), .RST(rst), .Q(\stack[6][34] )
         );
  DFF \stack_reg[7][34]  ( .D(n2357), .CLK(clk), .RST(rst), .Q(\stack[7][34] )
         );
  DFF \stack_reg[0][35]  ( .D(n2356), .CLK(clk), .RST(rst), .Q(o[35]) );
  DFF \stack_reg[1][35]  ( .D(n2355), .CLK(clk), .RST(rst), .Q(\stack[1][35] )
         );
  DFF \stack_reg[2][35]  ( .D(n2354), .CLK(clk), .RST(rst), .Q(\stack[2][35] )
         );
  DFF \stack_reg[3][35]  ( .D(n2353), .CLK(clk), .RST(rst), .Q(\stack[3][35] )
         );
  DFF \stack_reg[4][35]  ( .D(n2352), .CLK(clk), .RST(rst), .Q(\stack[4][35] )
         );
  DFF \stack_reg[5][35]  ( .D(n2351), .CLK(clk), .RST(rst), .Q(\stack[5][35] )
         );
  DFF \stack_reg[6][35]  ( .D(n2350), .CLK(clk), .RST(rst), .Q(\stack[6][35] )
         );
  DFF \stack_reg[7][35]  ( .D(n2349), .CLK(clk), .RST(rst), .Q(\stack[7][35] )
         );
  DFF \stack_reg[0][36]  ( .D(n2348), .CLK(clk), .RST(rst), .Q(o[36]) );
  DFF \stack_reg[1][36]  ( .D(n2347), .CLK(clk), .RST(rst), .Q(\stack[1][36] )
         );
  DFF \stack_reg[2][36]  ( .D(n2346), .CLK(clk), .RST(rst), .Q(\stack[2][36] )
         );
  DFF \stack_reg[3][36]  ( .D(n2345), .CLK(clk), .RST(rst), .Q(\stack[3][36] )
         );
  DFF \stack_reg[4][36]  ( .D(n2344), .CLK(clk), .RST(rst), .Q(\stack[4][36] )
         );
  DFF \stack_reg[5][36]  ( .D(n2343), .CLK(clk), .RST(rst), .Q(\stack[5][36] )
         );
  DFF \stack_reg[6][36]  ( .D(n2342), .CLK(clk), .RST(rst), .Q(\stack[6][36] )
         );
  DFF \stack_reg[7][36]  ( .D(n2341), .CLK(clk), .RST(rst), .Q(\stack[7][36] )
         );
  DFF \stack_reg[0][37]  ( .D(n2340), .CLK(clk), .RST(rst), .Q(o[37]) );
  DFF \stack_reg[1][37]  ( .D(n2339), .CLK(clk), .RST(rst), .Q(\stack[1][37] )
         );
  DFF \stack_reg[2][37]  ( .D(n2338), .CLK(clk), .RST(rst), .Q(\stack[2][37] )
         );
  DFF \stack_reg[3][37]  ( .D(n2337), .CLK(clk), .RST(rst), .Q(\stack[3][37] )
         );
  DFF \stack_reg[4][37]  ( .D(n2336), .CLK(clk), .RST(rst), .Q(\stack[4][37] )
         );
  DFF \stack_reg[5][37]  ( .D(n2335), .CLK(clk), .RST(rst), .Q(\stack[5][37] )
         );
  DFF \stack_reg[6][37]  ( .D(n2334), .CLK(clk), .RST(rst), .Q(\stack[6][37] )
         );
  DFF \stack_reg[7][37]  ( .D(n2333), .CLK(clk), .RST(rst), .Q(\stack[7][37] )
         );
  DFF \stack_reg[0][38]  ( .D(n2332), .CLK(clk), .RST(rst), .Q(o[38]) );
  DFF \stack_reg[1][38]  ( .D(n2331), .CLK(clk), .RST(rst), .Q(\stack[1][38] )
         );
  DFF \stack_reg[2][38]  ( .D(n2330), .CLK(clk), .RST(rst), .Q(\stack[2][38] )
         );
  DFF \stack_reg[3][38]  ( .D(n2329), .CLK(clk), .RST(rst), .Q(\stack[3][38] )
         );
  DFF \stack_reg[4][38]  ( .D(n2328), .CLK(clk), .RST(rst), .Q(\stack[4][38] )
         );
  DFF \stack_reg[5][38]  ( .D(n2327), .CLK(clk), .RST(rst), .Q(\stack[5][38] )
         );
  DFF \stack_reg[6][38]  ( .D(n2326), .CLK(clk), .RST(rst), .Q(\stack[6][38] )
         );
  DFF \stack_reg[7][38]  ( .D(n2325), .CLK(clk), .RST(rst), .Q(\stack[7][38] )
         );
  DFF \stack_reg[0][39]  ( .D(n2324), .CLK(clk), .RST(rst), .Q(o[39]) );
  DFF \stack_reg[1][39]  ( .D(n2323), .CLK(clk), .RST(rst), .Q(\stack[1][39] )
         );
  DFF \stack_reg[2][39]  ( .D(n2322), .CLK(clk), .RST(rst), .Q(\stack[2][39] )
         );
  DFF \stack_reg[3][39]  ( .D(n2321), .CLK(clk), .RST(rst), .Q(\stack[3][39] )
         );
  DFF \stack_reg[4][39]  ( .D(n2320), .CLK(clk), .RST(rst), .Q(\stack[4][39] )
         );
  DFF \stack_reg[5][39]  ( .D(n2319), .CLK(clk), .RST(rst), .Q(\stack[5][39] )
         );
  DFF \stack_reg[6][39]  ( .D(n2318), .CLK(clk), .RST(rst), .Q(\stack[6][39] )
         );
  DFF \stack_reg[7][39]  ( .D(n2317), .CLK(clk), .RST(rst), .Q(\stack[7][39] )
         );
  DFF \stack_reg[0][40]  ( .D(n2316), .CLK(clk), .RST(rst), .Q(o[40]) );
  DFF \stack_reg[1][40]  ( .D(n2315), .CLK(clk), .RST(rst), .Q(\stack[1][40] )
         );
  DFF \stack_reg[2][40]  ( .D(n2314), .CLK(clk), .RST(rst), .Q(\stack[2][40] )
         );
  DFF \stack_reg[3][40]  ( .D(n2313), .CLK(clk), .RST(rst), .Q(\stack[3][40] )
         );
  DFF \stack_reg[4][40]  ( .D(n2312), .CLK(clk), .RST(rst), .Q(\stack[4][40] )
         );
  DFF \stack_reg[5][40]  ( .D(n2311), .CLK(clk), .RST(rst), .Q(\stack[5][40] )
         );
  DFF \stack_reg[6][40]  ( .D(n2310), .CLK(clk), .RST(rst), .Q(\stack[6][40] )
         );
  DFF \stack_reg[7][40]  ( .D(n2309), .CLK(clk), .RST(rst), .Q(\stack[7][40] )
         );
  DFF \stack_reg[0][41]  ( .D(n2308), .CLK(clk), .RST(rst), .Q(o[41]) );
  DFF \stack_reg[1][41]  ( .D(n2307), .CLK(clk), .RST(rst), .Q(\stack[1][41] )
         );
  DFF \stack_reg[2][41]  ( .D(n2306), .CLK(clk), .RST(rst), .Q(\stack[2][41] )
         );
  DFF \stack_reg[3][41]  ( .D(n2305), .CLK(clk), .RST(rst), .Q(\stack[3][41] )
         );
  DFF \stack_reg[4][41]  ( .D(n2304), .CLK(clk), .RST(rst), .Q(\stack[4][41] )
         );
  DFF \stack_reg[5][41]  ( .D(n2303), .CLK(clk), .RST(rst), .Q(\stack[5][41] )
         );
  DFF \stack_reg[6][41]  ( .D(n2302), .CLK(clk), .RST(rst), .Q(\stack[6][41] )
         );
  DFF \stack_reg[7][41]  ( .D(n2301), .CLK(clk), .RST(rst), .Q(\stack[7][41] )
         );
  DFF \stack_reg[0][42]  ( .D(n2300), .CLK(clk), .RST(rst), .Q(o[42]) );
  DFF \stack_reg[1][42]  ( .D(n2299), .CLK(clk), .RST(rst), .Q(\stack[1][42] )
         );
  DFF \stack_reg[2][42]  ( .D(n2298), .CLK(clk), .RST(rst), .Q(\stack[2][42] )
         );
  DFF \stack_reg[3][42]  ( .D(n2297), .CLK(clk), .RST(rst), .Q(\stack[3][42] )
         );
  DFF \stack_reg[4][42]  ( .D(n2296), .CLK(clk), .RST(rst), .Q(\stack[4][42] )
         );
  DFF \stack_reg[5][42]  ( .D(n2295), .CLK(clk), .RST(rst), .Q(\stack[5][42] )
         );
  DFF \stack_reg[6][42]  ( .D(n2294), .CLK(clk), .RST(rst), .Q(\stack[6][42] )
         );
  DFF \stack_reg[7][42]  ( .D(n2293), .CLK(clk), .RST(rst), .Q(\stack[7][42] )
         );
  DFF \stack_reg[0][43]  ( .D(n2292), .CLK(clk), .RST(rst), .Q(o[43]) );
  DFF \stack_reg[1][43]  ( .D(n2291), .CLK(clk), .RST(rst), .Q(\stack[1][43] )
         );
  DFF \stack_reg[2][43]  ( .D(n2290), .CLK(clk), .RST(rst), .Q(\stack[2][43] )
         );
  DFF \stack_reg[3][43]  ( .D(n2289), .CLK(clk), .RST(rst), .Q(\stack[3][43] )
         );
  DFF \stack_reg[4][43]  ( .D(n2288), .CLK(clk), .RST(rst), .Q(\stack[4][43] )
         );
  DFF \stack_reg[5][43]  ( .D(n2287), .CLK(clk), .RST(rst), .Q(\stack[5][43] )
         );
  DFF \stack_reg[6][43]  ( .D(n2286), .CLK(clk), .RST(rst), .Q(\stack[6][43] )
         );
  DFF \stack_reg[7][43]  ( .D(n2285), .CLK(clk), .RST(rst), .Q(\stack[7][43] )
         );
  DFF \stack_reg[0][44]  ( .D(n2284), .CLK(clk), .RST(rst), .Q(o[44]) );
  DFF \stack_reg[1][44]  ( .D(n2283), .CLK(clk), .RST(rst), .Q(\stack[1][44] )
         );
  DFF \stack_reg[2][44]  ( .D(n2282), .CLK(clk), .RST(rst), .Q(\stack[2][44] )
         );
  DFF \stack_reg[3][44]  ( .D(n2281), .CLK(clk), .RST(rst), .Q(\stack[3][44] )
         );
  DFF \stack_reg[4][44]  ( .D(n2280), .CLK(clk), .RST(rst), .Q(\stack[4][44] )
         );
  DFF \stack_reg[5][44]  ( .D(n2279), .CLK(clk), .RST(rst), .Q(\stack[5][44] )
         );
  DFF \stack_reg[6][44]  ( .D(n2278), .CLK(clk), .RST(rst), .Q(\stack[6][44] )
         );
  DFF \stack_reg[7][44]  ( .D(n2277), .CLK(clk), .RST(rst), .Q(\stack[7][44] )
         );
  DFF \stack_reg[0][45]  ( .D(n2276), .CLK(clk), .RST(rst), .Q(o[45]) );
  DFF \stack_reg[1][45]  ( .D(n2275), .CLK(clk), .RST(rst), .Q(\stack[1][45] )
         );
  DFF \stack_reg[2][45]  ( .D(n2274), .CLK(clk), .RST(rst), .Q(\stack[2][45] )
         );
  DFF \stack_reg[3][45]  ( .D(n2273), .CLK(clk), .RST(rst), .Q(\stack[3][45] )
         );
  DFF \stack_reg[4][45]  ( .D(n2272), .CLK(clk), .RST(rst), .Q(\stack[4][45] )
         );
  DFF \stack_reg[5][45]  ( .D(n2271), .CLK(clk), .RST(rst), .Q(\stack[5][45] )
         );
  DFF \stack_reg[6][45]  ( .D(n2270), .CLK(clk), .RST(rst), .Q(\stack[6][45] )
         );
  DFF \stack_reg[7][45]  ( .D(n2269), .CLK(clk), .RST(rst), .Q(\stack[7][45] )
         );
  DFF \stack_reg[0][46]  ( .D(n2268), .CLK(clk), .RST(rst), .Q(o[46]) );
  DFF \stack_reg[1][46]  ( .D(n2267), .CLK(clk), .RST(rst), .Q(\stack[1][46] )
         );
  DFF \stack_reg[2][46]  ( .D(n2266), .CLK(clk), .RST(rst), .Q(\stack[2][46] )
         );
  DFF \stack_reg[3][46]  ( .D(n2265), .CLK(clk), .RST(rst), .Q(\stack[3][46] )
         );
  DFF \stack_reg[4][46]  ( .D(n2264), .CLK(clk), .RST(rst), .Q(\stack[4][46] )
         );
  DFF \stack_reg[5][46]  ( .D(n2263), .CLK(clk), .RST(rst), .Q(\stack[5][46] )
         );
  DFF \stack_reg[6][46]  ( .D(n2262), .CLK(clk), .RST(rst), .Q(\stack[6][46] )
         );
  DFF \stack_reg[7][46]  ( .D(n2261), .CLK(clk), .RST(rst), .Q(\stack[7][46] )
         );
  DFF \stack_reg[0][47]  ( .D(n2260), .CLK(clk), .RST(rst), .Q(o[47]) );
  DFF \stack_reg[1][47]  ( .D(n2259), .CLK(clk), .RST(rst), .Q(\stack[1][47] )
         );
  DFF \stack_reg[2][47]  ( .D(n2258), .CLK(clk), .RST(rst), .Q(\stack[2][47] )
         );
  DFF \stack_reg[3][47]  ( .D(n2257), .CLK(clk), .RST(rst), .Q(\stack[3][47] )
         );
  DFF \stack_reg[4][47]  ( .D(n2256), .CLK(clk), .RST(rst), .Q(\stack[4][47] )
         );
  DFF \stack_reg[5][47]  ( .D(n2255), .CLK(clk), .RST(rst), .Q(\stack[5][47] )
         );
  DFF \stack_reg[6][47]  ( .D(n2254), .CLK(clk), .RST(rst), .Q(\stack[6][47] )
         );
  DFF \stack_reg[7][47]  ( .D(n2253), .CLK(clk), .RST(rst), .Q(\stack[7][47] )
         );
  DFF \stack_reg[0][48]  ( .D(n2252), .CLK(clk), .RST(rst), .Q(o[48]) );
  DFF \stack_reg[1][48]  ( .D(n2251), .CLK(clk), .RST(rst), .Q(\stack[1][48] )
         );
  DFF \stack_reg[2][48]  ( .D(n2250), .CLK(clk), .RST(rst), .Q(\stack[2][48] )
         );
  DFF \stack_reg[3][48]  ( .D(n2249), .CLK(clk), .RST(rst), .Q(\stack[3][48] )
         );
  DFF \stack_reg[4][48]  ( .D(n2248), .CLK(clk), .RST(rst), .Q(\stack[4][48] )
         );
  DFF \stack_reg[5][48]  ( .D(n2247), .CLK(clk), .RST(rst), .Q(\stack[5][48] )
         );
  DFF \stack_reg[6][48]  ( .D(n2246), .CLK(clk), .RST(rst), .Q(\stack[6][48] )
         );
  DFF \stack_reg[7][48]  ( .D(n2245), .CLK(clk), .RST(rst), .Q(\stack[7][48] )
         );
  DFF \stack_reg[0][49]  ( .D(n2244), .CLK(clk), .RST(rst), .Q(o[49]) );
  DFF \stack_reg[1][49]  ( .D(n2243), .CLK(clk), .RST(rst), .Q(\stack[1][49] )
         );
  DFF \stack_reg[2][49]  ( .D(n2242), .CLK(clk), .RST(rst), .Q(\stack[2][49] )
         );
  DFF \stack_reg[3][49]  ( .D(n2241), .CLK(clk), .RST(rst), .Q(\stack[3][49] )
         );
  DFF \stack_reg[4][49]  ( .D(n2240), .CLK(clk), .RST(rst), .Q(\stack[4][49] )
         );
  DFF \stack_reg[5][49]  ( .D(n2239), .CLK(clk), .RST(rst), .Q(\stack[5][49] )
         );
  DFF \stack_reg[6][49]  ( .D(n2238), .CLK(clk), .RST(rst), .Q(\stack[6][49] )
         );
  DFF \stack_reg[7][49]  ( .D(n2237), .CLK(clk), .RST(rst), .Q(\stack[7][49] )
         );
  DFF \stack_reg[0][50]  ( .D(n2236), .CLK(clk), .RST(rst), .Q(o[50]) );
  DFF \stack_reg[1][50]  ( .D(n2235), .CLK(clk), .RST(rst), .Q(\stack[1][50] )
         );
  DFF \stack_reg[2][50]  ( .D(n2234), .CLK(clk), .RST(rst), .Q(\stack[2][50] )
         );
  DFF \stack_reg[3][50]  ( .D(n2233), .CLK(clk), .RST(rst), .Q(\stack[3][50] )
         );
  DFF \stack_reg[4][50]  ( .D(n2232), .CLK(clk), .RST(rst), .Q(\stack[4][50] )
         );
  DFF \stack_reg[5][50]  ( .D(n2231), .CLK(clk), .RST(rst), .Q(\stack[5][50] )
         );
  DFF \stack_reg[6][50]  ( .D(n2230), .CLK(clk), .RST(rst), .Q(\stack[6][50] )
         );
  DFF \stack_reg[7][50]  ( .D(n2229), .CLK(clk), .RST(rst), .Q(\stack[7][50] )
         );
  DFF \stack_reg[0][51]  ( .D(n2228), .CLK(clk), .RST(rst), .Q(o[51]) );
  DFF \stack_reg[1][51]  ( .D(n2227), .CLK(clk), .RST(rst), .Q(\stack[1][51] )
         );
  DFF \stack_reg[2][51]  ( .D(n2226), .CLK(clk), .RST(rst), .Q(\stack[2][51] )
         );
  DFF \stack_reg[3][51]  ( .D(n2225), .CLK(clk), .RST(rst), .Q(\stack[3][51] )
         );
  DFF \stack_reg[4][51]  ( .D(n2224), .CLK(clk), .RST(rst), .Q(\stack[4][51] )
         );
  DFF \stack_reg[5][51]  ( .D(n2223), .CLK(clk), .RST(rst), .Q(\stack[5][51] )
         );
  DFF \stack_reg[6][51]  ( .D(n2222), .CLK(clk), .RST(rst), .Q(\stack[6][51] )
         );
  DFF \stack_reg[7][51]  ( .D(n2221), .CLK(clk), .RST(rst), .Q(\stack[7][51] )
         );
  DFF \stack_reg[0][52]  ( .D(n2220), .CLK(clk), .RST(rst), .Q(o[52]) );
  DFF \stack_reg[1][52]  ( .D(n2219), .CLK(clk), .RST(rst), .Q(\stack[1][52] )
         );
  DFF \stack_reg[2][52]  ( .D(n2218), .CLK(clk), .RST(rst), .Q(\stack[2][52] )
         );
  DFF \stack_reg[3][52]  ( .D(n2217), .CLK(clk), .RST(rst), .Q(\stack[3][52] )
         );
  DFF \stack_reg[4][52]  ( .D(n2216), .CLK(clk), .RST(rst), .Q(\stack[4][52] )
         );
  DFF \stack_reg[5][52]  ( .D(n2215), .CLK(clk), .RST(rst), .Q(\stack[5][52] )
         );
  DFF \stack_reg[6][52]  ( .D(n2214), .CLK(clk), .RST(rst), .Q(\stack[6][52] )
         );
  DFF \stack_reg[7][52]  ( .D(n2213), .CLK(clk), .RST(rst), .Q(\stack[7][52] )
         );
  DFF \stack_reg[0][53]  ( .D(n2212), .CLK(clk), .RST(rst), .Q(o[53]) );
  DFF \stack_reg[1][53]  ( .D(n2211), .CLK(clk), .RST(rst), .Q(\stack[1][53] )
         );
  DFF \stack_reg[2][53]  ( .D(n2210), .CLK(clk), .RST(rst), .Q(\stack[2][53] )
         );
  DFF \stack_reg[3][53]  ( .D(n2209), .CLK(clk), .RST(rst), .Q(\stack[3][53] )
         );
  DFF \stack_reg[4][53]  ( .D(n2208), .CLK(clk), .RST(rst), .Q(\stack[4][53] )
         );
  DFF \stack_reg[5][53]  ( .D(n2207), .CLK(clk), .RST(rst), .Q(\stack[5][53] )
         );
  DFF \stack_reg[6][53]  ( .D(n2206), .CLK(clk), .RST(rst), .Q(\stack[6][53] )
         );
  DFF \stack_reg[7][53]  ( .D(n2205), .CLK(clk), .RST(rst), .Q(\stack[7][53] )
         );
  DFF \stack_reg[0][54]  ( .D(n2204), .CLK(clk), .RST(rst), .Q(o[54]) );
  DFF \stack_reg[1][54]  ( .D(n2203), .CLK(clk), .RST(rst), .Q(\stack[1][54] )
         );
  DFF \stack_reg[2][54]  ( .D(n2202), .CLK(clk), .RST(rst), .Q(\stack[2][54] )
         );
  DFF \stack_reg[3][54]  ( .D(n2201), .CLK(clk), .RST(rst), .Q(\stack[3][54] )
         );
  DFF \stack_reg[4][54]  ( .D(n2200), .CLK(clk), .RST(rst), .Q(\stack[4][54] )
         );
  DFF \stack_reg[5][54]  ( .D(n2199), .CLK(clk), .RST(rst), .Q(\stack[5][54] )
         );
  DFF \stack_reg[6][54]  ( .D(n2198), .CLK(clk), .RST(rst), .Q(\stack[6][54] )
         );
  DFF \stack_reg[7][54]  ( .D(n2197), .CLK(clk), .RST(rst), .Q(\stack[7][54] )
         );
  DFF \stack_reg[0][55]  ( .D(n2196), .CLK(clk), .RST(rst), .Q(o[55]) );
  DFF \stack_reg[1][55]  ( .D(n2195), .CLK(clk), .RST(rst), .Q(\stack[1][55] )
         );
  DFF \stack_reg[2][55]  ( .D(n2194), .CLK(clk), .RST(rst), .Q(\stack[2][55] )
         );
  DFF \stack_reg[3][55]  ( .D(n2193), .CLK(clk), .RST(rst), .Q(\stack[3][55] )
         );
  DFF \stack_reg[4][55]  ( .D(n2192), .CLK(clk), .RST(rst), .Q(\stack[4][55] )
         );
  DFF \stack_reg[5][55]  ( .D(n2191), .CLK(clk), .RST(rst), .Q(\stack[5][55] )
         );
  DFF \stack_reg[6][55]  ( .D(n2190), .CLK(clk), .RST(rst), .Q(\stack[6][55] )
         );
  DFF \stack_reg[7][55]  ( .D(n2189), .CLK(clk), .RST(rst), .Q(\stack[7][55] )
         );
  DFF \stack_reg[0][56]  ( .D(n2188), .CLK(clk), .RST(rst), .Q(o[56]) );
  DFF \stack_reg[1][56]  ( .D(n2187), .CLK(clk), .RST(rst), .Q(\stack[1][56] )
         );
  DFF \stack_reg[2][56]  ( .D(n2186), .CLK(clk), .RST(rst), .Q(\stack[2][56] )
         );
  DFF \stack_reg[3][56]  ( .D(n2185), .CLK(clk), .RST(rst), .Q(\stack[3][56] )
         );
  DFF \stack_reg[4][56]  ( .D(n2184), .CLK(clk), .RST(rst), .Q(\stack[4][56] )
         );
  DFF \stack_reg[5][56]  ( .D(n2183), .CLK(clk), .RST(rst), .Q(\stack[5][56] )
         );
  DFF \stack_reg[6][56]  ( .D(n2182), .CLK(clk), .RST(rst), .Q(\stack[6][56] )
         );
  DFF \stack_reg[7][56]  ( .D(n2181), .CLK(clk), .RST(rst), .Q(\stack[7][56] )
         );
  DFF \stack_reg[0][57]  ( .D(n2180), .CLK(clk), .RST(rst), .Q(o[57]) );
  DFF \stack_reg[1][57]  ( .D(n2179), .CLK(clk), .RST(rst), .Q(\stack[1][57] )
         );
  DFF \stack_reg[2][57]  ( .D(n2178), .CLK(clk), .RST(rst), .Q(\stack[2][57] )
         );
  DFF \stack_reg[3][57]  ( .D(n2177), .CLK(clk), .RST(rst), .Q(\stack[3][57] )
         );
  DFF \stack_reg[4][57]  ( .D(n2176), .CLK(clk), .RST(rst), .Q(\stack[4][57] )
         );
  DFF \stack_reg[5][57]  ( .D(n2175), .CLK(clk), .RST(rst), .Q(\stack[5][57] )
         );
  DFF \stack_reg[6][57]  ( .D(n2174), .CLK(clk), .RST(rst), .Q(\stack[6][57] )
         );
  DFF \stack_reg[7][57]  ( .D(n2173), .CLK(clk), .RST(rst), .Q(\stack[7][57] )
         );
  DFF \stack_reg[0][58]  ( .D(n2172), .CLK(clk), .RST(rst), .Q(o[58]) );
  DFF \stack_reg[1][58]  ( .D(n2171), .CLK(clk), .RST(rst), .Q(\stack[1][58] )
         );
  DFF \stack_reg[2][58]  ( .D(n2170), .CLK(clk), .RST(rst), .Q(\stack[2][58] )
         );
  DFF \stack_reg[3][58]  ( .D(n2169), .CLK(clk), .RST(rst), .Q(\stack[3][58] )
         );
  DFF \stack_reg[4][58]  ( .D(n2168), .CLK(clk), .RST(rst), .Q(\stack[4][58] )
         );
  DFF \stack_reg[5][58]  ( .D(n2167), .CLK(clk), .RST(rst), .Q(\stack[5][58] )
         );
  DFF \stack_reg[6][58]  ( .D(n2166), .CLK(clk), .RST(rst), .Q(\stack[6][58] )
         );
  DFF \stack_reg[7][58]  ( .D(n2165), .CLK(clk), .RST(rst), .Q(\stack[7][58] )
         );
  DFF \stack_reg[0][59]  ( .D(n2164), .CLK(clk), .RST(rst), .Q(o[59]) );
  DFF \stack_reg[1][59]  ( .D(n2163), .CLK(clk), .RST(rst), .Q(\stack[1][59] )
         );
  DFF \stack_reg[2][59]  ( .D(n2162), .CLK(clk), .RST(rst), .Q(\stack[2][59] )
         );
  DFF \stack_reg[3][59]  ( .D(n2161), .CLK(clk), .RST(rst), .Q(\stack[3][59] )
         );
  DFF \stack_reg[4][59]  ( .D(n2160), .CLK(clk), .RST(rst), .Q(\stack[4][59] )
         );
  DFF \stack_reg[5][59]  ( .D(n2159), .CLK(clk), .RST(rst), .Q(\stack[5][59] )
         );
  DFF \stack_reg[6][59]  ( .D(n2158), .CLK(clk), .RST(rst), .Q(\stack[6][59] )
         );
  DFF \stack_reg[7][59]  ( .D(n2157), .CLK(clk), .RST(rst), .Q(\stack[7][59] )
         );
  DFF \stack_reg[0][60]  ( .D(n2156), .CLK(clk), .RST(rst), .Q(o[60]) );
  DFF \stack_reg[1][60]  ( .D(n2155), .CLK(clk), .RST(rst), .Q(\stack[1][60] )
         );
  DFF \stack_reg[2][60]  ( .D(n2154), .CLK(clk), .RST(rst), .Q(\stack[2][60] )
         );
  DFF \stack_reg[3][60]  ( .D(n2153), .CLK(clk), .RST(rst), .Q(\stack[3][60] )
         );
  DFF \stack_reg[4][60]  ( .D(n2152), .CLK(clk), .RST(rst), .Q(\stack[4][60] )
         );
  DFF \stack_reg[5][60]  ( .D(n2151), .CLK(clk), .RST(rst), .Q(\stack[5][60] )
         );
  DFF \stack_reg[6][60]  ( .D(n2150), .CLK(clk), .RST(rst), .Q(\stack[6][60] )
         );
  DFF \stack_reg[7][60]  ( .D(n2149), .CLK(clk), .RST(rst), .Q(\stack[7][60] )
         );
  DFF \stack_reg[0][61]  ( .D(n2148), .CLK(clk), .RST(rst), .Q(o[61]) );
  DFF \stack_reg[1][61]  ( .D(n2147), .CLK(clk), .RST(rst), .Q(\stack[1][61] )
         );
  DFF \stack_reg[2][61]  ( .D(n2146), .CLK(clk), .RST(rst), .Q(\stack[2][61] )
         );
  DFF \stack_reg[3][61]  ( .D(n2145), .CLK(clk), .RST(rst), .Q(\stack[3][61] )
         );
  DFF \stack_reg[4][61]  ( .D(n2144), .CLK(clk), .RST(rst), .Q(\stack[4][61] )
         );
  DFF \stack_reg[5][61]  ( .D(n2143), .CLK(clk), .RST(rst), .Q(\stack[5][61] )
         );
  DFF \stack_reg[6][61]  ( .D(n2142), .CLK(clk), .RST(rst), .Q(\stack[6][61] )
         );
  DFF \stack_reg[7][61]  ( .D(n2141), .CLK(clk), .RST(rst), .Q(\stack[7][61] )
         );
  DFF \stack_reg[0][62]  ( .D(n2140), .CLK(clk), .RST(rst), .Q(o[62]) );
  DFF \stack_reg[1][62]  ( .D(n2139), .CLK(clk), .RST(rst), .Q(\stack[1][62] )
         );
  DFF \stack_reg[2][62]  ( .D(n2138), .CLK(clk), .RST(rst), .Q(\stack[2][62] )
         );
  DFF \stack_reg[3][62]  ( .D(n2137), .CLK(clk), .RST(rst), .Q(\stack[3][62] )
         );
  DFF \stack_reg[4][62]  ( .D(n2136), .CLK(clk), .RST(rst), .Q(\stack[4][62] )
         );
  DFF \stack_reg[5][62]  ( .D(n2135), .CLK(clk), .RST(rst), .Q(\stack[5][62] )
         );
  DFF \stack_reg[6][62]  ( .D(n2134), .CLK(clk), .RST(rst), .Q(\stack[6][62] )
         );
  DFF \stack_reg[7][62]  ( .D(n2133), .CLK(clk), .RST(rst), .Q(\stack[7][62] )
         );
  DFF \stack_reg[0][63]  ( .D(n2132), .CLK(clk), .RST(rst), .Q(o[63]) );
  DFF \stack_reg[1][63]  ( .D(n2131), .CLK(clk), .RST(rst), .Q(\stack[1][63] )
         );
  DFF \stack_reg[2][63]  ( .D(n2130), .CLK(clk), .RST(rst), .Q(\stack[2][63] )
         );
  DFF \stack_reg[3][63]  ( .D(n2129), .CLK(clk), .RST(rst), .Q(\stack[3][63] )
         );
  DFF \stack_reg[4][63]  ( .D(n2128), .CLK(clk), .RST(rst), .Q(\stack[4][63] )
         );
  DFF \stack_reg[5][63]  ( .D(n2127), .CLK(clk), .RST(rst), .Q(\stack[5][63] )
         );
  DFF \stack_reg[6][63]  ( .D(n2126), .CLK(clk), .RST(rst), .Q(\stack[6][63] )
         );
  DFF \stack_reg[7][63]  ( .D(n2125), .CLK(clk), .RST(rst), .Q(\stack[7][63] )
         );
  DFF \stack_reg[2][0]  ( .D(n2124), .CLK(clk), .RST(rst), .Q(\stack[2][0] )
         );
  DFF \stack_reg[3][0]  ( .D(n2123), .CLK(clk), .RST(rst), .Q(\stack[3][0] )
         );
  DFF \stack_reg[4][0]  ( .D(n2122), .CLK(clk), .RST(rst), .Q(\stack[4][0] )
         );
  DFF \stack_reg[5][0]  ( .D(n2121), .CLK(clk), .RST(rst), .Q(\stack[5][0] )
         );
  DFF \stack_reg[6][0]  ( .D(n2120), .CLK(clk), .RST(rst), .Q(\stack[6][0] )
         );
  DFF \stack_reg[7][0]  ( .D(n2119), .CLK(clk), .RST(rst), .Q(\stack[7][0] )
         );
  XOR \DP_OP_25_64_8855/U383  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_0 ), .Z(
        \DP_OP_25_64_8855/n656 ) );
  XOR \DP_OP_25_64_8855/U382  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_1 ), .Z(
        \DP_OP_25_64_8855/n655 ) );
  XOR \DP_OP_25_64_8855/U381  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_2 ), .Z(
        \DP_OP_25_64_8855/n654 ) );
  XOR \DP_OP_25_64_8855/U380  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_3 ), .Z(
        \DP_OP_25_64_8855/n653 ) );
  XOR \DP_OP_25_64_8855/U379  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_4 ), .Z(
        \DP_OP_25_64_8855/n652 ) );
  XOR \DP_OP_25_64_8855/U378  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_5 ), .Z(
        \DP_OP_25_64_8855/n651 ) );
  XOR \DP_OP_25_64_8855/U377  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_6 ), .Z(
        \DP_OP_25_64_8855/n650 ) );
  XOR \DP_OP_25_64_8855/U376  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_7 ), .Z(
        \DP_OP_25_64_8855/n649 ) );
  XOR \DP_OP_25_64_8855/U375  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_8 ), .Z(
        \DP_OP_25_64_8855/n648 ) );
  XOR \DP_OP_25_64_8855/U374  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_9 ), .Z(
        \DP_OP_25_64_8855/n647 ) );
  XOR \DP_OP_25_64_8855/U373  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_10 ), .Z(
        \DP_OP_25_64_8855/n646 ) );
  XOR \DP_OP_25_64_8855/U372  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_11 ), .Z(
        \DP_OP_25_64_8855/n645 ) );
  XOR \DP_OP_25_64_8855/U371  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_12 ), .Z(
        \DP_OP_25_64_8855/n644 ) );
  XOR \DP_OP_25_64_8855/U370  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_13 ), .Z(
        \DP_OP_25_64_8855/n643 ) );
  XOR \DP_OP_25_64_8855/U369  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_14 ), .Z(
        \DP_OP_25_64_8855/n642 ) );
  XOR \DP_OP_25_64_8855/U368  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_15 ), .Z(
        \DP_OP_25_64_8855/n641 ) );
  XOR \DP_OP_25_64_8855/U367  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_16 ), .Z(
        \DP_OP_25_64_8855/n640 ) );
  XOR \DP_OP_25_64_8855/U366  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_17 ), .Z(
        \DP_OP_25_64_8855/n639 ) );
  XOR \DP_OP_25_64_8855/U365  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_18 ), .Z(
        \DP_OP_25_64_8855/n638 ) );
  XOR \DP_OP_25_64_8855/U364  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_19 ), .Z(
        \DP_OP_25_64_8855/n637 ) );
  XOR \DP_OP_25_64_8855/U363  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_20 ), .Z(
        \DP_OP_25_64_8855/n636 ) );
  XOR \DP_OP_25_64_8855/U309  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_21 ), .Z(
        \DP_OP_25_64_8855/n635 ) );
  XOR \DP_OP_25_64_8855/U308  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_22 ), .Z(
        \DP_OP_25_64_8855/n634 ) );
  XOR \DP_OP_25_64_8855/U307  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_23 ), .Z(
        \DP_OP_25_64_8855/n633 ) );
  XOR \DP_OP_25_64_8855/U306  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_24 ), .Z(
        \DP_OP_25_64_8855/n632 ) );
  XOR \DP_OP_25_64_8855/U305  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_25 ), .Z(
        \DP_OP_25_64_8855/n631 ) );
  XOR \DP_OP_25_64_8855/U304  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_26 ), .Z(
        \DP_OP_25_64_8855/n630 ) );
  XOR \DP_OP_25_64_8855/U303  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_27 ), .Z(
        \DP_OP_25_64_8855/n629 ) );
  XOR \DP_OP_25_64_8855/U302  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_28 ), .Z(
        \DP_OP_25_64_8855/n628 ) );
  XOR \DP_OP_25_64_8855/U301  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_29 ), .Z(
        \DP_OP_25_64_8855/n627 ) );
  XOR \DP_OP_25_64_8855/U300  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_30 ), .Z(
        \DP_OP_25_64_8855/n626 ) );
  XOR \DP_OP_25_64_8855/U299  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_31 ), .Z(
        \DP_OP_25_64_8855/n625 ) );
  XOR \DP_OP_25_64_8855/U298  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_32 ), .Z(
        \DP_OP_25_64_8855/n624 ) );
  XOR \DP_OP_25_64_8855/U297  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_33 ), .Z(
        \DP_OP_25_64_8855/n623 ) );
  XOR \DP_OP_25_64_8855/U296  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_34 ), .Z(
        \DP_OP_25_64_8855/n622 ) );
  XOR \DP_OP_25_64_8855/U295  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_35 ), .Z(
        \DP_OP_25_64_8855/n621 ) );
  XOR \DP_OP_25_64_8855/U294  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_36 ), .Z(
        \DP_OP_25_64_8855/n620 ) );
  XOR \DP_OP_25_64_8855/U293  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_37 ), .Z(
        \DP_OP_25_64_8855/n619 ) );
  XOR \DP_OP_25_64_8855/U292  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_38 ), .Z(
        \DP_OP_25_64_8855/n618 ) );
  XOR \DP_OP_25_64_8855/U291  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_39 ), .Z(
        \DP_OP_25_64_8855/n617 ) );
  XOR \DP_OP_25_64_8855/U290  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_40 ), .Z(
        \DP_OP_25_64_8855/n616 ) );
  XOR \DP_OP_25_64_8855/U289  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_41 ), .Z(
        \DP_OP_25_64_8855/n615 ) );
  XOR \DP_OP_25_64_8855/U288  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_42 ), .Z(
        \DP_OP_25_64_8855/n614 ) );
  XOR \DP_OP_25_64_8855/U287  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_43 ), .Z(
        \DP_OP_25_64_8855/n613 ) );
  XOR \DP_OP_25_64_8855/U286  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_44 ), .Z(
        \DP_OP_25_64_8855/n612 ) );
  XOR \DP_OP_25_64_8855/U285  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_45 ), .Z(
        \DP_OP_25_64_8855/n611 ) );
  XOR \DP_OP_25_64_8855/U284  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_46 ), .Z(
        \DP_OP_25_64_8855/n610 ) );
  XOR \DP_OP_25_64_8855/U283  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_47 ), .Z(
        \DP_OP_25_64_8855/n609 ) );
  XOR \DP_OP_25_64_8855/U282  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_48 ), .Z(
        \DP_OP_25_64_8855/n608 ) );
  XOR \DP_OP_25_64_8855/U281  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_49 ), .Z(
        \DP_OP_25_64_8855/n607 ) );
  XOR \DP_OP_25_64_8855/U280  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_50 ), .Z(
        \DP_OP_25_64_8855/n606 ) );
  XOR \DP_OP_25_64_8855/U279  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_51 ), .Z(
        \DP_OP_25_64_8855/n605 ) );
  XOR \DP_OP_25_64_8855/U278  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_52 ), .Z(
        \DP_OP_25_64_8855/n604 ) );
  XOR \DP_OP_25_64_8855/U277  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_53 ), .Z(
        \DP_OP_25_64_8855/n603 ) );
  XOR \DP_OP_25_64_8855/U276  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_54 ), .Z(
        \DP_OP_25_64_8855/n602 ) );
  XOR \DP_OP_25_64_8855/U275  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_55 ), .Z(
        \DP_OP_25_64_8855/n601 ) );
  XOR \DP_OP_25_64_8855/U274  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_56 ), .Z(
        \DP_OP_25_64_8855/n600 ) );
  XOR \DP_OP_25_64_8855/U273  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_57 ), .Z(
        \DP_OP_25_64_8855/n599 ) );
  XOR \DP_OP_25_64_8855/U272  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_58 ), .Z(
        \DP_OP_25_64_8855/n598 ) );
  XOR \DP_OP_25_64_8855/U271  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_59 ), .Z(
        \DP_OP_25_64_8855/n597 ) );
  XOR \DP_OP_25_64_8855/U270  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_60 ), .Z(
        \DP_OP_25_64_8855/n596 ) );
  XOR \DP_OP_25_64_8855/U269  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_61 ), .Z(
        \DP_OP_25_64_8855/n595 ) );
  XOR \DP_OP_25_64_8855/U268  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_62 ), .Z(
        \DP_OP_25_64_8855/n594 ) );
  XOR \DP_OP_25_64_8855/U267  ( .A(\C1/Z_0 ), .B(\U1/RSOP_16/C3/Z_63 ), .Z(
        \DP_OP_25_64_8855/n593 ) );
  XOR \DP_OP_25_64_8855/U264  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_8855/n525 ) );
  XOR \DP_OP_25_64_8855/U263  ( .A(\DP_OP_25_64_8855/n525 ), .B(
        \DP_OP_25_64_8855/n656 ), .Z(\C3/DATA5_0 ) );
  XOR \DP_OP_25_64_8855/U209  ( .A(\DP_OP_25_64_8855/n655 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_8855/n524 ) );
  XOR \DP_OP_25_64_8855/U208  ( .A(\DP_OP_25_64_8855/n588 ), .B(
        \DP_OP_25_64_8855/n524 ), .Z(\C3/DATA5_1 ) );
  XOR \DP_OP_25_64_8855/U207  ( .A(\DP_OP_25_64_8855/n654 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_8855/n523 ) );
  XOR \DP_OP_25_64_8855/U206  ( .A(\DP_OP_25_64_8855/n587 ), .B(
        \DP_OP_25_64_8855/n523 ), .Z(\C3/DATA5_2 ) );
  XOR \DP_OP_25_64_8855/U205  ( .A(\DP_OP_25_64_8855/n653 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_8855/n522 ) );
  XOR \DP_OP_25_64_8855/U204  ( .A(\DP_OP_25_64_8855/n586 ), .B(
        \DP_OP_25_64_8855/n522 ), .Z(\C3/DATA5_3 ) );
  XOR \DP_OP_25_64_8855/U203  ( .A(\DP_OP_25_64_8855/n652 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_8855/n521 ) );
  XOR \DP_OP_25_64_8855/U202  ( .A(\DP_OP_25_64_8855/n585 ), .B(
        \DP_OP_25_64_8855/n521 ), .Z(\C3/DATA5_4 ) );
  XOR \DP_OP_25_64_8855/U201  ( .A(\DP_OP_25_64_8855/n651 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_8855/n520 ) );
  XOR \DP_OP_25_64_8855/U200  ( .A(\DP_OP_25_64_8855/n584 ), .B(
        \DP_OP_25_64_8855/n520 ), .Z(\C3/DATA5_5 ) );
  XOR \DP_OP_25_64_8855/U199  ( .A(\DP_OP_25_64_8855/n650 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_8855/n519 ) );
  XOR \DP_OP_25_64_8855/U198  ( .A(\DP_OP_25_64_8855/n583 ), .B(
        \DP_OP_25_64_8855/n519 ), .Z(\C3/DATA5_6 ) );
  XOR \DP_OP_25_64_8855/U197  ( .A(\DP_OP_25_64_8855/n649 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_8855/n518 ) );
  XOR \DP_OP_25_64_8855/U196  ( .A(\DP_OP_25_64_8855/n582 ), .B(
        \DP_OP_25_64_8855/n518 ), .Z(\C3/DATA5_7 ) );
  XOR \DP_OP_25_64_8855/U195  ( .A(\DP_OP_25_64_8855/n648 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_8855/n517 ) );
  XOR \DP_OP_25_64_8855/U194  ( .A(\DP_OP_25_64_8855/n581 ), .B(
        \DP_OP_25_64_8855/n517 ), .Z(\C3/DATA5_8 ) );
  XOR \DP_OP_25_64_8855/U193  ( .A(\DP_OP_25_64_8855/n647 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_8855/n516 ) );
  XOR \DP_OP_25_64_8855/U192  ( .A(\DP_OP_25_64_8855/n580 ), .B(
        \DP_OP_25_64_8855/n516 ), .Z(\C3/DATA5_9 ) );
  XOR \DP_OP_25_64_8855/U191  ( .A(\DP_OP_25_64_8855/n646 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_8855/n515 ) );
  XOR \DP_OP_25_64_8855/U190  ( .A(\DP_OP_25_64_8855/n579 ), .B(
        \DP_OP_25_64_8855/n515 ), .Z(\C3/DATA5_10 ) );
  XOR \DP_OP_25_64_8855/U189  ( .A(\DP_OP_25_64_8855/n645 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_8855/n514 ) );
  XOR \DP_OP_25_64_8855/U188  ( .A(\DP_OP_25_64_8855/n578 ), .B(
        \DP_OP_25_64_8855/n514 ), .Z(\C3/DATA5_11 ) );
  XOR \DP_OP_25_64_8855/U187  ( .A(\DP_OP_25_64_8855/n644 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_8855/n513 ) );
  XOR \DP_OP_25_64_8855/U186  ( .A(\DP_OP_25_64_8855/n577 ), .B(
        \DP_OP_25_64_8855/n513 ), .Z(\C3/DATA5_12 ) );
  XOR \DP_OP_25_64_8855/U185  ( .A(\DP_OP_25_64_8855/n643 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_8855/n512 ) );
  XOR \DP_OP_25_64_8855/U184  ( .A(\DP_OP_25_64_8855/n576 ), .B(
        \DP_OP_25_64_8855/n512 ), .Z(\C3/DATA5_13 ) );
  XOR \DP_OP_25_64_8855/U183  ( .A(\DP_OP_25_64_8855/n642 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_8855/n511 ) );
  XOR \DP_OP_25_64_8855/U182  ( .A(\DP_OP_25_64_8855/n575 ), .B(
        \DP_OP_25_64_8855/n511 ), .Z(\C3/DATA5_14 ) );
  XOR \DP_OP_25_64_8855/U181  ( .A(\DP_OP_25_64_8855/n641 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_8855/n510 ) );
  XOR \DP_OP_25_64_8855/U180  ( .A(\DP_OP_25_64_8855/n574 ), .B(
        \DP_OP_25_64_8855/n510 ), .Z(\C3/DATA5_15 ) );
  XOR \DP_OP_25_64_8855/U179  ( .A(\DP_OP_25_64_8855/n640 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_8855/n509 ) );
  XOR \DP_OP_25_64_8855/U178  ( .A(\DP_OP_25_64_8855/n573 ), .B(
        \DP_OP_25_64_8855/n509 ), .Z(\C3/DATA5_16 ) );
  XOR \DP_OP_25_64_8855/U177  ( .A(\DP_OP_25_64_8855/n639 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_8855/n508 ) );
  XOR \DP_OP_25_64_8855/U176  ( .A(\DP_OP_25_64_8855/n572 ), .B(
        \DP_OP_25_64_8855/n508 ), .Z(\C3/DATA5_17 ) );
  XOR \DP_OP_25_64_8855/U175  ( .A(\DP_OP_25_64_8855/n638 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_8855/n507 ) );
  XOR \DP_OP_25_64_8855/U174  ( .A(\DP_OP_25_64_8855/n571 ), .B(
        \DP_OP_25_64_8855/n507 ), .Z(\C3/DATA5_18 ) );
  XOR \DP_OP_25_64_8855/U173  ( .A(\DP_OP_25_64_8855/n637 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_8855/n506 ) );
  XOR \DP_OP_25_64_8855/U172  ( .A(\DP_OP_25_64_8855/n570 ), .B(
        \DP_OP_25_64_8855/n506 ), .Z(\C3/DATA5_19 ) );
  XOR \DP_OP_25_64_8855/U171  ( .A(\DP_OP_25_64_8855/n636 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_8855/n505 ) );
  XOR \DP_OP_25_64_8855/U170  ( .A(\DP_OP_25_64_8855/n569 ), .B(
        \DP_OP_25_64_8855/n505 ), .Z(\C3/DATA5_20 ) );
  XOR \DP_OP_25_64_8855/U169  ( .A(\DP_OP_25_64_8855/n635 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_8855/n504 ) );
  XOR \DP_OP_25_64_8855/U168  ( .A(\DP_OP_25_64_8855/n568 ), .B(
        \DP_OP_25_64_8855/n504 ), .Z(\C3/DATA5_21 ) );
  XOR \DP_OP_25_64_8855/U167  ( .A(\DP_OP_25_64_8855/n634 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_8855/n503 ) );
  XOR \DP_OP_25_64_8855/U166  ( .A(\DP_OP_25_64_8855/n567 ), .B(
        \DP_OP_25_64_8855/n503 ), .Z(\C3/DATA5_22 ) );
  XOR \DP_OP_25_64_8855/U165  ( .A(\DP_OP_25_64_8855/n633 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_8855/n502 ) );
  XOR \DP_OP_25_64_8855/U164  ( .A(\DP_OP_25_64_8855/n566 ), .B(
        \DP_OP_25_64_8855/n502 ), .Z(\C3/DATA5_23 ) );
  XOR \DP_OP_25_64_8855/U163  ( .A(\DP_OP_25_64_8855/n632 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_8855/n501 ) );
  XOR \DP_OP_25_64_8855/U109  ( .A(\DP_OP_25_64_8855/n565 ), .B(
        \DP_OP_25_64_8855/n501 ), .Z(\C3/DATA5_24 ) );
  XOR \DP_OP_25_64_8855/U108  ( .A(\DP_OP_25_64_8855/n631 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_8855/n500 ) );
  XOR \DP_OP_25_64_8855/U107  ( .A(\DP_OP_25_64_8855/n564 ), .B(
        \DP_OP_25_64_8855/n500 ), .Z(\C3/DATA5_25 ) );
  XOR \DP_OP_25_64_8855/U106  ( .A(\DP_OP_25_64_8855/n630 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_8855/n499 ) );
  XOR \DP_OP_25_64_8855/U105  ( .A(\DP_OP_25_64_8855/n563 ), .B(
        \DP_OP_25_64_8855/n499 ), .Z(\C3/DATA5_26 ) );
  XOR \DP_OP_25_64_8855/U104  ( .A(\DP_OP_25_64_8855/n629 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_8855/n498 ) );
  XOR \DP_OP_25_64_8855/U103  ( .A(\DP_OP_25_64_8855/n562 ), .B(
        \DP_OP_25_64_8855/n498 ), .Z(\C3/DATA5_27 ) );
  XOR \DP_OP_25_64_8855/U102  ( .A(\DP_OP_25_64_8855/n628 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_8855/n497 ) );
  XOR \DP_OP_25_64_8855/U101  ( .A(\DP_OP_25_64_8855/n561 ), .B(
        \DP_OP_25_64_8855/n497 ), .Z(\C3/DATA5_28 ) );
  XOR \DP_OP_25_64_8855/U100  ( .A(\DP_OP_25_64_8855/n627 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_8855/n496 ) );
  XOR \DP_OP_25_64_8855/U99  ( .A(\DP_OP_25_64_8855/n560 ), .B(
        \DP_OP_25_64_8855/n496 ), .Z(\C3/DATA5_29 ) );
  XOR \DP_OP_25_64_8855/U98  ( .A(\DP_OP_25_64_8855/n626 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_8855/n495 ) );
  XOR \DP_OP_25_64_8855/U97  ( .A(\DP_OP_25_64_8855/n559 ), .B(
        \DP_OP_25_64_8855/n495 ), .Z(\C3/DATA5_30 ) );
  XOR \DP_OP_25_64_8855/U96  ( .A(\DP_OP_25_64_8855/n625 ), .B(
        \U1/RSOP_16/C2/Z_31 ), .Z(\DP_OP_25_64_8855/n494 ) );
  XOR \DP_OP_25_64_8855/U95  ( .A(\DP_OP_25_64_8855/n558 ), .B(
        \DP_OP_25_64_8855/n494 ), .Z(\C3/DATA5_31 ) );
  XOR \DP_OP_25_64_8855/U94  ( .A(\DP_OP_25_64_8855/n624 ), .B(
        \U1/RSOP_16/C2/Z_32 ), .Z(\DP_OP_25_64_8855/n493 ) );
  XOR \DP_OP_25_64_8855/U93  ( .A(\DP_OP_25_64_8855/n557 ), .B(
        \DP_OP_25_64_8855/n493 ), .Z(\C3/DATA5_32 ) );
  XOR \DP_OP_25_64_8855/U92  ( .A(\DP_OP_25_64_8855/n623 ), .B(
        \U1/RSOP_16/C2/Z_33 ), .Z(\DP_OP_25_64_8855/n492 ) );
  XOR \DP_OP_25_64_8855/U91  ( .A(\DP_OP_25_64_8855/n556 ), .B(
        \DP_OP_25_64_8855/n492 ), .Z(\C3/DATA5_33 ) );
  XOR \DP_OP_25_64_8855/U90  ( .A(\DP_OP_25_64_8855/n622 ), .B(
        \U1/RSOP_16/C2/Z_34 ), .Z(\DP_OP_25_64_8855/n491 ) );
  XOR \DP_OP_25_64_8855/U89  ( .A(\DP_OP_25_64_8855/n555 ), .B(
        \DP_OP_25_64_8855/n491 ), .Z(\C3/DATA5_34 ) );
  XOR \DP_OP_25_64_8855/U88  ( .A(\DP_OP_25_64_8855/n621 ), .B(
        \U1/RSOP_16/C2/Z_35 ), .Z(\DP_OP_25_64_8855/n490 ) );
  XOR \DP_OP_25_64_8855/U87  ( .A(\DP_OP_25_64_8855/n554 ), .B(
        \DP_OP_25_64_8855/n490 ), .Z(\C3/DATA5_35 ) );
  XOR \DP_OP_25_64_8855/U86  ( .A(\DP_OP_25_64_8855/n620 ), .B(
        \U1/RSOP_16/C2/Z_36 ), .Z(\DP_OP_25_64_8855/n489 ) );
  XOR \DP_OP_25_64_8855/U85  ( .A(\DP_OP_25_64_8855/n553 ), .B(
        \DP_OP_25_64_8855/n489 ), .Z(\C3/DATA5_36 ) );
  XOR \DP_OP_25_64_8855/U84  ( .A(\DP_OP_25_64_8855/n619 ), .B(
        \U1/RSOP_16/C2/Z_37 ), .Z(\DP_OP_25_64_8855/n488 ) );
  XOR \DP_OP_25_64_8855/U83  ( .A(\DP_OP_25_64_8855/n552 ), .B(
        \DP_OP_25_64_8855/n488 ), .Z(\C3/DATA5_37 ) );
  XOR \DP_OP_25_64_8855/U82  ( .A(\DP_OP_25_64_8855/n618 ), .B(
        \U1/RSOP_16/C2/Z_38 ), .Z(\DP_OP_25_64_8855/n487 ) );
  XOR \DP_OP_25_64_8855/U81  ( .A(\DP_OP_25_64_8855/n551 ), .B(
        \DP_OP_25_64_8855/n487 ), .Z(\C3/DATA5_38 ) );
  XOR \DP_OP_25_64_8855/U80  ( .A(\DP_OP_25_64_8855/n617 ), .B(
        \U1/RSOP_16/C2/Z_39 ), .Z(\DP_OP_25_64_8855/n486 ) );
  XOR \DP_OP_25_64_8855/U79  ( .A(\DP_OP_25_64_8855/n550 ), .B(
        \DP_OP_25_64_8855/n486 ), .Z(\C3/DATA5_39 ) );
  XOR \DP_OP_25_64_8855/U78  ( .A(\DP_OP_25_64_8855/n616 ), .B(
        \U1/RSOP_16/C2/Z_40 ), .Z(\DP_OP_25_64_8855/n485 ) );
  XOR \DP_OP_25_64_8855/U77  ( .A(\DP_OP_25_64_8855/n549 ), .B(
        \DP_OP_25_64_8855/n485 ), .Z(\C3/DATA5_40 ) );
  XOR \DP_OP_25_64_8855/U76  ( .A(\DP_OP_25_64_8855/n615 ), .B(
        \U1/RSOP_16/C2/Z_41 ), .Z(\DP_OP_25_64_8855/n484 ) );
  XOR \DP_OP_25_64_8855/U75  ( .A(\DP_OP_25_64_8855/n548 ), .B(
        \DP_OP_25_64_8855/n484 ), .Z(\C3/DATA5_41 ) );
  XOR \DP_OP_25_64_8855/U74  ( .A(\DP_OP_25_64_8855/n614 ), .B(
        \U1/RSOP_16/C2/Z_42 ), .Z(\DP_OP_25_64_8855/n483 ) );
  XOR \DP_OP_25_64_8855/U73  ( .A(\DP_OP_25_64_8855/n547 ), .B(
        \DP_OP_25_64_8855/n483 ), .Z(\C3/DATA5_42 ) );
  XOR \DP_OP_25_64_8855/U72  ( .A(\DP_OP_25_64_8855/n613 ), .B(
        \U1/RSOP_16/C2/Z_43 ), .Z(\DP_OP_25_64_8855/n482 ) );
  XOR \DP_OP_25_64_8855/U71  ( .A(\DP_OP_25_64_8855/n546 ), .B(
        \DP_OP_25_64_8855/n482 ), .Z(\C3/DATA5_43 ) );
  XOR \DP_OP_25_64_8855/U70  ( .A(\DP_OP_25_64_8855/n612 ), .B(
        \U1/RSOP_16/C2/Z_44 ), .Z(\DP_OP_25_64_8855/n481 ) );
  XOR \DP_OP_25_64_8855/U69  ( .A(\DP_OP_25_64_8855/n545 ), .B(
        \DP_OP_25_64_8855/n481 ), .Z(\C3/DATA5_44 ) );
  XOR \DP_OP_25_64_8855/U68  ( .A(\DP_OP_25_64_8855/n611 ), .B(
        \U1/RSOP_16/C2/Z_45 ), .Z(\DP_OP_25_64_8855/n480 ) );
  XOR \DP_OP_25_64_8855/U67  ( .A(\DP_OP_25_64_8855/n544 ), .B(
        \DP_OP_25_64_8855/n480 ), .Z(\C3/DATA5_45 ) );
  XOR \DP_OP_25_64_8855/U66  ( .A(\DP_OP_25_64_8855/n610 ), .B(
        \U1/RSOP_16/C2/Z_46 ), .Z(\DP_OP_25_64_8855/n479 ) );
  XOR \DP_OP_25_64_8855/U65  ( .A(\DP_OP_25_64_8855/n543 ), .B(
        \DP_OP_25_64_8855/n479 ), .Z(\C3/DATA5_46 ) );
  XOR \DP_OP_25_64_8855/U64  ( .A(\DP_OP_25_64_8855/n609 ), .B(
        \U1/RSOP_16/C2/Z_47 ), .Z(\DP_OP_25_64_8855/n478 ) );
  XOR \DP_OP_25_64_8855/U63  ( .A(\DP_OP_25_64_8855/n542 ), .B(
        \DP_OP_25_64_8855/n478 ), .Z(\C3/DATA5_47 ) );
  XOR \DP_OP_25_64_8855/U62  ( .A(\DP_OP_25_64_8855/n608 ), .B(
        \U1/RSOP_16/C2/Z_48 ), .Z(\DP_OP_25_64_8855/n477 ) );
  XOR \DP_OP_25_64_8855/U61  ( .A(\DP_OP_25_64_8855/n541 ), .B(
        \DP_OP_25_64_8855/n477 ), .Z(\C3/DATA5_48 ) );
  XOR \DP_OP_25_64_8855/U60  ( .A(\DP_OP_25_64_8855/n607 ), .B(
        \U1/RSOP_16/C2/Z_49 ), .Z(\DP_OP_25_64_8855/n476 ) );
  XOR \DP_OP_25_64_8855/U59  ( .A(\DP_OP_25_64_8855/n540 ), .B(
        \DP_OP_25_64_8855/n476 ), .Z(\C3/DATA5_49 ) );
  XOR \DP_OP_25_64_8855/U58  ( .A(\DP_OP_25_64_8855/n606 ), .B(
        \U1/RSOP_16/C2/Z_50 ), .Z(\DP_OP_25_64_8855/n475 ) );
  XOR \DP_OP_25_64_8855/U57  ( .A(\DP_OP_25_64_8855/n539 ), .B(
        \DP_OP_25_64_8855/n475 ), .Z(\C3/DATA5_50 ) );
  XOR \DP_OP_25_64_8855/U56  ( .A(\DP_OP_25_64_8855/n605 ), .B(
        \U1/RSOP_16/C2/Z_51 ), .Z(\DP_OP_25_64_8855/n474 ) );
  XOR \DP_OP_25_64_8855/U55  ( .A(\DP_OP_25_64_8855/n538 ), .B(
        \DP_OP_25_64_8855/n474 ), .Z(\C3/DATA5_51 ) );
  XOR \DP_OP_25_64_8855/U54  ( .A(\DP_OP_25_64_8855/n604 ), .B(
        \U1/RSOP_16/C2/Z_52 ), .Z(\DP_OP_25_64_8855/n473 ) );
  XOR \DP_OP_25_64_8855/U53  ( .A(\DP_OP_25_64_8855/n537 ), .B(
        \DP_OP_25_64_8855/n473 ), .Z(\C3/DATA5_52 ) );
  XOR \DP_OP_25_64_8855/U52  ( .A(\DP_OP_25_64_8855/n603 ), .B(
        \U1/RSOP_16/C2/Z_53 ), .Z(\DP_OP_25_64_8855/n472 ) );
  XOR \DP_OP_25_64_8855/U51  ( .A(\DP_OP_25_64_8855/n536 ), .B(
        \DP_OP_25_64_8855/n472 ), .Z(\C3/DATA5_53 ) );
  XOR \DP_OP_25_64_8855/U50  ( .A(\DP_OP_25_64_8855/n602 ), .B(
        \U1/RSOP_16/C2/Z_54 ), .Z(\DP_OP_25_64_8855/n471 ) );
  XOR \DP_OP_25_64_8855/U49  ( .A(\DP_OP_25_64_8855/n535 ), .B(
        \DP_OP_25_64_8855/n471 ), .Z(\C3/DATA5_54 ) );
  XOR \DP_OP_25_64_8855/U48  ( .A(\DP_OP_25_64_8855/n601 ), .B(
        \U1/RSOP_16/C2/Z_55 ), .Z(\DP_OP_25_64_8855/n470 ) );
  XOR \DP_OP_25_64_8855/U47  ( .A(\DP_OP_25_64_8855/n534 ), .B(
        \DP_OP_25_64_8855/n470 ), .Z(\C3/DATA5_55 ) );
  XOR \DP_OP_25_64_8855/U46  ( .A(\DP_OP_25_64_8855/n600 ), .B(
        \U1/RSOP_16/C2/Z_56 ), .Z(\DP_OP_25_64_8855/n469 ) );
  XOR \DP_OP_25_64_8855/U45  ( .A(\DP_OP_25_64_8855/n533 ), .B(
        \DP_OP_25_64_8855/n469 ), .Z(\C3/DATA5_56 ) );
  XOR \DP_OP_25_64_8855/U44  ( .A(\DP_OP_25_64_8855/n599 ), .B(
        \U1/RSOP_16/C2/Z_57 ), .Z(\DP_OP_25_64_8855/n468 ) );
  XOR \DP_OP_25_64_8855/U43  ( .A(\DP_OP_25_64_8855/n532 ), .B(
        \DP_OP_25_64_8855/n468 ), .Z(\C3/DATA5_57 ) );
  XOR \DP_OP_25_64_8855/U42  ( .A(\DP_OP_25_64_8855/n598 ), .B(
        \U1/RSOP_16/C2/Z_58 ), .Z(\DP_OP_25_64_8855/n467 ) );
  XOR \DP_OP_25_64_8855/U41  ( .A(\DP_OP_25_64_8855/n531 ), .B(
        \DP_OP_25_64_8855/n467 ), .Z(\C3/DATA5_58 ) );
  XOR \DP_OP_25_64_8855/U40  ( .A(\DP_OP_25_64_8855/n597 ), .B(
        \U1/RSOP_16/C2/Z_59 ), .Z(\DP_OP_25_64_8855/n466 ) );
  XOR \DP_OP_25_64_8855/U30  ( .A(\DP_OP_25_64_8855/n530 ), .B(
        \DP_OP_25_64_8855/n466 ), .Z(\C3/DATA5_59 ) );
  XOR \DP_OP_25_64_8855/U20  ( .A(\DP_OP_25_64_8855/n596 ), .B(
        \U1/RSOP_16/C2/Z_60 ), .Z(\DP_OP_25_64_8855/n465 ) );
  XOR \DP_OP_25_64_8855/U10  ( .A(\DP_OP_25_64_8855/n529 ), .B(
        \DP_OP_25_64_8855/n465 ), .Z(\C3/DATA5_60 ) );
  XOR \DP_OP_25_64_8855/U9  ( .A(\DP_OP_25_64_8855/n595 ), .B(
        \U1/RSOP_16/C2/Z_61 ), .Z(\DP_OP_25_64_8855/n464 ) );
  XOR \DP_OP_25_64_8855/U8  ( .A(\DP_OP_25_64_8855/n528 ), .B(
        \DP_OP_25_64_8855/n464 ), .Z(\C3/DATA5_61 ) );
  XOR \DP_OP_25_64_8855/U7  ( .A(\DP_OP_25_64_8855/n594 ), .B(
        \U1/RSOP_16/C2/Z_62 ), .Z(\DP_OP_25_64_8855/n463 ) );
  XOR \DP_OP_25_64_8855/U6  ( .A(\DP_OP_25_64_8855/n527 ), .B(
        \DP_OP_25_64_8855/n463 ), .Z(\C3/DATA5_62 ) );
  XOR \DP_OP_25_64_8855/U5  ( .A(\DP_OP_25_64_8855/n593 ), .B(
        \U1/RSOP_16/C2/Z_63 ), .Z(\DP_OP_25_64_8855/n462 ) );
  XOR \DP_OP_25_64_8855/U4  ( .A(\DP_OP_25_64_8855/n526 ), .B(
        \DP_OP_25_64_8855/n462 ), .Z(\C3/DATA5_63 ) );
  NAND \DP_OP_25_64_8855/U162  ( .A(\DP_OP_25_64_8855/n594 ), .B(
        \U1/RSOP_16/C2/Z_62 ), .Z(\DP_OP_25_64_8855/n5 ) );
  NAND \DP_OP_25_64_8855/U262  ( .A(\DP_OP_25_64_8855/n527 ), .B(
        \DP_OP_25_64_8855/n463 ), .Z(\DP_OP_25_64_8855/n8 ) );
  NAND \DP_OP_25_64_8855/U362  ( .A(\DP_OP_25_64_8855/n5 ), .B(
        \DP_OP_25_64_8855/n8 ), .Z(\DP_OP_25_64_8855/n526 ) );
  NAND \DP_OP_25_64_8855/U161  ( .A(\DP_OP_25_64_8855/n595 ), .B(
        \U1/RSOP_16/C2/Z_61 ), .Z(\DP_OP_25_64_8855/n14 ) );
  NAND \DP_OP_25_64_8855/U261  ( .A(\DP_OP_25_64_8855/n528 ), .B(
        \DP_OP_25_64_8855/n464 ), .Z(\DP_OP_25_64_8855/n15 ) );
  NAND \DP_OP_25_64_8855/U361  ( .A(\DP_OP_25_64_8855/n14 ), .B(
        \DP_OP_25_64_8855/n15 ), .Z(\DP_OP_25_64_8855/n527 ) );
  NAND \DP_OP_25_64_8855/U160  ( .A(\DP_OP_25_64_8855/n596 ), .B(
        \U1/RSOP_16/C2/Z_60 ), .Z(\DP_OP_25_64_8855/n21 ) );
  NAND \DP_OP_25_64_8855/U260  ( .A(\DP_OP_25_64_8855/n529 ), .B(
        \DP_OP_25_64_8855/n465 ), .Z(\DP_OP_25_64_8855/n22 ) );
  NAND \DP_OP_25_64_8855/U360  ( .A(\DP_OP_25_64_8855/n21 ), .B(
        \DP_OP_25_64_8855/n22 ), .Z(\DP_OP_25_64_8855/n528 ) );
  NAND \DP_OP_25_64_8855/U159  ( .A(\DP_OP_25_64_8855/n597 ), .B(
        \U1/RSOP_16/C2/Z_59 ), .Z(\DP_OP_25_64_8855/n28 ) );
  NAND \DP_OP_25_64_8855/U259  ( .A(\DP_OP_25_64_8855/n530 ), .B(
        \DP_OP_25_64_8855/n466 ), .Z(\DP_OP_25_64_8855/n29 ) );
  NAND \DP_OP_25_64_8855/U359  ( .A(\DP_OP_25_64_8855/n28 ), .B(
        \DP_OP_25_64_8855/n29 ), .Z(\DP_OP_25_64_8855/n529 ) );
  NAND \DP_OP_25_64_8855/U158  ( .A(\DP_OP_25_64_8855/n598 ), .B(
        \U1/RSOP_16/C2/Z_58 ), .Z(\DP_OP_25_64_8855/n35 ) );
  NAND \DP_OP_25_64_8855/U258  ( .A(\DP_OP_25_64_8855/n531 ), .B(
        \DP_OP_25_64_8855/n467 ), .Z(\DP_OP_25_64_8855/n36 ) );
  NAND \DP_OP_25_64_8855/U358  ( .A(\DP_OP_25_64_8855/n35 ), .B(
        \DP_OP_25_64_8855/n36 ), .Z(\DP_OP_25_64_8855/n530 ) );
  NAND \DP_OP_25_64_8855/U157  ( .A(\DP_OP_25_64_8855/n599 ), .B(
        \U1/RSOP_16/C2/Z_57 ), .Z(\DP_OP_25_64_8855/n42 ) );
  NAND \DP_OP_25_64_8855/U257  ( .A(\DP_OP_25_64_8855/n532 ), .B(
        \DP_OP_25_64_8855/n468 ), .Z(\DP_OP_25_64_8855/n43 ) );
  NAND \DP_OP_25_64_8855/U357  ( .A(\DP_OP_25_64_8855/n42 ), .B(
        \DP_OP_25_64_8855/n43 ), .Z(\DP_OP_25_64_8855/n531 ) );
  NAND \DP_OP_25_64_8855/U156  ( .A(\DP_OP_25_64_8855/n600 ), .B(
        \U1/RSOP_16/C2/Z_56 ), .Z(\DP_OP_25_64_8855/n49 ) );
  NAND \DP_OP_25_64_8855/U256  ( .A(\DP_OP_25_64_8855/n533 ), .B(
        \DP_OP_25_64_8855/n469 ), .Z(\DP_OP_25_64_8855/n50 ) );
  NAND \DP_OP_25_64_8855/U356  ( .A(\DP_OP_25_64_8855/n49 ), .B(
        \DP_OP_25_64_8855/n50 ), .Z(\DP_OP_25_64_8855/n532 ) );
  NAND \DP_OP_25_64_8855/U155  ( .A(\DP_OP_25_64_8855/n601 ), .B(
        \U1/RSOP_16/C2/Z_55 ), .Z(\DP_OP_25_64_8855/n56 ) );
  NAND \DP_OP_25_64_8855/U255  ( .A(\DP_OP_25_64_8855/n534 ), .B(
        \DP_OP_25_64_8855/n470 ), .Z(\DP_OP_25_64_8855/n57 ) );
  NAND \DP_OP_25_64_8855/U355  ( .A(\DP_OP_25_64_8855/n56 ), .B(
        \DP_OP_25_64_8855/n57 ), .Z(\DP_OP_25_64_8855/n533 ) );
  NAND \DP_OP_25_64_8855/U154  ( .A(\DP_OP_25_64_8855/n602 ), .B(
        \U1/RSOP_16/C2/Z_54 ), .Z(\DP_OP_25_64_8855/n81 ) );
  NAND \DP_OP_25_64_8855/U254  ( .A(\DP_OP_25_64_8855/n535 ), .B(
        \DP_OP_25_64_8855/n471 ), .Z(\DP_OP_25_64_8855/n82 ) );
  NAND \DP_OP_25_64_8855/U354  ( .A(\DP_OP_25_64_8855/n81 ), .B(
        \DP_OP_25_64_8855/n82 ), .Z(\DP_OP_25_64_8855/n534 ) );
  NAND \DP_OP_25_64_8855/U153  ( .A(\DP_OP_25_64_8855/n603 ), .B(
        \U1/RSOP_16/C2/Z_53 ), .Z(\DP_OP_25_64_8855/n88 ) );
  NAND \DP_OP_25_64_8855/U253  ( .A(\DP_OP_25_64_8855/n536 ), .B(
        \DP_OP_25_64_8855/n472 ), .Z(\DP_OP_25_64_8855/n89 ) );
  NAND \DP_OP_25_64_8855/U353  ( .A(\DP_OP_25_64_8855/n88 ), .B(
        \DP_OP_25_64_8855/n89 ), .Z(\DP_OP_25_64_8855/n535 ) );
  NAND \DP_OP_25_64_8855/U152  ( .A(\DP_OP_25_64_8855/n604 ), .B(
        \U1/RSOP_16/C2/Z_52 ), .Z(\DP_OP_25_64_8855/n95 ) );
  NAND \DP_OP_25_64_8855/U252  ( .A(\DP_OP_25_64_8855/n537 ), .B(
        \DP_OP_25_64_8855/n473 ), .Z(\DP_OP_25_64_8855/n96 ) );
  NAND \DP_OP_25_64_8855/U352  ( .A(\DP_OP_25_64_8855/n95 ), .B(
        \DP_OP_25_64_8855/n96 ), .Z(\DP_OP_25_64_8855/n536 ) );
  NAND \DP_OP_25_64_8855/U151  ( .A(\DP_OP_25_64_8855/n605 ), .B(
        \U1/RSOP_16/C2/Z_51 ), .Z(\DP_OP_25_64_8855/n102 ) );
  NAND \DP_OP_25_64_8855/U251  ( .A(\DP_OP_25_64_8855/n538 ), .B(
        \DP_OP_25_64_8855/n474 ), .Z(\DP_OP_25_64_8855/n103 ) );
  NAND \DP_OP_25_64_8855/U351  ( .A(\DP_OP_25_64_8855/n102 ), .B(
        \DP_OP_25_64_8855/n103 ), .Z(\DP_OP_25_64_8855/n537 ) );
  NAND \DP_OP_25_64_8855/U150  ( .A(\DP_OP_25_64_8855/n606 ), .B(
        \U1/RSOP_16/C2/Z_50 ), .Z(\DP_OP_25_64_8855/n109 ) );
  NAND \DP_OP_25_64_8855/U250  ( .A(\DP_OP_25_64_8855/n539 ), .B(
        \DP_OP_25_64_8855/n475 ), .Z(\DP_OP_25_64_8855/n110 ) );
  NAND \DP_OP_25_64_8855/U350  ( .A(\DP_OP_25_64_8855/n109 ), .B(
        \DP_OP_25_64_8855/n110 ), .Z(\DP_OP_25_64_8855/n538 ) );
  NAND \DP_OP_25_64_8855/U149  ( .A(\DP_OP_25_64_8855/n607 ), .B(
        \U1/RSOP_16/C2/Z_49 ), .Z(\DP_OP_25_64_8855/n116 ) );
  NAND \DP_OP_25_64_8855/U249  ( .A(\DP_OP_25_64_8855/n540 ), .B(
        \DP_OP_25_64_8855/n476 ), .Z(\DP_OP_25_64_8855/n117 ) );
  NAND \DP_OP_25_64_8855/U349  ( .A(\DP_OP_25_64_8855/n116 ), .B(
        \DP_OP_25_64_8855/n117 ), .Z(\DP_OP_25_64_8855/n539 ) );
  NAND \DP_OP_25_64_8855/U148  ( .A(\DP_OP_25_64_8855/n608 ), .B(
        \U1/RSOP_16/C2/Z_48 ), .Z(\DP_OP_25_64_8855/n123 ) );
  NAND \DP_OP_25_64_8855/U248  ( .A(\DP_OP_25_64_8855/n541 ), .B(
        \DP_OP_25_64_8855/n477 ), .Z(\DP_OP_25_64_8855/n124 ) );
  NAND \DP_OP_25_64_8855/U348  ( .A(\DP_OP_25_64_8855/n123 ), .B(
        \DP_OP_25_64_8855/n124 ), .Z(\DP_OP_25_64_8855/n540 ) );
  NAND \DP_OP_25_64_8855/U147  ( .A(\DP_OP_25_64_8855/n609 ), .B(
        \U1/RSOP_16/C2/Z_47 ), .Z(\DP_OP_25_64_8855/n130 ) );
  NAND \DP_OP_25_64_8855/U247  ( .A(\DP_OP_25_64_8855/n542 ), .B(
        \DP_OP_25_64_8855/n478 ), .Z(\DP_OP_25_64_8855/n131 ) );
  NAND \DP_OP_25_64_8855/U347  ( .A(\DP_OP_25_64_8855/n130 ), .B(
        \DP_OP_25_64_8855/n131 ), .Z(\DP_OP_25_64_8855/n541 ) );
  NAND \DP_OP_25_64_8855/U146  ( .A(\DP_OP_25_64_8855/n610 ), .B(
        \U1/RSOP_16/C2/Z_46 ), .Z(\DP_OP_25_64_8855/n137 ) );
  NAND \DP_OP_25_64_8855/U246  ( .A(\DP_OP_25_64_8855/n543 ), .B(
        \DP_OP_25_64_8855/n479 ), .Z(\DP_OP_25_64_8855/n138 ) );
  NAND \DP_OP_25_64_8855/U346  ( .A(\DP_OP_25_64_8855/n137 ), .B(
        \DP_OP_25_64_8855/n138 ), .Z(\DP_OP_25_64_8855/n542 ) );
  NAND \DP_OP_25_64_8855/U145  ( .A(\DP_OP_25_64_8855/n611 ), .B(
        \U1/RSOP_16/C2/Z_45 ), .Z(\DP_OP_25_64_8855/n144 ) );
  NAND \DP_OP_25_64_8855/U245  ( .A(\DP_OP_25_64_8855/n544 ), .B(
        \DP_OP_25_64_8855/n480 ), .Z(\DP_OP_25_64_8855/n145 ) );
  NAND \DP_OP_25_64_8855/U345  ( .A(\DP_OP_25_64_8855/n144 ), .B(
        \DP_OP_25_64_8855/n145 ), .Z(\DP_OP_25_64_8855/n543 ) );
  NAND \DP_OP_25_64_8855/U144  ( .A(\DP_OP_25_64_8855/n612 ), .B(
        \U1/RSOP_16/C2/Z_44 ), .Z(\DP_OP_25_64_8855/n151 ) );
  NAND \DP_OP_25_64_8855/U244  ( .A(\DP_OP_25_64_8855/n545 ), .B(
        \DP_OP_25_64_8855/n481 ), .Z(\DP_OP_25_64_8855/n152 ) );
  NAND \DP_OP_25_64_8855/U344  ( .A(\DP_OP_25_64_8855/n151 ), .B(
        \DP_OP_25_64_8855/n152 ), .Z(\DP_OP_25_64_8855/n544 ) );
  NAND \DP_OP_25_64_8855/U143  ( .A(\DP_OP_25_64_8855/n613 ), .B(
        \U1/RSOP_16/C2/Z_43 ), .Z(\DP_OP_25_64_8855/n158 ) );
  NAND \DP_OP_25_64_8855/U243  ( .A(\DP_OP_25_64_8855/n546 ), .B(
        \DP_OP_25_64_8855/n482 ), .Z(\DP_OP_25_64_8855/n159 ) );
  NAND \DP_OP_25_64_8855/U343  ( .A(\DP_OP_25_64_8855/n158 ), .B(
        \DP_OP_25_64_8855/n159 ), .Z(\DP_OP_25_64_8855/n545 ) );
  NAND \DP_OP_25_64_8855/U142  ( .A(\DP_OP_25_64_8855/n614 ), .B(
        \U1/RSOP_16/C2/Z_42 ), .Z(\DP_OP_25_64_8855/n165 ) );
  NAND \DP_OP_25_64_8855/U242  ( .A(\DP_OP_25_64_8855/n547 ), .B(
        \DP_OP_25_64_8855/n483 ), .Z(\DP_OP_25_64_8855/n166 ) );
  NAND \DP_OP_25_64_8855/U342  ( .A(\DP_OP_25_64_8855/n165 ), .B(
        \DP_OP_25_64_8855/n166 ), .Z(\DP_OP_25_64_8855/n546 ) );
  NAND \DP_OP_25_64_8855/U141  ( .A(\DP_OP_25_64_8855/n615 ), .B(
        \U1/RSOP_16/C2/Z_41 ), .Z(\DP_OP_25_64_8855/n172 ) );
  NAND \DP_OP_25_64_8855/U241  ( .A(\DP_OP_25_64_8855/n548 ), .B(
        \DP_OP_25_64_8855/n484 ), .Z(\DP_OP_25_64_8855/n173 ) );
  NAND \DP_OP_25_64_8855/U341  ( .A(\DP_OP_25_64_8855/n172 ), .B(
        \DP_OP_25_64_8855/n173 ), .Z(\DP_OP_25_64_8855/n547 ) );
  NAND \DP_OP_25_64_8855/U140  ( .A(\DP_OP_25_64_8855/n616 ), .B(
        \U1/RSOP_16/C2/Z_40 ), .Z(\DP_OP_25_64_8855/n179 ) );
  NAND \DP_OP_25_64_8855/U240  ( .A(\DP_OP_25_64_8855/n549 ), .B(
        \DP_OP_25_64_8855/n485 ), .Z(\DP_OP_25_64_8855/n180 ) );
  NAND \DP_OP_25_64_8855/U340  ( .A(\DP_OP_25_64_8855/n179 ), .B(
        \DP_OP_25_64_8855/n180 ), .Z(\DP_OP_25_64_8855/n548 ) );
  NAND \DP_OP_25_64_8855/U139  ( .A(\DP_OP_25_64_8855/n617 ), .B(
        \U1/RSOP_16/C2/Z_39 ), .Z(\DP_OP_25_64_8855/n186 ) );
  NAND \DP_OP_25_64_8855/U239  ( .A(\DP_OP_25_64_8855/n550 ), .B(
        \DP_OP_25_64_8855/n486 ), .Z(\DP_OP_25_64_8855/n187 ) );
  NAND \DP_OP_25_64_8855/U339  ( .A(\DP_OP_25_64_8855/n186 ), .B(
        \DP_OP_25_64_8855/n187 ), .Z(\DP_OP_25_64_8855/n549 ) );
  NAND \DP_OP_25_64_8855/U138  ( .A(\DP_OP_25_64_8855/n618 ), .B(
        \U1/RSOP_16/C2/Z_38 ), .Z(\DP_OP_25_64_8855/n193 ) );
  NAND \DP_OP_25_64_8855/U238  ( .A(\DP_OP_25_64_8855/n551 ), .B(
        \DP_OP_25_64_8855/n487 ), .Z(\DP_OP_25_64_8855/n194 ) );
  NAND \DP_OP_25_64_8855/U338  ( .A(\DP_OP_25_64_8855/n193 ), .B(
        \DP_OP_25_64_8855/n194 ), .Z(\DP_OP_25_64_8855/n550 ) );
  NAND \DP_OP_25_64_8855/U137  ( .A(\DP_OP_25_64_8855/n619 ), .B(
        \U1/RSOP_16/C2/Z_37 ), .Z(\DP_OP_25_64_8855/n200 ) );
  NAND \DP_OP_25_64_8855/U237  ( .A(\DP_OP_25_64_8855/n552 ), .B(
        \DP_OP_25_64_8855/n488 ), .Z(\DP_OP_25_64_8855/n201 ) );
  NAND \DP_OP_25_64_8855/U337  ( .A(\DP_OP_25_64_8855/n200 ), .B(
        \DP_OP_25_64_8855/n201 ), .Z(\DP_OP_25_64_8855/n551 ) );
  NAND \DP_OP_25_64_8855/U136  ( .A(\DP_OP_25_64_8855/n620 ), .B(
        \U1/RSOP_16/C2/Z_36 ), .Z(\DP_OP_25_64_8855/n207 ) );
  NAND \DP_OP_25_64_8855/U236  ( .A(\DP_OP_25_64_8855/n553 ), .B(
        \DP_OP_25_64_8855/n489 ), .Z(\DP_OP_25_64_8855/n208 ) );
  NAND \DP_OP_25_64_8855/U336  ( .A(\DP_OP_25_64_8855/n207 ), .B(
        \DP_OP_25_64_8855/n208 ), .Z(\DP_OP_25_64_8855/n552 ) );
  NAND \DP_OP_25_64_8855/U135  ( .A(\DP_OP_25_64_8855/n621 ), .B(
        \U1/RSOP_16/C2/Z_35 ), .Z(\DP_OP_25_64_8855/n214 ) );
  NAND \DP_OP_25_64_8855/U235  ( .A(\DP_OP_25_64_8855/n554 ), .B(
        \DP_OP_25_64_8855/n490 ), .Z(\DP_OP_25_64_8855/n215 ) );
  NAND \DP_OP_25_64_8855/U335  ( .A(\DP_OP_25_64_8855/n214 ), .B(
        \DP_OP_25_64_8855/n215 ), .Z(\DP_OP_25_64_8855/n553 ) );
  NAND \DP_OP_25_64_8855/U134  ( .A(\DP_OP_25_64_8855/n622 ), .B(
        \U1/RSOP_16/C2/Z_34 ), .Z(\DP_OP_25_64_8855/n221 ) );
  NAND \DP_OP_25_64_8855/U234  ( .A(\DP_OP_25_64_8855/n555 ), .B(
        \DP_OP_25_64_8855/n491 ), .Z(\DP_OP_25_64_8855/n222 ) );
  NAND \DP_OP_25_64_8855/U334  ( .A(\DP_OP_25_64_8855/n221 ), .B(
        \DP_OP_25_64_8855/n222 ), .Z(\DP_OP_25_64_8855/n554 ) );
  NAND \DP_OP_25_64_8855/U133  ( .A(\DP_OP_25_64_8855/n623 ), .B(
        \U1/RSOP_16/C2/Z_33 ), .Z(\DP_OP_25_64_8855/n228 ) );
  NAND \DP_OP_25_64_8855/U233  ( .A(\DP_OP_25_64_8855/n556 ), .B(
        \DP_OP_25_64_8855/n492 ), .Z(\DP_OP_25_64_8855/n229 ) );
  NAND \DP_OP_25_64_8855/U333  ( .A(\DP_OP_25_64_8855/n228 ), .B(
        \DP_OP_25_64_8855/n229 ), .Z(\DP_OP_25_64_8855/n555 ) );
  NAND \DP_OP_25_64_8855/U132  ( .A(\DP_OP_25_64_8855/n624 ), .B(
        \U1/RSOP_16/C2/Z_32 ), .Z(\DP_OP_25_64_8855/n235 ) );
  NAND \DP_OP_25_64_8855/U232  ( .A(\DP_OP_25_64_8855/n557 ), .B(
        \DP_OP_25_64_8855/n493 ), .Z(\DP_OP_25_64_8855/n236 ) );
  NAND \DP_OP_25_64_8855/U332  ( .A(\DP_OP_25_64_8855/n235 ), .B(
        \DP_OP_25_64_8855/n236 ), .Z(\DP_OP_25_64_8855/n556 ) );
  NAND \DP_OP_25_64_8855/U131  ( .A(\DP_OP_25_64_8855/n625 ), .B(
        \U1/RSOP_16/C2/Z_31 ), .Z(\DP_OP_25_64_8855/n242 ) );
  NAND \DP_OP_25_64_8855/U231  ( .A(\DP_OP_25_64_8855/n558 ), .B(
        \DP_OP_25_64_8855/n494 ), .Z(\DP_OP_25_64_8855/n243 ) );
  NAND \DP_OP_25_64_8855/U331  ( .A(\DP_OP_25_64_8855/n242 ), .B(
        \DP_OP_25_64_8855/n243 ), .Z(\DP_OP_25_64_8855/n557 ) );
  NAND \DP_OP_25_64_8855/U130  ( .A(\DP_OP_25_64_8855/n626 ), .B(
        \U1/RSOP_16/C2/Z_30 ), .Z(\DP_OP_25_64_8855/n249 ) );
  NAND \DP_OP_25_64_8855/U230  ( .A(\DP_OP_25_64_8855/n559 ), .B(
        \DP_OP_25_64_8855/n495 ), .Z(\DP_OP_25_64_8855/n250 ) );
  NAND \DP_OP_25_64_8855/U330  ( .A(\DP_OP_25_64_8855/n249 ), .B(
        \DP_OP_25_64_8855/n250 ), .Z(\DP_OP_25_64_8855/n558 ) );
  NAND \DP_OP_25_64_8855/U129  ( .A(\DP_OP_25_64_8855/n627 ), .B(
        \U1/RSOP_16/C2/Z_29 ), .Z(\DP_OP_25_64_8855/n256 ) );
  NAND \DP_OP_25_64_8855/U229  ( .A(\DP_OP_25_64_8855/n560 ), .B(
        \DP_OP_25_64_8855/n496 ), .Z(\DP_OP_25_64_8855/n257 ) );
  NAND \DP_OP_25_64_8855/U329  ( .A(\DP_OP_25_64_8855/n256 ), .B(
        \DP_OP_25_64_8855/n257 ), .Z(\DP_OP_25_64_8855/n559 ) );
  NAND \DP_OP_25_64_8855/U128  ( .A(\DP_OP_25_64_8855/n628 ), .B(
        \U1/RSOP_16/C2/Z_28 ), .Z(\DP_OP_25_64_8855/n263 ) );
  NAND \DP_OP_25_64_8855/U228  ( .A(\DP_OP_25_64_8855/n561 ), .B(
        \DP_OP_25_64_8855/n497 ), .Z(\DP_OP_25_64_8855/n264 ) );
  NAND \DP_OP_25_64_8855/U328  ( .A(\DP_OP_25_64_8855/n263 ), .B(
        \DP_OP_25_64_8855/n264 ), .Z(\DP_OP_25_64_8855/n560 ) );
  NAND \DP_OP_25_64_8855/U127  ( .A(\DP_OP_25_64_8855/n629 ), .B(
        \U1/RSOP_16/C2/Z_27 ), .Z(\DP_OP_25_64_8855/n270 ) );
  NAND \DP_OP_25_64_8855/U227  ( .A(\DP_OP_25_64_8855/n562 ), .B(
        \DP_OP_25_64_8855/n498 ), .Z(\DP_OP_25_64_8855/n271 ) );
  NAND \DP_OP_25_64_8855/U327  ( .A(\DP_OP_25_64_8855/n270 ), .B(
        \DP_OP_25_64_8855/n271 ), .Z(\DP_OP_25_64_8855/n561 ) );
  NAND \DP_OP_25_64_8855/U126  ( .A(\DP_OP_25_64_8855/n630 ), .B(
        \U1/RSOP_16/C2/Z_26 ), .Z(\DP_OP_25_64_8855/n277 ) );
  NAND \DP_OP_25_64_8855/U226  ( .A(\DP_OP_25_64_8855/n563 ), .B(
        \DP_OP_25_64_8855/n499 ), .Z(\DP_OP_25_64_8855/n278 ) );
  NAND \DP_OP_25_64_8855/U326  ( .A(\DP_OP_25_64_8855/n277 ), .B(
        \DP_OP_25_64_8855/n278 ), .Z(\DP_OP_25_64_8855/n562 ) );
  NAND \DP_OP_25_64_8855/U125  ( .A(\DP_OP_25_64_8855/n631 ), .B(
        \U1/RSOP_16/C2/Z_25 ), .Z(\DP_OP_25_64_8855/n284 ) );
  NAND \DP_OP_25_64_8855/U225  ( .A(\DP_OP_25_64_8855/n564 ), .B(
        \DP_OP_25_64_8855/n500 ), .Z(\DP_OP_25_64_8855/n285 ) );
  NAND \DP_OP_25_64_8855/U325  ( .A(\DP_OP_25_64_8855/n284 ), .B(
        \DP_OP_25_64_8855/n285 ), .Z(\DP_OP_25_64_8855/n563 ) );
  NAND \DP_OP_25_64_8855/U124  ( .A(\DP_OP_25_64_8855/n632 ), .B(
        \U1/RSOP_16/C2/Z_24 ), .Z(\DP_OP_25_64_8855/n291 ) );
  NAND \DP_OP_25_64_8855/U224  ( .A(\DP_OP_25_64_8855/n565 ), .B(
        \DP_OP_25_64_8855/n501 ), .Z(\DP_OP_25_64_8855/n292 ) );
  NAND \DP_OP_25_64_8855/U324  ( .A(\DP_OP_25_64_8855/n291 ), .B(
        \DP_OP_25_64_8855/n292 ), .Z(\DP_OP_25_64_8855/n564 ) );
  NAND \DP_OP_25_64_8855/U123  ( .A(\DP_OP_25_64_8855/n633 ), .B(
        \U1/RSOP_16/C2/Z_23 ), .Z(\DP_OP_25_64_8855/n298 ) );
  NAND \DP_OP_25_64_8855/U223  ( .A(\DP_OP_25_64_8855/n566 ), .B(
        \DP_OP_25_64_8855/n502 ), .Z(\DP_OP_25_64_8855/n299 ) );
  NAND \DP_OP_25_64_8855/U323  ( .A(\DP_OP_25_64_8855/n298 ), .B(
        \DP_OP_25_64_8855/n299 ), .Z(\DP_OP_25_64_8855/n565 ) );
  NAND \DP_OP_25_64_8855/U122  ( .A(\DP_OP_25_64_8855/n634 ), .B(
        \U1/RSOP_16/C2/Z_22 ), .Z(\DP_OP_25_64_8855/n305 ) );
  NAND \DP_OP_25_64_8855/U222  ( .A(\DP_OP_25_64_8855/n567 ), .B(
        \DP_OP_25_64_8855/n503 ), .Z(\DP_OP_25_64_8855/n306 ) );
  NAND \DP_OP_25_64_8855/U322  ( .A(\DP_OP_25_64_8855/n305 ), .B(
        \DP_OP_25_64_8855/n306 ), .Z(\DP_OP_25_64_8855/n566 ) );
  NAND \DP_OP_25_64_8855/U121  ( .A(\DP_OP_25_64_8855/n635 ), .B(
        \U1/RSOP_16/C2/Z_21 ), .Z(\DP_OP_25_64_8855/n312 ) );
  NAND \DP_OP_25_64_8855/U221  ( .A(\DP_OP_25_64_8855/n568 ), .B(
        \DP_OP_25_64_8855/n504 ), .Z(\DP_OP_25_64_8855/n313 ) );
  NAND \DP_OP_25_64_8855/U321  ( .A(\DP_OP_25_64_8855/n312 ), .B(
        \DP_OP_25_64_8855/n313 ), .Z(\DP_OP_25_64_8855/n567 ) );
  NAND \DP_OP_25_64_8855/U120  ( .A(\DP_OP_25_64_8855/n636 ), .B(
        \U1/RSOP_16/C2/Z_20 ), .Z(\DP_OP_25_64_8855/n319 ) );
  NAND \DP_OP_25_64_8855/U220  ( .A(\DP_OP_25_64_8855/n569 ), .B(
        \DP_OP_25_64_8855/n505 ), .Z(\DP_OP_25_64_8855/n320 ) );
  NAND \DP_OP_25_64_8855/U320  ( .A(\DP_OP_25_64_8855/n319 ), .B(
        \DP_OP_25_64_8855/n320 ), .Z(\DP_OP_25_64_8855/n568 ) );
  NAND \DP_OP_25_64_8855/U119  ( .A(\DP_OP_25_64_8855/n637 ), .B(
        \U1/RSOP_16/C2/Z_19 ), .Z(\DP_OP_25_64_8855/n326 ) );
  NAND \DP_OP_25_64_8855/U219  ( .A(\DP_OP_25_64_8855/n570 ), .B(
        \DP_OP_25_64_8855/n506 ), .Z(\DP_OP_25_64_8855/n327 ) );
  NAND \DP_OP_25_64_8855/U319  ( .A(\DP_OP_25_64_8855/n326 ), .B(
        \DP_OP_25_64_8855/n327 ), .Z(\DP_OP_25_64_8855/n569 ) );
  NAND \DP_OP_25_64_8855/U118  ( .A(\DP_OP_25_64_8855/n638 ), .B(
        \U1/RSOP_16/C2/Z_18 ), .Z(\DP_OP_25_64_8855/n333 ) );
  NAND \DP_OP_25_64_8855/U218  ( .A(\DP_OP_25_64_8855/n571 ), .B(
        \DP_OP_25_64_8855/n507 ), .Z(\DP_OP_25_64_8855/n334 ) );
  NAND \DP_OP_25_64_8855/U318  ( .A(\DP_OP_25_64_8855/n333 ), .B(
        \DP_OP_25_64_8855/n334 ), .Z(\DP_OP_25_64_8855/n570 ) );
  NAND \DP_OP_25_64_8855/U117  ( .A(\DP_OP_25_64_8855/n639 ), .B(
        \U1/RSOP_16/C2/Z_17 ), .Z(\DP_OP_25_64_8855/n340 ) );
  NAND \DP_OP_25_64_8855/U217  ( .A(\DP_OP_25_64_8855/n572 ), .B(
        \DP_OP_25_64_8855/n508 ), .Z(\DP_OP_25_64_8855/n341 ) );
  NAND \DP_OP_25_64_8855/U317  ( .A(\DP_OP_25_64_8855/n340 ), .B(
        \DP_OP_25_64_8855/n341 ), .Z(\DP_OP_25_64_8855/n571 ) );
  NAND \DP_OP_25_64_8855/U116  ( .A(\DP_OP_25_64_8855/n640 ), .B(
        \U1/RSOP_16/C2/Z_16 ), .Z(\DP_OP_25_64_8855/n347 ) );
  NAND \DP_OP_25_64_8855/U216  ( .A(\DP_OP_25_64_8855/n573 ), .B(
        \DP_OP_25_64_8855/n509 ), .Z(\DP_OP_25_64_8855/n348 ) );
  NAND \DP_OP_25_64_8855/U316  ( .A(\DP_OP_25_64_8855/n347 ), .B(
        \DP_OP_25_64_8855/n348 ), .Z(\DP_OP_25_64_8855/n572 ) );
  NAND \DP_OP_25_64_8855/U115  ( .A(\DP_OP_25_64_8855/n641 ), .B(
        \U1/RSOP_16/C2/Z_15 ), .Z(\DP_OP_25_64_8855/n354 ) );
  NAND \DP_OP_25_64_8855/U215  ( .A(\DP_OP_25_64_8855/n574 ), .B(
        \DP_OP_25_64_8855/n510 ), .Z(\DP_OP_25_64_8855/n355 ) );
  NAND \DP_OP_25_64_8855/U315  ( .A(\DP_OP_25_64_8855/n354 ), .B(
        \DP_OP_25_64_8855/n355 ), .Z(\DP_OP_25_64_8855/n573 ) );
  NAND \DP_OP_25_64_8855/U114  ( .A(\DP_OP_25_64_8855/n642 ), .B(
        \U1/RSOP_16/C2/Z_14 ), .Z(\DP_OP_25_64_8855/n361 ) );
  NAND \DP_OP_25_64_8855/U214  ( .A(\DP_OP_25_64_8855/n575 ), .B(
        \DP_OP_25_64_8855/n511 ), .Z(\DP_OP_25_64_8855/n362 ) );
  NAND \DP_OP_25_64_8855/U314  ( .A(\DP_OP_25_64_8855/n361 ), .B(
        \DP_OP_25_64_8855/n362 ), .Z(\DP_OP_25_64_8855/n574 ) );
  NAND \DP_OP_25_64_8855/U113  ( .A(\DP_OP_25_64_8855/n643 ), .B(
        \U1/RSOP_16/C2/Z_13 ), .Z(\DP_OP_25_64_8855/n368 ) );
  NAND \DP_OP_25_64_8855/U213  ( .A(\DP_OP_25_64_8855/n576 ), .B(
        \DP_OP_25_64_8855/n512 ), .Z(\DP_OP_25_64_8855/n369 ) );
  NAND \DP_OP_25_64_8855/U313  ( .A(\DP_OP_25_64_8855/n368 ), .B(
        \DP_OP_25_64_8855/n369 ), .Z(\DP_OP_25_64_8855/n575 ) );
  NAND \DP_OP_25_64_8855/U112  ( .A(\DP_OP_25_64_8855/n644 ), .B(
        \U1/RSOP_16/C2/Z_12 ), .Z(\DP_OP_25_64_8855/n375 ) );
  NAND \DP_OP_25_64_8855/U212  ( .A(\DP_OP_25_64_8855/n577 ), .B(
        \DP_OP_25_64_8855/n513 ), .Z(\DP_OP_25_64_8855/n376 ) );
  NAND \DP_OP_25_64_8855/U312  ( .A(\DP_OP_25_64_8855/n375 ), .B(
        \DP_OP_25_64_8855/n376 ), .Z(\DP_OP_25_64_8855/n576 ) );
  NAND \DP_OP_25_64_8855/U111  ( .A(\DP_OP_25_64_8855/n645 ), .B(
        \U1/RSOP_16/C2/Z_11 ), .Z(\DP_OP_25_64_8855/n382 ) );
  NAND \DP_OP_25_64_8855/U211  ( .A(\DP_OP_25_64_8855/n578 ), .B(
        \DP_OP_25_64_8855/n514 ), .Z(\DP_OP_25_64_8855/n383 ) );
  NAND \DP_OP_25_64_8855/U311  ( .A(\DP_OP_25_64_8855/n382 ), .B(
        \DP_OP_25_64_8855/n383 ), .Z(\DP_OP_25_64_8855/n577 ) );
  NAND \DP_OP_25_64_8855/U110  ( .A(\DP_OP_25_64_8855/n646 ), .B(
        \U1/RSOP_16/C2/Z_10 ), .Z(\DP_OP_25_64_8855/n389 ) );
  NAND \DP_OP_25_64_8855/U210  ( .A(\DP_OP_25_64_8855/n579 ), .B(
        \DP_OP_25_64_8855/n515 ), .Z(\DP_OP_25_64_8855/n390 ) );
  NAND \DP_OP_25_64_8855/U310  ( .A(\DP_OP_25_64_8855/n389 ), .B(
        \DP_OP_25_64_8855/n390 ), .Z(\DP_OP_25_64_8855/n578 ) );
  NAND \DP_OP_25_64_8855/U19  ( .A(\DP_OP_25_64_8855/n647 ), .B(
        \U1/RSOP_16/C2/Z_9 ), .Z(\DP_OP_25_64_8855/n396 ) );
  NAND \DP_OP_25_64_8855/U29  ( .A(\DP_OP_25_64_8855/n580 ), .B(
        \DP_OP_25_64_8855/n516 ), .Z(\DP_OP_25_64_8855/n397 ) );
  NAND \DP_OP_25_64_8855/U39  ( .A(\DP_OP_25_64_8855/n396 ), .B(
        \DP_OP_25_64_8855/n397 ), .Z(\DP_OP_25_64_8855/n579 ) );
  NAND \DP_OP_25_64_8855/U18  ( .A(\DP_OP_25_64_8855/n648 ), .B(
        \U1/RSOP_16/C2/Z_8 ), .Z(\DP_OP_25_64_8855/n403 ) );
  NAND \DP_OP_25_64_8855/U28  ( .A(\DP_OP_25_64_8855/n581 ), .B(
        \DP_OP_25_64_8855/n517 ), .Z(\DP_OP_25_64_8855/n404 ) );
  NAND \DP_OP_25_64_8855/U38  ( .A(\DP_OP_25_64_8855/n403 ), .B(
        \DP_OP_25_64_8855/n404 ), .Z(\DP_OP_25_64_8855/n580 ) );
  NAND \DP_OP_25_64_8855/U17  ( .A(\DP_OP_25_64_8855/n649 ), .B(
        \U1/RSOP_16/C2/Z_7 ), .Z(\DP_OP_25_64_8855/n410 ) );
  NAND \DP_OP_25_64_8855/U27  ( .A(\DP_OP_25_64_8855/n582 ), .B(
        \DP_OP_25_64_8855/n518 ), .Z(\DP_OP_25_64_8855/n411 ) );
  NAND \DP_OP_25_64_8855/U37  ( .A(\DP_OP_25_64_8855/n410 ), .B(
        \DP_OP_25_64_8855/n411 ), .Z(\DP_OP_25_64_8855/n581 ) );
  NAND \DP_OP_25_64_8855/U16  ( .A(\DP_OP_25_64_8855/n650 ), .B(
        \U1/RSOP_16/C2/Z_6 ), .Z(\DP_OP_25_64_8855/n417 ) );
  NAND \DP_OP_25_64_8855/U26  ( .A(\DP_OP_25_64_8855/n583 ), .B(
        \DP_OP_25_64_8855/n519 ), .Z(\DP_OP_25_64_8855/n418 ) );
  NAND \DP_OP_25_64_8855/U36  ( .A(\DP_OP_25_64_8855/n417 ), .B(
        \DP_OP_25_64_8855/n418 ), .Z(\DP_OP_25_64_8855/n582 ) );
  NAND \DP_OP_25_64_8855/U15  ( .A(\DP_OP_25_64_8855/n651 ), .B(
        \U1/RSOP_16/C2/Z_5 ), .Z(\DP_OP_25_64_8855/n424 ) );
  NAND \DP_OP_25_64_8855/U25  ( .A(\DP_OP_25_64_8855/n584 ), .B(
        \DP_OP_25_64_8855/n520 ), .Z(\DP_OP_25_64_8855/n425 ) );
  NAND \DP_OP_25_64_8855/U35  ( .A(\DP_OP_25_64_8855/n424 ), .B(
        \DP_OP_25_64_8855/n425 ), .Z(\DP_OP_25_64_8855/n583 ) );
  NAND \DP_OP_25_64_8855/U14  ( .A(\DP_OP_25_64_8855/n652 ), .B(
        \U1/RSOP_16/C2/Z_4 ), .Z(\DP_OP_25_64_8855/n431 ) );
  NAND \DP_OP_25_64_8855/U24  ( .A(\DP_OP_25_64_8855/n585 ), .B(
        \DP_OP_25_64_8855/n521 ), .Z(\DP_OP_25_64_8855/n432 ) );
  NAND \DP_OP_25_64_8855/U34  ( .A(\DP_OP_25_64_8855/n431 ), .B(
        \DP_OP_25_64_8855/n432 ), .Z(\DP_OP_25_64_8855/n584 ) );
  NAND \DP_OP_25_64_8855/U13  ( .A(\DP_OP_25_64_8855/n653 ), .B(
        \U1/RSOP_16/C2/Z_3 ), .Z(\DP_OP_25_64_8855/n438 ) );
  NAND \DP_OP_25_64_8855/U23  ( .A(\DP_OP_25_64_8855/n586 ), .B(
        \DP_OP_25_64_8855/n522 ), .Z(\DP_OP_25_64_8855/n439 ) );
  NAND \DP_OP_25_64_8855/U33  ( .A(\DP_OP_25_64_8855/n438 ), .B(
        \DP_OP_25_64_8855/n439 ), .Z(\DP_OP_25_64_8855/n585 ) );
  NAND \DP_OP_25_64_8855/U12  ( .A(\DP_OP_25_64_8855/n654 ), .B(
        \U1/RSOP_16/C2/Z_2 ), .Z(\DP_OP_25_64_8855/n445 ) );
  NAND \DP_OP_25_64_8855/U22  ( .A(\DP_OP_25_64_8855/n587 ), .B(
        \DP_OP_25_64_8855/n523 ), .Z(\DP_OP_25_64_8855/n446 ) );
  NAND \DP_OP_25_64_8855/U32  ( .A(\DP_OP_25_64_8855/n445 ), .B(
        \DP_OP_25_64_8855/n446 ), .Z(\DP_OP_25_64_8855/n586 ) );
  NAND \DP_OP_25_64_8855/U11  ( .A(\DP_OP_25_64_8855/n655 ), .B(
        \U1/RSOP_16/C2/Z_1 ), .Z(\DP_OP_25_64_8855/n452 ) );
  NAND \DP_OP_25_64_8855/U21  ( .A(\DP_OP_25_64_8855/n588 ), .B(
        \DP_OP_25_64_8855/n524 ), .Z(\DP_OP_25_64_8855/n453 ) );
  NAND \DP_OP_25_64_8855/U31  ( .A(\DP_OP_25_64_8855/n452 ), .B(
        \DP_OP_25_64_8855/n453 ), .Z(\DP_OP_25_64_8855/n587 ) );
  NAND \DP_OP_25_64_8855/U1  ( .A(\U1/RSOP_16/C2/Z_0 ), .B(\C1/Z_0 ), .Z(
        \DP_OP_25_64_8855/n459 ) );
  NAND \DP_OP_25_64_8855/U2  ( .A(\DP_OP_25_64_8855/n525 ), .B(
        \DP_OP_25_64_8855/n656 ), .Z(\DP_OP_25_64_8855/n460 ) );
  NAND \DP_OP_25_64_8855/U3  ( .A(\DP_OP_25_64_8855/n459 ), .B(
        \DP_OP_25_64_8855/n460 ), .Z(\DP_OP_25_64_8855/n588 ) );
  XOR U2965 ( .A(n5835), .B(n5834), .Z(n5746) );
  XOR U2966 ( .A(n5845), .B(n5844), .Z(n5846) );
  XOR U2967 ( .A(n7951), .B(n7950), .Z(n7742) );
  XOR U2968 ( .A(n7485), .B(n7484), .Z(n7288) );
  XOR U2969 ( .A(n5198), .B(n5197), .Z(n5074) );
  XOR U2970 ( .A(n4901), .B(n4900), .Z(n4788) );
  XOR U2971 ( .A(n8948), .B(n8947), .Z(n8728) );
  XOR U2972 ( .A(n10058), .B(n10057), .Z(n9791) );
  XOR U2973 ( .A(n12514), .B(n12515), .Z(n13421) );
  XOR U2974 ( .A(n13320), .B(n13321), .Z(n13670) );
  XOR U2975 ( .A(n13272), .B(n13273), .Z(n13622) );
  XOR U2976 ( .A(n13148), .B(n17175), .Z(n13496) );
  XOR U2977 ( .A(n11256), .B(n11255), .Z(n10963) );
  XOR U2978 ( .A(n10659), .B(n10660), .Z(n12532) );
  XOR U2979 ( .A(n12539), .B(n12540), .Z(n13448) );
  XOR U2980 ( .A(n14140), .B(n14141), .Z(n14498) );
  XOR U2981 ( .A(n4851), .B(n4850), .Z(n4852) );
  XOR U2982 ( .A(n5148), .B(n5147), .Z(n5149) );
  XOR U2983 ( .A(n5488), .B(n5487), .Z(n5489) );
  XOR U2984 ( .A(n5592), .B(n5591), .Z(n5586) );
  XOR U2985 ( .A(n4348), .B(n4347), .Z(n4317) );
  XOR U2986 ( .A(n4120), .B(n4119), .Z(n4121) );
  XOR U2987 ( .A(n5839), .B(n5838), .Z(n5840) );
  XOR U2988 ( .A(n5174), .B(n5173), .Z(n5097) );
  XOR U2989 ( .A(n4543), .B(n4542), .Z(n4544) );
  XOR U2990 ( .A(n4134), .B(n4133), .Z(n4093) );
  XOR U2991 ( .A(n3903), .B(n3902), .Z(n3904) );
  XOR U2992 ( .A(n3753), .B(n3752), .Z(n3754) );
  XOR U2993 ( .A(n5851), .B(n5850), .Z(n5853) );
  XOR U2994 ( .A(n6223), .B(n6222), .Z(n6086) );
  XOR U2995 ( .A(n5508), .B(n5507), .Z(n5395) );
  XOR U2996 ( .A(n6618), .B(n6617), .Z(n6620) );
  XOR U2997 ( .A(n5190), .B(n5189), .Z(n5191) );
  XOR U2998 ( .A(n4619), .B(n4618), .Z(n4620) );
  XOR U2999 ( .A(n3943), .B(n3942), .Z(n3944) );
  XOR U3000 ( .A(n7943), .B(n7942), .Z(n7944) );
  XOR U3001 ( .A(n5859), .B(n5858), .Z(n5723) );
  XOR U3002 ( .A(n5388), .B(n5387), .Z(n5390) );
  XOR U3003 ( .A(n7287), .B(n7286), .Z(n7289) );
  XOR U3004 ( .A(n6626), .B(n6625), .Z(n6458) );
  XOR U3005 ( .A(n5716), .B(n5715), .Z(n5718) );
  XOR U3006 ( .A(n5382), .B(n5381), .Z(n5384) );
  XOR U3007 ( .A(n4152), .B(n4151), .Z(n4075) );
  XOR U3008 ( .A(n16907), .B(n3950), .Z(n3886) );
  XOR U3009 ( .A(n3306), .B(n3305), .Z(n3307) );
  XOR U3010 ( .A(n8988), .B(n8987), .Z(n8989) );
  XOR U3011 ( .A(n4381), .B(n4380), .Z(n4382) );
  XOR U3012 ( .A(n9220), .B(n9219), .Z(n9221) );
  XOR U3013 ( .A(n8447), .B(n8446), .Z(n8214) );
  XOR U3014 ( .A(n7957), .B(n7956), .Z(n7736) );
  XOR U3015 ( .A(n7049), .B(n7048), .Z(n6853) );
  XOR U3016 ( .A(n5204), .B(n5203), .Z(n5068) );
  XOR U3017 ( .A(n4907), .B(n4906), .Z(n4782) );
  XOR U3018 ( .A(n10046), .B(n10045), .Z(n9803) );
  XOR U3019 ( .A(n6636), .B(n6635), .Z(n6637) );
  XOR U3020 ( .A(n5875), .B(n5874), .Z(n5876) );
  XOR U3021 ( .A(n3783), .B(n3782), .Z(n3784) );
  XOR U3022 ( .A(n10062), .B(n10061), .Z(n10063) );
  XOR U3023 ( .A(n5532), .B(n5531), .Z(n12390) );
  XOR U3024 ( .A(n4164), .B(n4163), .Z(n12332) );
  XOR U3025 ( .A(n10644), .B(n10643), .Z(n10365) );
  XOR U3026 ( .A(n12462), .B(n12463), .Z(n13369) );
  XOR U3027 ( .A(n12346), .B(n12347), .Z(n13247) );
  XOR U3028 ( .A(n13332), .B(n13333), .Z(n13682) );
  XOR U3029 ( .A(n13308), .B(n13309), .Z(n13658) );
  XOR U3030 ( .A(n13296), .B(n13297), .Z(n13646) );
  XOR U3031 ( .A(n13260), .B(n13261), .Z(n13610) );
  XOR U3032 ( .A(n13212), .B(n13213), .Z(n13566) );
  XOR U3033 ( .A(n13146), .B(n13147), .Z(n13497) );
  XOR U3034 ( .A(n10962), .B(n10961), .Z(n10964) );
  XOR U3035 ( .A(n13672), .B(n13673), .Z(n14033) );
  XOR U3036 ( .A(n13624), .B(n13625), .Z(n13985) );
  XOR U3037 ( .A(n13590), .B(n13591), .Z(n13949) );
  XOR U3038 ( .A(n13544), .B(n13545), .Z(n13899) );
  XOR U3039 ( .A(n13490), .B(n13491), .Z(n13831) );
  XOR U3040 ( .A(n12537), .B(n12538), .Z(n13449) );
  XOR U3041 ( .A(n13794), .B(n13795), .Z(n14156) );
  XOR U3042 ( .A(n14152), .B(n14153), .Z(n14510) );
  XOR U3043 ( .A(n13772), .B(n13773), .Z(n14132) );
  XOR U3044 ( .A(n14128), .B(n14129), .Z(n14486) );
  XOR U3045 ( .A(n14116), .B(n14117), .Z(n14474) );
  XOR U3046 ( .A(n14104), .B(n14105), .Z(n14462) );
  XOR U3047 ( .A(n13890), .B(n13891), .Z(n14255) );
  XOR U3048 ( .A(n13876), .B(n13877), .Z(n14187) );
  XOR U3049 ( .A(n4715), .B(n4714), .Z(n4698) );
  XOR U3050 ( .A(n4847), .B(n4846), .Z(n4834) );
  XOR U3051 ( .A(n4583), .B(n4582), .Z(n4584) );
  XOR U3052 ( .A(n4987), .B(n4986), .Z(n4970) );
  XOR U3053 ( .A(n4997), .B(n4996), .Z(n4998) );
  XOR U3054 ( .A(n4863), .B(n4862), .Z(n4864) );
  XOR U3055 ( .A(n4459), .B(n4458), .Z(n4442) );
  XOR U3056 ( .A(n5160), .B(n5159), .Z(n5161) );
  XOR U3057 ( .A(n5120), .B(n5119), .Z(n5121) );
  XOR U3058 ( .A(n4823), .B(n4822), .Z(n4824) );
  XOR U3059 ( .A(n4340), .B(n4339), .Z(n4341) );
  XOR U3060 ( .A(n5108), .B(n5107), .Z(n5109) );
  XOR U3061 ( .A(n5482), .B(n5481), .Z(n5483) );
  XOR U3062 ( .A(n4595), .B(n4594), .Z(n4596) );
  XOR U3063 ( .A(n4222), .B(n4221), .Z(n4205) );
  XOR U3064 ( .A(n5654), .B(n5653), .Z(n5655) );
  XOR U3065 ( .A(n5412), .B(n5411), .Z(n5414) );
  XOR U3066 ( .A(n4555), .B(n4554), .Z(n4557) );
  XOR U3067 ( .A(n5829), .B(n5828), .Z(n5752) );
  XOR U3068 ( .A(n5923), .B(n5922), .Z(n5924) );
  XOR U3069 ( .A(n4352), .B(n4351), .Z(n4353) );
  XOR U3070 ( .A(n6209), .B(n6208), .Z(n6210) );
  XOR U3071 ( .A(n5660), .B(n5659), .Z(n5661) );
  XOR U3072 ( .A(n5406), .B(n5405), .Z(n5408) );
  XOR U3073 ( .A(n5096), .B(n5095), .Z(n5098) );
  XOR U3074 ( .A(n4811), .B(n4810), .Z(n4813) );
  XOR U3075 ( .A(n4128), .B(n4127), .Z(n4097) );
  XOR U3076 ( .A(n3925), .B(n3924), .Z(n3926) );
  XOR U3077 ( .A(n6097), .B(n6096), .Z(n6098) );
  XOR U3078 ( .A(n6596), .B(n6595), .Z(n6488) );
  XOR U3079 ( .A(n4607), .B(n4606), .Z(n4609) );
  XOR U3080 ( .A(n3835), .B(n3834), .Z(n3818) );
  XOR U3081 ( .A(n6790), .B(n6789), .Z(n6791) );
  XOR U3082 ( .A(n6091), .B(n6090), .Z(n6093) );
  XOR U3083 ( .A(n5666), .B(n5665), .Z(n5667) );
  XOR U3084 ( .A(n5400), .B(n5399), .Z(n5402) );
  XOR U3085 ( .A(n5090), .B(n16714), .Z(n5091) );
  XOR U3086 ( .A(n3739), .B(n3738), .Z(n3755) );
  XOR U3087 ( .A(n6882), .B(n6881), .Z(n6883) );
  XOR U3088 ( .A(n7095), .B(n7094), .Z(n7096) );
  XOR U3089 ( .A(n7029), .B(n7028), .Z(n7030) );
  XOR U3090 ( .A(n4138), .B(n4137), .Z(n4139) );
  XOR U3091 ( .A(n3937), .B(n3936), .Z(n3938) );
  XOR U3092 ( .A(n3665), .B(n3664), .Z(n3666) );
  XOR U3093 ( .A(n6870), .B(n6869), .Z(n6871) );
  XOR U3094 ( .A(n6085), .B(n6084), .Z(n6087) );
  XOR U3095 ( .A(n5672), .B(n5671), .Z(n5673) );
  XOR U3096 ( .A(n5394), .B(n5393), .Z(n5396) );
  XOR U3097 ( .A(n4799), .B(n4798), .Z(n4800) );
  XOR U3098 ( .A(n4615), .B(n4614), .Z(n4538) );
  XOR U3099 ( .A(n4086), .B(n4085), .Z(n4087) );
  XOR U3100 ( .A(n7311), .B(n7310), .Z(n7312) );
  XOR U3101 ( .A(n7471), .B(n7470), .Z(n7472) );
  XOR U3102 ( .A(n7539), .B(n7538), .Z(n7533) );
  XOR U3103 ( .A(n3765), .B(n3764), .Z(n3767) );
  XOR U3104 ( .A(n3517), .B(n3516), .Z(n3518) );
  XOR U3105 ( .A(n7927), .B(n7926), .Z(n7766) );
  XOR U3106 ( .A(n7709), .B(n7708), .Z(n7710) );
  XOR U3107 ( .A(n7479), .B(n7478), .Z(n7294) );
  XOR U3108 ( .A(n6269), .B(n6268), .Z(n6270) );
  XOR U3109 ( .A(n6079), .B(n6078), .Z(n6081) );
  XOR U3110 ( .A(n5684), .B(n5683), .Z(n5685) );
  XOR U3111 ( .A(n5192), .B(n5191), .Z(n5080) );
  XOR U3112 ( .A(n4505), .B(n4504), .Z(n4506) );
  XOR U3113 ( .A(n4048), .B(n4047), .Z(n4049) );
  XOR U3114 ( .A(n3891), .B(n3890), .Z(n3892) );
  XOR U3115 ( .A(n3725), .B(n3724), .Z(n3727) );
  XOR U3116 ( .A(n3481), .B(n3480), .Z(n3482) );
  XOR U3117 ( .A(n3302), .B(n3301), .Z(n3289) );
  XOR U3118 ( .A(n8225), .B(n8224), .Z(n8226) );
  XOR U3119 ( .A(n8423), .B(n8422), .Z(n8239) );
  XOR U3120 ( .A(n5863), .B(n5862), .Z(n5864) );
  XOR U3121 ( .A(n5518), .B(n5517), .Z(n5519) );
  XOR U3122 ( .A(n3617), .B(n3616), .Z(n3618) );
  XOR U3123 ( .A(n3428), .B(n3427), .Z(n3411) );
  XOR U3124 ( .A(n8681), .B(n8680), .Z(n8682) );
  XOR U3125 ( .A(n8219), .B(n8218), .Z(n8221) );
  XOR U3126 ( .A(n7715), .B(n7714), .Z(n7716) );
  XOR U3127 ( .A(n6654), .B(n6653), .Z(n6655) );
  XOR U3128 ( .A(n5045), .B(n5044), .Z(n5046) );
  XOR U3129 ( .A(n4787), .B(n4786), .Z(n4789) );
  XOR U3130 ( .A(n4262), .B(n4261), .Z(n4264) );
  XOR U3131 ( .A(n4074), .B(n4073), .Z(n4076) );
  XOR U3132 ( .A(n3719), .B(n3718), .Z(n3720) );
  XOR U3133 ( .A(n3577), .B(n3576), .Z(n3579) );
  XOR U3134 ( .A(n8693), .B(n8692), .Z(n8694) );
  XOR U3135 ( .A(n8946), .B(n8945), .Z(n8947) );
  XOR U3136 ( .A(n6630), .B(n6629), .Z(n6631) );
  XOR U3137 ( .A(n3493), .B(n3492), .Z(n3494) );
  XOR U3138 ( .A(n3235), .B(n3236), .Z(n3254) );
  XOR U3139 ( .A(n8990), .B(n8989), .Z(n9222) );
  XNOR U3140 ( .A(n9260), .B(n9259), .Z(n9483) );
  XOR U3141 ( .A(n8213), .B(n8212), .Z(n8215) );
  XOR U3142 ( .A(n7721), .B(n7720), .Z(n7722) );
  XOR U3143 ( .A(n7491), .B(n7490), .Z(n7282) );
  XOR U3144 ( .A(n5871), .B(n5870), .Z(n5711) );
  XOR U3145 ( .A(n5526), .B(n5525), .Z(n5377) );
  XOR U3146 ( .A(n5067), .B(n5066), .Z(n5069) );
  XOR U3147 ( .A(n5051), .B(n5050), .Z(n5052) );
  XOR U3148 ( .A(n4519), .B(n4518), .Z(n4521) );
  XOR U3149 ( .A(n4383), .B(n4382), .Z(n4283) );
  XOR U3150 ( .A(n4268), .B(n4267), .Z(n4269) );
  XOR U3151 ( .A(n4068), .B(n4067), .Z(n4070) );
  XOR U3152 ( .A(n4054), .B(n4053), .Z(n4055) );
  XOR U3153 ( .A(n3956), .B(n3955), .Z(n3880) );
  XOR U3154 ( .A(n3647), .B(n3646), .Z(n3648) );
  XOR U3155 ( .A(n3453), .B(n17020), .Z(n3455) );
  XOR U3156 ( .A(n3314), .B(n3313), .Z(n3286) );
  XOR U3157 ( .A(n9757), .B(n9756), .Z(n9758) );
  XOR U3158 ( .A(n7961), .B(n7960), .Z(n7962) );
  XOR U3159 ( .A(n3333), .B(n3334), .Z(n3355) );
  XOR U3160 ( .A(n10081), .B(n10080), .Z(n10082) );
  XOR U3161 ( .A(n7970), .B(n7971), .Z(n12473) );
  XOR U3162 ( .A(n7062), .B(n7063), .Z(n12449) );
  XOR U3163 ( .A(n7055), .B(n7054), .Z(n12436) );
  XOR U3164 ( .A(n6638), .B(n6637), .Z(n12424) );
  XOR U3165 ( .A(n6059), .B(n6058), .Z(n6060) );
  XOR U3166 ( .A(n5368), .B(n5367), .Z(n5369) );
  XOR U3167 ( .A(n5062), .B(n5063), .Z(n12378) );
  XOR U3168 ( .A(n5057), .B(n5056), .Z(n5058) );
  XOR U3169 ( .A(n4913), .B(n4912), .Z(n12366) );
  XOR U3170 ( .A(n4274), .B(n4273), .Z(n4275) );
  XOR U3171 ( .A(n3785), .B(n3784), .Z(n12310) );
  XOR U3172 ( .A(n3563), .B(n3562), .Z(n3564) );
  XOR U3173 ( .A(n3449), .B(n3450), .Z(n12231) );
  XOR U3174 ( .A(n10064), .B(n10063), .Z(n12506) );
  XOR U3175 ( .A(n10337), .B(n10336), .Z(n10338) );
  XOR U3176 ( .A(n12392), .B(n12393), .Z(n13295) );
  XOR U3177 ( .A(n12300), .B(n12301), .Z(n13201) );
  XOR U3178 ( .A(n12278), .B(n12279), .Z(n13177) );
  XOR U3179 ( .A(n12266), .B(n12267), .Z(n13167) );
  XOR U3180 ( .A(n12249), .B(n12250), .Z(n13130) );
  XOR U3181 ( .A(n10662), .B(n10661), .Z(n10663) );
  XOR U3182 ( .A(n13414), .B(n13415), .Z(n13765) );
  XOR U3183 ( .A(n12490), .B(n12491), .Z(n13396) );
  XOR U3184 ( .A(n13392), .B(n13393), .Z(n13742) );
  XOR U3185 ( .A(n13368), .B(n13369), .Z(n13718) );
  XOR U3186 ( .A(n13342), .B(n13343), .Z(n13695) );
  XOR U3187 ( .A(n13330), .B(n13331), .Z(n13683) );
  XOR U3188 ( .A(n12420), .B(n12421), .Z(n13324) );
  XOR U3189 ( .A(n12410), .B(n12411), .Z(n13312) );
  XOR U3190 ( .A(n12374), .B(n12375), .Z(n13276) );
  XOR U3191 ( .A(n12362), .B(n12363), .Z(n13264) );
  XOR U3192 ( .A(n12340), .B(n12341), .Z(n13240) );
  XOR U3193 ( .A(n13236), .B(n13237), .Z(n13588) );
  XOR U3194 ( .A(n13178), .B(n13179), .Z(n13475) );
  XOR U3195 ( .A(n13168), .B(n13169), .Z(n13520) );
  XOR U3196 ( .A(n11262), .B(n11261), .Z(n12531) );
  XOR U3197 ( .A(n11570), .B(n11569), .Z(n11571) );
  XOR U3198 ( .A(n12622), .B(n12621), .Z(n12620) );
  XOR U3199 ( .A(n13450), .B(n13451), .Z(n13793) );
  XOR U3200 ( .A(n13732), .B(n13733), .Z(n14091) );
  XOR U3201 ( .A(n13510), .B(n13511), .Z(n13867) );
  XOR U3202 ( .A(n13800), .B(n13801), .Z(n14163) );
  XOR U3203 ( .A(n14150), .B(n14151), .Z(n14511) );
  XOR U3204 ( .A(n13782), .B(n13783), .Z(n14144) );
  XOR U3205 ( .A(n14126), .B(n14127), .Z(n14487) );
  XOR U3206 ( .A(n13750), .B(n13751), .Z(n14108) );
  XOR U3207 ( .A(n14102), .B(n14103), .Z(n14463) );
  XOR U3208 ( .A(n14078), .B(n14079), .Z(n14441) );
  XOR U3209 ( .A(n14068), .B(n14069), .Z(n14428) );
  XOR U3210 ( .A(n14044), .B(n14045), .Z(n14404) );
  XOR U3211 ( .A(n13678), .B(n13679), .Z(n14036) );
  XOR U3212 ( .A(n14030), .B(n14031), .Z(n14393) );
  XOR U3213 ( .A(n14020), .B(n14021), .Z(n14380) );
  XOR U3214 ( .A(n14006), .B(n14007), .Z(n14369) );
  XOR U3215 ( .A(n13630), .B(n13631), .Z(n13988) );
  XOR U3216 ( .A(n13982), .B(n13983), .Z(n14347) );
  XOR U3217 ( .A(n13972), .B(n13973), .Z(n14334) );
  XOR U3218 ( .A(n13596), .B(n13597), .Z(n13952) );
  XOR U3219 ( .A(n13946), .B(n13947), .Z(n14313) );
  XOR U3220 ( .A(n13936), .B(n13937), .Z(n14300) );
  XOR U3221 ( .A(n13922), .B(n13923), .Z(n14289) );
  XOR U3222 ( .A(n13912), .B(n13913), .Z(n14185) );
  XOR U3223 ( .A(n13550), .B(n13551), .Z(n13905) );
  XOR U3224 ( .A(n13900), .B(n13901), .Z(n14266) );
  XOR U3225 ( .A(n13868), .B(n13869), .Z(n14232) );
  XOR U3226 ( .A(n13854), .B(n13855), .Z(n13857) );
  XOR U3227 ( .A(n13846), .B(n13847), .Z(n14208) );
  XOR U3228 ( .A(n14164), .B(n14165), .Z(n14177) );
  XOR U3229 ( .A(n11895), .B(n11894), .Z(n12543) );
  XOR U3230 ( .A(n13463), .B(n13464), .Z(n13804) );
  XOR U3231 ( .A(n14254), .B(n14255), .Z(n14257) );
  XOR U3232 ( .A(n14196), .B(n14197), .Z(n14199) );
  XNOR U3233 ( .A(n13124), .B(n13125), .Z(n13815) );
  XOR U3234 ( .A(n14244), .B(n14245), .Z(n14643) );
  XOR U3235 ( .A(n4579), .B(n4578), .Z(n4566) );
  XOR U3236 ( .A(n4857), .B(n4856), .Z(n4858) );
  XOR U3237 ( .A(n4969), .B(n4968), .Z(n4971) );
  XOR U3238 ( .A(n4719), .B(n4718), .Z(n4720) );
  XOR U3239 ( .A(n4978), .B(n4977), .Z(n4984) );
  XOR U3240 ( .A(n4963), .B(n4962), .Z(n4964) );
  XOR U3241 ( .A(n4589), .B(n4588), .Z(n4590) );
  XOR U3242 ( .A(n4324), .B(n4323), .Z(n4325) );
  XOR U3243 ( .A(n5150), .B(n5149), .Z(n5119) );
  XOR U3244 ( .A(n5156), .B(n5155), .Z(n5115) );
  XOR U3245 ( .A(n5003), .B(n5002), .Z(n5004) );
  XOR U3246 ( .A(n4865), .B(n4864), .Z(n4825) );
  XOR U3247 ( .A(n4116), .B(n4115), .Z(n4103) );
  XOR U3248 ( .A(n5430), .B(n5429), .Z(n5432) );
  XOR U3249 ( .A(n5424), .B(n5423), .Z(n5425) );
  XOR U3250 ( .A(n5268), .B(n5267), .Z(n5269) );
  XOR U3251 ( .A(n4731), .B(n4730), .Z(n4732) );
  XOR U3252 ( .A(n4465), .B(n4464), .Z(n4468) );
  XOR U3253 ( .A(n5484), .B(n5483), .Z(n5419) );
  XOR U3254 ( .A(n5584), .B(n5583), .Z(n5585) );
  XOR U3255 ( .A(n5650), .B(n5649), .Z(n5589) );
  XOR U3256 ( .A(n5102), .B(n5101), .Z(n5104) );
  XOR U3257 ( .A(n4817), .B(n4816), .Z(n4818) );
  XOR U3258 ( .A(n4737), .B(n4736), .Z(n4738) );
  XOR U3259 ( .A(n4318), .B(n4317), .Z(n4319) );
  XOR U3260 ( .A(n5656), .B(n5655), .Z(n5571) );
  XOR U3261 ( .A(n5931), .B(n5930), .Z(n5925) );
  XOR U3262 ( .A(n5494), .B(n5493), .Z(n5495) );
  XOR U3263 ( .A(n4228), .B(n4227), .Z(n4231) );
  XOR U3264 ( .A(n3909), .B(n3908), .Z(n3910) );
  XNOR U3265 ( .A(n6385), .B(n6384), .Z(n6335) );
  XOR U3266 ( .A(n5841), .B(n5840), .Z(n5740) );
  XOR U3267 ( .A(n4685), .B(n4684), .Z(n4686) );
  XOR U3268 ( .A(n4603), .B(n4602), .Z(n4551) );
  XOR U3269 ( .A(n4312), .B(n4311), .Z(n4313) );
  XOR U3270 ( .A(n4098), .B(n4097), .Z(n4099) );
  XOR U3271 ( .A(n6407), .B(n6406), .Z(n6408) );
  XOR U3272 ( .A(n3749), .B(n3748), .Z(n3736) );
  XNOR U3273 ( .A(n6099), .B(n6098), .Z(n6215) );
  XOR U3274 ( .A(n6600), .B(n6599), .Z(n6602) );
  XOR U3275 ( .A(n5566), .B(n5565), .Z(n5567) );
  XOR U3276 ( .A(n4881), .B(n4880), .Z(n4883) );
  XOR U3277 ( .A(n4026), .B(n4025), .Z(n4029) );
  XOR U3278 ( .A(n6023), .B(n6022), .Z(n6024) );
  XOR U3279 ( .A(n5734), .B(n5733), .Z(n5736) );
  XOR U3280 ( .A(n5180), .B(n5179), .Z(n5092) );
  XOR U3281 ( .A(n4487), .B(n4486), .Z(n4488) );
  XOR U3282 ( .A(n4306), .B(n4305), .Z(n4307) );
  XOR U3283 ( .A(n4092), .B(n4091), .Z(n4094) );
  XOR U3284 ( .A(n3674), .B(n3673), .Z(n3680) );
  XNOR U3285 ( .A(n6902), .B(n6901), .Z(n7006) );
  XOR U3286 ( .A(n3839), .B(n3838), .Z(n3840) );
  XOR U3287 ( .A(n6802), .B(n6801), .Z(n6803) );
  XOR U3288 ( .A(n7019), .B(n7018), .Z(n6884) );
  XOR U3289 ( .A(n7103), .B(n7102), .Z(n7097) );
  XOR U3290 ( .A(n6612), .B(n6611), .Z(n6614) );
  XOR U3291 ( .A(n6221), .B(n6220), .Z(n6222) );
  XOR U3292 ( .A(n4667), .B(n4666), .Z(n4669) );
  XOR U3293 ( .A(n3759), .B(n3758), .Z(n3760) );
  XOR U3294 ( .A(n7089), .B(n7088), .Z(n7090) );
  XOR U3295 ( .A(n7317), .B(n7316), .Z(n7319) );
  XOR U3296 ( .A(n7031), .B(n7030), .Z(n6872) );
  XOR U3297 ( .A(n5728), .B(n5727), .Z(n5729) );
  XOR U3298 ( .A(n5562), .B(n5561), .Z(n5674) );
  XOR U3299 ( .A(n4661), .B(n4660), .Z(n4662) );
  XOR U3300 ( .A(n4499), .B(n4498), .Z(n4500) );
  XOR U3301 ( .A(n4300), .B(n4299), .Z(n4301) );
  XOR U3302 ( .A(n4192), .B(n4191), .Z(n4193) );
  XOR U3303 ( .A(n3939), .B(n3938), .Z(n3898) );
  XOR U3304 ( .A(n3605), .B(n3604), .Z(n3606) );
  XOR U3305 ( .A(n7467), .B(n7466), .Z(n7306) );
  XOR U3306 ( .A(n7697), .B(n7696), .Z(n7698) );
  XOR U3307 ( .A(n8091), .B(n8090), .Z(n8093) );
  XNOR U3308 ( .A(n4801), .B(n4800), .Z(n4893) );
  XOR U3309 ( .A(n3687), .B(n3686), .Z(n3688) );
  XOR U3310 ( .A(n7299), .B(n7298), .Z(n7301) );
  XOR U3311 ( .A(n7531), .B(n7530), .Z(n7532) );
  XNOR U3312 ( .A(n8035), .B(n8034), .Z(n8103) );
  XOR U3313 ( .A(n5512), .B(n5511), .Z(n5513) );
  XOR U3314 ( .A(n4144), .B(n4143), .Z(n4145) );
  XOR U3315 ( .A(n3811), .B(n3810), .Z(n3812) );
  XOR U3316 ( .A(n7703), .B(n7702), .Z(n7704) );
  XOR U3317 ( .A(n7765), .B(n7764), .Z(n7767) );
  XOR U3318 ( .A(n7759), .B(n7758), .Z(n7761) );
  XOR U3319 ( .A(n8869), .B(n8868), .Z(n8871) );
  XOR U3320 ( .A(n6463), .B(n6462), .Z(n6464) );
  XOR U3321 ( .A(n6277), .B(n6276), .Z(n6271) );
  XOR U3322 ( .A(n6229), .B(n6228), .Z(n6080) );
  XOR U3323 ( .A(n4793), .B(n4792), .Z(n4794) );
  XOR U3324 ( .A(n4621), .B(n4620), .Z(n4532) );
  XOR U3325 ( .A(n3851), .B(n3850), .Z(n3852) );
  XNOR U3326 ( .A(n3519), .B(n3518), .Z(n3538) );
  XOR U3327 ( .A(n8181), .B(n8180), .Z(n8182) );
  XNOR U3328 ( .A(n8263), .B(n8262), .Z(n8403) );
  XOR U3329 ( .A(n8823), .B(n8822), .Z(n8825) );
  XOR U3330 ( .A(n8169), .B(n8168), .Z(n8170) );
  XOR U3331 ( .A(n8243), .B(n8242), .Z(n8245) );
  XOR U3332 ( .A(n8433), .B(n8432), .Z(n8435) );
  XOR U3333 ( .A(n8187), .B(n8186), .Z(n8188) );
  XOR U3334 ( .A(n7949), .B(n7948), .Z(n7950) );
  XOR U3335 ( .A(n7519), .B(n7518), .Z(n7520) );
  XOR U3336 ( .A(n7041), .B(n7040), .Z(n7043) );
  XOR U3337 ( .A(n5893), .B(n5892), .Z(n5894) );
  XOR U3338 ( .A(n5554), .B(n5553), .Z(n5555) );
  XOR U3339 ( .A(n5196), .B(n5195), .Z(n5197) );
  XOR U3340 ( .A(n4423), .B(n4422), .Z(n4424) );
  XOR U3341 ( .A(n4186), .B(n4185), .Z(n4187) );
  XOR U3342 ( .A(n3990), .B(n3989), .Z(n3991) );
  XOR U3343 ( .A(n3659), .B(n3658), .Z(n3660) );
  XOR U3344 ( .A(n3487), .B(n3486), .Z(n3488) );
  XOR U3345 ( .A(n3290), .B(n3289), .Z(n3291) );
  XOR U3346 ( .A(n8485), .B(n8484), .Z(n8486) );
  XOR U3347 ( .A(n9026), .B(n9025), .Z(n9149) );
  XOR U3348 ( .A(n7741), .B(n7740), .Z(n7743) );
  XOR U3349 ( .A(n6431), .B(n6430), .Z(n6432) );
  XOR U3350 ( .A(n6073), .B(n6072), .Z(n6075) );
  XOR U3351 ( .A(n6041), .B(n6040), .Z(n6042) );
  XOR U3352 ( .A(n5690), .B(n5689), .Z(n5691) );
  XOR U3353 ( .A(n5073), .B(n5072), .Z(n5075) );
  XOR U3354 ( .A(n4525), .B(n4524), .Z(n4527) );
  XOR U3355 ( .A(n4511), .B(n4510), .Z(n4512) );
  XOR U3356 ( .A(n4377), .B(n4376), .Z(n4289) );
  XOR U3357 ( .A(n3984), .B(n3983), .Z(n3985) );
  XOR U3358 ( .A(n3885), .B(n3884), .Z(n3887) );
  XOR U3359 ( .A(n3699), .B(n3698), .Z(n3700) );
  XOR U3360 ( .A(n3619), .B(n3618), .Z(n3578) );
  XOR U3361 ( .A(n8475), .B(n8474), .Z(n8695) );
  XOR U3362 ( .A(n8727), .B(n8726), .Z(n8729) );
  XNOR U3363 ( .A(n9569), .B(n9568), .Z(n9661) );
  XOR U3364 ( .A(n9927), .B(n9926), .Z(n9929) );
  XOR U3365 ( .A(n8942), .B(n8941), .Z(n8734) );
  XOR U3366 ( .A(n9198), .B(n9197), .Z(n9204) );
  XOR U3367 ( .A(n8958), .B(n8957), .Z(n8960) );
  XOR U3368 ( .A(n8445), .B(n8444), .Z(n8446) );
  XOR U3369 ( .A(n6832), .B(n6831), .Z(n6833) );
  XOR U3370 ( .A(n5869), .B(n5868), .Z(n5870) );
  XOR U3371 ( .A(n5524), .B(n5523), .Z(n5525) );
  XOR U3372 ( .A(n3511), .B(n3510), .Z(n3512) );
  XOR U3373 ( .A(n3434), .B(n3433), .Z(n3437) );
  XNOR U3374 ( .A(n10472), .B(n10471), .Z(n10464) );
  XOR U3375 ( .A(n9226), .B(n9225), .Z(n9227) );
  XOR U3376 ( .A(n8715), .B(n8714), .Z(n8717) );
  XOR U3377 ( .A(n7735), .B(n7734), .Z(n7737) );
  XOR U3378 ( .A(n7515), .B(n7514), .Z(n7723) );
  XOR U3379 ( .A(n7281), .B(n7280), .Z(n7283) );
  XOR U3380 ( .A(n7267), .B(n7266), .Z(n7268) );
  XOR U3381 ( .A(n6852), .B(n6851), .Z(n6854) );
  XOR U3382 ( .A(n6838), .B(n6837), .Z(n6839) );
  XOR U3383 ( .A(n6632), .B(n6631), .Z(n6452) );
  XOR U3384 ( .A(n6067), .B(n6066), .Z(n6068) );
  XOR U3385 ( .A(n4929), .B(n4928), .Z(n5053) );
  XOR U3386 ( .A(n4781), .B(n4780), .Z(n4783) );
  XOR U3387 ( .A(n4767), .B(n4766), .Z(n4768) );
  XOR U3388 ( .A(n4182), .B(n4181), .Z(n4270) );
  XOR U3389 ( .A(n4158), .B(n4157), .Z(n4069) );
  XOR U3390 ( .A(n3879), .B(n3878), .Z(n3881) );
  XOR U3391 ( .A(n3779), .B(n3778), .Z(n3714) );
  XOR U3392 ( .A(n3551), .B(n3550), .Z(n3552) );
  XOR U3393 ( .A(n3255), .B(n3256), .Z(n3337) );
  XNOR U3394 ( .A(n3266), .B(n3265), .Z(n3260) );
  XOR U3395 ( .A(n9745), .B(n9744), .Z(n9746) );
  XOR U3396 ( .A(n4056), .B(n4055), .Z(n3971) );
  XOR U3397 ( .A(n3649), .B(n3648), .Z(n3640) );
  XOR U3398 ( .A(n9769), .B(n9768), .Z(n9770) );
  XOR U3399 ( .A(n9501), .B(n9500), .Z(n9503) );
  XOR U3400 ( .A(n5542), .B(n5541), .Z(n5543) );
  XOR U3401 ( .A(n4405), .B(n4404), .Z(n4406) );
  XOR U3402 ( .A(n3629), .B(n3628), .Z(n3630) );
  XOR U3403 ( .A(n3499), .B(n3498), .Z(n3500) );
  XOR U3404 ( .A(n3351), .B(n3352), .Z(n3395) );
  XOR U3405 ( .A(n3327), .B(n3328), .Z(n3371) );
  XOR U3406 ( .A(n10050), .B(n10049), .Z(n10051) );
  XNOR U3407 ( .A(n10401), .B(n10400), .Z(n10612) );
  XOR U3408 ( .A(n9795), .B(n9794), .Z(n9796) );
  XOR U3409 ( .A(n8710), .B(n8711), .Z(n12224) );
  XOR U3410 ( .A(n8453), .B(n8452), .Z(n12472) );
  XOR U3411 ( .A(n7727), .B(n7726), .Z(n7728) );
  XOR U3412 ( .A(n6645), .B(n6646), .Z(n12437) );
  XOR U3413 ( .A(n6055), .B(n6054), .Z(n6061) );
  XOR U3414 ( .A(n5539), .B(n5540), .Z(n12403) );
  XOR U3415 ( .A(n5702), .B(n5701), .Z(n5703) );
  XOR U3416 ( .A(n5217), .B(n5218), .Z(n12391) );
  XOR U3417 ( .A(n5222), .B(n5221), .Z(n5370) );
  XOR U3418 ( .A(n5210), .B(n5209), .Z(n12379) );
  XOR U3419 ( .A(n4773), .B(n4772), .Z(n4774) );
  XOR U3420 ( .A(n4396), .B(n4397), .Z(n12228) );
  XOR U3421 ( .A(n4399), .B(n4398), .Z(n4400) );
  XOR U3422 ( .A(n4389), .B(n4388), .Z(n12344) );
  XOR U3423 ( .A(n4060), .B(n4059), .Z(n4061) );
  XOR U3424 ( .A(n3869), .B(n3868), .Z(n3870) );
  XOR U3425 ( .A(n3638), .B(n3639), .Z(n12311) );
  XOR U3426 ( .A(n3373), .B(n3374), .Z(n12253) );
  XOR U3427 ( .A(n9510), .B(n9511), .Z(n12507) );
  XOR U3428 ( .A(n10349), .B(n10348), .Z(n10350) );
  XOR U3429 ( .A(n10355), .B(n10354), .Z(n10356) );
  XOR U3430 ( .A(n10083), .B(n10082), .Z(n10339) );
  XOR U3431 ( .A(n10375), .B(n10374), .Z(n10377) );
  XNOR U3432 ( .A(n10389), .B(n10388), .Z(n10624) );
  XOR U3433 ( .A(n12005), .B(n12004), .Z(n12006) );
  XNOR U3434 ( .A(n12229), .B(n12230), .Z(n12323) );
  XOR U3435 ( .A(n3377), .B(n3378), .Z(n12260) );
  XOR U3436 ( .A(n10642), .B(n10641), .Z(n10643) );
  XOR U3437 ( .A(n7966), .B(n7967), .Z(n12467) );
  XOR U3438 ( .A(n12426), .B(n12427), .Z(n13333) );
  XOR U3439 ( .A(n4916), .B(n4917), .Z(n12373) );
  XOR U3440 ( .A(n4167), .B(n4168), .Z(n12339) );
  XOR U3441 ( .A(n12334), .B(n12335), .Z(n13237) );
  XOR U3442 ( .A(n3504), .B(n3505), .Z(n12293) );
  XOR U3443 ( .A(n3399), .B(n3400), .Z(n12283) );
  XOR U3444 ( .A(n3389), .B(n3390), .Z(n12271) );
  XOR U3445 ( .A(n12247), .B(n12248), .Z(n13131) );
  XOR U3446 ( .A(n12652), .B(n12651), .Z(n12650) );
  XOR U3447 ( .A(n10942), .B(n10941), .Z(n10943) );
  XOR U3448 ( .A(n13404), .B(n13405), .Z(n13470) );
  XOR U3449 ( .A(n12468), .B(n12469), .Z(n13372) );
  XOR U3450 ( .A(n13366), .B(n13367), .Z(n13719) );
  XOR U3451 ( .A(n12456), .B(n12457), .Z(n13360) );
  XOR U3452 ( .A(n13356), .B(n13357), .Z(n13706) );
  XOR U3453 ( .A(n12386), .B(n12387), .Z(n13288) );
  XOR U3454 ( .A(n13282), .B(n13283), .Z(n13635) );
  XOR U3455 ( .A(n12294), .B(n12295), .Z(n13126) );
  XOR U3456 ( .A(n13190), .B(n13191), .Z(n13543) );
  XOR U3457 ( .A(n12284), .B(n12285), .Z(n13183) );
  XOR U3458 ( .A(n13176), .B(n13177), .Z(n13476) );
  XOR U3459 ( .A(n12272), .B(n12273), .Z(n13128) );
  XOR U3460 ( .A(n13140), .B(n13141), .Z(n13143) );
  XNOR U3461 ( .A(n13471), .B(n13472), .Z(n13601) );
  XNOR U3462 ( .A(n12608), .B(n12607), .Z(n12971) );
  XOR U3463 ( .A(n13338), .B(n13339), .Z(n13689) );
  XOR U3464 ( .A(n13314), .B(n13315), .Z(n13665) );
  XOR U3465 ( .A(n13302), .B(n13303), .Z(n13653) );
  XOR U3466 ( .A(n13266), .B(n13267), .Z(n13617) );
  XOR U3467 ( .A(n13218), .B(n13219), .Z(n13573) );
  XOR U3468 ( .A(n13556), .B(n13557), .Z(n13911) );
  XOR U3469 ( .A(n13162), .B(n13163), .Z(n13515) );
  XOR U3470 ( .A(n11584), .B(n11583), .Z(n11585) );
  XOR U3471 ( .A(n13792), .B(n13793), .Z(n14157) );
  XOR U3472 ( .A(n13780), .B(n13781), .Z(n14145) );
  XOR U3473 ( .A(n13770), .B(n13771), .Z(n14133) );
  XOR U3474 ( .A(n13760), .B(n13761), .Z(n14120) );
  XOR U3475 ( .A(n13748), .B(n13749), .Z(n14109) );
  XOR U3476 ( .A(n13714), .B(n13715), .Z(n14072) );
  XOR U3477 ( .A(n13702), .B(n13703), .Z(n14060) );
  XOR U3478 ( .A(n13690), .B(n13691), .Z(n14048) );
  XOR U3479 ( .A(n13676), .B(n13677), .Z(n14037) );
  XOR U3480 ( .A(n13666), .B(n13667), .Z(n14024) );
  XOR U3481 ( .A(n13654), .B(n13655), .Z(n14012) );
  XOR U3482 ( .A(n13642), .B(n13643), .Z(n14000) );
  XOR U3483 ( .A(n13996), .B(n13997), .Z(n14181) );
  XOR U3484 ( .A(n13628), .B(n13629), .Z(n13989) );
  XOR U3485 ( .A(n13618), .B(n13619), .Z(n13976) );
  XOR U3486 ( .A(n13960), .B(n13961), .Z(n14183) );
  XOR U3487 ( .A(n13594), .B(n13595), .Z(n13953) );
  XOR U3488 ( .A(n13574), .B(n13575), .Z(n13928) );
  XOR U3489 ( .A(n13528), .B(n13529), .Z(n13883) );
  XOR U3490 ( .A(n13516), .B(n13517), .Z(n13828) );
  XOR U3491 ( .A(n13504), .B(n13505), .Z(n13860) );
  XOR U3492 ( .A(n11269), .B(n11270), .Z(n12544) );
  XOR U3493 ( .A(n11917), .B(n11916), .Z(n12208) );
  XNOR U3494 ( .A(n14176), .B(n14177), .Z(n14523) );
  XNOR U3495 ( .A(n14178), .B(n14179), .Z(n14453) );
  XOR U3496 ( .A(n13904), .B(n13905), .Z(n13907) );
  XOR U3497 ( .A(n13850), .B(n13851), .Z(n14215) );
  XOR U3498 ( .A(n12551), .B(n12552), .Z(n13461) );
  XOR U3499 ( .A(n14512), .B(n14513), .Z(n14535) );
  XOR U3500 ( .A(n14500), .B(n14501), .Z(n14537) );
  XOR U3501 ( .A(n14488), .B(n14489), .Z(n14539) );
  XOR U3502 ( .A(n14476), .B(n14477), .Z(n14541) );
  XOR U3503 ( .A(n14464), .B(n14465), .Z(n14543) );
  XOR U3504 ( .A(n14442), .B(n14443), .Z(n14547) );
  XOR U3505 ( .A(n14430), .B(n14431), .Z(n14549) );
  XOR U3506 ( .A(n14418), .B(n14419), .Z(n14551) );
  XOR U3507 ( .A(n14406), .B(n14407), .Z(n14553) );
  XOR U3508 ( .A(n14394), .B(n14395), .Z(n14555) );
  XOR U3509 ( .A(n14382), .B(n14383), .Z(n14557) );
  XOR U3510 ( .A(n14370), .B(n14371), .Z(n14559) );
  XOR U3511 ( .A(n14348), .B(n14349), .Z(n14563) );
  XOR U3512 ( .A(n14336), .B(n14337), .Z(n14565) );
  XOR U3513 ( .A(n14314), .B(n14315), .Z(n14569) );
  XOR U3514 ( .A(n14302), .B(n14303), .Z(n14571) );
  XOR U3515 ( .A(n14290), .B(n14291), .Z(n14573) );
  XOR U3516 ( .A(n14268), .B(n14269), .Z(n14577) );
  XOR U3517 ( .A(n14256), .B(n14257), .Z(n14579) );
  XOR U3518 ( .A(n14234), .B(n14235), .Z(n14581) );
  XOR U3519 ( .A(n14222), .B(n14223), .Z(n14621) );
  XOR U3520 ( .A(n14210), .B(n14211), .Z(n14583) );
  XOR U3521 ( .A(n14198), .B(n14199), .Z(n14585) );
  XOR U3522 ( .A(n14901), .B(n14900), .Z(n14899) );
  XOR U3523 ( .A(n14642), .B(n14643), .Z(n14645) );
  XOR U3524 ( .A(n4567), .B(n4566), .Z(n4568) );
  XOR U3525 ( .A(n4706), .B(n4705), .Z(n4712) );
  XOR U3526 ( .A(n4450), .B(n4449), .Z(n4456) );
  XOR U3527 ( .A(n4837), .B(n4836), .Z(n4853) );
  XOR U3528 ( .A(n4829), .B(n4828), .Z(n4830) );
  XOR U3529 ( .A(n4336), .B(n4335), .Z(n4323) );
  XOR U3530 ( .A(n4991), .B(n4990), .Z(n4992) );
  XOR U3531 ( .A(n5126), .B(n5125), .Z(n5127) );
  XOR U3532 ( .A(n4721), .B(n4720), .Z(n4724) );
  XOR U3533 ( .A(n5142), .B(n5141), .Z(n5143) );
  XOR U3534 ( .A(n5154), .B(n5153), .Z(n5155) );
  XOR U3535 ( .A(n4591), .B(n4590), .Z(n4560) );
  XOR U3536 ( .A(n4213), .B(n4212), .Z(n4219) );
  XOR U3537 ( .A(n5162), .B(n5161), .Z(n5110) );
  XOR U3538 ( .A(n5326), .B(n5325), .Z(n5327) );
  XOR U3539 ( .A(n5320), .B(n5319), .Z(n5322) );
  XOR U3540 ( .A(n4463), .B(n4462), .Z(n4464) );
  XOR U3541 ( .A(n5476), .B(n5475), .Z(n5477) );
  XOR U3542 ( .A(n5009), .B(n5008), .Z(n5011) );
  XOR U3543 ( .A(n4346), .B(n4345), .Z(n4347) );
  XOR U3544 ( .A(n4104), .B(n4103), .Z(n4105) );
  XOR U3545 ( .A(n5418), .B(n5417), .Z(n5420) );
  XOR U3546 ( .A(n5771), .B(n5770), .Z(n5815) );
  XOR U3547 ( .A(n5805), .B(n5804), .Z(n5775) );
  XOR U3548 ( .A(n5590), .B(n5589), .Z(n5591) );
  XOR U3549 ( .A(n5262), .B(n5261), .Z(n5263) );
  XOR U3550 ( .A(n5015), .B(n5014), .Z(n5016) );
  XOR U3551 ( .A(n4733), .B(n4732), .Z(n4739) );
  XOR U3552 ( .A(n4597), .B(n4596), .Z(n4556) );
  XOR U3553 ( .A(n5827), .B(n5826), .Z(n5828) );
  XOR U3554 ( .A(n4819), .B(n4818), .Z(n4874) );
  XOR U3555 ( .A(n4226), .B(n4225), .Z(n4227) );
  XOR U3556 ( .A(n4018), .B(n4017), .Z(n4020) );
  XOR U3557 ( .A(n5751), .B(n5750), .Z(n5753) );
  XOR U3558 ( .A(n5987), .B(n5986), .Z(n5989) );
  XOR U3559 ( .A(n5917), .B(n5916), .Z(n5918) );
  XOR U3560 ( .A(n5572), .B(n5571), .Z(n5573) );
  XOR U3561 ( .A(n5172), .B(n5171), .Z(n5173) );
  XOR U3562 ( .A(n4435), .B(n4434), .Z(n4436) );
  XOR U3563 ( .A(n4002), .B(n4001), .Z(n4004) );
  XOR U3564 ( .A(n6343), .B(n6342), .Z(n6373) );
  XOR U3565 ( .A(n6169), .B(n6168), .Z(n6139) );
  XOR U3566 ( .A(n6191), .B(n6190), .Z(n6193) );
  XOR U3567 ( .A(n6335), .B(n6334), .Z(n6337) );
  XNOR U3568 ( .A(n6546), .B(n6545), .Z(n6548) );
  XOR U3569 ( .A(n5911), .B(n5910), .Z(n5912) );
  XOR U3570 ( .A(n5739), .B(n16637), .Z(n5741) );
  XOR U3571 ( .A(n5496), .B(n5495), .Z(n5407) );
  XOR U3572 ( .A(n4549), .B(n4548), .Z(n4550) );
  XOR U3573 ( .A(n4475), .B(n4474), .Z(n4476) );
  XOR U3574 ( .A(n4354), .B(n4353), .Z(n4314) );
  XOR U3575 ( .A(n3826), .B(n3825), .Z(n3832) );
  XOR U3576 ( .A(n6109), .B(n6108), .Z(n6111) );
  XOR U3577 ( .A(n6415), .B(n6414), .Z(n6421) );
  XOR U3578 ( .A(n6576), .B(n6575), .Z(n6578) );
  XOR U3579 ( .A(n4687), .B(n4686), .Z(n4678) );
  XOR U3580 ( .A(n6594), .B(n6593), .Z(n6595) );
  XOR U3581 ( .A(n5250), .B(n5249), .Z(n5251) );
  XOR U3582 ( .A(n4951), .B(n4950), .Z(n4953) );
  XOR U3583 ( .A(n4238), .B(n4237), .Z(n4239) );
  XOR U3584 ( .A(n3817), .B(n3816), .Z(n3819) );
  XOR U3585 ( .A(n6481), .B(n6480), .Z(n6483) );
  XOR U3586 ( .A(n6666), .B(n6665), .Z(n6667) );
  XOR U3587 ( .A(n6964), .B(n6963), .Z(n6966) );
  XNOR U3588 ( .A(n7169), .B(n7168), .Z(n7201) );
  XNOR U3589 ( .A(n7189), .B(n7188), .Z(n7191) );
  XOR U3590 ( .A(n6475), .B(n6474), .Z(n6477) );
  XOR U3591 ( .A(n6293), .B(n6292), .Z(n6294) );
  XOR U3592 ( .A(n6217), .B(n6216), .Z(n6092) );
  XOR U3593 ( .A(n5568), .B(n5567), .Z(n5668) );
  XOR U3594 ( .A(n5338), .B(n5337), .Z(n5339) );
  XOR U3595 ( .A(n5027), .B(n5026), .Z(n5028) );
  XOR U3596 ( .A(n4244), .B(n4243), .Z(n4245) );
  XOR U3597 ( .A(n4030), .B(n4029), .Z(n4031) );
  XOR U3598 ( .A(n7017), .B(n7016), .Z(n7018) );
  XNOR U3599 ( .A(n6896), .B(n6895), .Z(n7012) );
  XNOR U3600 ( .A(n7383), .B(n7382), .Z(n7387) );
  XOR U3601 ( .A(n4489), .B(n4488), .Z(n4492) );
  XOR U3602 ( .A(n4308), .B(n4307), .Z(n4363) );
  XOR U3603 ( .A(n3905), .B(n3904), .Z(n3936) );
  XOR U3604 ( .A(n3595), .B(n3594), .Z(n3598) );
  XOR U3605 ( .A(n3681), .B(n3680), .Z(n3682) );
  XOR U3606 ( .A(n7025), .B(n7024), .Z(n6878) );
  XNOR U3607 ( .A(n7399), .B(n7398), .Z(n7401) );
  XOR U3608 ( .A(n7611), .B(n7610), .Z(n7655) );
  XOR U3609 ( .A(n5905), .B(n5904), .Z(n5906) );
  XOR U3610 ( .A(n5506), .B(n5505), .Z(n5507) );
  XOR U3611 ( .A(n5184), .B(n5183), .Z(n5186) );
  XOR U3612 ( .A(n4887), .B(n4886), .Z(n4889) );
  XOR U3613 ( .A(n4613), .B(n4612), .Z(n4614) );
  XOR U3614 ( .A(n7237), .B(n7236), .Z(n7238) );
  XOR U3615 ( .A(n7459), .B(n7458), .Z(n7461) );
  XOR U3616 ( .A(n7249), .B(n7248), .Z(n7250) );
  XOR U3617 ( .A(n6814), .B(n6813), .Z(n6815) );
  XOR U3618 ( .A(n6029), .B(n6028), .Z(n6030) );
  XOR U3619 ( .A(n4140), .B(n4139), .Z(n4088) );
  XOR U3620 ( .A(n3845), .B(n3844), .Z(n3846) );
  XOR U3621 ( .A(n3526), .B(n3525), .Z(n3532) );
  XOR U3622 ( .A(n7243), .B(n7242), .Z(n7244) );
  XOR U3623 ( .A(n7305), .B(n7304), .Z(n7307) );
  XNOR U3624 ( .A(n7871), .B(n7870), .Z(n7873) );
  XOR U3625 ( .A(n8075), .B(n8074), .Z(n8045) );
  XOR U3626 ( .A(n4194), .B(n4193), .Z(n4249) );
  XOR U3627 ( .A(n3471), .B(n3470), .Z(n3474) );
  XOR U3628 ( .A(n7925), .B(n7924), .Z(n7926) );
  XOR U3629 ( .A(n8103), .B(n8102), .Z(n8105) );
  XNOR U3630 ( .A(n7791), .B(n7790), .Z(n7907) );
  XOR U3631 ( .A(n8311), .B(n8310), .Z(n8305) );
  XOR U3632 ( .A(n7477), .B(n7476), .Z(n7478) );
  XOR U3633 ( .A(n7035), .B(n7034), .Z(n7037) );
  XOR U3634 ( .A(n6275), .B(n6274), .Z(n6276) );
  XOR U3635 ( .A(n5678), .B(n5677), .Z(n5679) );
  XOR U3636 ( .A(n4743), .B(n4742), .Z(n4744) );
  XOR U3637 ( .A(n4429), .B(n4428), .Z(n4431) );
  XOR U3638 ( .A(n4370), .B(n4369), .Z(n4371) );
  XOR U3639 ( .A(n4042), .B(n4041), .Z(n4044) );
  XOR U3640 ( .A(n3689), .B(n3688), .Z(n3692) );
  XOR U3641 ( .A(n7545), .B(n7544), .Z(n7705) );
  XOR U3642 ( .A(n7525), .B(n7524), .Z(n7526) );
  XOR U3643 ( .A(n7937), .B(n7936), .Z(n7939) );
  XOR U3644 ( .A(n8153), .B(n8152), .Z(n8159) );
  XOR U3645 ( .A(n7945), .B(n7944), .Z(n7748) );
  XOR U3646 ( .A(n7293), .B(n7292), .Z(n7295) );
  XOR U3647 ( .A(n6035), .B(n6034), .Z(n6036) );
  XOR U3648 ( .A(n5722), .B(n5721), .Z(n5724) );
  XOR U3649 ( .A(n5350), .B(n5349), .Z(n5351) );
  XOR U3650 ( .A(n5079), .B(n5078), .Z(n5081) );
  XOR U3651 ( .A(n4749), .B(n4748), .Z(n4750) );
  XOR U3652 ( .A(n4531), .B(n4530), .Z(n4533) );
  XOR U3653 ( .A(n4294), .B(n4293), .Z(n4296) );
  XOR U3654 ( .A(n4146), .B(n4145), .Z(n4081) );
  XOR U3655 ( .A(n3945), .B(n3944), .Z(n3893) );
  XOR U3656 ( .A(n3613), .B(n3612), .Z(n3582) );
  XOR U3657 ( .A(n7993), .B(n7992), .Z(n7987) );
  XNOR U3658 ( .A(n8257), .B(n8256), .Z(n8409) );
  XOR U3659 ( .A(n8529), .B(n8528), .Z(n8641) );
  XNOR U3660 ( .A(n8609), .B(n8608), .Z(n8611) );
  XNOR U3661 ( .A(n8813), .B(n8812), .Z(n8887) );
  XOR U3662 ( .A(n9072), .B(n9071), .Z(n9074) );
  XOR U3663 ( .A(n8829), .B(n8828), .Z(n8831) );
  XNOR U3664 ( .A(n6465), .B(n6464), .Z(n6624) );
  XNOR U3665 ( .A(n4795), .B(n4794), .Z(n4899) );
  XOR U3666 ( .A(n3426), .B(n3425), .Z(n3427) );
  XOR U3667 ( .A(n7999), .B(n7998), .Z(n8171) );
  XOR U3668 ( .A(n8427), .B(n8426), .Z(n8429) );
  XOR U3669 ( .A(n9066), .B(n9065), .Z(n9068) );
  XOR U3670 ( .A(n6233), .B(n6232), .Z(n6235) );
  XOR U3671 ( .A(n3857), .B(n3856), .Z(n3859) );
  XOR U3672 ( .A(n3410), .B(n3409), .Z(n3412) );
  XOR U3673 ( .A(n9044), .B(n9043), .Z(n9143) );
  XOR U3674 ( .A(n9020), .B(n9019), .Z(n9156) );
  XOR U3675 ( .A(n9585), .B(n9584), .Z(n9587) );
  XOR U3676 ( .A(n8441), .B(n8440), .Z(n8220) );
  XOR U3677 ( .A(n7521), .B(n7520), .Z(n7717) );
  XOR U3678 ( .A(n7261), .B(n7260), .Z(n7262) );
  XOR U3679 ( .A(n6858), .B(n6857), .Z(n6859) );
  XOR U3680 ( .A(n6662), .B(n6661), .Z(n6656) );
  XOR U3681 ( .A(n6427), .B(n6426), .Z(n6433) );
  XOR U3682 ( .A(n5556), .B(n5555), .Z(n5692) );
  XOR U3683 ( .A(n5520), .B(n5519), .Z(n5383) );
  XOR U3684 ( .A(n4935), .B(n4934), .Z(n5047) );
  XOR U3685 ( .A(n4761), .B(n4760), .Z(n4762) );
  XOR U3686 ( .A(n4425), .B(n4424), .Z(n4513) );
  XOR U3687 ( .A(n4288), .B(n4287), .Z(n4290) );
  XNOR U3688 ( .A(n4188), .B(n4187), .Z(n4263) );
  XOR U3689 ( .A(n3992), .B(n3991), .Z(n3986) );
  XOR U3690 ( .A(n3863), .B(n3862), .Z(n3864) );
  XOR U3691 ( .A(n3661), .B(n3660), .Z(n3701) );
  XOR U3692 ( .A(n3545), .B(n3544), .Z(n3546) );
  XOR U3693 ( .A(n3459), .B(n3458), .Z(n3460) );
  XOR U3694 ( .A(n3273), .B(n3272), .Z(n3279) );
  XOR U3695 ( .A(n8493), .B(n8492), .Z(n8677) );
  XOR U3696 ( .A(n8940), .B(n8939), .Z(n8941) );
  XOR U3697 ( .A(n9186), .B(n9185), .Z(n9192) );
  XOR U3698 ( .A(n9661), .B(n9660), .Z(n9663) );
  XNOR U3699 ( .A(n9597), .B(n9596), .Z(n9599) );
  XOR U3700 ( .A(n3721), .B(n3720), .Z(n3776) );
  XOR U3701 ( .A(n3233), .B(n3234), .Z(n3236) );
  XNOR U3702 ( .A(n8747), .B(n8746), .Z(n8934) );
  XOR U3703 ( .A(n8952), .B(n8951), .Z(n8953) );
  XOR U3704 ( .A(n9214), .B(n9213), .Z(n9215) );
  XOR U3705 ( .A(n9539), .B(n9538), .Z(n9687) );
  XOR U3706 ( .A(n9655), .B(n9654), .Z(n9657) );
  XNOR U3707 ( .A(n9675), .B(n9674), .Z(n9543) );
  XOR U3708 ( .A(n9897), .B(n9896), .Z(n9899) );
  XOR U3709 ( .A(n10195), .B(n10194), .Z(n10196) );
  XOR U3710 ( .A(n8721), .B(n8720), .Z(n8723) );
  XOR U3711 ( .A(n7979), .B(n7978), .Z(n7980) );
  XOR U3712 ( .A(n7489), .B(n7488), .Z(n7490) );
  XOR U3713 ( .A(n5887), .B(n5886), .Z(n5888) );
  XOR U3714 ( .A(n5226), .B(n5225), .Z(n5227) );
  XOR U3715 ( .A(n4905), .B(n4904), .Z(n4906) );
  XOR U3716 ( .A(n4631), .B(n4630), .Z(n4633) );
  XOR U3717 ( .A(n4156), .B(n4155), .Z(n4157) );
  XOR U3718 ( .A(n3954), .B(n3953), .Z(n3955) );
  XOR U3719 ( .A(n3623), .B(n3622), .Z(n3624) );
  XOR U3720 ( .A(n9208), .B(n9207), .Z(n9209) );
  XNOR U3721 ( .A(n9266), .B(n9265), .Z(n9477) );
  XOR U3722 ( .A(n9527), .B(n9526), .Z(n9699) );
  XOR U3723 ( .A(n9232), .B(n9231), .Z(n9233) );
  XOR U3724 ( .A(n8199), .B(n8198), .Z(n8200) );
  XOR U3725 ( .A(n6437), .B(n6436), .Z(n6438) );
  XOR U3726 ( .A(n6047), .B(n6046), .Z(n6048) );
  XOR U3727 ( .A(n5710), .B(n5709), .Z(n5712) );
  XOR U3728 ( .A(n5376), .B(n5375), .Z(n5378) );
  XOR U3729 ( .A(n5362), .B(n5361), .Z(n5363) );
  XOR U3730 ( .A(n3438), .B(n3437), .Z(n3439) );
  XOR U3731 ( .A(n3285), .B(n3286), .Z(n3349) );
  XOR U3732 ( .A(n3247), .B(n3248), .Z(n3250) );
  XOR U3733 ( .A(n9489), .B(n9488), .Z(n9491) );
  XOR U3734 ( .A(n9827), .B(n9826), .Z(n10026) );
  XOR U3735 ( .A(n10149), .B(n10148), .Z(n10272) );
  XOR U3736 ( .A(n10137), .B(n10136), .Z(n10130) );
  XOR U3737 ( .A(n10476), .B(n10475), .Z(n10478) );
  XOR U3738 ( .A(n10822), .B(n10821), .Z(n10823) );
  XNOR U3739 ( .A(n11100), .B(n11099), .Z(n11102) );
  XOR U3740 ( .A(n11112), .B(n11111), .Z(n11114) );
  XOR U3741 ( .A(n10546), .B(n10545), .Z(n10548) );
  XOR U3742 ( .A(n9246), .B(n9245), .Z(n9247) );
  XNOR U3743 ( .A(n6069), .B(n6068), .Z(n6245) );
  XOR U3744 ( .A(n3325), .B(n3326), .Z(n3328) );
  XOR U3745 ( .A(n9753), .B(n9752), .Z(n9759) );
  XOR U3746 ( .A(n9801), .B(n9800), .Z(n9802) );
  XOR U3747 ( .A(n10095), .B(n10094), .Z(n10303) );
  XOR U3748 ( .A(n10854), .B(n10853), .Z(n10858) );
  XOR U3749 ( .A(n10764), .B(n10763), .Z(n10766) );
  XOR U3750 ( .A(n10846), .B(n10845), .Z(n10848) );
  XOR U3751 ( .A(n8461), .B(n8460), .Z(n8462) );
  XOR U3752 ( .A(n7507), .B(n7506), .Z(n7508) );
  XOR U3753 ( .A(n7065), .B(n7064), .Z(n7066) );
  XOR U3754 ( .A(n6648), .B(n6647), .Z(n6649) );
  XOR U3755 ( .A(n5208), .B(n5207), .Z(n5209) );
  XOR U3756 ( .A(n4921), .B(n4920), .Z(n4922) );
  XOR U3757 ( .A(n4387), .B(n4386), .Z(n4388) );
  XOR U3758 ( .A(n4174), .B(n4173), .Z(n4175) );
  XOR U3759 ( .A(n3641), .B(n3640), .Z(n3642) );
  XOR U3760 ( .A(n3557), .B(n3556), .Z(n3559) );
  XOR U3761 ( .A(n3339), .B(n3340), .Z(n3381) );
  XOR U3762 ( .A(n3343), .B(n3344), .Z(n3346) );
  XOR U3763 ( .A(n9807), .B(n9806), .Z(n9808) );
  XOR U3764 ( .A(n10056), .B(n10055), .Z(n10057) );
  XOR U3765 ( .A(n10321), .B(n10320), .Z(n10327) );
  XOR U3766 ( .A(n11386), .B(n11385), .Z(n11388) );
  XOR U3767 ( .A(n11739), .B(n11738), .Z(n11741) );
  XOR U3768 ( .A(n8976), .B(n8975), .Z(n8977) );
  XOR U3769 ( .A(n8705), .B(n8704), .Z(n8706) );
  XOR U3770 ( .A(n8205), .B(n8204), .Z(n8206) );
  XOR U3771 ( .A(n7963), .B(n7962), .Z(n12460) );
  XOR U3772 ( .A(n7273), .B(n7272), .Z(n7274) );
  XOR U3773 ( .A(n6844), .B(n6843), .Z(n6845) );
  XOR U3774 ( .A(n6254), .B(n6255), .Z(n12425) );
  XOR U3775 ( .A(n5544), .B(n5543), .Z(n5704) );
  XOR U3776 ( .A(n4651), .B(n4650), .Z(n4775) );
  XOR U3777 ( .A(n4407), .B(n4406), .Z(n4401) );
  XOR U3778 ( .A(n4171), .B(n4172), .Z(n12345) );
  XOR U3779 ( .A(n3974), .B(n3973), .Z(n4062) );
  XOR U3780 ( .A(n3874), .B(n3875), .Z(n12230) );
  XOR U3781 ( .A(n3795), .B(n3794), .Z(n3871) );
  XOR U3782 ( .A(n3705), .B(n3704), .Z(n3706) );
  XOR U3783 ( .A(n3508), .B(n3509), .Z(n12299) );
  XOR U3784 ( .A(n3501), .B(n3500), .Z(n12232) );
  XOR U3785 ( .A(n3365), .B(n3366), .Z(n3368) );
  XOR U3786 ( .A(n10351), .B(n10350), .Z(n10357) );
  XNOR U3787 ( .A(n12023), .B(n12022), .Z(n12025) );
  XOR U3788 ( .A(n10075), .B(n10074), .Z(n10076) );
  XNOR U3789 ( .A(n12223), .B(n12224), .Z(n12485) );
  XOR U3790 ( .A(n12241), .B(n12242), .Z(n12244) );
  XOR U3791 ( .A(n10363), .B(n10362), .Z(n10364) );
  XNOR U3792 ( .A(n10395), .B(n10394), .Z(n10618) );
  XOR U3793 ( .A(n11012), .B(n11011), .Z(n11212) );
  XOR U3794 ( .A(n11506), .B(n11505), .Z(n11511) );
  XOR U3795 ( .A(n12011), .B(n12010), .Z(n12013) );
  XOR U3796 ( .A(n11691), .B(n11690), .Z(n11693) );
  XOR U3797 ( .A(n12861), .B(n12860), .Z(n12857) );
  XOR U3798 ( .A(n12838), .B(n12839), .Z(n12837) );
  XOR U3799 ( .A(n10638), .B(n10637), .Z(n10370) );
  XOR U3800 ( .A(n12508), .B(n12509), .Z(n13418) );
  XOR U3801 ( .A(n12496), .B(n12497), .Z(n13403) );
  XOR U3802 ( .A(n12474), .B(n12475), .Z(n13381) );
  XOR U3803 ( .A(n12450), .B(n12451), .Z(n13357) );
  XOR U3804 ( .A(n12438), .B(n12439), .Z(n13345) );
  XOR U3805 ( .A(n12414), .B(n12415), .Z(n13321) );
  XOR U3806 ( .A(n5880), .B(n5881), .Z(n12409) );
  XOR U3807 ( .A(n12404), .B(n12405), .Z(n13309) );
  XOR U3808 ( .A(n5213), .B(n5214), .Z(n12385) );
  XOR U3809 ( .A(n12368), .B(n12369), .Z(n13273) );
  XOR U3810 ( .A(n12356), .B(n12357), .Z(n13261) );
  XOR U3811 ( .A(n12312), .B(n12313), .Z(n13213) );
  XOR U3812 ( .A(n12255), .B(n12256), .Z(n13155) );
  XOR U3813 ( .A(n12259), .B(n12260), .Z(n12262) );
  XOR U3814 ( .A(n10948), .B(n10947), .Z(n10949) );
  XOR U3815 ( .A(n11322), .B(n11321), .Z(n11530) );
  XOR U3816 ( .A(n11975), .B(n11974), .Z(n11977) );
  XOR U3817 ( .A(n12875), .B(n12874), .Z(n12873) );
  XOR U3818 ( .A(n12893), .B(n12892), .Z(n12891) );
  XOR U3819 ( .A(n12520), .B(n12521), .Z(n13431) );
  XOR U3820 ( .A(n12454), .B(n12455), .Z(n13361) );
  XOR U3821 ( .A(n13354), .B(n13355), .Z(n13707) );
  XOR U3822 ( .A(n12418), .B(n12419), .Z(n13325) );
  XOR U3823 ( .A(n13318), .B(n13319), .Z(n13671) );
  XOR U3824 ( .A(n13306), .B(n13307), .Z(n13659) );
  XOR U3825 ( .A(n13294), .B(n13295), .Z(n13647) );
  XOR U3826 ( .A(n12372), .B(n12373), .Z(n13277) );
  XOR U3827 ( .A(n13270), .B(n13271), .Z(n13623) );
  XOR U3828 ( .A(n13258), .B(n13259), .Z(n13611) );
  XOR U3829 ( .A(n13248), .B(n13249), .Z(n13472) );
  XOR U3830 ( .A(n12338), .B(n12339), .Z(n13241) );
  XOR U3831 ( .A(n13234), .B(n13235), .Z(n13589) );
  XOR U3832 ( .A(n12328), .B(n12329), .Z(n13228) );
  XOR U3833 ( .A(n13224), .B(n13225), .Z(n13474) );
  XOR U3834 ( .A(n13210), .B(n13211), .Z(n13567) );
  XOR U3835 ( .A(n13198), .B(n13199), .Z(n13555) );
  XOR U3836 ( .A(n12292), .B(n12293), .Z(n13127) );
  XOR U3837 ( .A(n12270), .B(n12271), .Z(n13129) );
  XOR U3838 ( .A(n13166), .B(n13167), .Z(n13521) );
  XNOR U3839 ( .A(n10970), .B(n10969), .Z(n11254) );
  XOR U3840 ( .A(n12130), .B(n12129), .Z(n12136) );
  XOR U3841 ( .A(n13542), .B(n13543), .Z(n13545) );
  XOR U3842 ( .A(n13151), .B(n13152), .Z(n13503) );
  XOR U3843 ( .A(n13142), .B(n13143), .Z(n13493) );
  XOR U3844 ( .A(n13484), .B(n13485), .Z(n13487) );
  XOR U3845 ( .A(n11576), .B(n11575), .Z(n11577) );
  XNOR U3846 ( .A(n11604), .B(n11603), .Z(n11875) );
  XOR U3847 ( .A(n11935), .B(n11934), .Z(n12154) );
  XNOR U3848 ( .A(n12971), .B(n12970), .Z(n12969) );
  XOR U3849 ( .A(n12533), .B(n12534), .Z(n13445) );
  XOR U3850 ( .A(n13423), .B(n13424), .Z(n13771) );
  XOR U3851 ( .A(n13398), .B(n13399), .Z(n13749) );
  XOR U3852 ( .A(n13744), .B(n13745), .Z(n14105) );
  XOR U3853 ( .A(n13374), .B(n13375), .Z(n13724) );
  XOR U3854 ( .A(n13636), .B(n13637), .Z(n13995) );
  XOR U3855 ( .A(n13184), .B(n13185), .Z(n13536) );
  XOR U3856 ( .A(n13498), .B(n13499), .Z(n13855) );
  XOR U3857 ( .A(n13454), .B(n13455), .Z(n13799) );
  XNOR U3858 ( .A(n11586), .B(n11585), .Z(n11893) );
  XOR U3859 ( .A(n14138), .B(n14139), .Z(n14499) );
  XOR U3860 ( .A(n14114), .B(n14115), .Z(n14475) );
  XOR U3861 ( .A(n14092), .B(n14093), .Z(n14179) );
  XOR U3862 ( .A(n13726), .B(n13727), .Z(n14084) );
  XOR U3863 ( .A(n14080), .B(n14081), .Z(n14440) );
  XOR U3864 ( .A(n13700), .B(n13701), .Z(n14061) );
  XOR U3865 ( .A(n14054), .B(n14055), .Z(n14417) );
  XOR U3866 ( .A(n13688), .B(n13689), .Z(n14049) );
  XOR U3867 ( .A(n14042), .B(n14043), .Z(n14405) );
  XOR U3868 ( .A(n13664), .B(n13665), .Z(n14025) );
  XOR U3869 ( .A(n14018), .B(n14019), .Z(n14381) );
  XOR U3870 ( .A(n13652), .B(n13653), .Z(n14013) );
  XOR U3871 ( .A(n14008), .B(n14009), .Z(n14368) );
  XOR U3872 ( .A(n13640), .B(n13641), .Z(n14001) );
  XOR U3873 ( .A(n13616), .B(n13617), .Z(n13977) );
  XOR U3874 ( .A(n13970), .B(n13971), .Z(n14335) );
  XOR U3875 ( .A(n13606), .B(n13607), .Z(n13964) );
  XOR U3876 ( .A(n13584), .B(n13585), .Z(n13940) );
  XOR U3877 ( .A(n13934), .B(n13935), .Z(n14301) );
  XOR U3878 ( .A(n13572), .B(n13573), .Z(n13929) );
  XOR U3879 ( .A(n13924), .B(n13925), .Z(n14288) );
  XOR U3880 ( .A(n13562), .B(n13563), .Z(n13916) );
  XOR U3881 ( .A(n13538), .B(n13539), .Z(n13826) );
  XOR U3882 ( .A(n13878), .B(n13879), .Z(n14186) );
  XOR U3883 ( .A(n13514), .B(n13515), .Z(n13829) );
  XOR U3884 ( .A(n13866), .B(n13867), .Z(n14233) );
  XOR U3885 ( .A(n13806), .B(n13807), .Z(n14168) );
  XOR U3886 ( .A(n11911), .B(n11910), .Z(n12214) );
  XOR U3887 ( .A(n12572), .B(n12571), .Z(n13073) );
  XOR U3888 ( .A(n13882), .B(n13883), .Z(n13885) );
  XOR U3889 ( .A(n13839), .B(n13840), .Z(n13842) );
  XNOR U3890 ( .A(n13815), .B(n13814), .Z(n13811) );
  XOR U3891 ( .A(n12549), .B(n12550), .Z(n13462) );
  XOR U3892 ( .A(n14074), .B(n14075), .Z(n14435) );
  XOR U3893 ( .A(n14038), .B(n14039), .Z(n14399) );
  XOR U3894 ( .A(n13990), .B(n13991), .Z(n14353) );
  XOR U3895 ( .A(n13954), .B(n13955), .Z(n14319) );
  XOR U3896 ( .A(n13906), .B(n13907), .Z(n14273) );
  XOR U3897 ( .A(n13862), .B(n13863), .Z(n14227) );
  XOR U3898 ( .A(n14214), .B(n14215), .Z(n14217) );
  XOR U3899 ( .A(n14516), .B(n14517), .Z(n14881) );
  XOR U3900 ( .A(n14492), .B(n14493), .Z(n14861) );
  XOR U3901 ( .A(n14468), .B(n14469), .Z(n14841) );
  XOR U3902 ( .A(n14436), .B(n14437), .Z(n14810) );
  XOR U3903 ( .A(n14424), .B(n14425), .Z(n14800) );
  XOR U3904 ( .A(n14400), .B(n14401), .Z(n14780) );
  XOR U3905 ( .A(n14364), .B(n14365), .Z(n14750) );
  XOR U3906 ( .A(n14354), .B(n14355), .Z(n14740) );
  XOR U3907 ( .A(n14330), .B(n14331), .Z(n14720) );
  XOR U3908 ( .A(n14320), .B(n14321), .Z(n14710) );
  XOR U3909 ( .A(n14284), .B(n14285), .Z(n14680) );
  XOR U3910 ( .A(n14274), .B(n14275), .Z(n14670) );
  XOR U3911 ( .A(n14228), .B(n14229), .Z(n14628) );
  XOR U3912 ( .A(n14895), .B(n14894), .Z(n14960) );
  XOR U3913 ( .A(n14884), .B(n14885), .Z(n15036) );
  XOR U3914 ( .A(n14874), .B(n14875), .Z(n15112) );
  XOR U3915 ( .A(n14864), .B(n14865), .Z(n15188) );
  XOR U3916 ( .A(n14854), .B(n14855), .Z(n15264) );
  XOR U3917 ( .A(n14844), .B(n14845), .Z(n15340) );
  XOR U3918 ( .A(n14834), .B(n14835), .Z(n15416) );
  XOR U3919 ( .A(n14824), .B(n14825), .Z(n15492) );
  XOR U3920 ( .A(n14814), .B(n14815), .Z(n15568) );
  XOR U3921 ( .A(n14804), .B(n14805), .Z(n15644) );
  XOR U3922 ( .A(n14794), .B(n14795), .Z(n15720) );
  XOR U3923 ( .A(n14784), .B(n14785), .Z(n15796) );
  XOR U3924 ( .A(n14774), .B(n14775), .Z(n15872) );
  XOR U3925 ( .A(n14764), .B(n14765), .Z(n15947) );
  XOR U3926 ( .A(n14754), .B(n14755), .Z(n16023) );
  XOR U3927 ( .A(n14744), .B(n14745), .Z(n16099) );
  XOR U3928 ( .A(n14734), .B(n14735), .Z(n16176) );
  XOR U3929 ( .A(n14724), .B(n14725), .Z(n16253) );
  XOR U3930 ( .A(n14714), .B(n14715), .Z(n16331) );
  XOR U3931 ( .A(n14704), .B(n14705), .Z(n16408) );
  XOR U3932 ( .A(n14694), .B(n14695), .Z(n16484) );
  XOR U3933 ( .A(n14684), .B(n14685), .Z(n16562) );
  XOR U3934 ( .A(n14674), .B(n14675), .Z(n16639) );
  XOR U3935 ( .A(n14664), .B(n14665), .Z(n16716) );
  XOR U3936 ( .A(n14654), .B(n14655), .Z(n16792) );
  XOR U3937 ( .A(n14644), .B(n14645), .Z(n16870) );
  XOR U3938 ( .A(n14632), .B(n14633), .Z(n16947) );
  XOR U3939 ( .A(n14622), .B(n14623), .Z(n17024) );
  XOR U3940 ( .A(n14610), .B(n14611), .Z(n17101) );
  XOR U3941 ( .A(n14600), .B(n14601), .Z(n17179) );
  XOR U3942 ( .A(n4713), .B(n4712), .Z(n4714) );
  XOR U3943 ( .A(n4697), .B(n4696), .Z(n4699) );
  XOR U3944 ( .A(n4835), .B(n4834), .Z(n4836) );
  XOR U3945 ( .A(n4831), .B(n4830), .Z(n4862) );
  XOR U3946 ( .A(n4457), .B(n4456), .Z(n4458) );
  XOR U3947 ( .A(n4985), .B(n4984), .Z(n4986) );
  XOR U3948 ( .A(n4993), .B(n4992), .Z(n4996) );
  XOR U3949 ( .A(n4441), .B(n4440), .Z(n4443) );
  XOR U3950 ( .A(n5128), .B(n5127), .Z(n5144) );
  XOR U3951 ( .A(n5114), .B(n5113), .Z(n5116) );
  XOR U3952 ( .A(n4965), .B(n4964), .Z(n5005) );
  XOR U3953 ( .A(n4725), .B(n4724), .Z(n4726) );
  XOR U3954 ( .A(n4561), .B(n4560), .Z(n4562) );
  XOR U3955 ( .A(n5274), .B(n5273), .Z(n5275) );
  XOR U3956 ( .A(n5314), .B(n5313), .Z(n5315) );
  XOR U3957 ( .A(n5444), .B(n5443), .Z(n5460) );
  XOR U3958 ( .A(n4220), .B(n4219), .Z(n4221) );
  XOR U3959 ( .A(n5328), .B(n5327), .Z(n5267) );
  XOR U3960 ( .A(n5478), .B(n5477), .Z(n5426) );
  XOR U3961 ( .A(n5166), .B(n5165), .Z(n5167) );
  XOR U3962 ( .A(n4869), .B(n4868), .Z(n4871) );
  XOR U3963 ( .A(n4204), .B(n4203), .Z(n4206) );
  XOR U3964 ( .A(n5642), .B(n5641), .Z(n5644) );
  XOR U3965 ( .A(n5490), .B(n5489), .Z(n5413) );
  XOR U3966 ( .A(n4469), .B(n4468), .Z(n4470) );
  XOR U3967 ( .A(n4011), .B(n4010), .Z(n4017) );
  XOR U3968 ( .A(n5578), .B(n5577), .Z(n5580) );
  XOR U3969 ( .A(n5745), .B(n5744), .Z(n5747) );
  XOR U3970 ( .A(n5833), .B(n5832), .Z(n5834) );
  XOR U3971 ( .A(n5821), .B(n5820), .Z(n5823) );
  XOR U3972 ( .A(n5943), .B(n5942), .Z(n5983) );
  XOR U3973 ( .A(n5757), .B(n5756), .Z(n5759) );
  XOR U3974 ( .A(n5017), .B(n5016), .Z(n4956) );
  XOR U3975 ( .A(n4320), .B(n4319), .Z(n4351) );
  XOR U3976 ( .A(n3921), .B(n3920), .Z(n3908) );
  XNOR U3977 ( .A(n5995), .B(n5994), .Z(n5935) );
  XOR U3978 ( .A(n6185), .B(n6184), .Z(n6187) );
  XOR U3979 ( .A(n5256), .B(n5255), .Z(n5257) );
  XOR U3980 ( .A(n4691), .B(n4690), .Z(n4693) );
  XOR U3981 ( .A(n4601), .B(n4600), .Z(n4602) );
  XOR U3982 ( .A(n5929), .B(n5928), .Z(n5930) );
  XOR U3983 ( .A(n6103), .B(n6102), .Z(n6105) );
  XOR U3984 ( .A(n6117), .B(n6116), .Z(n6197) );
  XOR U3985 ( .A(n6203), .B(n6202), .Z(n6205) );
  XOR U3986 ( .A(n5574), .B(n5573), .Z(n5662) );
  XOR U3987 ( .A(n5332), .B(n5331), .Z(n5333) );
  XOR U3988 ( .A(n5021), .B(n5020), .Z(n5022) );
  XOR U3989 ( .A(n4877), .B(n4876), .Z(n4812) );
  XOR U3990 ( .A(n4232), .B(n4231), .Z(n4233) );
  XOR U3991 ( .A(n6419), .B(n6418), .Z(n6420) );
  XOR U3992 ( .A(n6307), .B(n6306), .Z(n6409) );
  XOR U3993 ( .A(n6377), .B(n6376), .Z(n6379) );
  XNOR U3994 ( .A(n6331), .B(n6330), .Z(n6323) );
  XNOR U3995 ( .A(n6397), .B(n6396), .Z(n6311) );
  XOR U3996 ( .A(n4024), .B(n4023), .Z(n4025) );
  XOR U3997 ( .A(n3833), .B(n3832), .Z(n3834) );
  XOR U3998 ( .A(n6486), .B(n16560), .Z(n6487) );
  NANDN U3999 ( .A(n6556), .B(n6555), .Z(n2964) );
  NANDN U4000 ( .A(n6724), .B(n6554), .Z(n2965) );
  NAND U4001 ( .A(n2964), .B(n2965), .Z(n6729) );
  XOR U4002 ( .A(n6970), .B(n6969), .Z(n6971) );
  XOR U4003 ( .A(n6017), .B(n6016), .Z(n6018) );
  XOR U4004 ( .A(n5500), .B(n5499), .Z(n5501) );
  XOR U4005 ( .A(n5178), .B(n5177), .Z(n5179) );
  XOR U4006 ( .A(n4679), .B(n4678), .Z(n4680) );
  XOR U4007 ( .A(n4481), .B(n4480), .Z(n4483) );
  XOR U4008 ( .A(n4358), .B(n4357), .Z(n4360) );
  XOR U4009 ( .A(n4132), .B(n4131), .Z(n4133) );
  XOR U4010 ( .A(n3931), .B(n3930), .Z(n3932) );
  XOR U4011 ( .A(n3737), .B(n3736), .Z(n3738) );
  XOR U4012 ( .A(n6492), .B(n6491), .Z(n6494) );
  XOR U4013 ( .A(n6668), .B(n6667), .Z(n6792) );
  XNOR U4014 ( .A(n6768), .B(n6767), .Z(n6684) );
  XOR U4015 ( .A(n7201), .B(n7200), .Z(n7203) );
  XOR U4016 ( .A(n5847), .B(n5846), .Z(n5735) );
  XOR U4017 ( .A(n4805), .B(n4804), .Z(n4807) );
  XOR U4018 ( .A(n4673), .B(n4672), .Z(n4674) );
  XOR U4019 ( .A(n6606), .B(n6605), .Z(n6608) );
  XOR U4020 ( .A(n6888), .B(n6887), .Z(n6890) );
  XOR U4021 ( .A(n7006), .B(n7005), .Z(n7008) );
  XOR U4022 ( .A(n7012), .B(n7011), .Z(n7013) );
  XOR U4023 ( .A(n7133), .B(n7132), .Z(n7221) );
  XOR U4024 ( .A(n7195), .B(n7194), .Z(n7197) );
  XOR U4025 ( .A(n7387), .B(n7386), .Z(n7389) );
  XOR U4026 ( .A(n5029), .B(n5028), .Z(n5032) );
  XOR U4027 ( .A(n4545), .B(n4544), .Z(n4612) );
  XOR U4028 ( .A(n6876), .B(n6875), .Z(n6877) );
  XOR U4029 ( .A(n7209), .B(n7208), .Z(n7149) );
  XOR U4030 ( .A(n7633), .B(n7632), .Z(n7637) );
  XOR U4031 ( .A(n7861), .B(n7860), .Z(n7843) );
  XOR U4032 ( .A(n6287), .B(n6286), .Z(n6288) );
  XOR U4033 ( .A(n5560), .B(n5559), .Z(n5561) );
  XOR U4034 ( .A(n5244), .B(n5243), .Z(n5245) );
  XOR U4035 ( .A(n4198), .B(n4197), .Z(n4200) );
  XOR U4036 ( .A(n3996), .B(n3995), .Z(n3997) );
  XOR U4037 ( .A(n3841), .B(n3840), .Z(n3844) );
  XOR U4038 ( .A(n3599), .B(n3598), .Z(n3600) );
  XOR U4039 ( .A(n3683), .B(n3682), .Z(n3667) );
  XOR U4040 ( .A(n7023), .B(n7022), .Z(n7024) );
  XOR U4041 ( .A(n7599), .B(n7598), .Z(n7663) );
  XOR U4042 ( .A(n7649), .B(n7648), .Z(n7651) );
  XOR U4043 ( .A(n6810), .B(n6809), .Z(n6816) );
  XOR U4044 ( .A(n6469), .B(n6468), .Z(n6471) );
  XOR U4045 ( .A(n6281), .B(n6280), .Z(n6282) );
  XOR U4046 ( .A(n5907), .B(n5906), .Z(n6031) );
  XOR U4047 ( .A(n5344), .B(n5343), .Z(n5345) );
  XOR U4048 ( .A(n5085), .B(n5084), .Z(n5087) );
  XOR U4049 ( .A(n5039), .B(n5038), .Z(n5040) );
  XOR U4050 ( .A(n4537), .B(n4536), .Z(n4539) );
  XOR U4051 ( .A(n4495), .B(n4494), .Z(n4501) );
  XOR U4052 ( .A(n4366), .B(n4365), .Z(n4302) );
  XOR U4053 ( .A(n4036), .B(n4035), .Z(n4037) );
  XOR U4054 ( .A(n3897), .B(n3896), .Z(n3899) );
  XOR U4055 ( .A(n3731), .B(n3730), .Z(n3732) );
  XOR U4056 ( .A(n7239), .B(n7238), .Z(n7245) );
  XOR U4057 ( .A(n7551), .B(n7550), .Z(n7699) );
  XOR U4058 ( .A(n7563), .B(n7562), .Z(n7687) );
  XOR U4059 ( .A(n8097), .B(n8096), .Z(n8099) );
  XNOR U4060 ( .A(n5730), .B(n5729), .Z(n5857) );
  XOR U4061 ( .A(n4663), .B(n4662), .Z(n4742) );
  XOR U4062 ( .A(n3533), .B(n3532), .Z(n3535) );
  XNOR U4063 ( .A(n7313), .B(n7312), .Z(n7465) );
  XOR U4064 ( .A(n7473), .B(n7472), .Z(n7300) );
  XOR U4065 ( .A(n7537), .B(n7536), .Z(n7538) );
  XOR U4066 ( .A(n7771), .B(n7770), .Z(n7773) );
  XOR U4067 ( .A(n7907), .B(n7906), .Z(n7909) );
  XOR U4068 ( .A(n8129), .B(n8128), .Z(n8135) );
  XOR U4069 ( .A(n8039), .B(n8038), .Z(n8041) );
  XOR U4070 ( .A(n8363), .B(n8362), .Z(n8315) );
  XOR U4071 ( .A(n8581), .B(n8580), .Z(n8563) );
  XOR U4072 ( .A(n7083), .B(n7082), .Z(n7084) );
  XOR U4073 ( .A(n6227), .B(n6226), .Z(n6228) );
  XOR U4074 ( .A(n4250), .B(n4249), .Z(n4251) );
  XOR U4075 ( .A(n3475), .B(n3474), .Z(n3476) );
  XNOR U4076 ( .A(n8111), .B(n8110), .Z(n8027) );
  XOR U4077 ( .A(n8275), .B(n8274), .Z(n8391) );
  XNOR U4078 ( .A(n8621), .B(n8620), .Z(n8623) );
  XNOR U4079 ( .A(n8551), .B(n8550), .Z(n8553) );
  XOR U4080 ( .A(n8859), .B(n8858), .Z(n8841) );
  XOR U4081 ( .A(n7747), .B(n7746), .Z(n7749) );
  XOR U4082 ( .A(n7527), .B(n7526), .Z(n7711) );
  XOR U4083 ( .A(n7255), .B(n7254), .Z(n7256) );
  XOR U4084 ( .A(n6864), .B(n6863), .Z(n6866) );
  XOR U4085 ( .A(n6826), .B(n6825), .Z(n6827) );
  XOR U4086 ( .A(n5680), .B(n5679), .Z(n5686) );
  XOR U4087 ( .A(n5514), .B(n5513), .Z(n5389) );
  XOR U4088 ( .A(n4939), .B(n4938), .Z(n4940) );
  XOR U4089 ( .A(n4256), .B(n4255), .Z(n4257) );
  XOR U4090 ( .A(n3813), .B(n3812), .Z(n3853) );
  XOR U4091 ( .A(n3693), .B(n3692), .Z(n3694) );
  XOR U4092 ( .A(n3583), .B(n3582), .Z(n3584) );
  XOR U4093 ( .A(n3419), .B(n3418), .Z(n3425) );
  XOR U4094 ( .A(n7931), .B(n7930), .Z(n7933) );
  XOR U4095 ( .A(n7753), .B(n7752), .Z(n7755) );
  XOR U4096 ( .A(n7997), .B(n7996), .Z(n7998) );
  XOR U4097 ( .A(n7985), .B(n7984), .Z(n7986) );
  XOR U4098 ( .A(n8177), .B(n8176), .Z(n8183) );
  XOR U4099 ( .A(n8403), .B(n8402), .Z(n8405) );
  XOR U4100 ( .A(n8409), .B(n8408), .Z(n8411) );
  XOR U4101 ( .A(n8541), .B(n8540), .Z(n8629) );
  XOR U4102 ( .A(n8523), .B(n8522), .Z(n8647) );
  XOR U4103 ( .A(n8835), .B(n8834), .Z(n8837) );
  XOR U4104 ( .A(n4507), .B(n4506), .Z(n4422) );
  XOR U4105 ( .A(n4050), .B(n4049), .Z(n3989) );
  XOR U4106 ( .A(n8237), .B(n8236), .Z(n8238) );
  XOR U4107 ( .A(n8499), .B(n8498), .Z(n8671) );
  XOR U4108 ( .A(n8881), .B(n8880), .Z(n8883) );
  XOR U4109 ( .A(n9050), .B(n9049), .Z(n9136) );
  XOR U4110 ( .A(n9359), .B(n9358), .Z(n9361) );
  XNOR U4111 ( .A(n9060), .B(n9059), .Z(n9062) );
  XOR U4112 ( .A(n9341), .B(n9340), .Z(n9343) );
  XOR U4113 ( .A(n9124), .B(n9123), .Z(n9126) );
  XOR U4114 ( .A(n7483), .B(n7482), .Z(n7484) );
  XOR U4115 ( .A(n6425), .B(n6424), .Z(n6426) );
  XOR U4116 ( .A(n5232), .B(n5231), .Z(n5233) );
  XOR U4117 ( .A(n4755), .B(n4754), .Z(n4756) );
  XOR U4118 ( .A(n4625), .B(n4624), .Z(n4627) );
  XOR U4119 ( .A(n4375), .B(n4374), .Z(n4376) );
  XOR U4120 ( .A(n4150), .B(n4149), .Z(n4151) );
  XOR U4121 ( .A(n3949), .B(n3948), .Z(n3950) );
  XOR U4122 ( .A(n3771), .B(n3770), .Z(n3773) );
  XOR U4123 ( .A(n3541), .B(n3540), .Z(n3544) );
  XOR U4124 ( .A(n8421), .B(n8420), .Z(n8422) );
  XOR U4125 ( .A(n8231), .B(n8230), .Z(n8233) );
  XNOR U4126 ( .A(n8227), .B(n8226), .Z(n8439) );
  XOR U4127 ( .A(n8687), .B(n8686), .Z(n8688) );
  XOR U4128 ( .A(n8487), .B(n8486), .Z(n8683) );
  XOR U4129 ( .A(n9038), .B(n9037), .Z(n9032) );
  XOR U4130 ( .A(n8193), .B(n8192), .Z(n8194) );
  XOR U4131 ( .A(n6457), .B(n6456), .Z(n6459) );
  XOR U4132 ( .A(n5895), .B(n5894), .Z(n6043) );
  XOR U4133 ( .A(n5865), .B(n5864), .Z(n5717) );
  XOR U4134 ( .A(n5356), .B(n5355), .Z(n5357) );
  XOR U4135 ( .A(n3489), .B(n3488), .Z(n3458) );
  XOR U4136 ( .A(n3292), .B(n3291), .Z(n3308) );
  XOR U4137 ( .A(n8739), .B(n8738), .Z(n8741) );
  XOR U4138 ( .A(n9008), .B(n9007), .Z(n9180) );
  XOR U4139 ( .A(n9014), .B(n9013), .Z(n9162) );
  XOR U4140 ( .A(n9649), .B(n9648), .Z(n9650) );
  XNOR U4141 ( .A(n6860), .B(n6859), .Z(n7047) );
  XOR U4142 ( .A(n3865), .B(n3864), .Z(n3804) );
  XOR U4143 ( .A(n3432), .B(n3431), .Z(n3433) );
  XOR U4144 ( .A(n3280), .B(n3279), .Z(n3282) );
  XOR U4145 ( .A(n8934), .B(n8933), .Z(n8936) );
  XOR U4146 ( .A(n8733), .B(n8732), .Z(n8735) );
  XOR U4147 ( .A(n9210), .B(n9209), .Z(n9216) );
  XOR U4148 ( .A(n9278), .B(n9277), .Z(n9465) );
  XOR U4149 ( .A(n9290), .B(n9289), .Z(n9453) );
  XOR U4150 ( .A(n9563), .B(n9562), .Z(n9555) );
  XNOR U4151 ( .A(n9543), .B(n9542), .Z(n9545) );
  XOR U4152 ( .A(n9921), .B(n9920), .Z(n9922) );
  XOR U4153 ( .A(n10201), .B(n10200), .Z(n10203) );
  XOR U4154 ( .A(n8954), .B(n8953), .Z(n8722) );
  XOR U4155 ( .A(n8467), .B(n8466), .Z(n8468) );
  XOR U4156 ( .A(n7955), .B(n7954), .Z(n7956) );
  XOR U4157 ( .A(n7513), .B(n7512), .Z(n7514) );
  XOR U4158 ( .A(n6239), .B(n6238), .Z(n6241) );
  XOR U4159 ( .A(n5548), .B(n5547), .Z(n5549) );
  XOR U4160 ( .A(n5202), .B(n5201), .Z(n5203) );
  XOR U4161 ( .A(n4927), .B(n4926), .Z(n4928) );
  XOR U4162 ( .A(n4417), .B(n4416), .Z(n4418) );
  XOR U4163 ( .A(n4180), .B(n4179), .Z(n4181) );
  XOR U4164 ( .A(n3978), .B(n3977), .Z(n3980) );
  XOR U4165 ( .A(n3653), .B(n3652), .Z(n3655) );
  XOR U4166 ( .A(n3264), .B(n3263), .Z(n3265) );
  XOR U4167 ( .A(n9252), .B(n9251), .Z(n9254) );
  XOR U4168 ( .A(n9477), .B(n9476), .Z(n9479) );
  XOR U4169 ( .A(n9711), .B(n9710), .Z(n9717) );
  XOR U4170 ( .A(n9533), .B(n9532), .Z(n9693) );
  XNOR U4171 ( .A(n9891), .B(n9890), .Z(n9893) );
  XNOR U4172 ( .A(n10161), .B(n10160), .Z(n10155) );
  XOR U4173 ( .A(n10482), .B(n10481), .Z(n10484) );
  XNOR U4174 ( .A(n10464), .B(n10463), .Z(n10466) );
  XOR U4175 ( .A(n9228), .B(n9227), .Z(n9234) );
  XOR U4176 ( .A(n8699), .B(n8698), .Z(n8700) );
  XOR U4177 ( .A(n7073), .B(n7072), .Z(n7269) );
  XOR U4178 ( .A(n6834), .B(n6833), .Z(n6840) );
  XOR U4179 ( .A(n6451), .B(n6450), .Z(n6453) );
  XOR U4180 ( .A(n6265), .B(n6264), .Z(n6439) );
  XOR U4181 ( .A(n5696), .B(n5695), .Z(n5697) );
  XOR U4182 ( .A(n4657), .B(n4656), .Z(n4769) );
  XOR U4183 ( .A(n4411), .B(n4410), .Z(n4412) );
  XOR U4184 ( .A(n4282), .B(n4281), .Z(n4284) );
  XOR U4185 ( .A(n3799), .B(n3798), .Z(n3800) );
  XOR U4186 ( .A(n3713), .B(n3712), .Z(n3715) );
  XOR U4187 ( .A(n3571), .B(n3570), .Z(n3572) );
  XOR U4188 ( .A(n3513), .B(n3512), .Z(n3553) );
  XOR U4189 ( .A(n3495), .B(n3494), .Z(n3454) );
  XOR U4190 ( .A(n3253), .B(n3254), .Z(n3338) );
  XOR U4191 ( .A(n9240), .B(n9239), .Z(n9242) );
  XOR U4192 ( .A(n9258), .B(n9257), .Z(n9259) );
  XNOR U4193 ( .A(n9248), .B(n9247), .Z(n9495) );
  XOR U4194 ( .A(n10125), .B(n10124), .Z(n10285) );
  XOR U4195 ( .A(n10143), .B(n10142), .Z(n10279) );
  XOR U4196 ( .A(n10770), .B(n10769), .Z(n10772) );
  XNOR U4197 ( .A(n10494), .B(n10493), .Z(n10496) );
  XNOR U4198 ( .A(n10458), .B(n10457), .Z(n10460) );
  XOR U4199 ( .A(n10830), .B(n10829), .Z(n10752) );
  XOR U4200 ( .A(n10758), .B(n10757), .Z(n10760) );
  XOR U4201 ( .A(n3249), .B(n3250), .Z(n3334) );
  XOR U4202 ( .A(n9765), .B(n9764), .Z(n9771) );
  XOR U4203 ( .A(n10044), .B(n10043), .Z(n10045) );
  XOR U4204 ( .A(n10746), .B(n10745), .Z(n10748) );
  XOR U4205 ( .A(n11134), .B(n11133), .Z(n11136) );
  XNOR U4206 ( .A(n11158), .B(n11157), .Z(n11160) );
  XOR U4207 ( .A(n11380), .B(n11379), .Z(n11381) );
  XOR U4208 ( .A(n8964), .B(n8963), .Z(n8966) );
  XOR U4209 ( .A(n8451), .B(n8450), .Z(n8452) );
  XOR U4210 ( .A(n7973), .B(n7972), .Z(n7974) );
  XOR U4211 ( .A(n7495), .B(n7494), .Z(n7497) );
  XOR U4212 ( .A(n7053), .B(n7052), .Z(n7054) );
  XOR U4213 ( .A(n6053), .B(n6052), .Z(n6054) );
  XOR U4214 ( .A(n5530), .B(n5529), .Z(n5531) );
  XOR U4215 ( .A(n5220), .B(n5219), .Z(n5221) );
  XOR U4216 ( .A(n4911), .B(n4910), .Z(n4912) );
  XOR U4217 ( .A(n4637), .B(n4636), .Z(n4639) );
  XOR U4218 ( .A(n4162), .B(n4161), .Z(n4163) );
  XOR U4219 ( .A(n3972), .B(n3971), .Z(n3973) );
  XOR U4220 ( .A(n3960), .B(n3959), .Z(n3962) );
  XOR U4221 ( .A(n3404), .B(n3403), .Z(n3405) );
  XOR U4222 ( .A(n3331), .B(n3332), .Z(n3356) );
  XOR U4223 ( .A(n9789), .B(n9788), .Z(n9790) );
  XOR U4224 ( .A(n9821), .B(n9820), .Z(n10032) );
  XOR U4225 ( .A(n10089), .B(n10088), .Z(n10333) );
  XOR U4226 ( .A(n10612), .B(n10611), .Z(n10614) );
  XNOR U4227 ( .A(n10734), .B(n10733), .Z(n10736) );
  XOR U4228 ( .A(n10419), .B(n10418), .Z(n10594) );
  XOR U4229 ( .A(n10740), .B(n10739), .Z(n10742) );
  XOR U4230 ( .A(n11184), .B(n11183), .Z(n11058) );
  XOR U4231 ( .A(n11088), .B(n11087), .Z(n11090) );
  XOR U4232 ( .A(n11070), .B(n11069), .Z(n11072) );
  XNOR U4233 ( .A(n11350), .B(n11349), .Z(n11352) );
  XNOR U4234 ( .A(n11076), .B(n11075), .Z(n11078) );
  XOR U4235 ( .A(n10052), .B(n10051), .Z(n9797) );
  XOR U4236 ( .A(n9781), .B(n9780), .Z(n9782) );
  XOR U4237 ( .A(n8973), .B(n8974), .Z(n12495) );
  XOR U4238 ( .A(n7504), .B(n7505), .Z(n12461) );
  XOR U4239 ( .A(n7509), .B(n7508), .Z(n7729) );
  XOR U4240 ( .A(n6443), .B(n6442), .Z(n6444) );
  XOR U4241 ( .A(n5884), .B(n5885), .Z(n12226) );
  XOR U4242 ( .A(n5877), .B(n5876), .Z(n12402) );
  XOR U4243 ( .A(n4923), .B(n4922), .Z(n5059) );
  XOR U4244 ( .A(n4646), .B(n4647), .Z(n12367) );
  XOR U4245 ( .A(n4176), .B(n4175), .Z(n4276) );
  XOR U4246 ( .A(n3969), .B(n3970), .Z(n12333) );
  XOR U4247 ( .A(n3643), .B(n3642), .Z(n3707) );
  XOR U4248 ( .A(n3631), .B(n3630), .Z(n12298) );
  XOR U4249 ( .A(n3444), .B(n3443), .Z(n3445) );
  XOR U4250 ( .A(n3393), .B(n3394), .Z(n12277) );
  XOR U4251 ( .A(n3345), .B(n3346), .Z(n3387) );
  XOR U4252 ( .A(n3383), .B(n3384), .Z(n12265) );
  XOR U4253 ( .A(n10343), .B(n10342), .Z(n10344) );
  XOR U4254 ( .A(n10624), .B(n10623), .Z(n10626) );
  XOR U4255 ( .A(n11470), .B(n11469), .Z(n11474) );
  XOR U4256 ( .A(n11733), .B(n11732), .Z(n11735) );
  XNOR U4257 ( .A(n11697), .B(n11696), .Z(n11699) );
  ANDN U4258 ( .B(n12051), .A(n12052), .Z(n12683) );
  XOR U4259 ( .A(n12779), .B(n12778), .Z(n12777) );
  XOR U4260 ( .A(n3565), .B(n3564), .Z(n3505) );
  XOR U4261 ( .A(n3367), .B(n3368), .Z(n12250) );
  XOR U4262 ( .A(n10649), .B(n10648), .Z(n10651) );
  XOR U4263 ( .A(n10618), .B(n10617), .Z(n10620) );
  XOR U4264 ( .A(n10636), .B(n10635), .Z(n10637) );
  XOR U4265 ( .A(n11006), .B(n11005), .Z(n11218) );
  XOR U4266 ( .A(n11334), .B(n11333), .Z(n11518) );
  XOR U4267 ( .A(n11817), .B(n11816), .Z(n11679) );
  XOR U4268 ( .A(n12842), .B(n12843), .Z(n12845) );
  XOR U4269 ( .A(n10369), .B(n10368), .Z(n10371) );
  XOR U4270 ( .A(n10067), .B(n10068), .Z(n12512) );
  XOR U4271 ( .A(n8456), .B(n8457), .Z(n12478) );
  XOR U4272 ( .A(n7058), .B(n7059), .Z(n12442) );
  XOR U4273 ( .A(n6641), .B(n6642), .Z(n12430) );
  XOR U4274 ( .A(n5535), .B(n5536), .Z(n12396) );
  XOR U4275 ( .A(n12380), .B(n12381), .Z(n13285) );
  XOR U4276 ( .A(n4392), .B(n4393), .Z(n12350) );
  XOR U4277 ( .A(n3788), .B(n3789), .Z(n12316) );
  XOR U4278 ( .A(n12288), .B(n12289), .Z(n13189) );
  XOR U4279 ( .A(n12243), .B(n12244), .Z(n13147) );
  XOR U4280 ( .A(n10944), .B(n10943), .Z(n10950) );
  XOR U4281 ( .A(n11316), .B(n11315), .Z(n11310) );
  XOR U4282 ( .A(n11663), .B(n11662), .Z(n11655) );
  XOR U4283 ( .A(n12106), .B(n12105), .Z(n12110) );
  XOR U4284 ( .A(n12001), .B(n12000), .Z(n11993) );
  XNOR U4285 ( .A(n11987), .B(n11986), .Z(n11989) );
  XOR U4286 ( .A(n12646), .B(n12645), .Z(n12643) );
  XOR U4287 ( .A(n11969), .B(n11968), .Z(n11970) );
  XNOR U4288 ( .A(n12658), .B(n12657), .Z(n12656) );
  XOR U4289 ( .A(n12502), .B(n12503), .Z(n13408) );
  XOR U4290 ( .A(n12488), .B(n12489), .Z(n13397) );
  XOR U4291 ( .A(n13390), .B(n13391), .Z(n13743) );
  XOR U4292 ( .A(n12480), .B(n12481), .Z(n13384) );
  XOR U4293 ( .A(n13378), .B(n13379), .Z(n13731) );
  XOR U4294 ( .A(n12466), .B(n12467), .Z(n13373) );
  XOR U4295 ( .A(n12444), .B(n12445), .Z(n13348) );
  XOR U4296 ( .A(n12432), .B(n12433), .Z(n13336) );
  XOR U4297 ( .A(n12408), .B(n12409), .Z(n13313) );
  XOR U4298 ( .A(n12398), .B(n12399), .Z(n13300) );
  XOR U4299 ( .A(n12384), .B(n12385), .Z(n13289) );
  XOR U4300 ( .A(n12360), .B(n12361), .Z(n13265) );
  XOR U4301 ( .A(n12352), .B(n12353), .Z(n13252) );
  XOR U4302 ( .A(n12326), .B(n12327), .Z(n13229) );
  XOR U4303 ( .A(n12318), .B(n12319), .Z(n13216) );
  XOR U4304 ( .A(n12306), .B(n12307), .Z(n13204) );
  XOR U4305 ( .A(n12261), .B(n12262), .Z(n13160) );
  XOR U4306 ( .A(n13156), .B(n13157), .Z(n13508) );
  XOR U4307 ( .A(n11260), .B(n11259), .Z(n11261) );
  XOR U4308 ( .A(n11286), .B(n11285), .Z(n11280) );
  XNOR U4309 ( .A(n11963), .B(n11962), .Z(n11965) );
  XOR U4310 ( .A(n11959), .B(n11958), .Z(n11952) );
  XOR U4311 ( .A(n12933), .B(n12932), .Z(n12929) );
  XOR U4312 ( .A(n10968), .B(n10967), .Z(n10969) );
  XNOR U4313 ( .A(n13469), .B(n13470), .Z(n13755) );
  XNOR U4314 ( .A(n13473), .B(n13474), .Z(n13579) );
  XOR U4315 ( .A(n13182), .B(n13183), .Z(n13185) );
  XOR U4316 ( .A(n11875), .B(n11874), .Z(n11877) );
  XOR U4317 ( .A(n11941), .B(n11940), .Z(n12148) );
  XOR U4318 ( .A(n12963), .B(n12962), .Z(n12989) );
  XNOR U4319 ( .A(n12628), .B(n12627), .Z(n12626) );
  XOR U4320 ( .A(n13788), .B(n13789), .Z(n14153) );
  XOR U4321 ( .A(n13776), .B(n13777), .Z(n14141) );
  XOR U4322 ( .A(n13766), .B(n13767), .Z(n14129) );
  XOR U4323 ( .A(n13720), .B(n13721), .Z(n14081) );
  XOR U4324 ( .A(n13362), .B(n13363), .Z(n13712) );
  XOR U4325 ( .A(n13708), .B(n13709), .Z(n14069) );
  XOR U4326 ( .A(n13696), .B(n13697), .Z(n14057) );
  XOR U4327 ( .A(n13684), .B(n13685), .Z(n14043) );
  XOR U4328 ( .A(n13326), .B(n13327), .Z(n13677) );
  XOR U4329 ( .A(n13660), .B(n13661), .Z(n14021) );
  XOR U4330 ( .A(n13648), .B(n13649), .Z(n14007) );
  XOR U4331 ( .A(n13278), .B(n13279), .Z(n13629) );
  XOR U4332 ( .A(n13612), .B(n13613), .Z(n13973) );
  XOR U4333 ( .A(n13242), .B(n13243), .Z(n13595) );
  XOR U4334 ( .A(n13568), .B(n13569), .Z(n13923) );
  XOR U4335 ( .A(n13194), .B(n13195), .Z(n13549) );
  XOR U4336 ( .A(n13532), .B(n13533), .Z(n13889) );
  XOR U4337 ( .A(n13172), .B(n13173), .Z(n13527) );
  XOR U4338 ( .A(n13522), .B(n13523), .Z(n13877) );
  XOR U4339 ( .A(n13502), .B(n13503), .Z(n13505) );
  XOR U4340 ( .A(n13492), .B(n13493), .Z(n13830) );
  XOR U4341 ( .A(n13486), .B(n13487), .Z(n13845) );
  XOR U4342 ( .A(n11265), .B(n11266), .Z(n12538) );
  XOR U4343 ( .A(n11592), .B(n11591), .Z(n11887) );
  XOR U4344 ( .A(n13738), .B(n13739), .Z(n14096) );
  XOR U4345 ( .A(n14066), .B(n14067), .Z(n14429) );
  XOR U4346 ( .A(n14032), .B(n14033), .Z(n14392) );
  XOR U4347 ( .A(n13984), .B(n13985), .Z(n14346) );
  XOR U4348 ( .A(n13948), .B(n13949), .Z(n14312) );
  XOR U4349 ( .A(n13898), .B(n13899), .Z(n14267) );
  XOR U4350 ( .A(n13856), .B(n13857), .Z(n14220) );
  XOR U4351 ( .A(n13059), .B(n13058), .Z(n13055) );
  XOR U4352 ( .A(n12545), .B(n12546), .Z(n13458) );
  XNOR U4353 ( .A(n14180), .B(n14181), .Z(n14359) );
  XNOR U4354 ( .A(n14182), .B(n14183), .Z(n14325) );
  XNOR U4355 ( .A(n14184), .B(n14185), .Z(n14279) );
  XOR U4356 ( .A(n11898), .B(n11899), .Z(n12550) );
  XOR U4357 ( .A(n14158), .B(n14159), .Z(n14517) );
  XOR U4358 ( .A(n14146), .B(n14147), .Z(n14504) );
  XOR U4359 ( .A(n14134), .B(n14135), .Z(n14493) );
  XOR U4360 ( .A(n14122), .B(n14123), .Z(n14480) );
  XOR U4361 ( .A(n14110), .B(n14111), .Z(n14469) );
  XOR U4362 ( .A(n14086), .B(n14087), .Z(n14446) );
  XOR U4363 ( .A(n14050), .B(n14051), .Z(n14410) );
  XOR U4364 ( .A(n14026), .B(n14027), .Z(n14386) );
  XOR U4365 ( .A(n14014), .B(n14015), .Z(n14374) );
  XOR U4366 ( .A(n13978), .B(n13979), .Z(n14340) );
  XOR U4367 ( .A(n13942), .B(n13943), .Z(n14306) );
  XOR U4368 ( .A(n13930), .B(n13931), .Z(n14294) );
  XOR U4369 ( .A(n13894), .B(n13895), .Z(n14261) );
  XOR U4370 ( .A(n13884), .B(n13885), .Z(n14248) );
  XOR U4371 ( .A(n13872), .B(n13873), .Z(n14239) );
  XOR U4372 ( .A(n13841), .B(n13842), .Z(n14202) );
  XOR U4373 ( .A(n12556), .B(n12555), .Z(n13125) );
  XOR U4374 ( .A(n14528), .B(n14529), .Z(n14890) );
  XOR U4375 ( .A(n14518), .B(n14519), .Z(n14880) );
  XOR U4376 ( .A(n14506), .B(n14507), .Z(n14870) );
  XOR U4377 ( .A(n14494), .B(n14495), .Z(n14860) );
  XOR U4378 ( .A(n14482), .B(n14483), .Z(n14850) );
  XOR U4379 ( .A(n14470), .B(n14471), .Z(n14840) );
  XOR U4380 ( .A(n14458), .B(n14459), .Z(n14830) );
  XOR U4381 ( .A(n14448), .B(n14449), .Z(n14820) );
  XOR U4382 ( .A(n14434), .B(n14435), .Z(n14811) );
  XOR U4383 ( .A(n14422), .B(n14423), .Z(n14801) );
  XOR U4384 ( .A(n14412), .B(n14413), .Z(n14790) );
  XOR U4385 ( .A(n14398), .B(n14399), .Z(n14781) );
  XOR U4386 ( .A(n14388), .B(n14389), .Z(n14770) );
  XOR U4387 ( .A(n14376), .B(n14377), .Z(n14760) );
  XOR U4388 ( .A(n14362), .B(n14363), .Z(n14751) );
  XOR U4389 ( .A(n14352), .B(n14353), .Z(n14741) );
  XOR U4390 ( .A(n14342), .B(n14343), .Z(n14730) );
  XOR U4391 ( .A(n14328), .B(n14329), .Z(n14721) );
  XOR U4392 ( .A(n14318), .B(n14319), .Z(n14711) );
  XOR U4393 ( .A(n14308), .B(n14309), .Z(n14700) );
  XOR U4394 ( .A(n14296), .B(n14297), .Z(n14690) );
  XOR U4395 ( .A(n14282), .B(n14283), .Z(n14681) );
  XOR U4396 ( .A(n14272), .B(n14273), .Z(n14671) );
  XOR U4397 ( .A(n14262), .B(n14263), .Z(n14660) );
  XOR U4398 ( .A(n14250), .B(n14251), .Z(n14650) );
  XOR U4399 ( .A(n14240), .B(n14241), .Z(n14638) );
  XOR U4400 ( .A(n14226), .B(n14227), .Z(n14629) );
  XOR U4401 ( .A(n14216), .B(n14217), .Z(n14616) );
  XOR U4402 ( .A(n14204), .B(n14205), .Z(n14606) );
  XOR U4403 ( .A(n14888), .B(n14889), .Z(n14998) );
  XOR U4404 ( .A(n14878), .B(n14879), .Z(n15074) );
  XOR U4405 ( .A(n14868), .B(n14869), .Z(n15150) );
  XOR U4406 ( .A(n14858), .B(n14859), .Z(n15226) );
  XOR U4407 ( .A(n14848), .B(n14849), .Z(n15302) );
  XOR U4408 ( .A(n14838), .B(n14839), .Z(n15378) );
  XOR U4409 ( .A(n14828), .B(n14829), .Z(n15454) );
  XOR U4410 ( .A(n14818), .B(n14819), .Z(n15530) );
  XOR U4411 ( .A(n14808), .B(n14809), .Z(n15606) );
  XOR U4412 ( .A(n14798), .B(n14799), .Z(n15682) );
  XOR U4413 ( .A(n14788), .B(n14789), .Z(n15758) );
  XOR U4414 ( .A(n14778), .B(n14779), .Z(n15834) );
  XOR U4415 ( .A(n14768), .B(n14769), .Z(n15910) );
  XOR U4416 ( .A(n14758), .B(n14759), .Z(n15986) );
  XOR U4417 ( .A(n14748), .B(n14749), .Z(n16062) );
  XOR U4418 ( .A(n14738), .B(n14739), .Z(n16137) );
  XOR U4419 ( .A(n14728), .B(n14729), .Z(n16214) );
  XOR U4420 ( .A(n14718), .B(n14719), .Z(n16292) );
  XOR U4421 ( .A(n14708), .B(n14709), .Z(n16370) );
  XOR U4422 ( .A(n14698), .B(n14699), .Z(n16446) );
  XOR U4423 ( .A(n14688), .B(n14689), .Z(n16523) );
  XOR U4424 ( .A(n14678), .B(n14679), .Z(n16600) );
  XOR U4425 ( .A(n14668), .B(n14669), .Z(n16677) );
  XOR U4426 ( .A(n14658), .B(n14659), .Z(n16754) );
  XOR U4427 ( .A(n14648), .B(n14649), .Z(n16831) );
  XOR U4428 ( .A(n14636), .B(n14637), .Z(n16910) );
  XOR U4429 ( .A(n14626), .B(n14627), .Z(n16985) );
  XOR U4430 ( .A(n14614), .B(n14615), .Z(n17062) );
  XOR U4431 ( .A(n14604), .B(n14605), .Z(n17140) );
  XOR U4432 ( .A(n14594), .B(n14595), .Z(n17218) );
  ANDN U4433 ( .B(opcode[0]), .A(opcode[1]), .Z(n3097) );
  ANDN U4434 ( .B(n3097), .A(opcode[2]), .Z(n3164) );
  ANDN U4435 ( .B(opcode[1]), .A(opcode[0]), .Z(n3163) );
  NANDN U4436 ( .A(opcode[2]), .B(n3163), .Z(n3096) );
  NANDN U4437 ( .A(n3164), .B(n3096), .Z(n3092) );
  AND U4438 ( .A(o[63]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_63 ) );
  AND U4439 ( .A(o[62]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_62 ) );
  AND U4440 ( .A(o[61]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_61 ) );
  AND U4441 ( .A(o[60]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_60 ) );
  AND U4442 ( .A(o[59]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_59 ) );
  AND U4443 ( .A(o[58]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_58 ) );
  AND U4444 ( .A(o[57]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_57 ) );
  AND U4445 ( .A(o[56]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_56 ) );
  AND U4446 ( .A(o[55]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_55 ) );
  AND U4447 ( .A(o[54]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_54 ) );
  AND U4448 ( .A(o[53]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_53 ) );
  AND U4449 ( .A(o[52]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_52 ) );
  AND U4450 ( .A(o[51]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_51 ) );
  AND U4451 ( .A(o[50]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_50 ) );
  AND U4452 ( .A(o[49]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_49 ) );
  AND U4453 ( .A(o[48]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_48 ) );
  AND U4454 ( .A(o[47]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_47 ) );
  AND U4455 ( .A(o[46]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_46 ) );
  AND U4456 ( .A(o[45]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_45 ) );
  AND U4457 ( .A(o[44]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_44 ) );
  AND U4458 ( .A(o[43]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_43 ) );
  AND U4459 ( .A(o[42]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_42 ) );
  AND U4460 ( .A(o[41]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_41 ) );
  AND U4461 ( .A(o[40]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_40 ) );
  AND U4462 ( .A(o[39]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_39 ) );
  AND U4463 ( .A(o[38]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_38 ) );
  AND U4464 ( .A(o[37]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_37 ) );
  AND U4465 ( .A(o[36]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_36 ) );
  AND U4466 ( .A(o[35]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_35 ) );
  AND U4467 ( .A(o[34]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_34 ) );
  AND U4468 ( .A(o[33]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_33 ) );
  AND U4469 ( .A(o[32]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_32 ) );
  AND U4470 ( .A(o[31]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_31 ) );
  AND U4471 ( .A(o[30]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_30 ) );
  AND U4472 ( .A(o[29]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_29 ) );
  AND U4473 ( .A(o[28]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_28 ) );
  AND U4474 ( .A(o[27]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_27 ) );
  AND U4475 ( .A(o[26]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_26 ) );
  AND U4476 ( .A(o[25]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_25 ) );
  AND U4477 ( .A(o[24]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_24 ) );
  AND U4478 ( .A(o[23]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_23 ) );
  AND U4479 ( .A(o[22]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_22 ) );
  AND U4480 ( .A(o[21]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_21 ) );
  AND U4481 ( .A(o[20]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_20 ) );
  AND U4482 ( .A(o[19]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_19 ) );
  AND U4483 ( .A(o[18]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_18 ) );
  AND U4484 ( .A(o[17]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_17 ) );
  AND U4485 ( .A(o[16]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_16 ) );
  AND U4486 ( .A(o[15]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_15 ) );
  AND U4487 ( .A(o[14]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_14 ) );
  AND U4488 ( .A(o[13]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_13 ) );
  AND U4489 ( .A(o[12]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_12 ) );
  AND U4490 ( .A(o[11]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_11 ) );
  AND U4491 ( .A(o[10]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_10 ) );
  AND U4492 ( .A(o[9]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_9 ) );
  AND U4493 ( .A(o[8]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_8 ) );
  AND U4494 ( .A(o[7]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_7 ) );
  AND U4495 ( .A(o[6]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_6 ) );
  AND U4496 ( .A(o[5]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_5 ) );
  AND U4497 ( .A(o[4]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_4 ) );
  AND U4498 ( .A(o[3]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_3 ) );
  AND U4499 ( .A(o[2]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_2 ) );
  AND U4500 ( .A(o[1]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_1 ) );
  AND U4501 ( .A(o[0]), .B(n3092), .Z(\U1/RSOP_16/C2/Z_0 ) );
  AND U4502 ( .A(n3097), .B(opcode[2]), .Z(n3095) );
  NAND U4503 ( .A(n3095), .B(o[63]), .Z(n2967) );
  NAND U4504 ( .A(\stack[1][63] ), .B(n3092), .Z(n2966) );
  NAND U4505 ( .A(n2967), .B(n2966), .Z(\U1/RSOP_16/C3/Z_63 ) );
  NAND U4506 ( .A(n3095), .B(o[62]), .Z(n2969) );
  NAND U4507 ( .A(\stack[1][62] ), .B(n3092), .Z(n2968) );
  NAND U4508 ( .A(n2969), .B(n2968), .Z(\U1/RSOP_16/C3/Z_62 ) );
  NAND U4509 ( .A(n3095), .B(o[61]), .Z(n2971) );
  NAND U4510 ( .A(\stack[1][61] ), .B(n3092), .Z(n2970) );
  NAND U4511 ( .A(n2971), .B(n2970), .Z(\U1/RSOP_16/C3/Z_61 ) );
  NAND U4512 ( .A(n3095), .B(o[60]), .Z(n2973) );
  NAND U4513 ( .A(\stack[1][60] ), .B(n3092), .Z(n2972) );
  NAND U4514 ( .A(n2973), .B(n2972), .Z(\U1/RSOP_16/C3/Z_60 ) );
  NAND U4515 ( .A(n3095), .B(o[59]), .Z(n2975) );
  NAND U4516 ( .A(\stack[1][59] ), .B(n3092), .Z(n2974) );
  NAND U4517 ( .A(n2975), .B(n2974), .Z(\U1/RSOP_16/C3/Z_59 ) );
  NAND U4518 ( .A(n3095), .B(o[58]), .Z(n2977) );
  NAND U4519 ( .A(\stack[1][58] ), .B(n3092), .Z(n2976) );
  NAND U4520 ( .A(n2977), .B(n2976), .Z(\U1/RSOP_16/C3/Z_58 ) );
  NAND U4521 ( .A(n3095), .B(o[57]), .Z(n2979) );
  NAND U4522 ( .A(\stack[1][57] ), .B(n3092), .Z(n2978) );
  NAND U4523 ( .A(n2979), .B(n2978), .Z(\U1/RSOP_16/C3/Z_57 ) );
  NAND U4524 ( .A(n3095), .B(o[56]), .Z(n2981) );
  NAND U4525 ( .A(\stack[1][56] ), .B(n3092), .Z(n2980) );
  NAND U4526 ( .A(n2981), .B(n2980), .Z(\U1/RSOP_16/C3/Z_56 ) );
  NAND U4527 ( .A(n3095), .B(o[55]), .Z(n2983) );
  NAND U4528 ( .A(\stack[1][55] ), .B(n3092), .Z(n2982) );
  NAND U4529 ( .A(n2983), .B(n2982), .Z(\U1/RSOP_16/C3/Z_55 ) );
  NAND U4530 ( .A(n3095), .B(o[54]), .Z(n2985) );
  NAND U4531 ( .A(\stack[1][54] ), .B(n3092), .Z(n2984) );
  NAND U4532 ( .A(n2985), .B(n2984), .Z(\U1/RSOP_16/C3/Z_54 ) );
  NAND U4533 ( .A(n3095), .B(o[53]), .Z(n2987) );
  NAND U4534 ( .A(\stack[1][53] ), .B(n3092), .Z(n2986) );
  NAND U4535 ( .A(n2987), .B(n2986), .Z(\U1/RSOP_16/C3/Z_53 ) );
  NAND U4536 ( .A(n3095), .B(o[52]), .Z(n2989) );
  NAND U4537 ( .A(\stack[1][52] ), .B(n3092), .Z(n2988) );
  NAND U4538 ( .A(n2989), .B(n2988), .Z(\U1/RSOP_16/C3/Z_52 ) );
  NAND U4539 ( .A(n3095), .B(o[51]), .Z(n2991) );
  NAND U4540 ( .A(\stack[1][51] ), .B(n3092), .Z(n2990) );
  NAND U4541 ( .A(n2991), .B(n2990), .Z(\U1/RSOP_16/C3/Z_51 ) );
  NAND U4542 ( .A(n3095), .B(o[50]), .Z(n2993) );
  NAND U4543 ( .A(\stack[1][50] ), .B(n3092), .Z(n2992) );
  NAND U4544 ( .A(n2993), .B(n2992), .Z(\U1/RSOP_16/C3/Z_50 ) );
  NAND U4545 ( .A(n3095), .B(o[49]), .Z(n2995) );
  NAND U4546 ( .A(\stack[1][49] ), .B(n3092), .Z(n2994) );
  NAND U4547 ( .A(n2995), .B(n2994), .Z(\U1/RSOP_16/C3/Z_49 ) );
  NAND U4548 ( .A(n3095), .B(o[48]), .Z(n2997) );
  NAND U4549 ( .A(\stack[1][48] ), .B(n3092), .Z(n2996) );
  NAND U4550 ( .A(n2997), .B(n2996), .Z(\U1/RSOP_16/C3/Z_48 ) );
  NAND U4551 ( .A(n3095), .B(o[47]), .Z(n2999) );
  NAND U4552 ( .A(\stack[1][47] ), .B(n3092), .Z(n2998) );
  NAND U4553 ( .A(n2999), .B(n2998), .Z(\U1/RSOP_16/C3/Z_47 ) );
  NAND U4554 ( .A(n3095), .B(o[46]), .Z(n3001) );
  NAND U4555 ( .A(\stack[1][46] ), .B(n3092), .Z(n3000) );
  NAND U4556 ( .A(n3001), .B(n3000), .Z(\U1/RSOP_16/C3/Z_46 ) );
  NAND U4557 ( .A(n3095), .B(o[45]), .Z(n3003) );
  NAND U4558 ( .A(\stack[1][45] ), .B(n3092), .Z(n3002) );
  NAND U4559 ( .A(n3003), .B(n3002), .Z(\U1/RSOP_16/C3/Z_45 ) );
  NAND U4560 ( .A(n3095), .B(o[44]), .Z(n3005) );
  NAND U4561 ( .A(\stack[1][44] ), .B(n3092), .Z(n3004) );
  NAND U4562 ( .A(n3005), .B(n3004), .Z(\U1/RSOP_16/C3/Z_44 ) );
  NAND U4563 ( .A(n3095), .B(o[43]), .Z(n3007) );
  NAND U4564 ( .A(\stack[1][43] ), .B(n3092), .Z(n3006) );
  NAND U4565 ( .A(n3007), .B(n3006), .Z(\U1/RSOP_16/C3/Z_43 ) );
  NAND U4566 ( .A(n3095), .B(o[42]), .Z(n3009) );
  NAND U4567 ( .A(\stack[1][42] ), .B(n3092), .Z(n3008) );
  NAND U4568 ( .A(n3009), .B(n3008), .Z(\U1/RSOP_16/C3/Z_42 ) );
  NAND U4569 ( .A(n3095), .B(o[41]), .Z(n3011) );
  NAND U4570 ( .A(\stack[1][41] ), .B(n3092), .Z(n3010) );
  NAND U4571 ( .A(n3011), .B(n3010), .Z(\U1/RSOP_16/C3/Z_41 ) );
  NAND U4572 ( .A(n3095), .B(o[40]), .Z(n3013) );
  NAND U4573 ( .A(\stack[1][40] ), .B(n3092), .Z(n3012) );
  NAND U4574 ( .A(n3013), .B(n3012), .Z(\U1/RSOP_16/C3/Z_40 ) );
  NAND U4575 ( .A(n3095), .B(o[39]), .Z(n3015) );
  NAND U4576 ( .A(\stack[1][39] ), .B(n3092), .Z(n3014) );
  NAND U4577 ( .A(n3015), .B(n3014), .Z(\U1/RSOP_16/C3/Z_39 ) );
  NAND U4578 ( .A(n3095), .B(o[38]), .Z(n3017) );
  NAND U4579 ( .A(\stack[1][38] ), .B(n3092), .Z(n3016) );
  NAND U4580 ( .A(n3017), .B(n3016), .Z(\U1/RSOP_16/C3/Z_38 ) );
  NAND U4581 ( .A(n3095), .B(o[37]), .Z(n3019) );
  NAND U4582 ( .A(\stack[1][37] ), .B(n3092), .Z(n3018) );
  NAND U4583 ( .A(n3019), .B(n3018), .Z(\U1/RSOP_16/C3/Z_37 ) );
  NAND U4584 ( .A(n3095), .B(o[36]), .Z(n3021) );
  NAND U4585 ( .A(\stack[1][36] ), .B(n3092), .Z(n3020) );
  NAND U4586 ( .A(n3021), .B(n3020), .Z(\U1/RSOP_16/C3/Z_36 ) );
  NAND U4587 ( .A(n3095), .B(o[35]), .Z(n3023) );
  NAND U4588 ( .A(\stack[1][35] ), .B(n3092), .Z(n3022) );
  NAND U4589 ( .A(n3023), .B(n3022), .Z(\U1/RSOP_16/C3/Z_35 ) );
  NAND U4590 ( .A(n3095), .B(o[34]), .Z(n3025) );
  NAND U4591 ( .A(\stack[1][34] ), .B(n3092), .Z(n3024) );
  NAND U4592 ( .A(n3025), .B(n3024), .Z(\U1/RSOP_16/C3/Z_34 ) );
  NAND U4593 ( .A(n3095), .B(o[33]), .Z(n3027) );
  NAND U4594 ( .A(\stack[1][33] ), .B(n3092), .Z(n3026) );
  NAND U4595 ( .A(n3027), .B(n3026), .Z(\U1/RSOP_16/C3/Z_33 ) );
  NAND U4596 ( .A(n3095), .B(o[32]), .Z(n3029) );
  NAND U4597 ( .A(\stack[1][32] ), .B(n3092), .Z(n3028) );
  NAND U4598 ( .A(n3029), .B(n3028), .Z(\U1/RSOP_16/C3/Z_32 ) );
  NAND U4599 ( .A(n3095), .B(o[31]), .Z(n3031) );
  NAND U4600 ( .A(\stack[1][31] ), .B(n3092), .Z(n3030) );
  NAND U4601 ( .A(n3031), .B(n3030), .Z(\U1/RSOP_16/C3/Z_31 ) );
  NAND U4602 ( .A(n3095), .B(o[30]), .Z(n3033) );
  NAND U4603 ( .A(\stack[1][30] ), .B(n3092), .Z(n3032) );
  NAND U4604 ( .A(n3033), .B(n3032), .Z(\U1/RSOP_16/C3/Z_30 ) );
  NAND U4605 ( .A(n3095), .B(o[29]), .Z(n3035) );
  NAND U4606 ( .A(\stack[1][29] ), .B(n3092), .Z(n3034) );
  NAND U4607 ( .A(n3035), .B(n3034), .Z(\U1/RSOP_16/C3/Z_29 ) );
  NAND U4608 ( .A(n3095), .B(o[28]), .Z(n3037) );
  NAND U4609 ( .A(\stack[1][28] ), .B(n3092), .Z(n3036) );
  NAND U4610 ( .A(n3037), .B(n3036), .Z(\U1/RSOP_16/C3/Z_28 ) );
  NAND U4611 ( .A(n3095), .B(o[27]), .Z(n3039) );
  NAND U4612 ( .A(\stack[1][27] ), .B(n3092), .Z(n3038) );
  NAND U4613 ( .A(n3039), .B(n3038), .Z(\U1/RSOP_16/C3/Z_27 ) );
  NAND U4614 ( .A(n3095), .B(o[26]), .Z(n3041) );
  NAND U4615 ( .A(\stack[1][26] ), .B(n3092), .Z(n3040) );
  NAND U4616 ( .A(n3041), .B(n3040), .Z(\U1/RSOP_16/C3/Z_26 ) );
  NAND U4617 ( .A(n3095), .B(o[25]), .Z(n3043) );
  NAND U4618 ( .A(\stack[1][25] ), .B(n3092), .Z(n3042) );
  NAND U4619 ( .A(n3043), .B(n3042), .Z(\U1/RSOP_16/C3/Z_25 ) );
  NAND U4620 ( .A(n3095), .B(o[24]), .Z(n3045) );
  NAND U4621 ( .A(\stack[1][24] ), .B(n3092), .Z(n3044) );
  NAND U4622 ( .A(n3045), .B(n3044), .Z(\U1/RSOP_16/C3/Z_24 ) );
  NAND U4623 ( .A(n3095), .B(o[23]), .Z(n3047) );
  NAND U4624 ( .A(\stack[1][23] ), .B(n3092), .Z(n3046) );
  NAND U4625 ( .A(n3047), .B(n3046), .Z(\U1/RSOP_16/C3/Z_23 ) );
  NAND U4626 ( .A(n3095), .B(o[22]), .Z(n3049) );
  NAND U4627 ( .A(\stack[1][22] ), .B(n3092), .Z(n3048) );
  NAND U4628 ( .A(n3049), .B(n3048), .Z(\U1/RSOP_16/C3/Z_22 ) );
  NAND U4629 ( .A(n3095), .B(o[21]), .Z(n3051) );
  NAND U4630 ( .A(\stack[1][21] ), .B(n3092), .Z(n3050) );
  NAND U4631 ( .A(n3051), .B(n3050), .Z(\U1/RSOP_16/C3/Z_21 ) );
  NAND U4632 ( .A(n3095), .B(o[20]), .Z(n3053) );
  NAND U4633 ( .A(\stack[1][20] ), .B(n3092), .Z(n3052) );
  NAND U4634 ( .A(n3053), .B(n3052), .Z(\U1/RSOP_16/C3/Z_20 ) );
  NAND U4635 ( .A(n3095), .B(o[19]), .Z(n3055) );
  NAND U4636 ( .A(\stack[1][19] ), .B(n3092), .Z(n3054) );
  NAND U4637 ( .A(n3055), .B(n3054), .Z(\U1/RSOP_16/C3/Z_19 ) );
  NAND U4638 ( .A(n3095), .B(o[18]), .Z(n3057) );
  NAND U4639 ( .A(\stack[1][18] ), .B(n3092), .Z(n3056) );
  NAND U4640 ( .A(n3057), .B(n3056), .Z(\U1/RSOP_16/C3/Z_18 ) );
  NAND U4641 ( .A(n3095), .B(o[17]), .Z(n3059) );
  NAND U4642 ( .A(\stack[1][17] ), .B(n3092), .Z(n3058) );
  NAND U4643 ( .A(n3059), .B(n3058), .Z(\U1/RSOP_16/C3/Z_17 ) );
  NAND U4644 ( .A(n3095), .B(o[16]), .Z(n3061) );
  NAND U4645 ( .A(\stack[1][16] ), .B(n3092), .Z(n3060) );
  NAND U4646 ( .A(n3061), .B(n3060), .Z(\U1/RSOP_16/C3/Z_16 ) );
  NAND U4647 ( .A(n3095), .B(o[15]), .Z(n3063) );
  NAND U4648 ( .A(\stack[1][15] ), .B(n3092), .Z(n3062) );
  NAND U4649 ( .A(n3063), .B(n3062), .Z(\U1/RSOP_16/C3/Z_15 ) );
  NAND U4650 ( .A(n3095), .B(o[14]), .Z(n3065) );
  NAND U4651 ( .A(\stack[1][14] ), .B(n3092), .Z(n3064) );
  NAND U4652 ( .A(n3065), .B(n3064), .Z(\U1/RSOP_16/C3/Z_14 ) );
  NAND U4653 ( .A(n3095), .B(o[13]), .Z(n3067) );
  NAND U4654 ( .A(\stack[1][13] ), .B(n3092), .Z(n3066) );
  NAND U4655 ( .A(n3067), .B(n3066), .Z(\U1/RSOP_16/C3/Z_13 ) );
  NAND U4656 ( .A(n3095), .B(o[12]), .Z(n3069) );
  NAND U4657 ( .A(\stack[1][12] ), .B(n3092), .Z(n3068) );
  NAND U4658 ( .A(n3069), .B(n3068), .Z(\U1/RSOP_16/C3/Z_12 ) );
  NAND U4659 ( .A(n3095), .B(o[11]), .Z(n3071) );
  NAND U4660 ( .A(\stack[1][11] ), .B(n3092), .Z(n3070) );
  NAND U4661 ( .A(n3071), .B(n3070), .Z(\U1/RSOP_16/C3/Z_11 ) );
  NAND U4662 ( .A(n3095), .B(o[10]), .Z(n3073) );
  NAND U4663 ( .A(\stack[1][10] ), .B(n3092), .Z(n3072) );
  NAND U4664 ( .A(n3073), .B(n3072), .Z(\U1/RSOP_16/C3/Z_10 ) );
  NAND U4665 ( .A(n3095), .B(o[9]), .Z(n3075) );
  NAND U4666 ( .A(\stack[1][9] ), .B(n3092), .Z(n3074) );
  NAND U4667 ( .A(n3075), .B(n3074), .Z(\U1/RSOP_16/C3/Z_9 ) );
  NAND U4668 ( .A(n3095), .B(o[8]), .Z(n3077) );
  NAND U4669 ( .A(\stack[1][8] ), .B(n3092), .Z(n3076) );
  NAND U4670 ( .A(n3077), .B(n3076), .Z(\U1/RSOP_16/C3/Z_8 ) );
  NAND U4671 ( .A(n3095), .B(o[7]), .Z(n3079) );
  NAND U4672 ( .A(\stack[1][7] ), .B(n3092), .Z(n3078) );
  NAND U4673 ( .A(n3079), .B(n3078), .Z(\U1/RSOP_16/C3/Z_7 ) );
  NAND U4674 ( .A(n3095), .B(o[6]), .Z(n3081) );
  NAND U4675 ( .A(\stack[1][6] ), .B(n3092), .Z(n3080) );
  NAND U4676 ( .A(n3081), .B(n3080), .Z(\U1/RSOP_16/C3/Z_6 ) );
  NAND U4677 ( .A(n3095), .B(o[5]), .Z(n3083) );
  NAND U4678 ( .A(\stack[1][5] ), .B(n3092), .Z(n3082) );
  NAND U4679 ( .A(n3083), .B(n3082), .Z(\U1/RSOP_16/C3/Z_5 ) );
  NAND U4680 ( .A(n3095), .B(o[4]), .Z(n3085) );
  NAND U4681 ( .A(\stack[1][4] ), .B(n3092), .Z(n3084) );
  NAND U4682 ( .A(n3085), .B(n3084), .Z(\U1/RSOP_16/C3/Z_4 ) );
  NAND U4683 ( .A(n3095), .B(o[3]), .Z(n3087) );
  NAND U4684 ( .A(\stack[1][3] ), .B(n3092), .Z(n3086) );
  NAND U4685 ( .A(n3087), .B(n3086), .Z(\U1/RSOP_16/C3/Z_3 ) );
  NAND U4686 ( .A(n3095), .B(o[2]), .Z(n3089) );
  NAND U4687 ( .A(\stack[1][2] ), .B(n3092), .Z(n3088) );
  NAND U4688 ( .A(n3089), .B(n3088), .Z(\U1/RSOP_16/C3/Z_2 ) );
  NAND U4689 ( .A(n3095), .B(o[1]), .Z(n3091) );
  NAND U4690 ( .A(\stack[1][1] ), .B(n3092), .Z(n3090) );
  NAND U4691 ( .A(n3091), .B(n3090), .Z(\U1/RSOP_16/C3/Z_1 ) );
  NAND U4692 ( .A(n3095), .B(o[0]), .Z(n3094) );
  NAND U4693 ( .A(\stack[1][0] ), .B(n3092), .Z(n3093) );
  NAND U4694 ( .A(n3094), .B(n3093), .Z(\U1/RSOP_16/C3/Z_0 ) );
  NANDN U4695 ( .A(n3095), .B(n3096), .Z(\C1/Z_0 ) );
  NANDN U4696 ( .A(n3097), .B(n3096), .Z(n3161) );
  NAND U4697 ( .A(\C3/DATA5_63 ), .B(n3161), .Z(n3098) );
  AND U4698 ( .A(n14923), .B(n3098), .Z(n14929) );
  NAND U4699 ( .A(\C3/DATA5_36 ), .B(n3161), .Z(n3099) );
  AND U4700 ( .A(n15946), .B(n3099), .Z(n15951) );
  NAND U4701 ( .A(\C3/DATA5_34 ), .B(n3161), .Z(n3100) );
  AND U4702 ( .A(n16022), .B(n3100), .Z(n16027) );
  NAND U4703 ( .A(\C3/DATA5_32 ), .B(n3161), .Z(n3101) );
  AND U4704 ( .A(n16098), .B(n3101), .Z(n16103) );
  NAND U4705 ( .A(\C3/DATA5_31 ), .B(n3161), .Z(n3102) );
  AND U4706 ( .A(n16136), .B(n3102), .Z(n16141) );
  NAND U4707 ( .A(\C3/DATA5_30 ), .B(n3161), .Z(n3103) );
  AND U4708 ( .A(n16175), .B(n3103), .Z(n16180) );
  NAND U4709 ( .A(\C3/DATA5_29 ), .B(n3161), .Z(n3104) );
  AND U4710 ( .A(n16213), .B(n3104), .Z(n16218) );
  NAND U4711 ( .A(\C3/DATA5_28 ), .B(n3161), .Z(n3105) );
  AND U4712 ( .A(n16252), .B(n3105), .Z(n16257) );
  NAND U4713 ( .A(\C3/DATA5_27 ), .B(n3161), .Z(n3106) );
  AND U4714 ( .A(n16291), .B(n3106), .Z(n16296) );
  NAND U4715 ( .A(\C3/DATA5_26 ), .B(n3161), .Z(n3107) );
  AND U4716 ( .A(n16330), .B(n3107), .Z(n16335) );
  NAND U4717 ( .A(\C3/DATA5_25 ), .B(n3161), .Z(n3108) );
  AND U4718 ( .A(n16369), .B(n3108), .Z(n16374) );
  NAND U4719 ( .A(\C3/DATA5_24 ), .B(n3161), .Z(n3109) );
  AND U4720 ( .A(n16407), .B(n3109), .Z(n16412) );
  NAND U4721 ( .A(\C3/DATA5_23 ), .B(n3161), .Z(n3110) );
  AND U4722 ( .A(n16445), .B(n3110), .Z(n16450) );
  NAND U4723 ( .A(\C3/DATA5_22 ), .B(n3161), .Z(n3111) );
  AND U4724 ( .A(n16483), .B(n3111), .Z(n16488) );
  NAND U4725 ( .A(\C3/DATA5_21 ), .B(n3161), .Z(n3112) );
  AND U4726 ( .A(n16522), .B(n3112), .Z(n16527) );
  NAND U4727 ( .A(\C3/DATA5_20 ), .B(n3161), .Z(n3113) );
  AND U4728 ( .A(n16561), .B(n3113), .Z(n16566) );
  NAND U4729 ( .A(\C3/DATA5_19 ), .B(n3161), .Z(n3114) );
  AND U4730 ( .A(n16599), .B(n3114), .Z(n16604) );
  NAND U4731 ( .A(\C3/DATA5_18 ), .B(n3161), .Z(n3115) );
  AND U4732 ( .A(n16638), .B(n3115), .Z(n16643) );
  NAND U4733 ( .A(\C3/DATA5_17 ), .B(n3161), .Z(n3116) );
  AND U4734 ( .A(n16676), .B(n3116), .Z(n16681) );
  NAND U4735 ( .A(\C3/DATA5_16 ), .B(n3161), .Z(n3117) );
  AND U4736 ( .A(n16715), .B(n3117), .Z(n16720) );
  NAND U4737 ( .A(\C3/DATA5_15 ), .B(n3161), .Z(n3118) );
  AND U4738 ( .A(n16753), .B(n3118), .Z(n16758) );
  NAND U4739 ( .A(\C3/DATA5_14 ), .B(n3161), .Z(n3119) );
  AND U4740 ( .A(n16791), .B(n3119), .Z(n16796) );
  NAND U4741 ( .A(\C3/DATA5_13 ), .B(n3161), .Z(n3120) );
  AND U4742 ( .A(n16830), .B(n3120), .Z(n16835) );
  NAND U4743 ( .A(\C3/DATA5_12 ), .B(n3161), .Z(n3121) );
  AND U4744 ( .A(n16869), .B(n3121), .Z(n16874) );
  NAND U4745 ( .A(\C3/DATA5_10 ), .B(n3161), .Z(n3122) );
  AND U4746 ( .A(n16946), .B(n3122), .Z(n16951) );
  NAND U4747 ( .A(\C3/DATA5_9 ), .B(n3161), .Z(n3123) );
  AND U4748 ( .A(n16984), .B(n3123), .Z(n16989) );
  NAND U4749 ( .A(\C3/DATA5_8 ), .B(n3161), .Z(n3124) );
  AND U4750 ( .A(n17023), .B(n3124), .Z(n17028) );
  NAND U4751 ( .A(\C3/DATA5_7 ), .B(n3161), .Z(n3125) );
  AND U4752 ( .A(n17061), .B(n3125), .Z(n17066) );
  NAND U4753 ( .A(\C3/DATA5_6 ), .B(n3161), .Z(n3126) );
  AND U4754 ( .A(n17100), .B(n3126), .Z(n17105) );
  NAND U4755 ( .A(\C3/DATA5_5 ), .B(n3161), .Z(n3127) );
  AND U4756 ( .A(n17139), .B(n3127), .Z(n17144) );
  NAND U4757 ( .A(\C3/DATA5_4 ), .B(n3161), .Z(n3128) );
  AND U4758 ( .A(n17178), .B(n3128), .Z(n17183) );
  NAND U4759 ( .A(\C3/DATA5_3 ), .B(n3161), .Z(n3129) );
  AND U4760 ( .A(n17217), .B(n3129), .Z(n17222) );
  NAND U4761 ( .A(\C3/DATA5_2 ), .B(n3161), .Z(n3130) );
  AND U4762 ( .A(n17255), .B(n3130), .Z(n17256) );
  NAND U4763 ( .A(\C3/DATA5_1 ), .B(n3161), .Z(n3131) );
  AND U4764 ( .A(n17302), .B(n3131), .Z(n17303) );
  NAND U4765 ( .A(\C3/DATA5_0 ), .B(n3161), .Z(n3132) );
  AND U4766 ( .A(n17312), .B(n3132), .Z(n17323) );
  NAND U4767 ( .A(\C3/DATA5_62 ), .B(n3161), .Z(n3133) );
  NAND U4768 ( .A(n14967), .B(n3133), .Z(n2140) );
  NAND U4769 ( .A(\C3/DATA5_61 ), .B(n3161), .Z(n3134) );
  NAND U4770 ( .A(n15005), .B(n3134), .Z(n2148) );
  NAND U4771 ( .A(\C3/DATA5_60 ), .B(n3161), .Z(n3135) );
  NAND U4772 ( .A(n15043), .B(n3135), .Z(n2156) );
  NAND U4773 ( .A(\C3/DATA5_59 ), .B(n3161), .Z(n3136) );
  NAND U4774 ( .A(n15081), .B(n3136), .Z(n2164) );
  NAND U4775 ( .A(\C3/DATA5_58 ), .B(n3161), .Z(n3137) );
  NAND U4776 ( .A(n15119), .B(n3137), .Z(n2172) );
  NAND U4777 ( .A(\C3/DATA5_57 ), .B(n3161), .Z(n3138) );
  NAND U4778 ( .A(n15157), .B(n3138), .Z(n2180) );
  NAND U4779 ( .A(\C3/DATA5_56 ), .B(n3161), .Z(n3139) );
  NAND U4780 ( .A(n15195), .B(n3139), .Z(n2188) );
  NAND U4781 ( .A(\C3/DATA5_55 ), .B(n3161), .Z(n3140) );
  NAND U4782 ( .A(n15233), .B(n3140), .Z(n2196) );
  NAND U4783 ( .A(\C3/DATA5_54 ), .B(n3161), .Z(n3141) );
  NAND U4784 ( .A(n15271), .B(n3141), .Z(n2204) );
  NAND U4785 ( .A(\C3/DATA5_53 ), .B(n3161), .Z(n3142) );
  NAND U4786 ( .A(n15309), .B(n3142), .Z(n2212) );
  NAND U4787 ( .A(\C3/DATA5_52 ), .B(n3161), .Z(n3143) );
  NAND U4788 ( .A(n15347), .B(n3143), .Z(n2220) );
  NAND U4789 ( .A(\C3/DATA5_51 ), .B(n3161), .Z(n3144) );
  NAND U4790 ( .A(n15385), .B(n3144), .Z(n2228) );
  NAND U4791 ( .A(\C3/DATA5_50 ), .B(n3161), .Z(n3145) );
  NAND U4792 ( .A(n15423), .B(n3145), .Z(n2236) );
  NAND U4793 ( .A(\C3/DATA5_49 ), .B(n3161), .Z(n3146) );
  NAND U4794 ( .A(n15461), .B(n3146), .Z(n2244) );
  NAND U4795 ( .A(\C3/DATA5_48 ), .B(n3161), .Z(n3147) );
  NAND U4796 ( .A(n15499), .B(n3147), .Z(n2252) );
  NAND U4797 ( .A(\C3/DATA5_47 ), .B(n3161), .Z(n3148) );
  NAND U4798 ( .A(n15537), .B(n3148), .Z(n2260) );
  NAND U4799 ( .A(\C3/DATA5_46 ), .B(n3161), .Z(n3149) );
  NAND U4800 ( .A(n15575), .B(n3149), .Z(n2268) );
  NAND U4801 ( .A(\C3/DATA5_45 ), .B(n3161), .Z(n3150) );
  NAND U4802 ( .A(n15613), .B(n3150), .Z(n2276) );
  NAND U4803 ( .A(\C3/DATA5_44 ), .B(n3161), .Z(n3151) );
  NAND U4804 ( .A(n15651), .B(n3151), .Z(n2284) );
  NAND U4805 ( .A(\C3/DATA5_43 ), .B(n3161), .Z(n3152) );
  NAND U4806 ( .A(n15689), .B(n3152), .Z(n2292) );
  NAND U4807 ( .A(\C3/DATA5_42 ), .B(n3161), .Z(n3153) );
  NAND U4808 ( .A(n15727), .B(n3153), .Z(n2300) );
  NAND U4809 ( .A(\C3/DATA5_41 ), .B(n3161), .Z(n3154) );
  NAND U4810 ( .A(n15765), .B(n3154), .Z(n2308) );
  NAND U4811 ( .A(\C3/DATA5_40 ), .B(n3161), .Z(n3155) );
  NAND U4812 ( .A(n15803), .B(n3155), .Z(n2316) );
  NAND U4813 ( .A(\C3/DATA5_39 ), .B(n3161), .Z(n3156) );
  NAND U4814 ( .A(n15841), .B(n3156), .Z(n2324) );
  NAND U4815 ( .A(\C3/DATA5_38 ), .B(n3161), .Z(n3157) );
  NAND U4816 ( .A(n15879), .B(n3157), .Z(n2332) );
  NAND U4817 ( .A(\C3/DATA5_37 ), .B(n3161), .Z(n3158) );
  NAND U4818 ( .A(n15917), .B(n3158), .Z(n2340) );
  NAND U4819 ( .A(\C3/DATA5_35 ), .B(n3161), .Z(n3159) );
  NAND U4820 ( .A(n15993), .B(n3159), .Z(n2356) );
  NAND U4821 ( .A(\C3/DATA5_33 ), .B(n3161), .Z(n3160) );
  NAND U4822 ( .A(n16069), .B(n3160), .Z(n2372) );
  NAND U4823 ( .A(\C3/DATA5_11 ), .B(n3161), .Z(n3162) );
  NAND U4824 ( .A(n16917), .B(n3162), .Z(n2548) );
  ANDN U4825 ( .B(opcode[2]), .A(opcode[0]), .Z(n3167) );
  ANDN U4826 ( .B(n3167), .A(opcode[1]), .Z(n17311) );
  NAND U4827 ( .A(\stack[6][0] ), .B(n17311), .Z(n3166) );
  NANDN U4828 ( .A(n17311), .B(\stack[7][0] ), .Z(n3165) );
  NAND U4829 ( .A(n3166), .B(n3165), .Z(n2119) );
  AND U4830 ( .A(n17311), .B(\stack[5][0] ), .Z(n3171) );
  OR U4831 ( .A(opcode[1]), .B(n3164), .Z(n17305) );
  NOR U4832 ( .A(n17305), .B(n3167), .Z(n17308) );
  NAND U4833 ( .A(n17308), .B(\stack[6][0] ), .Z(n3169) );
  NAND U4834 ( .A(n17305), .B(\stack[7][0] ), .Z(n3168) );
  AND U4835 ( .A(n3169), .B(n3168), .Z(n3170) );
  NANDN U4836 ( .A(n3171), .B(n3170), .Z(n2120) );
  NAND U4837 ( .A(\stack[4][0] ), .B(n17311), .Z(n3173) );
  NAND U4838 ( .A(n17305), .B(\stack[6][0] ), .Z(n3172) );
  AND U4839 ( .A(n3173), .B(n3172), .Z(n3175) );
  NAND U4840 ( .A(n17308), .B(\stack[5][0] ), .Z(n3174) );
  NAND U4841 ( .A(n3175), .B(n3174), .Z(n2121) );
  NAND U4842 ( .A(\stack[3][0] ), .B(n17311), .Z(n3177) );
  NAND U4843 ( .A(n17305), .B(\stack[5][0] ), .Z(n3176) );
  AND U4844 ( .A(n3177), .B(n3176), .Z(n3179) );
  NAND U4845 ( .A(n17308), .B(\stack[4][0] ), .Z(n3178) );
  NAND U4846 ( .A(n3179), .B(n3178), .Z(n2122) );
  NAND U4847 ( .A(\stack[2][0] ), .B(n17311), .Z(n3181) );
  NAND U4848 ( .A(n17305), .B(\stack[4][0] ), .Z(n3180) );
  AND U4849 ( .A(n3181), .B(n3180), .Z(n3183) );
  NAND U4850 ( .A(n17308), .B(\stack[3][0] ), .Z(n3182) );
  NAND U4851 ( .A(n3183), .B(n3182), .Z(n2123) );
  NAND U4852 ( .A(n17311), .B(\stack[1][0] ), .Z(n3185) );
  NAND U4853 ( .A(n17305), .B(\stack[3][0] ), .Z(n3184) );
  AND U4854 ( .A(n3185), .B(n3184), .Z(n3187) );
  NAND U4855 ( .A(n17308), .B(\stack[2][0] ), .Z(n3186) );
  NAND U4856 ( .A(n3187), .B(n3186), .Z(n2124) );
  NAND U4857 ( .A(\stack[6][63] ), .B(n17311), .Z(n3189) );
  NANDN U4858 ( .A(n17311), .B(\stack[7][63] ), .Z(n3188) );
  NAND U4859 ( .A(n3189), .B(n3188), .Z(n2125) );
  NAND U4860 ( .A(\stack[5][63] ), .B(n17311), .Z(n3191) );
  NAND U4861 ( .A(n17305), .B(\stack[7][63] ), .Z(n3190) );
  AND U4862 ( .A(n3191), .B(n3190), .Z(n3193) );
  NAND U4863 ( .A(n17308), .B(\stack[6][63] ), .Z(n3192) );
  NAND U4864 ( .A(n3193), .B(n3192), .Z(n2126) );
  NAND U4865 ( .A(\stack[4][63] ), .B(n17311), .Z(n3195) );
  NAND U4866 ( .A(n17305), .B(\stack[6][63] ), .Z(n3194) );
  AND U4867 ( .A(n3195), .B(n3194), .Z(n3197) );
  NAND U4868 ( .A(n17308), .B(\stack[5][63] ), .Z(n3196) );
  NAND U4869 ( .A(n3197), .B(n3196), .Z(n2127) );
  NAND U4870 ( .A(\stack[3][63] ), .B(n17311), .Z(n3199) );
  NAND U4871 ( .A(n17305), .B(\stack[5][63] ), .Z(n3198) );
  AND U4872 ( .A(n3199), .B(n3198), .Z(n3201) );
  NAND U4873 ( .A(n17308), .B(\stack[4][63] ), .Z(n3200) );
  NAND U4874 ( .A(n3201), .B(n3200), .Z(n2128) );
  NAND U4875 ( .A(\stack[2][63] ), .B(n17311), .Z(n3203) );
  NAND U4876 ( .A(n17305), .B(\stack[4][63] ), .Z(n3202) );
  AND U4877 ( .A(n3203), .B(n3202), .Z(n3205) );
  NAND U4878 ( .A(n17308), .B(\stack[3][63] ), .Z(n3204) );
  NAND U4879 ( .A(n3205), .B(n3204), .Z(n2129) );
  NAND U4880 ( .A(n17311), .B(\stack[1][63] ), .Z(n3207) );
  NAND U4881 ( .A(n17305), .B(\stack[3][63] ), .Z(n3206) );
  AND U4882 ( .A(n3207), .B(n3206), .Z(n3209) );
  NAND U4883 ( .A(n17308), .B(\stack[2][63] ), .Z(n3208) );
  NAND U4884 ( .A(n3209), .B(n3208), .Z(n2130) );
  NAND U4885 ( .A(n17311), .B(o[63]), .Z(n3211) );
  NAND U4886 ( .A(n17305), .B(\stack[2][63] ), .Z(n3210) );
  AND U4887 ( .A(n3211), .B(n3210), .Z(n3213) );
  NAND U4888 ( .A(\stack[1][63] ), .B(n17308), .Z(n3212) );
  NAND U4889 ( .A(n3213), .B(n3212), .Z(n2131) );
  AND U4890 ( .A(opcode[1]), .B(opcode[0]), .Z(n17314) );
  NANDN U4891 ( .A(opcode[2]), .B(n17314), .Z(n17294) );
  AND U4892 ( .A(\stack[1][5] ), .B(o[57]), .Z(n13124) );
  NAND U4893 ( .A(\stack[1][6] ), .B(o[50]), .Z(n10071) );
  NAND U4894 ( .A(\stack[1][6] ), .B(o[46]), .Z(n8973) );
  NAND U4895 ( .A(\stack[1][6] ), .B(o[44]), .Z(n8710) );
  NAND U4896 ( .A(\stack[1][6] ), .B(o[38]), .Z(n7062) );
  NAND U4897 ( .A(\stack[1][6] ), .B(o[32]), .Z(n5884) );
  NAND U4898 ( .A(\stack[1][6] ), .B(o[22]), .Z(n4396) );
  NAND U4899 ( .A(\stack[1][6] ), .B(o[16]), .Z(n3874) );
  NAND U4900 ( .A(\stack[1][6] ), .B(o[12]), .Z(n3508) );
  AND U4901 ( .A(o[10]), .B(\stack[1][6] ), .Z(n3449) );
  AND U4902 ( .A(\stack[1][8] ), .B(o[7]), .Z(n3406) );
  AND U4903 ( .A(\stack[1][8] ), .B(o[5]), .Z(n3259) );
  AND U4904 ( .A(\stack[1][12] ), .B(o[1]), .Z(n3269) );
  NAND U4905 ( .A(n3269), .B(o[0]), .Z(n3214) );
  XNOR U4906 ( .A(o[2]), .B(n3214), .Z(n3215) );
  AND U4907 ( .A(\stack[1][11] ), .B(n3215), .Z(n3272) );
  NAND U4908 ( .A(\stack[1][13] ), .B(o[0]), .Z(n3216) );
  XNOR U4909 ( .A(n3269), .B(n3216), .Z(n3273) );
  AND U4910 ( .A(o[0]), .B(\stack[1][10] ), .Z(n3217) );
  AND U4911 ( .A(o[1]), .B(\stack[1][11] ), .Z(n3222) );
  AND U4912 ( .A(n3217), .B(n3222), .Z(n3218) );
  NAND U4913 ( .A(o[2]), .B(n3218), .Z(n3224) );
  NAND U4914 ( .A(n3222), .B(o[0]), .Z(n3219) );
  XNOR U4915 ( .A(o[2]), .B(n3219), .Z(n3220) );
  AND U4916 ( .A(\stack[1][10] ), .B(n3220), .Z(n3233) );
  NAND U4917 ( .A(\stack[1][12] ), .B(o[0]), .Z(n3221) );
  XNOR U4918 ( .A(n3222), .B(n3221), .Z(n3234) );
  NAND U4919 ( .A(n3233), .B(n3234), .Z(n3223) );
  NAND U4920 ( .A(n3224), .B(n3223), .Z(n3280) );
  AND U4921 ( .A(o[3]), .B(\stack[1][10] ), .Z(n3281) );
  XNOR U4922 ( .A(n3282), .B(n3281), .Z(n3266) );
  AND U4923 ( .A(o[0]), .B(\stack[1][9] ), .Z(n3225) );
  AND U4924 ( .A(o[1]), .B(\stack[1][10] ), .Z(n3230) );
  AND U4925 ( .A(n3225), .B(n3230), .Z(n3226) );
  NAND U4926 ( .A(o[2]), .B(n3226), .Z(n3232) );
  NAND U4927 ( .A(n3230), .B(o[0]), .Z(n3227) );
  XNOR U4928 ( .A(o[2]), .B(n3227), .Z(n3228) );
  AND U4929 ( .A(\stack[1][9] ), .B(n3228), .Z(n3247) );
  NAND U4930 ( .A(\stack[1][11] ), .B(o[0]), .Z(n3229) );
  XNOR U4931 ( .A(n3230), .B(n3229), .Z(n3248) );
  NAND U4932 ( .A(n3247), .B(n3248), .Z(n3231) );
  NAND U4933 ( .A(n3232), .B(n3231), .Z(n3235) );
  NAND U4934 ( .A(n3235), .B(n3236), .Z(n3238) );
  AND U4935 ( .A(o[3]), .B(\stack[1][9] ), .Z(n3253) );
  NAND U4936 ( .A(n3253), .B(n3254), .Z(n3237) );
  AND U4937 ( .A(n3238), .B(n3237), .Z(n3263) );
  NAND U4938 ( .A(o[4]), .B(\stack[1][9] ), .Z(n3264) );
  NAND U4939 ( .A(n3259), .B(n3260), .Z(n3262) );
  AND U4940 ( .A(o[0]), .B(\stack[1][8] ), .Z(n3239) );
  AND U4941 ( .A(o[1]), .B(\stack[1][9] ), .Z(n3244) );
  AND U4942 ( .A(n3239), .B(n3244), .Z(n3240) );
  NAND U4943 ( .A(o[2]), .B(n3240), .Z(n3246) );
  NAND U4944 ( .A(n3244), .B(o[0]), .Z(n3241) );
  XNOR U4945 ( .A(o[2]), .B(n3241), .Z(n3242) );
  AND U4946 ( .A(\stack[1][8] ), .B(n3242), .Z(n3325) );
  NAND U4947 ( .A(\stack[1][10] ), .B(o[0]), .Z(n3243) );
  XNOR U4948 ( .A(n3244), .B(n3243), .Z(n3326) );
  NAND U4949 ( .A(n3325), .B(n3326), .Z(n3245) );
  NAND U4950 ( .A(n3246), .B(n3245), .Z(n3249) );
  NAND U4951 ( .A(n3249), .B(n3250), .Z(n3252) );
  AND U4952 ( .A(o[3]), .B(\stack[1][8] ), .Z(n3333) );
  NAND U4953 ( .A(n3333), .B(n3334), .Z(n3251) );
  NAND U4954 ( .A(n3252), .B(n3251), .Z(n3255) );
  AND U4955 ( .A(o[4]), .B(\stack[1][8] ), .Z(n3256) );
  NAND U4956 ( .A(n3255), .B(n3256), .Z(n3258) );
  NAND U4957 ( .A(n3338), .B(n3337), .Z(n3257) );
  NAND U4958 ( .A(n3258), .B(n3257), .Z(n3343) );
  XOR U4959 ( .A(n3260), .B(n3259), .Z(n3344) );
  NAND U4960 ( .A(n3343), .B(n3344), .Z(n3261) );
  NAND U4961 ( .A(n3262), .B(n3261), .Z(n3285) );
  NAND U4962 ( .A(n3264), .B(n3263), .Z(n3268) );
  NAND U4963 ( .A(n3266), .B(n3265), .Z(n3267) );
  AND U4964 ( .A(n3268), .B(n3267), .Z(n3312) );
  AND U4965 ( .A(o[0]), .B(\stack[1][11] ), .Z(n3270) );
  AND U4966 ( .A(n3270), .B(n3269), .Z(n3271) );
  NAND U4967 ( .A(o[2]), .B(n3271), .Z(n3275) );
  NAND U4968 ( .A(n3273), .B(n3272), .Z(n3274) );
  NAND U4969 ( .A(n3275), .B(n3274), .Z(n3290) );
  AND U4970 ( .A(o[1]), .B(\stack[1][13] ), .Z(n3298) );
  NAND U4971 ( .A(\stack[1][14] ), .B(o[0]), .Z(n3276) );
  XNOR U4972 ( .A(n3298), .B(n3276), .Z(n3301) );
  NAND U4973 ( .A(n3298), .B(o[0]), .Z(n3277) );
  XNOR U4974 ( .A(o[2]), .B(n3277), .Z(n3278) );
  AND U4975 ( .A(\stack[1][12] ), .B(n3278), .Z(n3302) );
  AND U4976 ( .A(o[3]), .B(\stack[1][11] ), .Z(n3292) );
  AND U4977 ( .A(o[4]), .B(\stack[1][10] ), .Z(n3305) );
  NAND U4978 ( .A(n3280), .B(n3279), .Z(n3284) );
  NAND U4979 ( .A(n3282), .B(n3281), .Z(n3283) );
  NAND U4980 ( .A(n3284), .B(n3283), .Z(n3306) );
  XOR U4981 ( .A(n3308), .B(n3307), .Z(n3311) );
  XOR U4982 ( .A(n3312), .B(n3311), .Z(n3313) );
  AND U4983 ( .A(o[5]), .B(\stack[1][9] ), .Z(n3314) );
  NAND U4984 ( .A(n3285), .B(n3286), .Z(n3288) );
  AND U4985 ( .A(\stack[1][8] ), .B(o[6]), .Z(n3350) );
  NAND U4986 ( .A(n3350), .B(n3349), .Z(n3287) );
  NAND U4987 ( .A(n3288), .B(n3287), .Z(n3404) );
  AND U4988 ( .A(o[6]), .B(\stack[1][9] ), .Z(n3440) );
  NAND U4989 ( .A(n3290), .B(n3289), .Z(n3294) );
  NAND U4990 ( .A(n3292), .B(n3291), .Z(n3293) );
  NAND U4991 ( .A(n3294), .B(n3293), .Z(n3410) );
  AND U4992 ( .A(o[4]), .B(\stack[1][11] ), .Z(n3409) );
  AND U4993 ( .A(o[1]), .B(\stack[1][14] ), .Z(n3415) );
  NAND U4994 ( .A(\stack[1][15] ), .B(o[0]), .Z(n3295) );
  XNOR U4995 ( .A(n3415), .B(n3295), .Z(n3418) );
  NAND U4996 ( .A(n3415), .B(o[0]), .Z(n3296) );
  XNOR U4997 ( .A(o[2]), .B(n3296), .Z(n3297) );
  AND U4998 ( .A(\stack[1][13] ), .B(n3297), .Z(n3419) );
  AND U4999 ( .A(o[0]), .B(\stack[1][12] ), .Z(n3299) );
  AND U5000 ( .A(n3299), .B(n3298), .Z(n3300) );
  NAND U5001 ( .A(o[2]), .B(n3300), .Z(n3304) );
  NAND U5002 ( .A(n3302), .B(n3301), .Z(n3303) );
  NAND U5003 ( .A(n3304), .B(n3303), .Z(n3426) );
  AND U5004 ( .A(o[3]), .B(\stack[1][12] ), .Z(n3428) );
  XOR U5005 ( .A(n3412), .B(n3411), .Z(n3431) );
  AND U5006 ( .A(o[5]), .B(\stack[1][10] ), .Z(n3432) );
  NAND U5007 ( .A(n3306), .B(n3305), .Z(n3310) );
  NAND U5008 ( .A(n3308), .B(n3307), .Z(n3309) );
  NAND U5009 ( .A(n3310), .B(n3309), .Z(n3434) );
  NAND U5010 ( .A(n3312), .B(n3311), .Z(n3316) );
  NAND U5011 ( .A(n3314), .B(n3313), .Z(n3315) );
  NAND U5012 ( .A(n3316), .B(n3315), .Z(n3438) );
  XOR U5013 ( .A(n3440), .B(n3439), .Z(n3403) );
  XOR U5014 ( .A(n3406), .B(n3405), .Z(n3446) );
  AND U5015 ( .A(\stack[1][7] ), .B(o[8]), .Z(n3443) );
  AND U5016 ( .A(o[0]), .B(\stack[1][7] ), .Z(n3317) );
  AND U5017 ( .A(\stack[1][8] ), .B(o[1]), .Z(n3320) );
  AND U5018 ( .A(n3317), .B(n3320), .Z(n3318) );
  NAND U5019 ( .A(o[2]), .B(n3318), .Z(n3324) );
  NAND U5020 ( .A(\stack[1][9] ), .B(o[0]), .Z(n3319) );
  XNOR U5021 ( .A(n3320), .B(n3319), .Z(n3365) );
  NAND U5022 ( .A(n3320), .B(o[0]), .Z(n3321) );
  XNOR U5023 ( .A(o[2]), .B(n3321), .Z(n3322) );
  AND U5024 ( .A(\stack[1][7] ), .B(n3322), .Z(n3366) );
  NAND U5025 ( .A(n3365), .B(n3366), .Z(n3323) );
  NAND U5026 ( .A(n3324), .B(n3323), .Z(n3327) );
  NAND U5027 ( .A(n3327), .B(n3328), .Z(n3330) );
  AND U5028 ( .A(o[3]), .B(\stack[1][7] ), .Z(n3372) );
  NAND U5029 ( .A(n3372), .B(n3371), .Z(n3329) );
  NAND U5030 ( .A(n3330), .B(n3329), .Z(n3331) );
  AND U5031 ( .A(o[4]), .B(\stack[1][7] ), .Z(n3332) );
  NAND U5032 ( .A(n3331), .B(n3332), .Z(n3336) );
  NAND U5033 ( .A(n3356), .B(n3355), .Z(n3335) );
  NAND U5034 ( .A(n3336), .B(n3335), .Z(n3339) );
  XOR U5035 ( .A(n3338), .B(n3337), .Z(n3340) );
  NAND U5036 ( .A(n3339), .B(n3340), .Z(n3342) );
  AND U5037 ( .A(\stack[1][7] ), .B(o[5]), .Z(n3382) );
  NAND U5038 ( .A(n3382), .B(n3381), .Z(n3341) );
  NAND U5039 ( .A(n3342), .B(n3341), .Z(n3345) );
  NAND U5040 ( .A(n3345), .B(n3346), .Z(n3348) );
  AND U5041 ( .A(\stack[1][7] ), .B(o[6]), .Z(n3388) );
  NAND U5042 ( .A(n3388), .B(n3387), .Z(n3347) );
  NAND U5043 ( .A(n3348), .B(n3347), .Z(n3351) );
  XOR U5044 ( .A(n3350), .B(n3349), .Z(n3352) );
  NAND U5045 ( .A(n3351), .B(n3352), .Z(n3354) );
  AND U5046 ( .A(\stack[1][7] ), .B(o[7]), .Z(n3396) );
  NAND U5047 ( .A(n3396), .B(n3395), .Z(n3353) );
  NAND U5048 ( .A(n3354), .B(n3353), .Z(n3444) );
  XNOR U5049 ( .A(n3446), .B(n3445), .Z(n3399) );
  AND U5050 ( .A(\stack[1][6] ), .B(o[5]), .Z(n3377) );
  XOR U5051 ( .A(n3356), .B(n3355), .Z(n3378) );
  NAND U5052 ( .A(n3377), .B(n3378), .Z(n3380) );
  AND U5053 ( .A(o[0]), .B(\stack[1][6] ), .Z(n3357) );
  AND U5054 ( .A(o[1]), .B(\stack[1][7] ), .Z(n3362) );
  AND U5055 ( .A(n3357), .B(n3362), .Z(n3358) );
  NAND U5056 ( .A(o[2]), .B(n3358), .Z(n3364) );
  NAND U5057 ( .A(n3362), .B(o[0]), .Z(n3359) );
  XNOR U5058 ( .A(o[2]), .B(n3359), .Z(n3360) );
  AND U5059 ( .A(\stack[1][6] ), .B(n3360), .Z(n12241) );
  NAND U5060 ( .A(\stack[1][8] ), .B(o[0]), .Z(n3361) );
  XNOR U5061 ( .A(n3362), .B(n3361), .Z(n12242) );
  NAND U5062 ( .A(n12241), .B(n12242), .Z(n3363) );
  NAND U5063 ( .A(n3364), .B(n3363), .Z(n3367) );
  NAND U5064 ( .A(n3367), .B(n3368), .Z(n3370) );
  AND U5065 ( .A(\stack[1][6] ), .B(o[3]), .Z(n12249) );
  NAND U5066 ( .A(n12249), .B(n12250), .Z(n3369) );
  NAND U5067 ( .A(n3370), .B(n3369), .Z(n3373) );
  AND U5068 ( .A(\stack[1][6] ), .B(o[4]), .Z(n3374) );
  NAND U5069 ( .A(n3373), .B(n3374), .Z(n3376) );
  XOR U5070 ( .A(n3372), .B(n3371), .Z(n12254) );
  NAND U5071 ( .A(n12254), .B(n12253), .Z(n3375) );
  NAND U5072 ( .A(n3376), .B(n3375), .Z(n12259) );
  NAND U5073 ( .A(n12259), .B(n12260), .Z(n3379) );
  NAND U5074 ( .A(n3380), .B(n3379), .Z(n3383) );
  XOR U5075 ( .A(n3382), .B(n3381), .Z(n3384) );
  NAND U5076 ( .A(n3383), .B(n3384), .Z(n3386) );
  AND U5077 ( .A(\stack[1][6] ), .B(o[6]), .Z(n17097) );
  NAND U5078 ( .A(n17097), .B(n12265), .Z(n3385) );
  NAND U5079 ( .A(n3386), .B(n3385), .Z(n3389) );
  XOR U5080 ( .A(n3388), .B(n3387), .Z(n3390) );
  NAND U5081 ( .A(n3389), .B(n3390), .Z(n3392) );
  AND U5082 ( .A(\stack[1][6] ), .B(o[7]), .Z(n12270) );
  NAND U5083 ( .A(n12270), .B(n12271), .Z(n3391) );
  NAND U5084 ( .A(n3392), .B(n3391), .Z(n3393) );
  AND U5085 ( .A(\stack[1][6] ), .B(o[8]), .Z(n3394) );
  NAND U5086 ( .A(n3393), .B(n3394), .Z(n3398) );
  XOR U5087 ( .A(n3396), .B(n3395), .Z(n12276) );
  NAND U5088 ( .A(n12277), .B(n12276), .Z(n3397) );
  AND U5089 ( .A(n3398), .B(n3397), .Z(n3400) );
  NAND U5090 ( .A(n3399), .B(n3400), .Z(n3402) );
  NAND U5091 ( .A(\stack[1][6] ), .B(o[9]), .Z(n12282) );
  NAND U5092 ( .A(n12283), .B(n12282), .Z(n3401) );
  AND U5093 ( .A(n3402), .B(n3401), .Z(n3450) );
  NAND U5094 ( .A(n3449), .B(n3450), .Z(n3452) );
  AND U5095 ( .A(\stack[1][8] ), .B(o[8]), .Z(n17020) );
  NAND U5096 ( .A(n3404), .B(n3403), .Z(n3408) );
  NAND U5097 ( .A(n3406), .B(n3405), .Z(n3407) );
  NAND U5098 ( .A(n3408), .B(n3407), .Z(n3453) );
  AND U5099 ( .A(o[6]), .B(\stack[1][10] ), .Z(n3461) );
  NAND U5100 ( .A(n3410), .B(n3409), .Z(n3414) );
  NAND U5101 ( .A(n3412), .B(n3411), .Z(n3413) );
  NAND U5102 ( .A(n3414), .B(n3413), .Z(n3487) );
  AND U5103 ( .A(o[3]), .B(\stack[1][13] ), .Z(n3477) );
  AND U5104 ( .A(o[0]), .B(\stack[1][13] ), .Z(n3416) );
  AND U5105 ( .A(n3416), .B(n3415), .Z(n3417) );
  NAND U5106 ( .A(o[2]), .B(n3417), .Z(n3421) );
  NAND U5107 ( .A(n3419), .B(n3418), .Z(n3420) );
  NAND U5108 ( .A(n3421), .B(n3420), .Z(n3475) );
  AND U5109 ( .A(o[1]), .B(\stack[1][15] ), .Z(n3467) );
  NAND U5110 ( .A(\stack[1][16] ), .B(o[0]), .Z(n3422) );
  XNOR U5111 ( .A(n3467), .B(n3422), .Z(n3470) );
  NAND U5112 ( .A(n3467), .B(o[0]), .Z(n3423) );
  XNOR U5113 ( .A(o[2]), .B(n3423), .Z(n3424) );
  AND U5114 ( .A(\stack[1][14] ), .B(n3424), .Z(n3471) );
  XOR U5115 ( .A(n3477), .B(n3476), .Z(n3483) );
  AND U5116 ( .A(o[4]), .B(\stack[1][12] ), .Z(n3480) );
  NAND U5117 ( .A(n3426), .B(n3425), .Z(n3430) );
  NAND U5118 ( .A(n3428), .B(n3427), .Z(n3429) );
  NAND U5119 ( .A(n3430), .B(n3429), .Z(n3481) );
  XOR U5120 ( .A(n3483), .B(n3482), .Z(n3486) );
  AND U5121 ( .A(o[5]), .B(\stack[1][11] ), .Z(n3489) );
  NAND U5122 ( .A(n3432), .B(n3431), .Z(n3436) );
  NAND U5123 ( .A(n3434), .B(n3433), .Z(n3435) );
  NAND U5124 ( .A(n3436), .B(n3435), .Z(n3459) );
  XOR U5125 ( .A(n3461), .B(n3460), .Z(n3492) );
  NAND U5126 ( .A(n3438), .B(n3437), .Z(n3442) );
  NAND U5127 ( .A(n3440), .B(n3439), .Z(n3441) );
  NAND U5128 ( .A(n3442), .B(n3441), .Z(n3493) );
  AND U5129 ( .A(\stack[1][9] ), .B(o[7]), .Z(n3495) );
  XOR U5130 ( .A(n3455), .B(n3454), .Z(n3498) );
  NAND U5131 ( .A(n3444), .B(n3443), .Z(n3448) );
  NAND U5132 ( .A(n3446), .B(n3445), .Z(n3447) );
  NAND U5133 ( .A(n3448), .B(n3447), .Z(n3499) );
  AND U5134 ( .A(\stack[1][7] ), .B(o[9]), .Z(n3501) );
  NAND U5135 ( .A(n12232), .B(n12231), .Z(n3451) );
  NAND U5136 ( .A(n3452), .B(n3451), .Z(n3504) );
  NAND U5137 ( .A(n3453), .B(n17020), .Z(n3457) );
  NAND U5138 ( .A(n3455), .B(n3454), .Z(n3456) );
  AND U5139 ( .A(n3457), .B(n3456), .Z(n3556) );
  NAND U5140 ( .A(n3459), .B(n3458), .Z(n3463) );
  NAND U5141 ( .A(n3461), .B(n3460), .Z(n3462) );
  NAND U5142 ( .A(n3463), .B(n3462), .Z(n3511) );
  AND U5143 ( .A(o[6]), .B(\stack[1][11] ), .Z(n3547) );
  AND U5144 ( .A(o[1]), .B(\stack[1][16] ), .Z(n3522) );
  NAND U5145 ( .A(\stack[1][17] ), .B(o[0]), .Z(n3464) );
  XNOR U5146 ( .A(n3522), .B(n3464), .Z(n3525) );
  NAND U5147 ( .A(n3522), .B(o[0]), .Z(n3465) );
  XNOR U5148 ( .A(o[2]), .B(n3465), .Z(n3466) );
  AND U5149 ( .A(\stack[1][15] ), .B(n3466), .Z(n3526) );
  AND U5150 ( .A(o[0]), .B(\stack[1][14] ), .Z(n3468) );
  AND U5151 ( .A(n3468), .B(n3467), .Z(n3469) );
  NAND U5152 ( .A(o[2]), .B(n3469), .Z(n3473) );
  NAND U5153 ( .A(n3471), .B(n3470), .Z(n3472) );
  NAND U5154 ( .A(n3473), .B(n3472), .Z(n3533) );
  AND U5155 ( .A(o[3]), .B(\stack[1][14] ), .Z(n3534) );
  XNOR U5156 ( .A(n3535), .B(n3534), .Z(n3519) );
  NAND U5157 ( .A(n3475), .B(n3474), .Z(n3479) );
  NAND U5158 ( .A(n3477), .B(n3476), .Z(n3478) );
  AND U5159 ( .A(n3479), .B(n3478), .Z(n3516) );
  NAND U5160 ( .A(o[4]), .B(\stack[1][13] ), .Z(n3517) );
  AND U5161 ( .A(o[5]), .B(\stack[1][12] ), .Z(n3539) );
  XOR U5162 ( .A(n3538), .B(n3539), .Z(n3540) );
  NAND U5163 ( .A(n3481), .B(n3480), .Z(n3485) );
  NAND U5164 ( .A(n3483), .B(n3482), .Z(n3484) );
  NAND U5165 ( .A(n3485), .B(n3484), .Z(n3541) );
  NAND U5166 ( .A(n3487), .B(n3486), .Z(n3491) );
  NAND U5167 ( .A(n3489), .B(n3488), .Z(n3490) );
  NAND U5168 ( .A(n3491), .B(n3490), .Z(n3545) );
  XOR U5169 ( .A(n3547), .B(n3546), .Z(n3510) );
  AND U5170 ( .A(o[7]), .B(\stack[1][10] ), .Z(n3513) );
  AND U5171 ( .A(\stack[1][9] ), .B(o[8]), .Z(n3550) );
  NAND U5172 ( .A(n3493), .B(n3492), .Z(n3497) );
  NAND U5173 ( .A(n3495), .B(n3494), .Z(n3496) );
  NAND U5174 ( .A(n3497), .B(n3496), .Z(n3551) );
  XNOR U5175 ( .A(n3553), .B(n3552), .Z(n3557) );
  NAND U5176 ( .A(\stack[1][8] ), .B(o[9]), .Z(n3558) );
  XNOR U5177 ( .A(n3559), .B(n3558), .Z(n3565) );
  AND U5178 ( .A(o[10]), .B(\stack[1][7] ), .Z(n3562) );
  NAND U5179 ( .A(n3499), .B(n3498), .Z(n3503) );
  NAND U5180 ( .A(n3501), .B(n3500), .Z(n3502) );
  NAND U5181 ( .A(n3503), .B(n3502), .Z(n3563) );
  NAND U5182 ( .A(n3504), .B(n3505), .Z(n3507) );
  AND U5183 ( .A(\stack[1][6] ), .B(o[11]), .Z(n12292) );
  NAND U5184 ( .A(n12292), .B(n12293), .Z(n3506) );
  AND U5185 ( .A(n3507), .B(n3506), .Z(n3509) );
  NAND U5186 ( .A(n3508), .B(n3509), .Z(n3569) );
  NAND U5187 ( .A(\stack[1][7] ), .B(o[11]), .Z(n3631) );
  AND U5188 ( .A(\stack[1][9] ), .B(o[9]), .Z(n3625) );
  NAND U5189 ( .A(n3511), .B(n3510), .Z(n3515) );
  NAND U5190 ( .A(n3513), .B(n3512), .Z(n3514) );
  NAND U5191 ( .A(n3515), .B(n3514), .Z(n3577) );
  AND U5192 ( .A(o[8]), .B(\stack[1][10] ), .Z(n3576) );
  AND U5193 ( .A(o[6]), .B(\stack[1][12] ), .Z(n3585) );
  NAND U5194 ( .A(n3517), .B(n3516), .Z(n3521) );
  NAND U5195 ( .A(n3519), .B(n3518), .Z(n3520) );
  AND U5196 ( .A(n3521), .B(n3520), .Z(n3611) );
  AND U5197 ( .A(o[3]), .B(\stack[1][15] ), .Z(n3601) );
  AND U5198 ( .A(o[0]), .B(\stack[1][15] ), .Z(n3523) );
  AND U5199 ( .A(n3523), .B(n3522), .Z(n3524) );
  NAND U5200 ( .A(o[2]), .B(n3524), .Z(n3528) );
  NAND U5201 ( .A(n3526), .B(n3525), .Z(n3527) );
  NAND U5202 ( .A(n3528), .B(n3527), .Z(n3599) );
  AND U5203 ( .A(o[1]), .B(\stack[1][17] ), .Z(n3591) );
  NAND U5204 ( .A(\stack[1][18] ), .B(o[0]), .Z(n3529) );
  XNOR U5205 ( .A(n3591), .B(n3529), .Z(n3594) );
  NAND U5206 ( .A(n3591), .B(o[0]), .Z(n3530) );
  XNOR U5207 ( .A(o[2]), .B(n3530), .Z(n3531) );
  AND U5208 ( .A(\stack[1][16] ), .B(n3531), .Z(n3595) );
  XOR U5209 ( .A(n3601), .B(n3600), .Z(n3607) );
  AND U5210 ( .A(o[4]), .B(\stack[1][14] ), .Z(n3604) );
  NAND U5211 ( .A(n3533), .B(n3532), .Z(n3537) );
  NAND U5212 ( .A(n3535), .B(n3534), .Z(n3536) );
  NAND U5213 ( .A(n3537), .B(n3536), .Z(n3605) );
  XOR U5214 ( .A(n3607), .B(n3606), .Z(n3610) );
  XOR U5215 ( .A(n3611), .B(n3610), .Z(n3612) );
  AND U5216 ( .A(o[5]), .B(\stack[1][13] ), .Z(n3613) );
  NAND U5217 ( .A(n3539), .B(n3538), .Z(n3543) );
  NAND U5218 ( .A(n3541), .B(n3540), .Z(n3542) );
  NAND U5219 ( .A(n3543), .B(n3542), .Z(n3583) );
  XOR U5220 ( .A(n3585), .B(n3584), .Z(n3616) );
  NAND U5221 ( .A(n3545), .B(n3544), .Z(n3549) );
  NAND U5222 ( .A(n3547), .B(n3546), .Z(n3548) );
  NAND U5223 ( .A(n3549), .B(n3548), .Z(n3617) );
  AND U5224 ( .A(o[7]), .B(\stack[1][11] ), .Z(n3619) );
  XOR U5225 ( .A(n3579), .B(n3578), .Z(n3622) );
  NAND U5226 ( .A(n3551), .B(n3550), .Z(n3555) );
  NAND U5227 ( .A(n3553), .B(n3552), .Z(n3554) );
  NAND U5228 ( .A(n3555), .B(n3554), .Z(n3623) );
  XOR U5229 ( .A(n3625), .B(n3624), .Z(n3573) );
  AND U5230 ( .A(o[10]), .B(\stack[1][8] ), .Z(n3570) );
  NAND U5231 ( .A(n3557), .B(n3556), .Z(n3561) );
  NAND U5232 ( .A(n3559), .B(n3558), .Z(n3560) );
  AND U5233 ( .A(n3561), .B(n3560), .Z(n3571) );
  XNOR U5234 ( .A(n3573), .B(n3572), .Z(n3629) );
  NAND U5235 ( .A(n3563), .B(n3562), .Z(n3567) );
  NAND U5236 ( .A(n3565), .B(n3564), .Z(n3566) );
  AND U5237 ( .A(n3567), .B(n3566), .Z(n3628) );
  NAND U5238 ( .A(n12299), .B(n12298), .Z(n3568) );
  AND U5239 ( .A(n3569), .B(n3568), .Z(n3635) );
  NAND U5240 ( .A(n3571), .B(n3570), .Z(n3575) );
  NAND U5241 ( .A(n3573), .B(n3572), .Z(n3574) );
  NAND U5242 ( .A(n3575), .B(n3574), .Z(n3641) );
  NAND U5243 ( .A(n3577), .B(n3576), .Z(n3581) );
  NAND U5244 ( .A(n3579), .B(n3578), .Z(n3580) );
  AND U5245 ( .A(n3581), .B(n3580), .Z(n3652) );
  NAND U5246 ( .A(n3583), .B(n3582), .Z(n3587) );
  NAND U5247 ( .A(n3585), .B(n3584), .Z(n3586) );
  NAND U5248 ( .A(n3587), .B(n3586), .Z(n3659) );
  AND U5249 ( .A(o[6]), .B(\stack[1][13] ), .Z(n3695) );
  AND U5250 ( .A(\stack[1][18] ), .B(o[1]), .Z(n3670) );
  NAND U5251 ( .A(n3670), .B(o[0]), .Z(n3588) );
  XNOR U5252 ( .A(o[2]), .B(n3588), .Z(n3589) );
  AND U5253 ( .A(\stack[1][17] ), .B(n3589), .Z(n3673) );
  NAND U5254 ( .A(\stack[1][19] ), .B(o[0]), .Z(n3590) );
  XNOR U5255 ( .A(n3670), .B(n3590), .Z(n3674) );
  AND U5256 ( .A(o[0]), .B(\stack[1][16] ), .Z(n3592) );
  AND U5257 ( .A(n3592), .B(n3591), .Z(n3593) );
  NAND U5258 ( .A(o[2]), .B(n3593), .Z(n3597) );
  NAND U5259 ( .A(n3595), .B(n3594), .Z(n3596) );
  NAND U5260 ( .A(n3597), .B(n3596), .Z(n3681) );
  AND U5261 ( .A(o[3]), .B(\stack[1][16] ), .Z(n3683) );
  NAND U5262 ( .A(n3599), .B(n3598), .Z(n3603) );
  NAND U5263 ( .A(n3601), .B(n3600), .Z(n3602) );
  NAND U5264 ( .A(n3603), .B(n3602), .Z(n3665) );
  AND U5265 ( .A(o[4]), .B(\stack[1][15] ), .Z(n3664) );
  XOR U5266 ( .A(n3667), .B(n3666), .Z(n3686) );
  AND U5267 ( .A(o[5]), .B(\stack[1][14] ), .Z(n3687) );
  NAND U5268 ( .A(n3605), .B(n3604), .Z(n3609) );
  NAND U5269 ( .A(n3607), .B(n3606), .Z(n3608) );
  NAND U5270 ( .A(n3609), .B(n3608), .Z(n3689) );
  NAND U5271 ( .A(n3611), .B(n3610), .Z(n3615) );
  NAND U5272 ( .A(n3613), .B(n3612), .Z(n3614) );
  NAND U5273 ( .A(n3615), .B(n3614), .Z(n3693) );
  XOR U5274 ( .A(n3695), .B(n3694), .Z(n3658) );
  AND U5275 ( .A(o[7]), .B(\stack[1][12] ), .Z(n3661) );
  AND U5276 ( .A(o[8]), .B(\stack[1][11] ), .Z(n3698) );
  NAND U5277 ( .A(n3617), .B(n3616), .Z(n3621) );
  NAND U5278 ( .A(n3619), .B(n3618), .Z(n3620) );
  NAND U5279 ( .A(n3621), .B(n3620), .Z(n3699) );
  XNOR U5280 ( .A(n3701), .B(n3700), .Z(n3653) );
  NAND U5281 ( .A(\stack[1][10] ), .B(o[9]), .Z(n3654) );
  XNOR U5282 ( .A(n3655), .B(n3654), .Z(n3649) );
  AND U5283 ( .A(o[10]), .B(\stack[1][9] ), .Z(n3646) );
  NAND U5284 ( .A(n3623), .B(n3622), .Z(n3627) );
  NAND U5285 ( .A(n3625), .B(n3624), .Z(n3626) );
  NAND U5286 ( .A(n3627), .B(n3626), .Z(n3647) );
  AND U5287 ( .A(\stack[1][8] ), .B(o[11]), .Z(n3643) );
  AND U5288 ( .A(\stack[1][7] ), .B(o[12]), .Z(n3704) );
  NAND U5289 ( .A(n3629), .B(n3628), .Z(n3633) );
  NAND U5290 ( .A(n3631), .B(n3630), .Z(n3632) );
  AND U5291 ( .A(n3633), .B(n3632), .Z(n3705) );
  XOR U5292 ( .A(n3707), .B(n3706), .Z(n3634) );
  NAND U5293 ( .A(n3635), .B(n3634), .Z(n3637) );
  AND U5294 ( .A(\stack[1][6] ), .B(o[13]), .Z(n12305) );
  XOR U5295 ( .A(n3635), .B(n3634), .Z(n12304) );
  NAND U5296 ( .A(n12305), .B(n12304), .Z(n3636) );
  NAND U5297 ( .A(n3637), .B(n3636), .Z(n3638) );
  AND U5298 ( .A(\stack[1][6] ), .B(o[14]), .Z(n3639) );
  NAND U5299 ( .A(n3638), .B(n3639), .Z(n3711) );
  NAND U5300 ( .A(n3641), .B(n3640), .Z(n3645) );
  NAND U5301 ( .A(n3643), .B(n3642), .Z(n3644) );
  AND U5302 ( .A(n3645), .B(n3644), .Z(n3712) );
  NAND U5303 ( .A(\stack[1][8] ), .B(o[12]), .Z(n3713) );
  NAND U5304 ( .A(n3647), .B(n3646), .Z(n3651) );
  NAND U5305 ( .A(n3649), .B(n3648), .Z(n3650) );
  AND U5306 ( .A(n3651), .B(n3650), .Z(n3777) );
  NAND U5307 ( .A(o[10]), .B(\stack[1][10] ), .Z(n3719) );
  NAND U5308 ( .A(n3653), .B(n3652), .Z(n3657) );
  NAND U5309 ( .A(n3655), .B(n3654), .Z(n3656) );
  NAND U5310 ( .A(n3657), .B(n3656), .Z(n3718) );
  NAND U5311 ( .A(n3659), .B(n3658), .Z(n3663) );
  NAND U5312 ( .A(n3661), .B(n3660), .Z(n3662) );
  AND U5313 ( .A(n3663), .B(n3662), .Z(n3724) );
  NAND U5314 ( .A(o[8]), .B(\stack[1][12] ), .Z(n3725) );
  AND U5315 ( .A(o[6]), .B(\stack[1][14] ), .Z(n3733) );
  AND U5316 ( .A(o[5]), .B(\stack[1][15] ), .Z(n3761) );
  NAND U5317 ( .A(n3665), .B(n3664), .Z(n3669) );
  NAND U5318 ( .A(n3667), .B(n3666), .Z(n3668) );
  NAND U5319 ( .A(n3669), .B(n3668), .Z(n3759) );
  AND U5320 ( .A(o[0]), .B(\stack[1][17] ), .Z(n3671) );
  AND U5321 ( .A(n3671), .B(n3670), .Z(n3672) );
  NAND U5322 ( .A(o[2]), .B(n3672), .Z(n3676) );
  NAND U5323 ( .A(n3674), .B(n3673), .Z(n3675) );
  NAND U5324 ( .A(n3676), .B(n3675), .Z(n3737) );
  AND U5325 ( .A(o[1]), .B(\stack[1][19] ), .Z(n3745) );
  NAND U5326 ( .A(\stack[1][20] ), .B(o[0]), .Z(n3677) );
  XNOR U5327 ( .A(n3745), .B(n3677), .Z(n3748) );
  NAND U5328 ( .A(n3745), .B(o[0]), .Z(n3678) );
  XNOR U5329 ( .A(o[2]), .B(n3678), .Z(n3679) );
  AND U5330 ( .A(\stack[1][18] ), .B(n3679), .Z(n3749) );
  AND U5331 ( .A(o[3]), .B(\stack[1][17] ), .Z(n3739) );
  AND U5332 ( .A(o[4]), .B(\stack[1][16] ), .Z(n3752) );
  NAND U5333 ( .A(n3681), .B(n3680), .Z(n3685) );
  NAND U5334 ( .A(n3683), .B(n3682), .Z(n3684) );
  NAND U5335 ( .A(n3685), .B(n3684), .Z(n3753) );
  XOR U5336 ( .A(n3755), .B(n3754), .Z(n3758) );
  XOR U5337 ( .A(n3761), .B(n3760), .Z(n3730) );
  NAND U5338 ( .A(n3687), .B(n3686), .Z(n3691) );
  NAND U5339 ( .A(n3689), .B(n3688), .Z(n3690) );
  NAND U5340 ( .A(n3691), .B(n3690), .Z(n3731) );
  XOR U5341 ( .A(n3733), .B(n3732), .Z(n3764) );
  NAND U5342 ( .A(n3693), .B(n3692), .Z(n3697) );
  NAND U5343 ( .A(n3695), .B(n3694), .Z(n3696) );
  NAND U5344 ( .A(n3697), .B(n3696), .Z(n3765) );
  AND U5345 ( .A(o[7]), .B(\stack[1][13] ), .Z(n3766) );
  XNOR U5346 ( .A(n3767), .B(n3766), .Z(n3726) );
  XNOR U5347 ( .A(n3727), .B(n3726), .Z(n3771) );
  NAND U5348 ( .A(n3699), .B(n3698), .Z(n3703) );
  NAND U5349 ( .A(n3701), .B(n3700), .Z(n3702) );
  NAND U5350 ( .A(n3703), .B(n3702), .Z(n3770) );
  AND U5351 ( .A(\stack[1][11] ), .B(o[9]), .Z(n3772) );
  XNOR U5352 ( .A(n3773), .B(n3772), .Z(n3721) );
  XOR U5353 ( .A(n3777), .B(n3776), .Z(n3778) );
  NAND U5354 ( .A(\stack[1][9] ), .B(o[11]), .Z(n3779) );
  XNOR U5355 ( .A(n3715), .B(n3714), .Z(n3783) );
  NAND U5356 ( .A(n3705), .B(n3704), .Z(n3709) );
  NAND U5357 ( .A(n3707), .B(n3706), .Z(n3708) );
  NAND U5358 ( .A(n3709), .B(n3708), .Z(n3782) );
  AND U5359 ( .A(\stack[1][7] ), .B(o[13]), .Z(n3785) );
  NAND U5360 ( .A(n12311), .B(n12310), .Z(n3710) );
  NAND U5361 ( .A(n3711), .B(n3710), .Z(n3788) );
  NAND U5362 ( .A(n3713), .B(n3712), .Z(n3717) );
  NAND U5363 ( .A(n3715), .B(n3714), .Z(n3716) );
  AND U5364 ( .A(n3717), .B(n3716), .Z(n3793) );
  AND U5365 ( .A(\stack[1][10] ), .B(o[11]), .Z(n3807) );
  NAND U5366 ( .A(n3719), .B(n3718), .Z(n3723) );
  NAND U5367 ( .A(n3721), .B(n3720), .Z(n3722) );
  AND U5368 ( .A(n3723), .B(n3722), .Z(n3805) );
  NAND U5369 ( .A(n3725), .B(n3724), .Z(n3729) );
  NAND U5370 ( .A(n3727), .B(n3726), .Z(n3728) );
  NAND U5371 ( .A(n3729), .B(n3728), .Z(n3857) );
  NAND U5372 ( .A(n3731), .B(n3730), .Z(n3735) );
  NAND U5373 ( .A(n3733), .B(n3732), .Z(n3734) );
  NAND U5374 ( .A(n3735), .B(n3734), .Z(n3811) );
  AND U5375 ( .A(o[6]), .B(\stack[1][15] ), .Z(n3847) );
  NAND U5376 ( .A(n3737), .B(n3736), .Z(n3741) );
  NAND U5377 ( .A(n3739), .B(n3738), .Z(n3740) );
  NAND U5378 ( .A(n3741), .B(n3740), .Z(n3817) );
  AND U5379 ( .A(o[4]), .B(\stack[1][17] ), .Z(n3816) );
  AND U5380 ( .A(o[1]), .B(\stack[1][20] ), .Z(n3822) );
  NAND U5381 ( .A(\stack[1][21] ), .B(o[0]), .Z(n3742) );
  XNOR U5382 ( .A(n3822), .B(n3742), .Z(n3825) );
  NAND U5383 ( .A(n3822), .B(o[0]), .Z(n3743) );
  XNOR U5384 ( .A(o[2]), .B(n3743), .Z(n3744) );
  AND U5385 ( .A(\stack[1][19] ), .B(n3744), .Z(n3826) );
  AND U5386 ( .A(o[0]), .B(\stack[1][18] ), .Z(n3746) );
  AND U5387 ( .A(n3746), .B(n3745), .Z(n3747) );
  NAND U5388 ( .A(o[2]), .B(n3747), .Z(n3751) );
  NAND U5389 ( .A(n3749), .B(n3748), .Z(n3750) );
  NAND U5390 ( .A(n3751), .B(n3750), .Z(n3833) );
  AND U5391 ( .A(o[3]), .B(\stack[1][18] ), .Z(n3835) );
  XOR U5392 ( .A(n3819), .B(n3818), .Z(n3838) );
  AND U5393 ( .A(o[5]), .B(\stack[1][16] ), .Z(n3839) );
  NAND U5394 ( .A(n3753), .B(n3752), .Z(n3757) );
  NAND U5395 ( .A(n3755), .B(n3754), .Z(n3756) );
  NAND U5396 ( .A(n3757), .B(n3756), .Z(n3841) );
  NAND U5397 ( .A(n3759), .B(n3758), .Z(n3763) );
  NAND U5398 ( .A(n3761), .B(n3760), .Z(n3762) );
  NAND U5399 ( .A(n3763), .B(n3762), .Z(n3845) );
  XOR U5400 ( .A(n3847), .B(n3846), .Z(n3810) );
  AND U5401 ( .A(o[7]), .B(\stack[1][14] ), .Z(n3813) );
  AND U5402 ( .A(o[8]), .B(\stack[1][13] ), .Z(n3850) );
  NAND U5403 ( .A(n3765), .B(n3764), .Z(n3769) );
  NAND U5404 ( .A(n3767), .B(n3766), .Z(n3768) );
  NAND U5405 ( .A(n3769), .B(n3768), .Z(n3851) );
  XNOR U5406 ( .A(n3853), .B(n3852), .Z(n3856) );
  NAND U5407 ( .A(o[9]), .B(\stack[1][12] ), .Z(n3858) );
  XNOR U5408 ( .A(n3859), .B(n3858), .Z(n3865) );
  AND U5409 ( .A(o[10]), .B(\stack[1][11] ), .Z(n3862) );
  NAND U5410 ( .A(n3771), .B(n3770), .Z(n3775) );
  NAND U5411 ( .A(n3773), .B(n3772), .Z(n3774) );
  NAND U5412 ( .A(n3775), .B(n3774), .Z(n3863) );
  XOR U5413 ( .A(n3805), .B(n3804), .Z(n3806) );
  XOR U5414 ( .A(n3807), .B(n3806), .Z(n3801) );
  AND U5415 ( .A(\stack[1][9] ), .B(o[12]), .Z(n3798) );
  NAND U5416 ( .A(n3777), .B(n3776), .Z(n3781) );
  NAND U5417 ( .A(n3779), .B(n3778), .Z(n3780) );
  AND U5418 ( .A(n3781), .B(n3780), .Z(n3799) );
  XOR U5419 ( .A(n3801), .B(n3800), .Z(n3792) );
  XOR U5420 ( .A(n3793), .B(n3792), .Z(n3794) );
  AND U5421 ( .A(\stack[1][8] ), .B(o[13]), .Z(n3795) );
  AND U5422 ( .A(\stack[1][7] ), .B(o[14]), .Z(n3868) );
  NAND U5423 ( .A(n3783), .B(n3782), .Z(n3787) );
  NAND U5424 ( .A(n3785), .B(n3784), .Z(n3786) );
  NAND U5425 ( .A(n3787), .B(n3786), .Z(n3869) );
  XOR U5426 ( .A(n3871), .B(n3870), .Z(n3789) );
  NAND U5427 ( .A(n3788), .B(n3789), .Z(n3791) );
  AND U5428 ( .A(\stack[1][6] ), .B(o[15]), .Z(n12317) );
  NAND U5429 ( .A(n12317), .B(n12316), .Z(n3790) );
  AND U5430 ( .A(n3791), .B(n3790), .Z(n3875) );
  NAND U5431 ( .A(n3874), .B(n3875), .Z(n3877) );
  NAND U5432 ( .A(n3793), .B(n3792), .Z(n3797) );
  NAND U5433 ( .A(n3795), .B(n3794), .Z(n3796) );
  NAND U5434 ( .A(n3797), .B(n3796), .Z(n3879) );
  AND U5435 ( .A(\stack[1][8] ), .B(o[14]), .Z(n3878) );
  NAND U5436 ( .A(n3799), .B(n3798), .Z(n3803) );
  NAND U5437 ( .A(n3801), .B(n3800), .Z(n3802) );
  NAND U5438 ( .A(n3803), .B(n3802), .Z(n3954) );
  NAND U5439 ( .A(n3805), .B(n3804), .Z(n3809) );
  NAND U5440 ( .A(n3807), .B(n3806), .Z(n3808) );
  AND U5441 ( .A(n3809), .B(n3808), .Z(n3884) );
  NAND U5442 ( .A(\stack[1][10] ), .B(o[12]), .Z(n3885) );
  NAND U5443 ( .A(\stack[1][11] ), .B(o[11]), .Z(n16907) );
  NAND U5444 ( .A(n3811), .B(n3810), .Z(n3815) );
  NAND U5445 ( .A(n3813), .B(n3812), .Z(n3814) );
  NAND U5446 ( .A(n3815), .B(n3814), .Z(n3897) );
  AND U5447 ( .A(o[8]), .B(\stack[1][14] ), .Z(n3896) );
  AND U5448 ( .A(o[5]), .B(\stack[1][17] ), .Z(n3933) );
  NAND U5449 ( .A(n3817), .B(n3816), .Z(n3821) );
  NAND U5450 ( .A(n3819), .B(n3818), .Z(n3820) );
  NAND U5451 ( .A(n3821), .B(n3820), .Z(n3931) );
  AND U5452 ( .A(o[3]), .B(\stack[1][19] ), .Z(n3911) );
  AND U5453 ( .A(o[0]), .B(\stack[1][19] ), .Z(n3823) );
  AND U5454 ( .A(n3823), .B(n3822), .Z(n3824) );
  NAND U5455 ( .A(o[2]), .B(n3824), .Z(n3828) );
  NAND U5456 ( .A(n3826), .B(n3825), .Z(n3827) );
  NAND U5457 ( .A(n3828), .B(n3827), .Z(n3909) );
  AND U5458 ( .A(o[1]), .B(\stack[1][21] ), .Z(n3917) );
  NAND U5459 ( .A(\stack[1][22] ), .B(o[0]), .Z(n3829) );
  XNOR U5460 ( .A(n3917), .B(n3829), .Z(n3920) );
  NAND U5461 ( .A(n3917), .B(o[0]), .Z(n3830) );
  XNOR U5462 ( .A(o[2]), .B(n3830), .Z(n3831) );
  AND U5463 ( .A(\stack[1][20] ), .B(n3831), .Z(n3921) );
  XOR U5464 ( .A(n3911), .B(n3910), .Z(n3927) );
  AND U5465 ( .A(o[4]), .B(\stack[1][18] ), .Z(n3924) );
  NAND U5466 ( .A(n3833), .B(n3832), .Z(n3837) );
  NAND U5467 ( .A(n3835), .B(n3834), .Z(n3836) );
  NAND U5468 ( .A(n3837), .B(n3836), .Z(n3925) );
  XOR U5469 ( .A(n3927), .B(n3926), .Z(n3930) );
  XOR U5470 ( .A(n3933), .B(n3932), .Z(n3902) );
  NAND U5471 ( .A(n3839), .B(n3838), .Z(n3843) );
  NAND U5472 ( .A(n3841), .B(n3840), .Z(n3842) );
  NAND U5473 ( .A(n3843), .B(n3842), .Z(n3903) );
  AND U5474 ( .A(o[6]), .B(\stack[1][16] ), .Z(n3905) );
  NAND U5475 ( .A(n3845), .B(n3844), .Z(n3849) );
  NAND U5476 ( .A(n3847), .B(n3846), .Z(n3848) );
  NAND U5477 ( .A(n3849), .B(n3848), .Z(n3937) );
  AND U5478 ( .A(o[7]), .B(\stack[1][15] ), .Z(n3939) );
  XOR U5479 ( .A(n3899), .B(n3898), .Z(n3942) );
  NAND U5480 ( .A(n3851), .B(n3850), .Z(n3855) );
  NAND U5481 ( .A(n3853), .B(n3852), .Z(n3854) );
  NAND U5482 ( .A(n3855), .B(n3854), .Z(n3943) );
  AND U5483 ( .A(o[9]), .B(\stack[1][13] ), .Z(n3945) );
  NAND U5484 ( .A(n3857), .B(n3856), .Z(n3861) );
  NAND U5485 ( .A(n3859), .B(n3858), .Z(n3860) );
  AND U5486 ( .A(n3861), .B(n3860), .Z(n3890) );
  AND U5487 ( .A(o[10]), .B(\stack[1][12] ), .Z(n3891) );
  XNOR U5488 ( .A(n3893), .B(n3892), .Z(n3949) );
  NAND U5489 ( .A(n3863), .B(n3862), .Z(n3867) );
  NAND U5490 ( .A(n3865), .B(n3864), .Z(n3866) );
  AND U5491 ( .A(n3867), .B(n3866), .Z(n3948) );
  XNOR U5492 ( .A(n3887), .B(n3886), .Z(n3953) );
  AND U5493 ( .A(\stack[1][9] ), .B(o[13]), .Z(n3956) );
  XOR U5494 ( .A(n3881), .B(n3880), .Z(n3959) );
  NAND U5495 ( .A(n3869), .B(n3868), .Z(n3873) );
  NAND U5496 ( .A(n3871), .B(n3870), .Z(n3872) );
  NAND U5497 ( .A(n3873), .B(n3872), .Z(n3960) );
  AND U5498 ( .A(\stack[1][7] ), .B(o[15]), .Z(n3961) );
  XNOR U5499 ( .A(n3962), .B(n3961), .Z(n12229) );
  NAND U5500 ( .A(n12229), .B(n12230), .Z(n3876) );
  AND U5501 ( .A(n3877), .B(n3876), .Z(n3966) );
  NAND U5502 ( .A(n3879), .B(n3878), .Z(n3883) );
  NAND U5503 ( .A(n3881), .B(n3880), .Z(n3882) );
  NAND U5504 ( .A(n3883), .B(n3882), .Z(n3972) );
  NAND U5505 ( .A(n3885), .B(n3884), .Z(n3889) );
  NAND U5506 ( .A(n3887), .B(n3886), .Z(n3888) );
  NAND U5507 ( .A(n3889), .B(n3888), .Z(n3978) );
  NAND U5508 ( .A(n3891), .B(n3890), .Z(n3895) );
  NAND U5509 ( .A(n3893), .B(n3892), .Z(n3894) );
  NAND U5510 ( .A(n3895), .B(n3894), .Z(n3990) );
  NAND U5511 ( .A(n3897), .B(n3896), .Z(n3901) );
  NAND U5512 ( .A(n3899), .B(n3898), .Z(n3900) );
  AND U5513 ( .A(n3901), .B(n3900), .Z(n4041) );
  AND U5514 ( .A(o[7]), .B(\stack[1][16] ), .Z(n3998) );
  NAND U5515 ( .A(n3903), .B(n3902), .Z(n3907) );
  NAND U5516 ( .A(n3905), .B(n3904), .Z(n3906) );
  NAND U5517 ( .A(n3907), .B(n3906), .Z(n3996) );
  AND U5518 ( .A(o[6]), .B(\stack[1][17] ), .Z(n4032) );
  NAND U5519 ( .A(n3909), .B(n3908), .Z(n3913) );
  NAND U5520 ( .A(n3911), .B(n3910), .Z(n3912) );
  AND U5521 ( .A(n3913), .B(n3912), .Z(n4001) );
  NAND U5522 ( .A(o[4]), .B(\stack[1][19] ), .Z(n4002) );
  AND U5523 ( .A(\stack[1][22] ), .B(o[1]), .Z(n4007) );
  NAND U5524 ( .A(n4007), .B(o[0]), .Z(n3914) );
  XNOR U5525 ( .A(o[2]), .B(n3914), .Z(n3915) );
  AND U5526 ( .A(\stack[1][21] ), .B(n3915), .Z(n4010) );
  NAND U5527 ( .A(\stack[1][23] ), .B(o[0]), .Z(n3916) );
  XNOR U5528 ( .A(n4007), .B(n3916), .Z(n4011) );
  AND U5529 ( .A(o[0]), .B(\stack[1][20] ), .Z(n3918) );
  AND U5530 ( .A(n3918), .B(n3917), .Z(n3919) );
  NAND U5531 ( .A(o[2]), .B(n3919), .Z(n3923) );
  NAND U5532 ( .A(n3921), .B(n3920), .Z(n3922) );
  NAND U5533 ( .A(n3923), .B(n3922), .Z(n4018) );
  AND U5534 ( .A(o[3]), .B(\stack[1][20] ), .Z(n4019) );
  XNOR U5535 ( .A(n4020), .B(n4019), .Z(n4003) );
  XNOR U5536 ( .A(n4004), .B(n4003), .Z(n4024) );
  AND U5537 ( .A(o[5]), .B(\stack[1][18] ), .Z(n4023) );
  NAND U5538 ( .A(n3925), .B(n3924), .Z(n3929) );
  NAND U5539 ( .A(n3927), .B(n3926), .Z(n3928) );
  NAND U5540 ( .A(n3929), .B(n3928), .Z(n4026) );
  NAND U5541 ( .A(n3931), .B(n3930), .Z(n3935) );
  NAND U5542 ( .A(n3933), .B(n3932), .Z(n3934) );
  NAND U5543 ( .A(n3935), .B(n3934), .Z(n4030) );
  XOR U5544 ( .A(n4032), .B(n4031), .Z(n3995) );
  XOR U5545 ( .A(n3998), .B(n3997), .Z(n4038) );
  AND U5546 ( .A(o[8]), .B(\stack[1][15] ), .Z(n4035) );
  NAND U5547 ( .A(n3937), .B(n3936), .Z(n3941) );
  NAND U5548 ( .A(n3939), .B(n3938), .Z(n3940) );
  NAND U5549 ( .A(n3941), .B(n3940), .Z(n4036) );
  XNOR U5550 ( .A(n4038), .B(n4037), .Z(n4042) );
  NAND U5551 ( .A(o[9]), .B(\stack[1][14] ), .Z(n4043) );
  XNOR U5552 ( .A(n4044), .B(n4043), .Z(n4050) );
  AND U5553 ( .A(o[10]), .B(\stack[1][13] ), .Z(n4047) );
  NAND U5554 ( .A(n3943), .B(n3942), .Z(n3947) );
  NAND U5555 ( .A(n3945), .B(n3944), .Z(n3946) );
  NAND U5556 ( .A(n3947), .B(n3946), .Z(n4048) );
  AND U5557 ( .A(\stack[1][12] ), .B(o[11]), .Z(n3992) );
  AND U5558 ( .A(\stack[1][11] ), .B(o[12]), .Z(n3983) );
  NAND U5559 ( .A(n3949), .B(n3948), .Z(n3952) );
  NAND U5560 ( .A(n16907), .B(n3950), .Z(n3951) );
  AND U5561 ( .A(n3952), .B(n3951), .Z(n3984) );
  XNOR U5562 ( .A(n3986), .B(n3985), .Z(n3977) );
  NAND U5563 ( .A(\stack[1][10] ), .B(o[13]), .Z(n3979) );
  XNOR U5564 ( .A(n3980), .B(n3979), .Z(n4056) );
  AND U5565 ( .A(\stack[1][9] ), .B(o[14]), .Z(n4053) );
  NAND U5566 ( .A(n3954), .B(n3953), .Z(n3958) );
  NAND U5567 ( .A(n3956), .B(n3955), .Z(n3957) );
  NAND U5568 ( .A(n3958), .B(n3957), .Z(n4054) );
  AND U5569 ( .A(\stack[1][8] ), .B(o[15]), .Z(n3974) );
  AND U5570 ( .A(\stack[1][7] ), .B(o[16]), .Z(n4059) );
  NAND U5571 ( .A(n3960), .B(n3959), .Z(n3964) );
  NAND U5572 ( .A(n3962), .B(n3961), .Z(n3963) );
  NAND U5573 ( .A(n3964), .B(n3963), .Z(n4060) );
  XOR U5574 ( .A(n4062), .B(n4061), .Z(n3965) );
  NAND U5575 ( .A(n3966), .B(n3965), .Z(n3968) );
  AND U5576 ( .A(\stack[1][6] ), .B(o[17]), .Z(n12326) );
  XOR U5577 ( .A(n3966), .B(n3965), .Z(n12327) );
  NAND U5578 ( .A(n12326), .B(n12327), .Z(n3967) );
  NAND U5579 ( .A(n3968), .B(n3967), .Z(n3969) );
  AND U5580 ( .A(\stack[1][6] ), .B(o[18]), .Z(n3970) );
  NAND U5581 ( .A(n3969), .B(n3970), .Z(n4066) );
  NAND U5582 ( .A(n3972), .B(n3971), .Z(n3976) );
  NAND U5583 ( .A(n3974), .B(n3973), .Z(n3975) );
  NAND U5584 ( .A(n3976), .B(n3975), .Z(n4068) );
  AND U5585 ( .A(\stack[1][8] ), .B(o[16]), .Z(n4067) );
  NAND U5586 ( .A(n3978), .B(n3977), .Z(n3982) );
  NAND U5587 ( .A(n3980), .B(n3979), .Z(n3981) );
  AND U5588 ( .A(n3982), .B(n3981), .Z(n4073) );
  AND U5589 ( .A(\stack[1][10] ), .B(o[14]), .Z(n4074) );
  NAND U5590 ( .A(n3984), .B(n3983), .Z(n3988) );
  NAND U5591 ( .A(n3986), .B(n3985), .Z(n3987) );
  NAND U5592 ( .A(n3988), .B(n3987), .Z(n4150) );
  NAND U5593 ( .A(\stack[1][12] ), .B(o[12]), .Z(n4080) );
  IV U5594 ( .A(n4080), .Z(n16868) );
  NAND U5595 ( .A(n3990), .B(n3989), .Z(n3994) );
  NAND U5596 ( .A(n3992), .B(n3991), .Z(n3993) );
  AND U5597 ( .A(n3994), .B(n3993), .Z(n4079) );
  XNOR U5598 ( .A(n16868), .B(n4079), .Z(n4082) );
  NAND U5599 ( .A(n3996), .B(n3995), .Z(n4000) );
  NAND U5600 ( .A(n3998), .B(n3997), .Z(n3999) );
  NAND U5601 ( .A(n4000), .B(n3999), .Z(n4092) );
  AND U5602 ( .A(o[8]), .B(\stack[1][16] ), .Z(n4091) );
  AND U5603 ( .A(o[6]), .B(\stack[1][18] ), .Z(n4100) );
  NAND U5604 ( .A(n4002), .B(n4001), .Z(n4006) );
  NAND U5605 ( .A(n4004), .B(n4003), .Z(n4005) );
  AND U5606 ( .A(n4006), .B(n4005), .Z(n4126) );
  AND U5607 ( .A(o[3]), .B(\stack[1][21] ), .Z(n4106) );
  AND U5608 ( .A(o[0]), .B(\stack[1][21] ), .Z(n4008) );
  AND U5609 ( .A(n4008), .B(n4007), .Z(n4009) );
  NAND U5610 ( .A(o[2]), .B(n4009), .Z(n4013) );
  NAND U5611 ( .A(n4011), .B(n4010), .Z(n4012) );
  NAND U5612 ( .A(n4013), .B(n4012), .Z(n4104) );
  AND U5613 ( .A(o[1]), .B(\stack[1][23] ), .Z(n4112) );
  NAND U5614 ( .A(\stack[1][24] ), .B(o[0]), .Z(n4014) );
  XNOR U5615 ( .A(n4112), .B(n4014), .Z(n4115) );
  NAND U5616 ( .A(n4112), .B(o[0]), .Z(n4015) );
  XNOR U5617 ( .A(o[2]), .B(n4015), .Z(n4016) );
  AND U5618 ( .A(\stack[1][22] ), .B(n4016), .Z(n4116) );
  XOR U5619 ( .A(n4106), .B(n4105), .Z(n4122) );
  AND U5620 ( .A(o[4]), .B(\stack[1][20] ), .Z(n4119) );
  NAND U5621 ( .A(n4018), .B(n4017), .Z(n4022) );
  NAND U5622 ( .A(n4020), .B(n4019), .Z(n4021) );
  NAND U5623 ( .A(n4022), .B(n4021), .Z(n4120) );
  XOR U5624 ( .A(n4122), .B(n4121), .Z(n4125) );
  XOR U5625 ( .A(n4126), .B(n4125), .Z(n4127) );
  AND U5626 ( .A(o[5]), .B(\stack[1][19] ), .Z(n4128) );
  NAND U5627 ( .A(n4024), .B(n4023), .Z(n4028) );
  NAND U5628 ( .A(n4026), .B(n4025), .Z(n4027) );
  NAND U5629 ( .A(n4028), .B(n4027), .Z(n4098) );
  XOR U5630 ( .A(n4100), .B(n4099), .Z(n4131) );
  NAND U5631 ( .A(n4030), .B(n4029), .Z(n4034) );
  NAND U5632 ( .A(n4032), .B(n4031), .Z(n4033) );
  NAND U5633 ( .A(n4034), .B(n4033), .Z(n4132) );
  AND U5634 ( .A(o[7]), .B(\stack[1][17] ), .Z(n4134) );
  XOR U5635 ( .A(n4094), .B(n4093), .Z(n4137) );
  NAND U5636 ( .A(n4036), .B(n4035), .Z(n4040) );
  NAND U5637 ( .A(n4038), .B(n4037), .Z(n4039) );
  NAND U5638 ( .A(n4040), .B(n4039), .Z(n4138) );
  AND U5639 ( .A(o[9]), .B(\stack[1][15] ), .Z(n4140) );
  NAND U5640 ( .A(n4042), .B(n4041), .Z(n4046) );
  NAND U5641 ( .A(n4044), .B(n4043), .Z(n4045) );
  AND U5642 ( .A(n4046), .B(n4045), .Z(n4085) );
  AND U5643 ( .A(o[10]), .B(\stack[1][14] ), .Z(n4086) );
  XNOR U5644 ( .A(n4088), .B(n4087), .Z(n4144) );
  NAND U5645 ( .A(n4048), .B(n4047), .Z(n4052) );
  NAND U5646 ( .A(n4050), .B(n4049), .Z(n4051) );
  AND U5647 ( .A(n4052), .B(n4051), .Z(n4143) );
  NAND U5648 ( .A(\stack[1][13] ), .B(o[11]), .Z(n4146) );
  XNOR U5649 ( .A(n4082), .B(n4081), .Z(n4149) );
  AND U5650 ( .A(\stack[1][11] ), .B(o[13]), .Z(n4152) );
  XOR U5651 ( .A(n4076), .B(n4075), .Z(n4155) );
  NAND U5652 ( .A(n4054), .B(n4053), .Z(n4058) );
  NAND U5653 ( .A(n4056), .B(n4055), .Z(n4057) );
  NAND U5654 ( .A(n4058), .B(n4057), .Z(n4156) );
  AND U5655 ( .A(\stack[1][9] ), .B(o[15]), .Z(n4158) );
  XOR U5656 ( .A(n4070), .B(n4069), .Z(n4161) );
  NAND U5657 ( .A(n4060), .B(n4059), .Z(n4064) );
  NAND U5658 ( .A(n4062), .B(n4061), .Z(n4063) );
  NAND U5659 ( .A(n4064), .B(n4063), .Z(n4162) );
  AND U5660 ( .A(\stack[1][7] ), .B(o[17]), .Z(n4164) );
  NAND U5661 ( .A(n12333), .B(n12332), .Z(n4065) );
  NAND U5662 ( .A(n4066), .B(n4065), .Z(n4167) );
  NAND U5663 ( .A(n4068), .B(n4067), .Z(n4072) );
  NAND U5664 ( .A(n4070), .B(n4069), .Z(n4071) );
  NAND U5665 ( .A(n4072), .B(n4071), .Z(n4174) );
  NAND U5666 ( .A(n4074), .B(n4073), .Z(n4078) );
  NAND U5667 ( .A(n4076), .B(n4075), .Z(n4077) );
  NAND U5668 ( .A(n4078), .B(n4077), .Z(n4180) );
  NAND U5669 ( .A(\stack[1][12] ), .B(o[13]), .Z(n4188) );
  NAND U5670 ( .A(n4080), .B(n4079), .Z(n4084) );
  NAND U5671 ( .A(n4082), .B(n4081), .Z(n4083) );
  NAND U5672 ( .A(n4084), .B(n4083), .Z(n4186) );
  AND U5673 ( .A(o[11]), .B(\stack[1][14] ), .Z(n4252) );
  NAND U5674 ( .A(n4086), .B(n4085), .Z(n4090) );
  NAND U5675 ( .A(n4088), .B(n4087), .Z(n4089) );
  NAND U5676 ( .A(n4090), .B(n4089), .Z(n4250) );
  NAND U5677 ( .A(n4092), .B(n4091), .Z(n4096) );
  NAND U5678 ( .A(n4094), .B(n4093), .Z(n4095) );
  AND U5679 ( .A(n4096), .B(n4095), .Z(n4197) );
  AND U5680 ( .A(o[7]), .B(\stack[1][18] ), .Z(n4240) );
  NAND U5681 ( .A(n4098), .B(n4097), .Z(n4102) );
  NAND U5682 ( .A(n4100), .B(n4099), .Z(n4101) );
  NAND U5683 ( .A(n4102), .B(n4101), .Z(n4238) );
  AND U5684 ( .A(o[6]), .B(\stack[1][19] ), .Z(n4234) );
  NAND U5685 ( .A(n4104), .B(n4103), .Z(n4108) );
  NAND U5686 ( .A(n4106), .B(n4105), .Z(n4107) );
  NAND U5687 ( .A(n4108), .B(n4107), .Z(n4204) );
  AND U5688 ( .A(o[4]), .B(\stack[1][21] ), .Z(n4203) );
  AND U5689 ( .A(o[1]), .B(\stack[1][24] ), .Z(n4209) );
  NAND U5690 ( .A(\stack[1][25] ), .B(o[0]), .Z(n4109) );
  XNOR U5691 ( .A(n4209), .B(n4109), .Z(n4212) );
  NAND U5692 ( .A(n4209), .B(o[0]), .Z(n4110) );
  XNOR U5693 ( .A(o[2]), .B(n4110), .Z(n4111) );
  AND U5694 ( .A(\stack[1][23] ), .B(n4111), .Z(n4213) );
  AND U5695 ( .A(o[0]), .B(\stack[1][22] ), .Z(n4113) );
  AND U5696 ( .A(n4113), .B(n4112), .Z(n4114) );
  NAND U5697 ( .A(o[2]), .B(n4114), .Z(n4118) );
  NAND U5698 ( .A(n4116), .B(n4115), .Z(n4117) );
  NAND U5699 ( .A(n4118), .B(n4117), .Z(n4220) );
  AND U5700 ( .A(o[3]), .B(\stack[1][22] ), .Z(n4222) );
  XOR U5701 ( .A(n4206), .B(n4205), .Z(n4225) );
  AND U5702 ( .A(o[5]), .B(\stack[1][20] ), .Z(n4226) );
  NAND U5703 ( .A(n4120), .B(n4119), .Z(n4124) );
  NAND U5704 ( .A(n4122), .B(n4121), .Z(n4123) );
  NAND U5705 ( .A(n4124), .B(n4123), .Z(n4228) );
  NAND U5706 ( .A(n4126), .B(n4125), .Z(n4130) );
  NAND U5707 ( .A(n4128), .B(n4127), .Z(n4129) );
  NAND U5708 ( .A(n4130), .B(n4129), .Z(n4232) );
  XOR U5709 ( .A(n4234), .B(n4233), .Z(n4237) );
  XOR U5710 ( .A(n4240), .B(n4239), .Z(n4246) );
  AND U5711 ( .A(o[8]), .B(\stack[1][17] ), .Z(n4243) );
  NAND U5712 ( .A(n4132), .B(n4131), .Z(n4136) );
  NAND U5713 ( .A(n4134), .B(n4133), .Z(n4135) );
  NAND U5714 ( .A(n4136), .B(n4135), .Z(n4244) );
  XNOR U5715 ( .A(n4246), .B(n4245), .Z(n4198) );
  NAND U5716 ( .A(o[9]), .B(\stack[1][16] ), .Z(n4199) );
  XNOR U5717 ( .A(n4200), .B(n4199), .Z(n4194) );
  AND U5718 ( .A(o[10]), .B(\stack[1][15] ), .Z(n4191) );
  NAND U5719 ( .A(n4138), .B(n4137), .Z(n4142) );
  NAND U5720 ( .A(n4140), .B(n4139), .Z(n4141) );
  NAND U5721 ( .A(n4142), .B(n4141), .Z(n4192) );
  XOR U5722 ( .A(n4252), .B(n4251), .Z(n4258) );
  AND U5723 ( .A(\stack[1][13] ), .B(o[12]), .Z(n4255) );
  NAND U5724 ( .A(n4144), .B(n4143), .Z(n4148) );
  NAND U5725 ( .A(n4146), .B(n4145), .Z(n4147) );
  AND U5726 ( .A(n4148), .B(n4147), .Z(n4256) );
  XNOR U5727 ( .A(n4258), .B(n4257), .Z(n4185) );
  AND U5728 ( .A(\stack[1][11] ), .B(o[14]), .Z(n4261) );
  NAND U5729 ( .A(n4150), .B(n4149), .Z(n4154) );
  NAND U5730 ( .A(n4152), .B(n4151), .Z(n4153) );
  NAND U5731 ( .A(n4154), .B(n4153), .Z(n4262) );
  XOR U5732 ( .A(n4263), .B(n4264), .Z(n4179) );
  AND U5733 ( .A(\stack[1][10] ), .B(o[15]), .Z(n4182) );
  AND U5734 ( .A(\stack[1][9] ), .B(o[16]), .Z(n4267) );
  NAND U5735 ( .A(n4156), .B(n4155), .Z(n4160) );
  NAND U5736 ( .A(n4158), .B(n4157), .Z(n4159) );
  NAND U5737 ( .A(n4160), .B(n4159), .Z(n4268) );
  XOR U5738 ( .A(n4270), .B(n4269), .Z(n4173) );
  AND U5739 ( .A(\stack[1][8] ), .B(o[17]), .Z(n4176) );
  AND U5740 ( .A(\stack[1][7] ), .B(o[18]), .Z(n4273) );
  NAND U5741 ( .A(n4162), .B(n4161), .Z(n4166) );
  NAND U5742 ( .A(n4164), .B(n4163), .Z(n4165) );
  NAND U5743 ( .A(n4166), .B(n4165), .Z(n4274) );
  XOR U5744 ( .A(n4276), .B(n4275), .Z(n4168) );
  NAND U5745 ( .A(n4167), .B(n4168), .Z(n4170) );
  AND U5746 ( .A(\stack[1][6] ), .B(o[19]), .Z(n12338) );
  NAND U5747 ( .A(n12338), .B(n12339), .Z(n4169) );
  NAND U5748 ( .A(n4170), .B(n4169), .Z(n4171) );
  AND U5749 ( .A(\stack[1][6] ), .B(o[20]), .Z(n4172) );
  NAND U5750 ( .A(n4171), .B(n4172), .Z(n4280) );
  NAND U5751 ( .A(n4174), .B(n4173), .Z(n4178) );
  NAND U5752 ( .A(n4176), .B(n4175), .Z(n4177) );
  NAND U5753 ( .A(n4178), .B(n4177), .Z(n4282) );
  AND U5754 ( .A(\stack[1][8] ), .B(o[18]), .Z(n4281) );
  NAND U5755 ( .A(n4180), .B(n4179), .Z(n4184) );
  NAND U5756 ( .A(n4182), .B(n4181), .Z(n4183) );
  NAND U5757 ( .A(n4184), .B(n4183), .Z(n4288) );
  AND U5758 ( .A(\stack[1][10] ), .B(o[16]), .Z(n4287) );
  NAND U5759 ( .A(n4186), .B(n4185), .Z(n4190) );
  NAND U5760 ( .A(n4188), .B(n4187), .Z(n4189) );
  AND U5761 ( .A(n4190), .B(n4189), .Z(n4293) );
  AND U5762 ( .A(\stack[1][12] ), .B(o[14]), .Z(n4294) );
  AND U5763 ( .A(\stack[1][13] ), .B(o[13]), .Z(n16829) );
  NAND U5764 ( .A(n4192), .B(n4191), .Z(n4196) );
  NAND U5765 ( .A(n4194), .B(n4193), .Z(n4195) );
  AND U5766 ( .A(n4196), .B(n4195), .Z(n4364) );
  NAND U5767 ( .A(n4198), .B(n4197), .Z(n4202) );
  NAND U5768 ( .A(n4200), .B(n4199), .Z(n4201) );
  NAND U5769 ( .A(n4202), .B(n4201), .Z(n4306) );
  NAND U5770 ( .A(o[10]), .B(\stack[1][16] ), .Z(n4305) );
  NAND U5771 ( .A(n4204), .B(n4203), .Z(n4208) );
  NAND U5772 ( .A(n4206), .B(n4205), .Z(n4207) );
  NAND U5773 ( .A(n4208), .B(n4207), .Z(n4346) );
  AND U5774 ( .A(o[3]), .B(\stack[1][23] ), .Z(n4326) );
  AND U5775 ( .A(o[0]), .B(\stack[1][23] ), .Z(n4210) );
  AND U5776 ( .A(n4210), .B(n4209), .Z(n4211) );
  NAND U5777 ( .A(o[2]), .B(n4211), .Z(n4215) );
  NAND U5778 ( .A(n4213), .B(n4212), .Z(n4214) );
  NAND U5779 ( .A(n4215), .B(n4214), .Z(n4324) );
  AND U5780 ( .A(o[1]), .B(\stack[1][25] ), .Z(n4332) );
  NAND U5781 ( .A(\stack[1][26] ), .B(o[0]), .Z(n4216) );
  XNOR U5782 ( .A(n4332), .B(n4216), .Z(n4335) );
  NAND U5783 ( .A(n4332), .B(o[0]), .Z(n4217) );
  XNOR U5784 ( .A(o[2]), .B(n4217), .Z(n4218) );
  AND U5785 ( .A(\stack[1][24] ), .B(n4218), .Z(n4336) );
  XOR U5786 ( .A(n4326), .B(n4325), .Z(n4342) );
  AND U5787 ( .A(o[4]), .B(\stack[1][22] ), .Z(n4339) );
  NAND U5788 ( .A(n4220), .B(n4219), .Z(n4224) );
  NAND U5789 ( .A(n4222), .B(n4221), .Z(n4223) );
  NAND U5790 ( .A(n4224), .B(n4223), .Z(n4340) );
  XOR U5791 ( .A(n4342), .B(n4341), .Z(n4345) );
  AND U5792 ( .A(o[5]), .B(\stack[1][21] ), .Z(n4348) );
  NAND U5793 ( .A(n4226), .B(n4225), .Z(n4230) );
  NAND U5794 ( .A(n4228), .B(n4227), .Z(n4229) );
  NAND U5795 ( .A(n4230), .B(n4229), .Z(n4318) );
  AND U5796 ( .A(o[6]), .B(\stack[1][20] ), .Z(n4320) );
  NAND U5797 ( .A(n4232), .B(n4231), .Z(n4236) );
  NAND U5798 ( .A(n4234), .B(n4233), .Z(n4235) );
  NAND U5799 ( .A(n4236), .B(n4235), .Z(n4352) );
  AND U5800 ( .A(o[7]), .B(\stack[1][19] ), .Z(n4354) );
  NAND U5801 ( .A(n4238), .B(n4237), .Z(n4242) );
  NAND U5802 ( .A(n4240), .B(n4239), .Z(n4241) );
  NAND U5803 ( .A(n4242), .B(n4241), .Z(n4312) );
  AND U5804 ( .A(o[8]), .B(\stack[1][18] ), .Z(n4311) );
  XOR U5805 ( .A(n4314), .B(n4313), .Z(n4357) );
  NAND U5806 ( .A(n4244), .B(n4243), .Z(n4248) );
  NAND U5807 ( .A(n4246), .B(n4245), .Z(n4247) );
  NAND U5808 ( .A(n4248), .B(n4247), .Z(n4358) );
  AND U5809 ( .A(o[9]), .B(\stack[1][17] ), .Z(n4359) );
  XNOR U5810 ( .A(n4360), .B(n4359), .Z(n4308) );
  XOR U5811 ( .A(n4364), .B(n4363), .Z(n4365) );
  NAND U5812 ( .A(o[11]), .B(\stack[1][15] ), .Z(n4366) );
  NAND U5813 ( .A(n4250), .B(n4249), .Z(n4254) );
  NAND U5814 ( .A(n4252), .B(n4251), .Z(n4253) );
  AND U5815 ( .A(n4254), .B(n4253), .Z(n4299) );
  NAND U5816 ( .A(o[12]), .B(\stack[1][14] ), .Z(n4300) );
  XNOR U5817 ( .A(n4302), .B(n4301), .Z(n4370) );
  NAND U5818 ( .A(n4256), .B(n4255), .Z(n4260) );
  NAND U5819 ( .A(n4258), .B(n4257), .Z(n4259) );
  NAND U5820 ( .A(n4260), .B(n4259), .Z(n4369) );
  XOR U5821 ( .A(n16829), .B(n4371), .Z(n4295) );
  XOR U5822 ( .A(n4296), .B(n4295), .Z(n4374) );
  NAND U5823 ( .A(n4262), .B(n4261), .Z(n4266) );
  NAND U5824 ( .A(n4264), .B(n4263), .Z(n4265) );
  NAND U5825 ( .A(n4266), .B(n4265), .Z(n4375) );
  AND U5826 ( .A(\stack[1][11] ), .B(o[15]), .Z(n4377) );
  XOR U5827 ( .A(n4290), .B(n4289), .Z(n4380) );
  NAND U5828 ( .A(n4268), .B(n4267), .Z(n4272) );
  NAND U5829 ( .A(n4270), .B(n4269), .Z(n4271) );
  NAND U5830 ( .A(n4272), .B(n4271), .Z(n4381) );
  AND U5831 ( .A(\stack[1][9] ), .B(o[17]), .Z(n4383) );
  XOR U5832 ( .A(n4284), .B(n4283), .Z(n4386) );
  NAND U5833 ( .A(n4274), .B(n4273), .Z(n4278) );
  NAND U5834 ( .A(n4276), .B(n4275), .Z(n4277) );
  NAND U5835 ( .A(n4278), .B(n4277), .Z(n4387) );
  AND U5836 ( .A(\stack[1][7] ), .B(o[19]), .Z(n4389) );
  NAND U5837 ( .A(n12345), .B(n12344), .Z(n4279) );
  NAND U5838 ( .A(n4280), .B(n4279), .Z(n4392) );
  NAND U5839 ( .A(n4282), .B(n4281), .Z(n4286) );
  NAND U5840 ( .A(n4284), .B(n4283), .Z(n4285) );
  NAND U5841 ( .A(n4286), .B(n4285), .Z(n4405) );
  AND U5842 ( .A(\stack[1][10] ), .B(o[17]), .Z(n4419) );
  NAND U5843 ( .A(n4288), .B(n4287), .Z(n4292) );
  NAND U5844 ( .A(n4290), .B(n4289), .Z(n4291) );
  NAND U5845 ( .A(n4292), .B(n4291), .Z(n4417) );
  NAND U5846 ( .A(n4294), .B(n4293), .Z(n4298) );
  NAND U5847 ( .A(n4296), .B(n4295), .Z(n4297) );
  NAND U5848 ( .A(n4298), .B(n4297), .Z(n4423) );
  NAND U5849 ( .A(n4300), .B(n4299), .Z(n4304) );
  NAND U5850 ( .A(n4302), .B(n4301), .Z(n4303) );
  NAND U5851 ( .A(n4304), .B(n4303), .Z(n4429) );
  NAND U5852 ( .A(n4306), .B(n4305), .Z(n4310) );
  NAND U5853 ( .A(n4308), .B(n4307), .Z(n4309) );
  AND U5854 ( .A(n4310), .B(n4309), .Z(n4493) );
  NAND U5855 ( .A(n4312), .B(n4311), .Z(n4316) );
  NAND U5856 ( .A(n4314), .B(n4313), .Z(n4315) );
  AND U5857 ( .A(n4316), .B(n4315), .Z(n4480) );
  AND U5858 ( .A(o[7]), .B(\stack[1][20] ), .Z(n4437) );
  NAND U5859 ( .A(n4318), .B(n4317), .Z(n4322) );
  NAND U5860 ( .A(n4320), .B(n4319), .Z(n4321) );
  NAND U5861 ( .A(n4322), .B(n4321), .Z(n4435) );
  AND U5862 ( .A(o[6]), .B(\stack[1][21] ), .Z(n4471) );
  NAND U5863 ( .A(n4324), .B(n4323), .Z(n4328) );
  NAND U5864 ( .A(n4326), .B(n4325), .Z(n4327) );
  NAND U5865 ( .A(n4328), .B(n4327), .Z(n4441) );
  AND U5866 ( .A(o[4]), .B(\stack[1][23] ), .Z(n4440) );
  AND U5867 ( .A(o[1]), .B(\stack[1][26] ), .Z(n4446) );
  NAND U5868 ( .A(\stack[1][27] ), .B(o[0]), .Z(n4329) );
  XNOR U5869 ( .A(n4446), .B(n4329), .Z(n4449) );
  NAND U5870 ( .A(n4446), .B(o[0]), .Z(n4330) );
  XNOR U5871 ( .A(o[2]), .B(n4330), .Z(n4331) );
  AND U5872 ( .A(\stack[1][25] ), .B(n4331), .Z(n4450) );
  AND U5873 ( .A(o[0]), .B(\stack[1][24] ), .Z(n4333) );
  AND U5874 ( .A(n4333), .B(n4332), .Z(n4334) );
  NAND U5875 ( .A(o[2]), .B(n4334), .Z(n4338) );
  NAND U5876 ( .A(n4336), .B(n4335), .Z(n4337) );
  NAND U5877 ( .A(n4338), .B(n4337), .Z(n4457) );
  AND U5878 ( .A(o[3]), .B(\stack[1][24] ), .Z(n4459) );
  XOR U5879 ( .A(n4443), .B(n4442), .Z(n4462) );
  AND U5880 ( .A(o[5]), .B(\stack[1][22] ), .Z(n4463) );
  NAND U5881 ( .A(n4340), .B(n4339), .Z(n4344) );
  NAND U5882 ( .A(n4342), .B(n4341), .Z(n4343) );
  NAND U5883 ( .A(n4344), .B(n4343), .Z(n4465) );
  NAND U5884 ( .A(n4346), .B(n4345), .Z(n4350) );
  NAND U5885 ( .A(n4348), .B(n4347), .Z(n4349) );
  NAND U5886 ( .A(n4350), .B(n4349), .Z(n4469) );
  XOR U5887 ( .A(n4471), .B(n4470), .Z(n4434) );
  XOR U5888 ( .A(n4437), .B(n4436), .Z(n4477) );
  AND U5889 ( .A(o[8]), .B(\stack[1][19] ), .Z(n4474) );
  NAND U5890 ( .A(n4352), .B(n4351), .Z(n4356) );
  NAND U5891 ( .A(n4354), .B(n4353), .Z(n4355) );
  NAND U5892 ( .A(n4356), .B(n4355), .Z(n4475) );
  XNOR U5893 ( .A(n4477), .B(n4476), .Z(n4481) );
  NAND U5894 ( .A(o[9]), .B(\stack[1][18] ), .Z(n4482) );
  XNOR U5895 ( .A(n4483), .B(n4482), .Z(n4489) );
  AND U5896 ( .A(o[10]), .B(\stack[1][17] ), .Z(n4486) );
  NAND U5897 ( .A(n4358), .B(n4357), .Z(n4362) );
  NAND U5898 ( .A(n4360), .B(n4359), .Z(n4361) );
  NAND U5899 ( .A(n4362), .B(n4361), .Z(n4487) );
  XOR U5900 ( .A(n4493), .B(n4492), .Z(n4494) );
  AND U5901 ( .A(o[11]), .B(\stack[1][16] ), .Z(n4495) );
  AND U5902 ( .A(o[12]), .B(\stack[1][15] ), .Z(n4498) );
  NAND U5903 ( .A(n4364), .B(n4363), .Z(n4368) );
  NAND U5904 ( .A(n4366), .B(n4365), .Z(n4367) );
  AND U5905 ( .A(n4368), .B(n4367), .Z(n4499) );
  XNOR U5906 ( .A(n4501), .B(n4500), .Z(n4428) );
  NAND U5907 ( .A(\stack[1][14] ), .B(o[13]), .Z(n4430) );
  XNOR U5908 ( .A(n4431), .B(n4430), .Z(n4507) );
  AND U5909 ( .A(\stack[1][13] ), .B(o[14]), .Z(n4504) );
  NAND U5910 ( .A(n4370), .B(n4369), .Z(n4373) );
  NAND U5911 ( .A(n16829), .B(n4371), .Z(n4372) );
  NAND U5912 ( .A(n4373), .B(n4372), .Z(n4505) );
  AND U5913 ( .A(\stack[1][12] ), .B(o[15]), .Z(n4425) );
  AND U5914 ( .A(\stack[1][11] ), .B(o[16]), .Z(n4510) );
  NAND U5915 ( .A(n4375), .B(n4374), .Z(n4379) );
  NAND U5916 ( .A(n4377), .B(n4376), .Z(n4378) );
  NAND U5917 ( .A(n4379), .B(n4378), .Z(n4511) );
  XOR U5918 ( .A(n4513), .B(n4512), .Z(n4416) );
  XOR U5919 ( .A(n4419), .B(n4418), .Z(n4413) );
  AND U5920 ( .A(\stack[1][9] ), .B(o[18]), .Z(n4410) );
  NAND U5921 ( .A(n4381), .B(n4380), .Z(n4385) );
  NAND U5922 ( .A(n4383), .B(n4382), .Z(n4384) );
  NAND U5923 ( .A(n4385), .B(n4384), .Z(n4411) );
  XOR U5924 ( .A(n4413), .B(n4412), .Z(n4404) );
  AND U5925 ( .A(\stack[1][8] ), .B(o[19]), .Z(n4407) );
  AND U5926 ( .A(\stack[1][7] ), .B(o[20]), .Z(n4398) );
  NAND U5927 ( .A(n4387), .B(n4386), .Z(n4391) );
  NAND U5928 ( .A(n4389), .B(n4388), .Z(n4390) );
  NAND U5929 ( .A(n4391), .B(n4390), .Z(n4399) );
  XOR U5930 ( .A(n4401), .B(n4400), .Z(n4393) );
  NAND U5931 ( .A(n4392), .B(n4393), .Z(n4395) );
  AND U5932 ( .A(\stack[1][6] ), .B(o[21]), .Z(n12351) );
  NAND U5933 ( .A(n12351), .B(n12350), .Z(n4394) );
  AND U5934 ( .A(n4395), .B(n4394), .Z(n4397) );
  NAND U5935 ( .A(n4396), .B(n4397), .Z(n4517) );
  NAND U5936 ( .A(n4399), .B(n4398), .Z(n4403) );
  NAND U5937 ( .A(n4401), .B(n4400), .Z(n4402) );
  NAND U5938 ( .A(n4403), .B(n4402), .Z(n4637) );
  NAND U5939 ( .A(n4405), .B(n4404), .Z(n4409) );
  NAND U5940 ( .A(n4407), .B(n4406), .Z(n4408) );
  AND U5941 ( .A(n4409), .B(n4408), .Z(n4518) );
  NAND U5942 ( .A(\stack[1][8] ), .B(o[20]), .Z(n4519) );
  NAND U5943 ( .A(n4411), .B(n4410), .Z(n4415) );
  NAND U5944 ( .A(n4413), .B(n4412), .Z(n4414) );
  NAND U5945 ( .A(n4415), .B(n4414), .Z(n4631) );
  NAND U5946 ( .A(n4417), .B(n4416), .Z(n4421) );
  NAND U5947 ( .A(n4419), .B(n4418), .Z(n4420) );
  AND U5948 ( .A(n4421), .B(n4420), .Z(n4524) );
  NAND U5949 ( .A(\stack[1][10] ), .B(o[18]), .Z(n4525) );
  NAND U5950 ( .A(n4423), .B(n4422), .Z(n4427) );
  NAND U5951 ( .A(n4425), .B(n4424), .Z(n4426) );
  NAND U5952 ( .A(n4427), .B(n4426), .Z(n4531) );
  AND U5953 ( .A(\stack[1][12] ), .B(o[16]), .Z(n4530) );
  AND U5954 ( .A(\stack[1][14] ), .B(o[14]), .Z(n4536) );
  NAND U5955 ( .A(n4429), .B(n4428), .Z(n4433) );
  NAND U5956 ( .A(n4431), .B(n4430), .Z(n4432) );
  AND U5957 ( .A(n4433), .B(n4432), .Z(n4537) );
  NAND U5958 ( .A(n4435), .B(n4434), .Z(n4439) );
  NAND U5959 ( .A(n4437), .B(n4436), .Z(n4438) );
  NAND U5960 ( .A(n4439), .B(n4438), .Z(n4555) );
  AND U5961 ( .A(o[8]), .B(\stack[1][20] ), .Z(n4554) );
  AND U5962 ( .A(o[6]), .B(\stack[1][22] ), .Z(n4563) );
  NAND U5963 ( .A(n4441), .B(n4440), .Z(n4445) );
  NAND U5964 ( .A(n4443), .B(n4442), .Z(n4444) );
  NAND U5965 ( .A(n4445), .B(n4444), .Z(n4589) );
  AND U5966 ( .A(o[3]), .B(\stack[1][25] ), .Z(n4569) );
  AND U5967 ( .A(o[0]), .B(\stack[1][25] ), .Z(n4447) );
  AND U5968 ( .A(n4447), .B(n4446), .Z(n4448) );
  NAND U5969 ( .A(o[2]), .B(n4448), .Z(n4452) );
  NAND U5970 ( .A(n4450), .B(n4449), .Z(n4451) );
  NAND U5971 ( .A(n4452), .B(n4451), .Z(n4567) );
  AND U5972 ( .A(o[1]), .B(\stack[1][27] ), .Z(n4575) );
  NAND U5973 ( .A(\stack[1][28] ), .B(o[0]), .Z(n4453) );
  XNOR U5974 ( .A(n4575), .B(n4453), .Z(n4578) );
  NAND U5975 ( .A(n4575), .B(o[0]), .Z(n4454) );
  XNOR U5976 ( .A(o[2]), .B(n4454), .Z(n4455) );
  AND U5977 ( .A(\stack[1][26] ), .B(n4455), .Z(n4579) );
  XOR U5978 ( .A(n4569), .B(n4568), .Z(n4585) );
  AND U5979 ( .A(o[4]), .B(\stack[1][24] ), .Z(n4582) );
  NAND U5980 ( .A(n4457), .B(n4456), .Z(n4461) );
  NAND U5981 ( .A(n4459), .B(n4458), .Z(n4460) );
  NAND U5982 ( .A(n4461), .B(n4460), .Z(n4583) );
  XOR U5983 ( .A(n4585), .B(n4584), .Z(n4588) );
  AND U5984 ( .A(o[5]), .B(\stack[1][23] ), .Z(n4591) );
  NAND U5985 ( .A(n4463), .B(n4462), .Z(n4467) );
  NAND U5986 ( .A(n4465), .B(n4464), .Z(n4466) );
  NAND U5987 ( .A(n4467), .B(n4466), .Z(n4561) );
  XOR U5988 ( .A(n4563), .B(n4562), .Z(n4594) );
  NAND U5989 ( .A(n4469), .B(n4468), .Z(n4473) );
  NAND U5990 ( .A(n4471), .B(n4470), .Z(n4472) );
  NAND U5991 ( .A(n4473), .B(n4472), .Z(n4595) );
  AND U5992 ( .A(o[7]), .B(\stack[1][21] ), .Z(n4597) );
  XOR U5993 ( .A(n4557), .B(n4556), .Z(n4600) );
  NAND U5994 ( .A(n4475), .B(n4474), .Z(n4479) );
  NAND U5995 ( .A(n4477), .B(n4476), .Z(n4478) );
  NAND U5996 ( .A(n4479), .B(n4478), .Z(n4601) );
  AND U5997 ( .A(o[9]), .B(\stack[1][19] ), .Z(n4603) );
  NAND U5998 ( .A(n4481), .B(n4480), .Z(n4485) );
  NAND U5999 ( .A(n4483), .B(n4482), .Z(n4484) );
  AND U6000 ( .A(n4485), .B(n4484), .Z(n4548) );
  AND U6001 ( .A(o[10]), .B(\stack[1][18] ), .Z(n4549) );
  XNOR U6002 ( .A(n4551), .B(n4550), .Z(n4607) );
  NAND U6003 ( .A(n4487), .B(n4486), .Z(n4491) );
  NAND U6004 ( .A(n4489), .B(n4488), .Z(n4490) );
  AND U6005 ( .A(n4491), .B(n4490), .Z(n4606) );
  NAND U6006 ( .A(o[11]), .B(\stack[1][17] ), .Z(n4608) );
  XNOR U6007 ( .A(n4609), .B(n4608), .Z(n4545) );
  NAND U6008 ( .A(n4493), .B(n4492), .Z(n4497) );
  NAND U6009 ( .A(n4495), .B(n4494), .Z(n4496) );
  NAND U6010 ( .A(n4497), .B(n4496), .Z(n4543) );
  AND U6011 ( .A(o[12]), .B(\stack[1][16] ), .Z(n4542) );
  NAND U6012 ( .A(n4499), .B(n4498), .Z(n4503) );
  NAND U6013 ( .A(n4501), .B(n4500), .Z(n4502) );
  NAND U6014 ( .A(n4503), .B(n4502), .Z(n4613) );
  AND U6015 ( .A(\stack[1][15] ), .B(o[13]), .Z(n4615) );
  XOR U6016 ( .A(n4539), .B(n4538), .Z(n4618) );
  NAND U6017 ( .A(n4505), .B(n4504), .Z(n4509) );
  NAND U6018 ( .A(n4507), .B(n4506), .Z(n4508) );
  NAND U6019 ( .A(n4509), .B(n4508), .Z(n4619) );
  AND U6020 ( .A(\stack[1][13] ), .B(o[15]), .Z(n4621) );
  XOR U6021 ( .A(n4533), .B(n4532), .Z(n4624) );
  NAND U6022 ( .A(n4511), .B(n4510), .Z(n4515) );
  NAND U6023 ( .A(n4513), .B(n4512), .Z(n4514) );
  NAND U6024 ( .A(n4515), .B(n4514), .Z(n4625) );
  AND U6025 ( .A(\stack[1][11] ), .B(o[17]), .Z(n4626) );
  XNOR U6026 ( .A(n4627), .B(n4626), .Z(n4526) );
  XNOR U6027 ( .A(n4527), .B(n4526), .Z(n4630) );
  AND U6028 ( .A(\stack[1][9] ), .B(o[19]), .Z(n4632) );
  XNOR U6029 ( .A(n4633), .B(n4632), .Z(n4520) );
  XNOR U6030 ( .A(n4521), .B(n4520), .Z(n4636) );
  AND U6031 ( .A(\stack[1][7] ), .B(o[21]), .Z(n4638) );
  XNOR U6032 ( .A(n4639), .B(n4638), .Z(n12227) );
  NAND U6033 ( .A(n12228), .B(n12227), .Z(n4516) );
  AND U6034 ( .A(n4517), .B(n4516), .Z(n4643) );
  NAND U6035 ( .A(n4519), .B(n4518), .Z(n4523) );
  NAND U6036 ( .A(n4521), .B(n4520), .Z(n4522) );
  AND U6037 ( .A(n4523), .B(n4522), .Z(n4649) );
  NAND U6038 ( .A(n4525), .B(n4524), .Z(n4529) );
  NAND U6039 ( .A(n4527), .B(n4526), .Z(n4528) );
  AND U6040 ( .A(n4529), .B(n4528), .Z(n4655) );
  AND U6041 ( .A(\stack[1][12] ), .B(o[17]), .Z(n4757) );
  NAND U6042 ( .A(n4531), .B(n4530), .Z(n4535) );
  NAND U6043 ( .A(n4533), .B(n4532), .Z(n4534) );
  NAND U6044 ( .A(n4535), .B(n4534), .Z(n4755) );
  AND U6045 ( .A(\stack[1][14] ), .B(o[15]), .Z(n4745) );
  NAND U6046 ( .A(n4537), .B(n4536), .Z(n4541) );
  NAND U6047 ( .A(n4539), .B(n4538), .Z(n4540) );
  NAND U6048 ( .A(n4541), .B(n4540), .Z(n4743) );
  NAND U6049 ( .A(n4543), .B(n4542), .Z(n4547) );
  NAND U6050 ( .A(n4545), .B(n4544), .Z(n4546) );
  AND U6051 ( .A(n4547), .B(n4546), .Z(n4666) );
  AND U6052 ( .A(o[11]), .B(\stack[1][18] ), .Z(n4681) );
  NAND U6053 ( .A(n4549), .B(n4548), .Z(n4553) );
  NAND U6054 ( .A(n4551), .B(n4550), .Z(n4552) );
  NAND U6055 ( .A(n4553), .B(n4552), .Z(n4679) );
  NAND U6056 ( .A(n4555), .B(n4554), .Z(n4559) );
  NAND U6057 ( .A(n4557), .B(n4556), .Z(n4558) );
  AND U6058 ( .A(n4559), .B(n4558), .Z(n4690) );
  NAND U6059 ( .A(n4561), .B(n4560), .Z(n4565) );
  NAND U6060 ( .A(n4563), .B(n4562), .Z(n4564) );
  NAND U6061 ( .A(n4565), .B(n4564), .Z(n4731) );
  AND U6062 ( .A(o[6]), .B(\stack[1][23] ), .Z(n4727) );
  NAND U6063 ( .A(n4567), .B(n4566), .Z(n4571) );
  NAND U6064 ( .A(n4569), .B(n4568), .Z(n4570) );
  NAND U6065 ( .A(n4571), .B(n4570), .Z(n4697) );
  AND U6066 ( .A(o[4]), .B(\stack[1][25] ), .Z(n4696) );
  AND U6067 ( .A(o[1]), .B(\stack[1][28] ), .Z(n4702) );
  NAND U6068 ( .A(\stack[1][29] ), .B(o[0]), .Z(n4572) );
  XNOR U6069 ( .A(n4702), .B(n4572), .Z(n4705) );
  NAND U6070 ( .A(n4702), .B(o[0]), .Z(n4573) );
  XNOR U6071 ( .A(o[2]), .B(n4573), .Z(n4574) );
  AND U6072 ( .A(\stack[1][27] ), .B(n4574), .Z(n4706) );
  AND U6073 ( .A(o[0]), .B(\stack[1][26] ), .Z(n4576) );
  AND U6074 ( .A(n4576), .B(n4575), .Z(n4577) );
  NAND U6075 ( .A(o[2]), .B(n4577), .Z(n4581) );
  NAND U6076 ( .A(n4579), .B(n4578), .Z(n4580) );
  NAND U6077 ( .A(n4581), .B(n4580), .Z(n4713) );
  AND U6078 ( .A(o[3]), .B(\stack[1][26] ), .Z(n4715) );
  XOR U6079 ( .A(n4699), .B(n4698), .Z(n4718) );
  AND U6080 ( .A(o[5]), .B(\stack[1][24] ), .Z(n4719) );
  NAND U6081 ( .A(n4583), .B(n4582), .Z(n4587) );
  NAND U6082 ( .A(n4585), .B(n4584), .Z(n4586) );
  NAND U6083 ( .A(n4587), .B(n4586), .Z(n4721) );
  NAND U6084 ( .A(n4589), .B(n4588), .Z(n4593) );
  NAND U6085 ( .A(n4591), .B(n4590), .Z(n4592) );
  NAND U6086 ( .A(n4593), .B(n4592), .Z(n4725) );
  XOR U6087 ( .A(n4727), .B(n4726), .Z(n4730) );
  AND U6088 ( .A(o[7]), .B(\stack[1][22] ), .Z(n4733) );
  AND U6089 ( .A(o[8]), .B(\stack[1][21] ), .Z(n4736) );
  NAND U6090 ( .A(n4595), .B(n4594), .Z(n4599) );
  NAND U6091 ( .A(n4597), .B(n4596), .Z(n4598) );
  NAND U6092 ( .A(n4599), .B(n4598), .Z(n4737) );
  XNOR U6093 ( .A(n4739), .B(n4738), .Z(n4691) );
  NAND U6094 ( .A(o[9]), .B(\stack[1][20] ), .Z(n4692) );
  XNOR U6095 ( .A(n4693), .B(n4692), .Z(n4687) );
  AND U6096 ( .A(o[10]), .B(\stack[1][19] ), .Z(n4684) );
  NAND U6097 ( .A(n4601), .B(n4600), .Z(n4605) );
  NAND U6098 ( .A(n4603), .B(n4602), .Z(n4604) );
  NAND U6099 ( .A(n4605), .B(n4604), .Z(n4685) );
  XOR U6100 ( .A(n4681), .B(n4680), .Z(n4675) );
  AND U6101 ( .A(o[12]), .B(\stack[1][17] ), .Z(n4672) );
  NAND U6102 ( .A(n4607), .B(n4606), .Z(n4611) );
  NAND U6103 ( .A(n4609), .B(n4608), .Z(n4610) );
  AND U6104 ( .A(n4611), .B(n4610), .Z(n4673) );
  XNOR U6105 ( .A(n4675), .B(n4674), .Z(n4667) );
  NAND U6106 ( .A(o[13]), .B(\stack[1][16] ), .Z(n4668) );
  XNOR U6107 ( .A(n4669), .B(n4668), .Z(n4663) );
  AND U6108 ( .A(\stack[1][15] ), .B(o[14]), .Z(n4660) );
  NAND U6109 ( .A(n4613), .B(n4612), .Z(n4617) );
  NAND U6110 ( .A(n4615), .B(n4614), .Z(n4616) );
  NAND U6111 ( .A(n4617), .B(n4616), .Z(n4661) );
  XOR U6112 ( .A(n4745), .B(n4744), .Z(n4751) );
  AND U6113 ( .A(\stack[1][13] ), .B(o[16]), .Z(n4748) );
  NAND U6114 ( .A(n4619), .B(n4618), .Z(n4623) );
  NAND U6115 ( .A(n4621), .B(n4620), .Z(n4622) );
  NAND U6116 ( .A(n4623), .B(n4622), .Z(n4749) );
  XOR U6117 ( .A(n4751), .B(n4750), .Z(n4754) );
  XOR U6118 ( .A(n4757), .B(n4756), .Z(n4763) );
  AND U6119 ( .A(\stack[1][11] ), .B(o[18]), .Z(n4760) );
  NAND U6120 ( .A(n4625), .B(n4624), .Z(n4629) );
  NAND U6121 ( .A(n4627), .B(n4626), .Z(n4628) );
  NAND U6122 ( .A(n4629), .B(n4628), .Z(n4761) );
  XOR U6123 ( .A(n4763), .B(n4762), .Z(n4654) );
  XOR U6124 ( .A(n4655), .B(n4654), .Z(n4656) );
  AND U6125 ( .A(\stack[1][10] ), .B(o[19]), .Z(n4657) );
  AND U6126 ( .A(\stack[1][9] ), .B(o[20]), .Z(n4766) );
  NAND U6127 ( .A(n4631), .B(n4630), .Z(n4635) );
  NAND U6128 ( .A(n4633), .B(n4632), .Z(n4634) );
  NAND U6129 ( .A(n4635), .B(n4634), .Z(n4767) );
  XOR U6130 ( .A(n4769), .B(n4768), .Z(n4648) );
  XOR U6131 ( .A(n4649), .B(n4648), .Z(n4650) );
  AND U6132 ( .A(\stack[1][8] ), .B(o[21]), .Z(n4651) );
  AND U6133 ( .A(\stack[1][7] ), .B(o[22]), .Z(n4772) );
  NAND U6134 ( .A(n4637), .B(n4636), .Z(n4641) );
  NAND U6135 ( .A(n4639), .B(n4638), .Z(n4640) );
  NAND U6136 ( .A(n4641), .B(n4640), .Z(n4773) );
  XOR U6137 ( .A(n4775), .B(n4774), .Z(n4642) );
  NAND U6138 ( .A(n4643), .B(n4642), .Z(n4645) );
  AND U6139 ( .A(\stack[1][6] ), .B(o[23]), .Z(n12360) );
  XOR U6140 ( .A(n4643), .B(n4642), .Z(n12361) );
  NAND U6141 ( .A(n12360), .B(n12361), .Z(n4644) );
  NAND U6142 ( .A(n4645), .B(n4644), .Z(n4646) );
  AND U6143 ( .A(\stack[1][6] ), .B(o[24]), .Z(n4647) );
  NAND U6144 ( .A(n4646), .B(n4647), .Z(n4779) );
  NAND U6145 ( .A(n4649), .B(n4648), .Z(n4653) );
  NAND U6146 ( .A(n4651), .B(n4650), .Z(n4652) );
  NAND U6147 ( .A(n4653), .B(n4652), .Z(n4781) );
  AND U6148 ( .A(\stack[1][8] ), .B(o[22]), .Z(n4780) );
  NAND U6149 ( .A(n4655), .B(n4654), .Z(n4659) );
  NAND U6150 ( .A(n4657), .B(n4656), .Z(n4658) );
  NAND U6151 ( .A(n4659), .B(n4658), .Z(n4787) );
  AND U6152 ( .A(\stack[1][10] ), .B(o[20]), .Z(n4786) );
  NAND U6153 ( .A(n4661), .B(n4660), .Z(n4665) );
  NAND U6154 ( .A(n4663), .B(n4662), .Z(n4664) );
  NAND U6155 ( .A(n4665), .B(n4664), .Z(n4887) );
  NAND U6156 ( .A(n4667), .B(n4666), .Z(n4671) );
  NAND U6157 ( .A(n4669), .B(n4668), .Z(n4670) );
  NAND U6158 ( .A(n4671), .B(n4670), .Z(n4805) );
  NAND U6159 ( .A(o[14]), .B(\stack[1][16] ), .Z(n4804) );
  NAND U6160 ( .A(n4673), .B(n4672), .Z(n4677) );
  NAND U6161 ( .A(n4675), .B(n4674), .Z(n4676) );
  NAND U6162 ( .A(n4677), .B(n4676), .Z(n4881) );
  NAND U6163 ( .A(n4679), .B(n4678), .Z(n4683) );
  NAND U6164 ( .A(n4681), .B(n4680), .Z(n4682) );
  AND U6165 ( .A(n4683), .B(n4682), .Z(n4810) );
  NAND U6166 ( .A(o[12]), .B(\stack[1][18] ), .Z(n4811) );
  NAND U6167 ( .A(n4685), .B(n4684), .Z(n4689) );
  NAND U6168 ( .A(n4687), .B(n4686), .Z(n4688) );
  AND U6169 ( .A(n4689), .B(n4688), .Z(n4875) );
  NAND U6170 ( .A(n4691), .B(n4690), .Z(n4695) );
  NAND U6171 ( .A(n4693), .B(n4692), .Z(n4694) );
  NAND U6172 ( .A(n4695), .B(n4694), .Z(n4817) );
  NAND U6173 ( .A(o[10]), .B(\stack[1][20] ), .Z(n4816) );
  AND U6174 ( .A(o[5]), .B(\stack[1][25] ), .Z(n4859) );
  NAND U6175 ( .A(n4697), .B(n4696), .Z(n4701) );
  NAND U6176 ( .A(n4699), .B(n4698), .Z(n4700) );
  NAND U6177 ( .A(n4701), .B(n4700), .Z(n4857) );
  AND U6178 ( .A(o[0]), .B(\stack[1][27] ), .Z(n4703) );
  AND U6179 ( .A(n4703), .B(n4702), .Z(n4704) );
  NAND U6180 ( .A(o[2]), .B(n4704), .Z(n4708) );
  NAND U6181 ( .A(n4706), .B(n4705), .Z(n4707) );
  NAND U6182 ( .A(n4708), .B(n4707), .Z(n4835) );
  AND U6183 ( .A(o[1]), .B(\stack[1][29] ), .Z(n4843) );
  NAND U6184 ( .A(\stack[1][30] ), .B(o[0]), .Z(n4709) );
  XNOR U6185 ( .A(n4843), .B(n4709), .Z(n4846) );
  NAND U6186 ( .A(n4843), .B(o[0]), .Z(n4710) );
  XNOR U6187 ( .A(o[2]), .B(n4710), .Z(n4711) );
  AND U6188 ( .A(\stack[1][28] ), .B(n4711), .Z(n4847) );
  AND U6189 ( .A(o[3]), .B(\stack[1][27] ), .Z(n4837) );
  AND U6190 ( .A(o[4]), .B(\stack[1][26] ), .Z(n4850) );
  NAND U6191 ( .A(n4713), .B(n4712), .Z(n4717) );
  NAND U6192 ( .A(n4715), .B(n4714), .Z(n4716) );
  NAND U6193 ( .A(n4717), .B(n4716), .Z(n4851) );
  XOR U6194 ( .A(n4853), .B(n4852), .Z(n4856) );
  XOR U6195 ( .A(n4859), .B(n4858), .Z(n4828) );
  NAND U6196 ( .A(n4719), .B(n4718), .Z(n4723) );
  NAND U6197 ( .A(n4721), .B(n4720), .Z(n4722) );
  NAND U6198 ( .A(n4723), .B(n4722), .Z(n4829) );
  AND U6199 ( .A(o[6]), .B(\stack[1][24] ), .Z(n4831) );
  NAND U6200 ( .A(n4725), .B(n4724), .Z(n4729) );
  NAND U6201 ( .A(n4727), .B(n4726), .Z(n4728) );
  NAND U6202 ( .A(n4729), .B(n4728), .Z(n4863) );
  AND U6203 ( .A(o[7]), .B(\stack[1][23] ), .Z(n4865) );
  NAND U6204 ( .A(n4731), .B(n4730), .Z(n4735) );
  NAND U6205 ( .A(n4733), .B(n4732), .Z(n4734) );
  NAND U6206 ( .A(n4735), .B(n4734), .Z(n4823) );
  AND U6207 ( .A(o[8]), .B(\stack[1][22] ), .Z(n4822) );
  XOR U6208 ( .A(n4825), .B(n4824), .Z(n4868) );
  NAND U6209 ( .A(n4737), .B(n4736), .Z(n4741) );
  NAND U6210 ( .A(n4739), .B(n4738), .Z(n4740) );
  NAND U6211 ( .A(n4741), .B(n4740), .Z(n4869) );
  AND U6212 ( .A(o[9]), .B(\stack[1][21] ), .Z(n4870) );
  XNOR U6213 ( .A(n4871), .B(n4870), .Z(n4819) );
  XOR U6214 ( .A(n4875), .B(n4874), .Z(n4876) );
  NAND U6215 ( .A(o[11]), .B(\stack[1][19] ), .Z(n4877) );
  XNOR U6216 ( .A(n4813), .B(n4812), .Z(n4880) );
  AND U6217 ( .A(o[13]), .B(\stack[1][17] ), .Z(n4882) );
  XNOR U6218 ( .A(n4883), .B(n4882), .Z(n4806) );
  XNOR U6219 ( .A(n4807), .B(n4806), .Z(n4886) );
  AND U6220 ( .A(\stack[1][15] ), .B(o[15]), .Z(n4888) );
  XNOR U6221 ( .A(n4889), .B(n4888), .Z(n4801) );
  NAND U6222 ( .A(n4743), .B(n4742), .Z(n4747) );
  NAND U6223 ( .A(n4745), .B(n4744), .Z(n4746) );
  AND U6224 ( .A(n4747), .B(n4746), .Z(n4798) );
  NAND U6225 ( .A(\stack[1][14] ), .B(o[16]), .Z(n4799) );
  NAND U6226 ( .A(n4749), .B(n4748), .Z(n4753) );
  NAND U6227 ( .A(n4751), .B(n4750), .Z(n4752) );
  NAND U6228 ( .A(n4753), .B(n4752), .Z(n4892) );
  XOR U6229 ( .A(n4893), .B(n4892), .Z(n4895) );
  AND U6230 ( .A(\stack[1][13] ), .B(o[17]), .Z(n4894) );
  XNOR U6231 ( .A(n4895), .B(n4894), .Z(n4795) );
  NAND U6232 ( .A(n4755), .B(n4754), .Z(n4759) );
  NAND U6233 ( .A(n4757), .B(n4756), .Z(n4758) );
  AND U6234 ( .A(n4759), .B(n4758), .Z(n4792) );
  NAND U6235 ( .A(\stack[1][12] ), .B(o[18]), .Z(n4793) );
  NAND U6236 ( .A(n4761), .B(n4760), .Z(n4765) );
  NAND U6237 ( .A(n4763), .B(n4762), .Z(n4764) );
  NAND U6238 ( .A(n4765), .B(n4764), .Z(n4898) );
  XOR U6239 ( .A(n4899), .B(n4898), .Z(n4900) );
  AND U6240 ( .A(\stack[1][11] ), .B(o[19]), .Z(n4901) );
  XOR U6241 ( .A(n4789), .B(n4788), .Z(n4904) );
  NAND U6242 ( .A(n4767), .B(n4766), .Z(n4771) );
  NAND U6243 ( .A(n4769), .B(n4768), .Z(n4770) );
  NAND U6244 ( .A(n4771), .B(n4770), .Z(n4905) );
  AND U6245 ( .A(\stack[1][9] ), .B(o[21]), .Z(n4907) );
  XOR U6246 ( .A(n4783), .B(n4782), .Z(n4910) );
  NAND U6247 ( .A(n4773), .B(n4772), .Z(n4777) );
  NAND U6248 ( .A(n4775), .B(n4774), .Z(n4776) );
  NAND U6249 ( .A(n4777), .B(n4776), .Z(n4911) );
  AND U6250 ( .A(\stack[1][7] ), .B(o[23]), .Z(n4913) );
  NAND U6251 ( .A(n12367), .B(n12366), .Z(n4778) );
  NAND U6252 ( .A(n4779), .B(n4778), .Z(n4916) );
  NAND U6253 ( .A(n4781), .B(n4780), .Z(n4785) );
  NAND U6254 ( .A(n4783), .B(n4782), .Z(n4784) );
  NAND U6255 ( .A(n4785), .B(n4784), .Z(n4921) );
  NAND U6256 ( .A(n4787), .B(n4786), .Z(n4791) );
  NAND U6257 ( .A(n4789), .B(n4788), .Z(n4790) );
  NAND U6258 ( .A(n4791), .B(n4790), .Z(n4927) );
  NAND U6259 ( .A(n4793), .B(n4792), .Z(n4797) );
  NAND U6260 ( .A(n4795), .B(n4794), .Z(n4796) );
  AND U6261 ( .A(n4797), .B(n4796), .Z(n4933) );
  AND U6262 ( .A(\stack[1][14] ), .B(o[17]), .Z(n4947) );
  NAND U6263 ( .A(n4799), .B(n4798), .Z(n4803) );
  NAND U6264 ( .A(n4801), .B(n4800), .Z(n4802) );
  AND U6265 ( .A(n4803), .B(n4802), .Z(n4945) );
  AND U6266 ( .A(\stack[1][16] ), .B(o[15]), .Z(n5035) );
  NAND U6267 ( .A(n4805), .B(n4804), .Z(n4809) );
  NAND U6268 ( .A(n4807), .B(n4806), .Z(n4808) );
  AND U6269 ( .A(n4809), .B(n4808), .Z(n5033) );
  NAND U6270 ( .A(n4811), .B(n4810), .Z(n4815) );
  NAND U6271 ( .A(n4813), .B(n4812), .Z(n4814) );
  NAND U6272 ( .A(n4815), .B(n4814), .Z(n4951) );
  AND U6273 ( .A(o[11]), .B(\stack[1][20] ), .Z(n4959) );
  NAND U6274 ( .A(n4817), .B(n4816), .Z(n4821) );
  NAND U6275 ( .A(n4819), .B(n4818), .Z(n4820) );
  AND U6276 ( .A(n4821), .B(n4820), .Z(n4957) );
  NAND U6277 ( .A(n4823), .B(n4822), .Z(n4827) );
  NAND U6278 ( .A(n4825), .B(n4824), .Z(n4826) );
  AND U6279 ( .A(n4827), .B(n4826), .Z(n5008) );
  NAND U6280 ( .A(n4829), .B(n4828), .Z(n4833) );
  NAND U6281 ( .A(n4831), .B(n4830), .Z(n4832) );
  NAND U6282 ( .A(n4833), .B(n4832), .Z(n4963) );
  AND U6283 ( .A(o[6]), .B(\stack[1][25] ), .Z(n4999) );
  NAND U6284 ( .A(n4835), .B(n4834), .Z(n4839) );
  NAND U6285 ( .A(n4837), .B(n4836), .Z(n4838) );
  NAND U6286 ( .A(n4839), .B(n4838), .Z(n4969) );
  AND U6287 ( .A(o[4]), .B(\stack[1][27] ), .Z(n4968) );
  AND U6288 ( .A(o[1]), .B(\stack[1][30] ), .Z(n4974) );
  NAND U6289 ( .A(\stack[1][31] ), .B(o[0]), .Z(n4840) );
  XNOR U6290 ( .A(n4974), .B(n4840), .Z(n4977) );
  NAND U6291 ( .A(n4974), .B(o[0]), .Z(n4841) );
  XNOR U6292 ( .A(o[2]), .B(n4841), .Z(n4842) );
  AND U6293 ( .A(\stack[1][29] ), .B(n4842), .Z(n4978) );
  AND U6294 ( .A(o[0]), .B(\stack[1][28] ), .Z(n4844) );
  AND U6295 ( .A(n4844), .B(n4843), .Z(n4845) );
  NAND U6296 ( .A(o[2]), .B(n4845), .Z(n4849) );
  NAND U6297 ( .A(n4847), .B(n4846), .Z(n4848) );
  NAND U6298 ( .A(n4849), .B(n4848), .Z(n4985) );
  AND U6299 ( .A(o[3]), .B(\stack[1][28] ), .Z(n4987) );
  XOR U6300 ( .A(n4971), .B(n4970), .Z(n4990) );
  AND U6301 ( .A(o[5]), .B(\stack[1][26] ), .Z(n4991) );
  NAND U6302 ( .A(n4851), .B(n4850), .Z(n4855) );
  NAND U6303 ( .A(n4853), .B(n4852), .Z(n4854) );
  NAND U6304 ( .A(n4855), .B(n4854), .Z(n4993) );
  NAND U6305 ( .A(n4857), .B(n4856), .Z(n4861) );
  NAND U6306 ( .A(n4859), .B(n4858), .Z(n4860) );
  NAND U6307 ( .A(n4861), .B(n4860), .Z(n4997) );
  XOR U6308 ( .A(n4999), .B(n4998), .Z(n4962) );
  AND U6309 ( .A(o[7]), .B(\stack[1][24] ), .Z(n4965) );
  AND U6310 ( .A(o[8]), .B(\stack[1][23] ), .Z(n5002) );
  NAND U6311 ( .A(n4863), .B(n4862), .Z(n4867) );
  NAND U6312 ( .A(n4865), .B(n4864), .Z(n4866) );
  NAND U6313 ( .A(n4867), .B(n4866), .Z(n5003) );
  XNOR U6314 ( .A(n5005), .B(n5004), .Z(n5009) );
  NAND U6315 ( .A(o[9]), .B(\stack[1][22] ), .Z(n5010) );
  XNOR U6316 ( .A(n5011), .B(n5010), .Z(n5017) );
  AND U6317 ( .A(o[10]), .B(\stack[1][21] ), .Z(n5014) );
  NAND U6318 ( .A(n4869), .B(n4868), .Z(n4873) );
  NAND U6319 ( .A(n4871), .B(n4870), .Z(n4872) );
  NAND U6320 ( .A(n4873), .B(n4872), .Z(n5015) );
  XOR U6321 ( .A(n4957), .B(n4956), .Z(n4958) );
  XOR U6322 ( .A(n4959), .B(n4958), .Z(n5023) );
  AND U6323 ( .A(o[12]), .B(\stack[1][19] ), .Z(n5020) );
  NAND U6324 ( .A(n4875), .B(n4874), .Z(n4879) );
  NAND U6325 ( .A(n4877), .B(n4876), .Z(n4878) );
  AND U6326 ( .A(n4879), .B(n4878), .Z(n5021) );
  XNOR U6327 ( .A(n5023), .B(n5022), .Z(n4950) );
  NAND U6328 ( .A(o[13]), .B(\stack[1][18] ), .Z(n4952) );
  XNOR U6329 ( .A(n4953), .B(n4952), .Z(n5029) );
  AND U6330 ( .A(o[14]), .B(\stack[1][17] ), .Z(n5026) );
  NAND U6331 ( .A(n4881), .B(n4880), .Z(n4885) );
  NAND U6332 ( .A(n4883), .B(n4882), .Z(n4884) );
  NAND U6333 ( .A(n4885), .B(n4884), .Z(n5027) );
  XOR U6334 ( .A(n5033), .B(n5032), .Z(n5034) );
  XOR U6335 ( .A(n5035), .B(n5034), .Z(n5041) );
  AND U6336 ( .A(\stack[1][15] ), .B(o[16]), .Z(n5038) );
  NAND U6337 ( .A(n4887), .B(n4886), .Z(n4891) );
  NAND U6338 ( .A(n4889), .B(n4888), .Z(n4890) );
  NAND U6339 ( .A(n4891), .B(n4890), .Z(n5039) );
  XOR U6340 ( .A(n5041), .B(n5040), .Z(n4944) );
  XOR U6341 ( .A(n4945), .B(n4944), .Z(n4946) );
  XOR U6342 ( .A(n4947), .B(n4946), .Z(n4941) );
  AND U6343 ( .A(\stack[1][13] ), .B(o[18]), .Z(n4938) );
  NAND U6344 ( .A(n4893), .B(n4892), .Z(n4897) );
  NAND U6345 ( .A(n4895), .B(n4894), .Z(n4896) );
  NAND U6346 ( .A(n4897), .B(n4896), .Z(n4939) );
  XOR U6347 ( .A(n4941), .B(n4940), .Z(n4932) );
  XOR U6348 ( .A(n4933), .B(n4932), .Z(n4934) );
  AND U6349 ( .A(\stack[1][12] ), .B(o[19]), .Z(n4935) );
  AND U6350 ( .A(\stack[1][11] ), .B(o[20]), .Z(n5044) );
  NAND U6351 ( .A(n4899), .B(n4898), .Z(n4903) );
  NAND U6352 ( .A(n4901), .B(n4900), .Z(n4902) );
  NAND U6353 ( .A(n4903), .B(n4902), .Z(n5045) );
  XOR U6354 ( .A(n5047), .B(n5046), .Z(n4926) );
  AND U6355 ( .A(\stack[1][10] ), .B(o[21]), .Z(n4929) );
  AND U6356 ( .A(\stack[1][9] ), .B(o[22]), .Z(n5050) );
  NAND U6357 ( .A(n4905), .B(n4904), .Z(n4909) );
  NAND U6358 ( .A(n4907), .B(n4906), .Z(n4908) );
  NAND U6359 ( .A(n4909), .B(n4908), .Z(n5051) );
  XOR U6360 ( .A(n5053), .B(n5052), .Z(n4920) );
  AND U6361 ( .A(\stack[1][8] ), .B(o[23]), .Z(n4923) );
  AND U6362 ( .A(\stack[1][7] ), .B(o[24]), .Z(n5056) );
  NAND U6363 ( .A(n4911), .B(n4910), .Z(n4915) );
  NAND U6364 ( .A(n4913), .B(n4912), .Z(n4914) );
  NAND U6365 ( .A(n4915), .B(n4914), .Z(n5057) );
  XOR U6366 ( .A(n5059), .B(n5058), .Z(n4917) );
  NAND U6367 ( .A(n4916), .B(n4917), .Z(n4919) );
  AND U6368 ( .A(\stack[1][6] ), .B(o[25]), .Z(n12372) );
  NAND U6369 ( .A(n12372), .B(n12373), .Z(n4918) );
  NAND U6370 ( .A(n4919), .B(n4918), .Z(n5062) );
  AND U6371 ( .A(\stack[1][6] ), .B(o[26]), .Z(n5063) );
  NAND U6372 ( .A(n5062), .B(n5063), .Z(n5065) );
  NAND U6373 ( .A(n4921), .B(n4920), .Z(n4925) );
  NAND U6374 ( .A(n4923), .B(n4922), .Z(n4924) );
  NAND U6375 ( .A(n4925), .B(n4924), .Z(n5067) );
  AND U6376 ( .A(\stack[1][8] ), .B(o[24]), .Z(n5066) );
  NAND U6377 ( .A(n4927), .B(n4926), .Z(n4931) );
  NAND U6378 ( .A(n4929), .B(n4928), .Z(n4930) );
  NAND U6379 ( .A(n4931), .B(n4930), .Z(n5073) );
  AND U6380 ( .A(\stack[1][10] ), .B(o[22]), .Z(n5072) );
  NAND U6381 ( .A(n4933), .B(n4932), .Z(n4937) );
  NAND U6382 ( .A(n4935), .B(n4934), .Z(n4936) );
  NAND U6383 ( .A(n4937), .B(n4936), .Z(n5079) );
  AND U6384 ( .A(\stack[1][12] ), .B(o[20]), .Z(n5078) );
  NAND U6385 ( .A(n4939), .B(n4938), .Z(n4943) );
  NAND U6386 ( .A(n4941), .B(n4940), .Z(n4942) );
  NAND U6387 ( .A(n4943), .B(n4942), .Z(n5190) );
  NAND U6388 ( .A(n4945), .B(n4944), .Z(n4949) );
  NAND U6389 ( .A(n4947), .B(n4946), .Z(n4948) );
  AND U6390 ( .A(n4949), .B(n4948), .Z(n5084) );
  NAND U6391 ( .A(\stack[1][14] ), .B(o[18]), .Z(n5085) );
  NAND U6392 ( .A(n4951), .B(n4950), .Z(n4955) );
  NAND U6393 ( .A(n4953), .B(n4952), .Z(n4954) );
  AND U6394 ( .A(n4955), .B(n4954), .Z(n5095) );
  AND U6395 ( .A(o[14]), .B(\stack[1][18] ), .Z(n5096) );
  NAND U6396 ( .A(n4957), .B(n4956), .Z(n4961) );
  NAND U6397 ( .A(n4959), .B(n4958), .Z(n4960) );
  NAND U6398 ( .A(n4961), .B(n4960), .Z(n5102) );
  AND U6399 ( .A(o[12]), .B(\stack[1][20] ), .Z(n5101) );
  AND U6400 ( .A(o[11]), .B(\stack[1][21] ), .Z(n5168) );
  NAND U6401 ( .A(n4963), .B(n4962), .Z(n4967) );
  NAND U6402 ( .A(n4965), .B(n4964), .Z(n4966) );
  NAND U6403 ( .A(n4967), .B(n4966), .Z(n5114) );
  AND U6404 ( .A(o[8]), .B(\stack[1][24] ), .Z(n5113) );
  AND U6405 ( .A(o[6]), .B(\stack[1][26] ), .Z(n5122) );
  NAND U6406 ( .A(n4969), .B(n4968), .Z(n4973) );
  NAND U6407 ( .A(n4971), .B(n4970), .Z(n4972) );
  NAND U6408 ( .A(n4973), .B(n4972), .Z(n5148) );
  AND U6409 ( .A(o[0]), .B(\stack[1][29] ), .Z(n4975) );
  AND U6410 ( .A(n4975), .B(n4974), .Z(n4976) );
  NAND U6411 ( .A(o[2]), .B(n4976), .Z(n4980) );
  NAND U6412 ( .A(n4978), .B(n4977), .Z(n4979) );
  NAND U6413 ( .A(n4980), .B(n4979), .Z(n5126) );
  AND U6414 ( .A(o[1]), .B(\stack[1][31] ), .Z(n5134) );
  NAND U6415 ( .A(\stack[1][32] ), .B(o[0]), .Z(n4981) );
  XNOR U6416 ( .A(n5134), .B(n4981), .Z(n5138) );
  NAND U6417 ( .A(n5134), .B(o[0]), .Z(n4982) );
  XNOR U6418 ( .A(o[2]), .B(n4982), .Z(n4983) );
  AND U6419 ( .A(\stack[1][30] ), .B(n4983), .Z(n5137) );
  XOR U6420 ( .A(n5138), .B(n5137), .Z(n5125) );
  AND U6421 ( .A(o[3]), .B(\stack[1][29] ), .Z(n5128) );
  AND U6422 ( .A(o[4]), .B(\stack[1][28] ), .Z(n5141) );
  NAND U6423 ( .A(n4985), .B(n4984), .Z(n4989) );
  NAND U6424 ( .A(n4987), .B(n4986), .Z(n4988) );
  NAND U6425 ( .A(n4989), .B(n4988), .Z(n5142) );
  XOR U6426 ( .A(n5144), .B(n5143), .Z(n5147) );
  AND U6427 ( .A(o[5]), .B(\stack[1][27] ), .Z(n5150) );
  NAND U6428 ( .A(n4991), .B(n4990), .Z(n4995) );
  NAND U6429 ( .A(n4993), .B(n4992), .Z(n4994) );
  NAND U6430 ( .A(n4995), .B(n4994), .Z(n5120) );
  XOR U6431 ( .A(n5122), .B(n5121), .Z(n5153) );
  NAND U6432 ( .A(n4997), .B(n4996), .Z(n5001) );
  NAND U6433 ( .A(n4999), .B(n4998), .Z(n5000) );
  NAND U6434 ( .A(n5001), .B(n5000), .Z(n5154) );
  AND U6435 ( .A(o[7]), .B(\stack[1][25] ), .Z(n5156) );
  XOR U6436 ( .A(n5116), .B(n5115), .Z(n5159) );
  NAND U6437 ( .A(n5003), .B(n5002), .Z(n5007) );
  NAND U6438 ( .A(n5005), .B(n5004), .Z(n5006) );
  NAND U6439 ( .A(n5007), .B(n5006), .Z(n5160) );
  AND U6440 ( .A(o[9]), .B(\stack[1][23] ), .Z(n5162) );
  NAND U6441 ( .A(n5009), .B(n5008), .Z(n5013) );
  NAND U6442 ( .A(n5011), .B(n5010), .Z(n5012) );
  AND U6443 ( .A(n5013), .B(n5012), .Z(n5107) );
  AND U6444 ( .A(o[10]), .B(\stack[1][22] ), .Z(n5108) );
  XOR U6445 ( .A(n5110), .B(n5109), .Z(n5165) );
  NAND U6446 ( .A(n5015), .B(n5014), .Z(n5019) );
  NAND U6447 ( .A(n5017), .B(n5016), .Z(n5018) );
  NAND U6448 ( .A(n5019), .B(n5018), .Z(n5166) );
  XOR U6449 ( .A(n5168), .B(n5167), .Z(n5103) );
  XOR U6450 ( .A(n5104), .B(n5103), .Z(n5171) );
  NAND U6451 ( .A(n5021), .B(n5020), .Z(n5025) );
  NAND U6452 ( .A(n5023), .B(n5022), .Z(n5024) );
  NAND U6453 ( .A(n5025), .B(n5024), .Z(n5172) );
  AND U6454 ( .A(o[13]), .B(\stack[1][19] ), .Z(n5174) );
  XOR U6455 ( .A(n5098), .B(n5097), .Z(n5177) );
  NAND U6456 ( .A(n5027), .B(n5026), .Z(n5031) );
  NAND U6457 ( .A(n5029), .B(n5028), .Z(n5030) );
  NAND U6458 ( .A(n5031), .B(n5030), .Z(n5178) );
  AND U6459 ( .A(\stack[1][17] ), .B(o[15]), .Z(n5180) );
  AND U6460 ( .A(\stack[1][16] ), .B(o[16]), .Z(n16714) );
  NAND U6461 ( .A(n5033), .B(n5032), .Z(n5037) );
  NAND U6462 ( .A(n5035), .B(n5034), .Z(n5036) );
  NAND U6463 ( .A(n5037), .B(n5036), .Z(n5090) );
  XOR U6464 ( .A(n5092), .B(n5091), .Z(n5183) );
  NAND U6465 ( .A(n5039), .B(n5038), .Z(n5043) );
  NAND U6466 ( .A(n5041), .B(n5040), .Z(n5042) );
  NAND U6467 ( .A(n5043), .B(n5042), .Z(n5184) );
  AND U6468 ( .A(\stack[1][15] ), .B(o[17]), .Z(n5185) );
  XNOR U6469 ( .A(n5186), .B(n5185), .Z(n5086) );
  XNOR U6470 ( .A(n5087), .B(n5086), .Z(n5189) );
  AND U6471 ( .A(\stack[1][13] ), .B(o[19]), .Z(n5192) );
  XOR U6472 ( .A(n5081), .B(n5080), .Z(n5195) );
  NAND U6473 ( .A(n5045), .B(n5044), .Z(n5049) );
  NAND U6474 ( .A(n5047), .B(n5046), .Z(n5048) );
  NAND U6475 ( .A(n5049), .B(n5048), .Z(n5196) );
  AND U6476 ( .A(\stack[1][11] ), .B(o[21]), .Z(n5198) );
  XOR U6477 ( .A(n5075), .B(n5074), .Z(n5201) );
  NAND U6478 ( .A(n5051), .B(n5050), .Z(n5055) );
  NAND U6479 ( .A(n5053), .B(n5052), .Z(n5054) );
  NAND U6480 ( .A(n5055), .B(n5054), .Z(n5202) );
  AND U6481 ( .A(\stack[1][9] ), .B(o[23]), .Z(n5204) );
  XOR U6482 ( .A(n5069), .B(n5068), .Z(n5207) );
  NAND U6483 ( .A(n5057), .B(n5056), .Z(n5061) );
  NAND U6484 ( .A(n5059), .B(n5058), .Z(n5060) );
  NAND U6485 ( .A(n5061), .B(n5060), .Z(n5208) );
  AND U6486 ( .A(\stack[1][7] ), .B(o[25]), .Z(n5210) );
  NAND U6487 ( .A(n12379), .B(n12378), .Z(n5064) );
  NAND U6488 ( .A(n5065), .B(n5064), .Z(n5213) );
  NAND U6489 ( .A(n5067), .B(n5066), .Z(n5071) );
  NAND U6490 ( .A(n5069), .B(n5068), .Z(n5070) );
  NAND U6491 ( .A(n5071), .B(n5070), .Z(n5220) );
  AND U6492 ( .A(\stack[1][10] ), .B(o[23]), .Z(n5228) );
  NAND U6493 ( .A(n5073), .B(n5072), .Z(n5077) );
  NAND U6494 ( .A(n5075), .B(n5074), .Z(n5076) );
  NAND U6495 ( .A(n5077), .B(n5076), .Z(n5226) );
  AND U6496 ( .A(\stack[1][12] ), .B(o[21]), .Z(n5234) );
  NAND U6497 ( .A(n5079), .B(n5078), .Z(n5083) );
  NAND U6498 ( .A(n5081), .B(n5080), .Z(n5082) );
  NAND U6499 ( .A(n5083), .B(n5082), .Z(n5232) );
  AND U6500 ( .A(\stack[1][14] ), .B(o[19]), .Z(n5240) );
  NAND U6501 ( .A(n5085), .B(n5084), .Z(n5089) );
  NAND U6502 ( .A(n5087), .B(n5086), .Z(n5088) );
  AND U6503 ( .A(n5089), .B(n5088), .Z(n5238) );
  AND U6504 ( .A(\stack[1][16] ), .B(o[17]), .Z(n5246) );
  NAND U6505 ( .A(n5090), .B(n16714), .Z(n5094) );
  NAND U6506 ( .A(n5092), .B(n5091), .Z(n5093) );
  NAND U6507 ( .A(n5094), .B(n5093), .Z(n5244) );
  AND U6508 ( .A(o[15]), .B(\stack[1][18] ), .Z(n5252) );
  NAND U6509 ( .A(n5096), .B(n5095), .Z(n5100) );
  NAND U6510 ( .A(n5098), .B(n5097), .Z(n5099) );
  NAND U6511 ( .A(n5100), .B(n5099), .Z(n5250) );
  AND U6512 ( .A(o[13]), .B(\stack[1][20] ), .Z(n5258) );
  NAND U6513 ( .A(n5102), .B(n5101), .Z(n5106) );
  NAND U6514 ( .A(n5104), .B(n5103), .Z(n5105) );
  NAND U6515 ( .A(n5106), .B(n5105), .Z(n5256) );
  AND U6516 ( .A(o[11]), .B(\stack[1][22] ), .Z(n5270) );
  NAND U6517 ( .A(n5108), .B(n5107), .Z(n5112) );
  NAND U6518 ( .A(n5110), .B(n5109), .Z(n5111) );
  NAND U6519 ( .A(n5112), .B(n5111), .Z(n5268) );
  NAND U6520 ( .A(n5114), .B(n5113), .Z(n5118) );
  NAND U6521 ( .A(n5116), .B(n5115), .Z(n5117) );
  AND U6522 ( .A(n5118), .B(n5117), .Z(n5319) );
  AND U6523 ( .A(o[7]), .B(\stack[1][26] ), .Z(n5276) );
  NAND U6524 ( .A(n5120), .B(n5119), .Z(n5124) );
  NAND U6525 ( .A(n5122), .B(n5121), .Z(n5123) );
  NAND U6526 ( .A(n5124), .B(n5123), .Z(n5274) );
  AND U6527 ( .A(o[6]), .B(\stack[1][27] ), .Z(n5310) );
  NAND U6528 ( .A(n5126), .B(n5125), .Z(n5130) );
  NAND U6529 ( .A(n5128), .B(n5127), .Z(n5129) );
  NAND U6530 ( .A(n5130), .B(n5129), .Z(n5279) );
  AND U6531 ( .A(o[4]), .B(\stack[1][29] ), .Z(n5280) );
  XOR U6532 ( .A(n5279), .B(n5280), .Z(n5282) );
  AND U6533 ( .A(o[1]), .B(\stack[1][32] ), .Z(n5285) );
  NAND U6534 ( .A(\stack[1][33] ), .B(o[0]), .Z(n5131) );
  XNOR U6535 ( .A(n5285), .B(n5131), .Z(n5289) );
  NAND U6536 ( .A(n5285), .B(o[0]), .Z(n5132) );
  XNOR U6537 ( .A(o[2]), .B(n5132), .Z(n5133) );
  AND U6538 ( .A(\stack[1][31] ), .B(n5133), .Z(n5288) );
  XOR U6539 ( .A(n5289), .B(n5288), .Z(n5296) );
  AND U6540 ( .A(o[0]), .B(\stack[1][30] ), .Z(n5135) );
  AND U6541 ( .A(n5135), .B(n5134), .Z(n5136) );
  NAND U6542 ( .A(o[2]), .B(n5136), .Z(n5140) );
  NAND U6543 ( .A(n5138), .B(n5137), .Z(n5139) );
  NAND U6544 ( .A(n5140), .B(n5139), .Z(n5295) );
  XOR U6545 ( .A(n5296), .B(n5295), .Z(n5298) );
  AND U6546 ( .A(o[3]), .B(\stack[1][30] ), .Z(n5297) );
  XOR U6547 ( .A(n5298), .B(n5297), .Z(n5281) );
  XOR U6548 ( .A(n5282), .B(n5281), .Z(n5302) );
  AND U6549 ( .A(o[5]), .B(\stack[1][28] ), .Z(n5301) );
  XOR U6550 ( .A(n5302), .B(n5301), .Z(n5304) );
  NAND U6551 ( .A(n5142), .B(n5141), .Z(n5146) );
  NAND U6552 ( .A(n5144), .B(n5143), .Z(n5145) );
  NAND U6553 ( .A(n5146), .B(n5145), .Z(n5303) );
  XOR U6554 ( .A(n5304), .B(n5303), .Z(n5308) );
  NAND U6555 ( .A(n5148), .B(n5147), .Z(n5152) );
  NAND U6556 ( .A(n5150), .B(n5149), .Z(n5151) );
  NAND U6557 ( .A(n5152), .B(n5151), .Z(n5307) );
  XOR U6558 ( .A(n5308), .B(n5307), .Z(n5309) );
  XOR U6559 ( .A(n5310), .B(n5309), .Z(n5273) );
  XOR U6560 ( .A(n5276), .B(n5275), .Z(n5316) );
  AND U6561 ( .A(o[8]), .B(\stack[1][25] ), .Z(n5313) );
  NAND U6562 ( .A(n5154), .B(n5153), .Z(n5158) );
  NAND U6563 ( .A(n5156), .B(n5155), .Z(n5157) );
  NAND U6564 ( .A(n5158), .B(n5157), .Z(n5314) );
  XNOR U6565 ( .A(n5316), .B(n5315), .Z(n5320) );
  NAND U6566 ( .A(o[9]), .B(\stack[1][24] ), .Z(n5321) );
  XNOR U6567 ( .A(n5322), .B(n5321), .Z(n5328) );
  AND U6568 ( .A(o[10]), .B(\stack[1][23] ), .Z(n5325) );
  NAND U6569 ( .A(n5160), .B(n5159), .Z(n5164) );
  NAND U6570 ( .A(n5162), .B(n5161), .Z(n5163) );
  NAND U6571 ( .A(n5164), .B(n5163), .Z(n5326) );
  XOR U6572 ( .A(n5270), .B(n5269), .Z(n5264) );
  AND U6573 ( .A(o[12]), .B(\stack[1][21] ), .Z(n5261) );
  NAND U6574 ( .A(n5166), .B(n5165), .Z(n5170) );
  NAND U6575 ( .A(n5168), .B(n5167), .Z(n5169) );
  NAND U6576 ( .A(n5170), .B(n5169), .Z(n5262) );
  XOR U6577 ( .A(n5264), .B(n5263), .Z(n5255) );
  XOR U6578 ( .A(n5258), .B(n5257), .Z(n5334) );
  AND U6579 ( .A(o[14]), .B(\stack[1][19] ), .Z(n5331) );
  NAND U6580 ( .A(n5172), .B(n5171), .Z(n5176) );
  NAND U6581 ( .A(n5174), .B(n5173), .Z(n5175) );
  NAND U6582 ( .A(n5176), .B(n5175), .Z(n5332) );
  XOR U6583 ( .A(n5334), .B(n5333), .Z(n5249) );
  XOR U6584 ( .A(n5252), .B(n5251), .Z(n5340) );
  AND U6585 ( .A(\stack[1][17] ), .B(o[16]), .Z(n5337) );
  NAND U6586 ( .A(n5178), .B(n5177), .Z(n5182) );
  NAND U6587 ( .A(n5180), .B(n5179), .Z(n5181) );
  NAND U6588 ( .A(n5182), .B(n5181), .Z(n5338) );
  XOR U6589 ( .A(n5340), .B(n5339), .Z(n5243) );
  XOR U6590 ( .A(n5246), .B(n5245), .Z(n5346) );
  AND U6591 ( .A(\stack[1][15] ), .B(o[18]), .Z(n5343) );
  NAND U6592 ( .A(n5184), .B(n5183), .Z(n5188) );
  NAND U6593 ( .A(n5186), .B(n5185), .Z(n5187) );
  NAND U6594 ( .A(n5188), .B(n5187), .Z(n5344) );
  XOR U6595 ( .A(n5346), .B(n5345), .Z(n5237) );
  XOR U6596 ( .A(n5238), .B(n5237), .Z(n5239) );
  XOR U6597 ( .A(n5240), .B(n5239), .Z(n5352) );
  AND U6598 ( .A(\stack[1][13] ), .B(o[20]), .Z(n5349) );
  NAND U6599 ( .A(n5190), .B(n5189), .Z(n5194) );
  NAND U6600 ( .A(n5192), .B(n5191), .Z(n5193) );
  NAND U6601 ( .A(n5194), .B(n5193), .Z(n5350) );
  XOR U6602 ( .A(n5352), .B(n5351), .Z(n5231) );
  XOR U6603 ( .A(n5234), .B(n5233), .Z(n5358) );
  AND U6604 ( .A(\stack[1][11] ), .B(o[22]), .Z(n5355) );
  NAND U6605 ( .A(n5196), .B(n5195), .Z(n5200) );
  NAND U6606 ( .A(n5198), .B(n5197), .Z(n5199) );
  NAND U6607 ( .A(n5200), .B(n5199), .Z(n5356) );
  XOR U6608 ( .A(n5358), .B(n5357), .Z(n5225) );
  XOR U6609 ( .A(n5228), .B(n5227), .Z(n5364) );
  AND U6610 ( .A(\stack[1][9] ), .B(o[24]), .Z(n5361) );
  NAND U6611 ( .A(n5202), .B(n5201), .Z(n5206) );
  NAND U6612 ( .A(n5204), .B(n5203), .Z(n5205) );
  NAND U6613 ( .A(n5206), .B(n5205), .Z(n5362) );
  XOR U6614 ( .A(n5364), .B(n5363), .Z(n5219) );
  AND U6615 ( .A(\stack[1][8] ), .B(o[25]), .Z(n5222) );
  AND U6616 ( .A(\stack[1][7] ), .B(o[26]), .Z(n5367) );
  NAND U6617 ( .A(n5208), .B(n5207), .Z(n5212) );
  NAND U6618 ( .A(n5210), .B(n5209), .Z(n5211) );
  NAND U6619 ( .A(n5212), .B(n5211), .Z(n5368) );
  XOR U6620 ( .A(n5370), .B(n5369), .Z(n5214) );
  NAND U6621 ( .A(n5213), .B(n5214), .Z(n5216) );
  AND U6622 ( .A(\stack[1][6] ), .B(o[27]), .Z(n12384) );
  NAND U6623 ( .A(n12384), .B(n12385), .Z(n5215) );
  NAND U6624 ( .A(n5216), .B(n5215), .Z(n5217) );
  AND U6625 ( .A(\stack[1][6] ), .B(o[28]), .Z(n5218) );
  NAND U6626 ( .A(n5217), .B(n5218), .Z(n5374) );
  NAND U6627 ( .A(n5220), .B(n5219), .Z(n5224) );
  NAND U6628 ( .A(n5222), .B(n5221), .Z(n5223) );
  NAND U6629 ( .A(n5224), .B(n5223), .Z(n5376) );
  AND U6630 ( .A(\stack[1][8] ), .B(o[26]), .Z(n5375) );
  NAND U6631 ( .A(n5226), .B(n5225), .Z(n5230) );
  NAND U6632 ( .A(n5228), .B(n5227), .Z(n5229) );
  NAND U6633 ( .A(n5230), .B(n5229), .Z(n5382) );
  AND U6634 ( .A(\stack[1][10] ), .B(o[24]), .Z(n5381) );
  NAND U6635 ( .A(n5232), .B(n5231), .Z(n5236) );
  NAND U6636 ( .A(n5234), .B(n5233), .Z(n5235) );
  NAND U6637 ( .A(n5236), .B(n5235), .Z(n5388) );
  AND U6638 ( .A(\stack[1][12] ), .B(o[22]), .Z(n5387) );
  NAND U6639 ( .A(n5238), .B(n5237), .Z(n5242) );
  NAND U6640 ( .A(n5240), .B(n5239), .Z(n5241) );
  NAND U6641 ( .A(n5242), .B(n5241), .Z(n5394) );
  AND U6642 ( .A(\stack[1][14] ), .B(o[20]), .Z(n5393) );
  NAND U6643 ( .A(n5244), .B(n5243), .Z(n5248) );
  NAND U6644 ( .A(n5246), .B(n5245), .Z(n5247) );
  NAND U6645 ( .A(n5248), .B(n5247), .Z(n5400) );
  AND U6646 ( .A(\stack[1][16] ), .B(o[18]), .Z(n5399) );
  AND U6647 ( .A(\stack[1][17] ), .B(o[17]), .Z(n5502) );
  NAND U6648 ( .A(n5250), .B(n5249), .Z(n5254) );
  NAND U6649 ( .A(n5252), .B(n5251), .Z(n5253) );
  NAND U6650 ( .A(n5254), .B(n5253), .Z(n5406) );
  AND U6651 ( .A(o[16]), .B(\stack[1][18] ), .Z(n5405) );
  NAND U6652 ( .A(n5256), .B(n5255), .Z(n5260) );
  NAND U6653 ( .A(n5258), .B(n5257), .Z(n5259) );
  NAND U6654 ( .A(n5260), .B(n5259), .Z(n5412) );
  AND U6655 ( .A(o[14]), .B(\stack[1][20] ), .Z(n5411) );
  NAND U6656 ( .A(n5262), .B(n5261), .Z(n5266) );
  NAND U6657 ( .A(n5264), .B(n5263), .Z(n5265) );
  NAND U6658 ( .A(n5266), .B(n5265), .Z(n5488) );
  NAND U6659 ( .A(n5268), .B(n5267), .Z(n5272) );
  NAND U6660 ( .A(n5270), .B(n5269), .Z(n5271) );
  AND U6661 ( .A(n5272), .B(n5271), .Z(n5417) );
  NAND U6662 ( .A(o[12]), .B(\stack[1][22] ), .Z(n5418) );
  NAND U6663 ( .A(n5274), .B(n5273), .Z(n5278) );
  NAND U6664 ( .A(n5276), .B(n5275), .Z(n5277) );
  NAND U6665 ( .A(n5278), .B(n5277), .Z(n5430) );
  AND U6666 ( .A(o[8]), .B(\stack[1][26] ), .Z(n5429) );
  AND U6667 ( .A(o[6]), .B(\stack[1][28] ), .Z(n5438) );
  NAND U6668 ( .A(n5280), .B(n5279), .Z(n5284) );
  NAND U6669 ( .A(n5282), .B(n5281), .Z(n5283) );
  NAND U6670 ( .A(n5284), .B(n5283), .Z(n5463) );
  AND U6671 ( .A(o[3]), .B(\stack[1][31] ), .Z(n5443) );
  AND U6672 ( .A(o[0]), .B(\stack[1][31] ), .Z(n5286) );
  AND U6673 ( .A(n5286), .B(n5285), .Z(n5287) );
  NAND U6674 ( .A(o[2]), .B(n5287), .Z(n5291) );
  NAND U6675 ( .A(n5289), .B(n5288), .Z(n5290) );
  NAND U6676 ( .A(n5291), .B(n5290), .Z(n5441) );
  AND U6677 ( .A(o[1]), .B(\stack[1][33] ), .Z(n5450) );
  NAND U6678 ( .A(\stack[1][34] ), .B(o[0]), .Z(n5292) );
  XNOR U6679 ( .A(n5450), .B(n5292), .Z(n5454) );
  NAND U6680 ( .A(n5450), .B(o[0]), .Z(n5293) );
  XNOR U6681 ( .A(o[2]), .B(n5293), .Z(n5294) );
  AND U6682 ( .A(\stack[1][32] ), .B(n5294), .Z(n5453) );
  XOR U6683 ( .A(n5454), .B(n5453), .Z(n5442) );
  XOR U6684 ( .A(n5441), .B(n5442), .Z(n5444) );
  AND U6685 ( .A(o[4]), .B(\stack[1][30] ), .Z(n5458) );
  NAND U6686 ( .A(n5296), .B(n5295), .Z(n5300) );
  NAND U6687 ( .A(n5298), .B(n5297), .Z(n5299) );
  NAND U6688 ( .A(n5300), .B(n5299), .Z(n5457) );
  XOR U6689 ( .A(n5458), .B(n5457), .Z(n5459) );
  XOR U6690 ( .A(n5460), .B(n5459), .Z(n5464) );
  XOR U6691 ( .A(n5463), .B(n5464), .Z(n5466) );
  AND U6692 ( .A(o[5]), .B(\stack[1][29] ), .Z(n5465) );
  XOR U6693 ( .A(n5466), .B(n5465), .Z(n5436) );
  NAND U6694 ( .A(n5302), .B(n5301), .Z(n5306) );
  NAND U6695 ( .A(n5304), .B(n5303), .Z(n5305) );
  NAND U6696 ( .A(n5306), .B(n5305), .Z(n5435) );
  XOR U6697 ( .A(n5436), .B(n5435), .Z(n5437) );
  XOR U6698 ( .A(n5438), .B(n5437), .Z(n5470) );
  NAND U6699 ( .A(n5308), .B(n5307), .Z(n5312) );
  NAND U6700 ( .A(n5310), .B(n5309), .Z(n5311) );
  NAND U6701 ( .A(n5312), .B(n5311), .Z(n5469) );
  XOR U6702 ( .A(n5470), .B(n5469), .Z(n5472) );
  AND U6703 ( .A(o[7]), .B(\stack[1][27] ), .Z(n5471) );
  XOR U6704 ( .A(n5472), .B(n5471), .Z(n5431) );
  XOR U6705 ( .A(n5432), .B(n5431), .Z(n5475) );
  NAND U6706 ( .A(n5314), .B(n5313), .Z(n5318) );
  NAND U6707 ( .A(n5316), .B(n5315), .Z(n5317) );
  NAND U6708 ( .A(n5318), .B(n5317), .Z(n5476) );
  AND U6709 ( .A(o[9]), .B(\stack[1][25] ), .Z(n5478) );
  NAND U6710 ( .A(n5320), .B(n5319), .Z(n5324) );
  NAND U6711 ( .A(n5322), .B(n5321), .Z(n5323) );
  AND U6712 ( .A(n5324), .B(n5323), .Z(n5423) );
  AND U6713 ( .A(o[10]), .B(\stack[1][24] ), .Z(n5424) );
  XNOR U6714 ( .A(n5426), .B(n5425), .Z(n5482) );
  NAND U6715 ( .A(n5326), .B(n5325), .Z(n5330) );
  NAND U6716 ( .A(n5328), .B(n5327), .Z(n5329) );
  AND U6717 ( .A(n5330), .B(n5329), .Z(n5481) );
  NAND U6718 ( .A(o[11]), .B(\stack[1][23] ), .Z(n5484) );
  XNOR U6719 ( .A(n5420), .B(n5419), .Z(n5487) );
  AND U6720 ( .A(o[13]), .B(\stack[1][21] ), .Z(n5490) );
  XOR U6721 ( .A(n5414), .B(n5413), .Z(n5493) );
  NAND U6722 ( .A(n5332), .B(n5331), .Z(n5336) );
  NAND U6723 ( .A(n5334), .B(n5333), .Z(n5335) );
  NAND U6724 ( .A(n5336), .B(n5335), .Z(n5494) );
  AND U6725 ( .A(o[15]), .B(\stack[1][19] ), .Z(n5496) );
  XOR U6726 ( .A(n5408), .B(n5407), .Z(n5499) );
  NAND U6727 ( .A(n5338), .B(n5337), .Z(n5342) );
  NAND U6728 ( .A(n5340), .B(n5339), .Z(n5341) );
  NAND U6729 ( .A(n5342), .B(n5341), .Z(n5500) );
  XOR U6730 ( .A(n5502), .B(n5501), .Z(n5401) );
  XOR U6731 ( .A(n5402), .B(n5401), .Z(n5505) );
  NAND U6732 ( .A(n5344), .B(n5343), .Z(n5348) );
  NAND U6733 ( .A(n5346), .B(n5345), .Z(n5347) );
  NAND U6734 ( .A(n5348), .B(n5347), .Z(n5506) );
  AND U6735 ( .A(\stack[1][15] ), .B(o[19]), .Z(n5508) );
  XOR U6736 ( .A(n5396), .B(n5395), .Z(n5511) );
  NAND U6737 ( .A(n5350), .B(n5349), .Z(n5354) );
  NAND U6738 ( .A(n5352), .B(n5351), .Z(n5353) );
  NAND U6739 ( .A(n5354), .B(n5353), .Z(n5512) );
  AND U6740 ( .A(\stack[1][13] ), .B(o[21]), .Z(n5514) );
  XOR U6741 ( .A(n5390), .B(n5389), .Z(n5517) );
  NAND U6742 ( .A(n5356), .B(n5355), .Z(n5360) );
  NAND U6743 ( .A(n5358), .B(n5357), .Z(n5359) );
  NAND U6744 ( .A(n5360), .B(n5359), .Z(n5518) );
  AND U6745 ( .A(\stack[1][11] ), .B(o[23]), .Z(n5520) );
  XOR U6746 ( .A(n5384), .B(n5383), .Z(n5523) );
  NAND U6747 ( .A(n5362), .B(n5361), .Z(n5366) );
  NAND U6748 ( .A(n5364), .B(n5363), .Z(n5365) );
  NAND U6749 ( .A(n5366), .B(n5365), .Z(n5524) );
  AND U6750 ( .A(\stack[1][9] ), .B(o[25]), .Z(n5526) );
  XOR U6751 ( .A(n5378), .B(n5377), .Z(n5529) );
  NAND U6752 ( .A(n5368), .B(n5367), .Z(n5372) );
  NAND U6753 ( .A(n5370), .B(n5369), .Z(n5371) );
  NAND U6754 ( .A(n5372), .B(n5371), .Z(n5530) );
  AND U6755 ( .A(\stack[1][7] ), .B(o[27]), .Z(n5532) );
  NAND U6756 ( .A(n12391), .B(n12390), .Z(n5373) );
  NAND U6757 ( .A(n5374), .B(n5373), .Z(n5535) );
  NAND U6758 ( .A(n5376), .B(n5375), .Z(n5380) );
  NAND U6759 ( .A(n5378), .B(n5377), .Z(n5379) );
  NAND U6760 ( .A(n5380), .B(n5379), .Z(n5542) );
  AND U6761 ( .A(\stack[1][10] ), .B(o[25]), .Z(n5550) );
  NAND U6762 ( .A(n5382), .B(n5381), .Z(n5386) );
  NAND U6763 ( .A(n5384), .B(n5383), .Z(n5385) );
  NAND U6764 ( .A(n5386), .B(n5385), .Z(n5548) );
  NAND U6765 ( .A(n5388), .B(n5387), .Z(n5392) );
  NAND U6766 ( .A(n5390), .B(n5389), .Z(n5391) );
  NAND U6767 ( .A(n5392), .B(n5391), .Z(n5554) );
  NAND U6768 ( .A(n5394), .B(n5393), .Z(n5398) );
  NAND U6769 ( .A(n5396), .B(n5395), .Z(n5397) );
  NAND U6770 ( .A(n5398), .B(n5397), .Z(n5678) );
  NAND U6771 ( .A(n5400), .B(n5399), .Z(n5404) );
  NAND U6772 ( .A(n5402), .B(n5401), .Z(n5403) );
  NAND U6773 ( .A(n5404), .B(n5403), .Z(n5560) );
  NAND U6774 ( .A(n5406), .B(n5405), .Z(n5410) );
  NAND U6775 ( .A(n5408), .B(n5407), .Z(n5409) );
  NAND U6776 ( .A(n5410), .B(n5409), .Z(n5566) );
  NAND U6777 ( .A(n5412), .B(n5411), .Z(n5416) );
  NAND U6778 ( .A(n5414), .B(n5413), .Z(n5415) );
  NAND U6779 ( .A(n5416), .B(n5415), .Z(n5572) );
  NAND U6780 ( .A(n5418), .B(n5417), .Z(n5422) );
  NAND U6781 ( .A(n5420), .B(n5419), .Z(n5421) );
  NAND U6782 ( .A(n5422), .B(n5421), .Z(n5578) );
  NAND U6783 ( .A(n5424), .B(n5423), .Z(n5428) );
  NAND U6784 ( .A(n5426), .B(n5425), .Z(n5427) );
  NAND U6785 ( .A(n5428), .B(n5427), .Z(n5590) );
  NAND U6786 ( .A(n5430), .B(n5429), .Z(n5434) );
  NAND U6787 ( .A(n5432), .B(n5431), .Z(n5433) );
  AND U6788 ( .A(n5434), .B(n5433), .Z(n5641) );
  NAND U6789 ( .A(n5436), .B(n5435), .Z(n5440) );
  NAND U6790 ( .A(n5438), .B(n5437), .Z(n5439) );
  NAND U6791 ( .A(n5440), .B(n5439), .Z(n5629) );
  AND U6792 ( .A(o[6]), .B(\stack[1][29] ), .Z(n5626) );
  NAND U6793 ( .A(n5442), .B(n5441), .Z(n5446) );
  NAND U6794 ( .A(n5444), .B(n5443), .Z(n5445) );
  NAND U6795 ( .A(n5446), .B(n5445), .Z(n5595) );
  AND U6796 ( .A(o[4]), .B(\stack[1][31] ), .Z(n5596) );
  XOR U6797 ( .A(n5595), .B(n5596), .Z(n5598) );
  AND U6798 ( .A(o[1]), .B(\stack[1][34] ), .Z(n5601) );
  NAND U6799 ( .A(\stack[1][35] ), .B(o[0]), .Z(n5447) );
  XNOR U6800 ( .A(n5601), .B(n5447), .Z(n5605) );
  NAND U6801 ( .A(n5601), .B(o[0]), .Z(n5448) );
  XNOR U6802 ( .A(o[2]), .B(n5448), .Z(n5449) );
  AND U6803 ( .A(\stack[1][33] ), .B(n5449), .Z(n5604) );
  XOR U6804 ( .A(n5605), .B(n5604), .Z(n5612) );
  AND U6805 ( .A(o[0]), .B(\stack[1][32] ), .Z(n5451) );
  AND U6806 ( .A(n5451), .B(n5450), .Z(n5452) );
  NAND U6807 ( .A(o[2]), .B(n5452), .Z(n5456) );
  NAND U6808 ( .A(n5454), .B(n5453), .Z(n5455) );
  NAND U6809 ( .A(n5456), .B(n5455), .Z(n5611) );
  XOR U6810 ( .A(n5612), .B(n5611), .Z(n5614) );
  AND U6811 ( .A(o[3]), .B(\stack[1][32] ), .Z(n5613) );
  XOR U6812 ( .A(n5614), .B(n5613), .Z(n5597) );
  XOR U6813 ( .A(n5598), .B(n5597), .Z(n5618) );
  AND U6814 ( .A(o[5]), .B(\stack[1][30] ), .Z(n5617) );
  XOR U6815 ( .A(n5618), .B(n5617), .Z(n5620) );
  NAND U6816 ( .A(n5458), .B(n5457), .Z(n5462) );
  NAND U6817 ( .A(n5460), .B(n5459), .Z(n5461) );
  NAND U6818 ( .A(n5462), .B(n5461), .Z(n5619) );
  XOR U6819 ( .A(n5620), .B(n5619), .Z(n5624) );
  NAND U6820 ( .A(n5464), .B(n5463), .Z(n5468) );
  NAND U6821 ( .A(n5466), .B(n5465), .Z(n5467) );
  NAND U6822 ( .A(n5468), .B(n5467), .Z(n5623) );
  XOR U6823 ( .A(n5624), .B(n5623), .Z(n5625) );
  XOR U6824 ( .A(n5626), .B(n5625), .Z(n5630) );
  XOR U6825 ( .A(n5629), .B(n5630), .Z(n5632) );
  AND U6826 ( .A(o[7]), .B(\stack[1][28] ), .Z(n5631) );
  XOR U6827 ( .A(n5632), .B(n5631), .Z(n5638) );
  AND U6828 ( .A(o[8]), .B(\stack[1][27] ), .Z(n5636) );
  NAND U6829 ( .A(n5470), .B(n5469), .Z(n5474) );
  NAND U6830 ( .A(n5472), .B(n5471), .Z(n5473) );
  NAND U6831 ( .A(n5474), .B(n5473), .Z(n5635) );
  XOR U6832 ( .A(n5636), .B(n5635), .Z(n5637) );
  XNOR U6833 ( .A(n5638), .B(n5637), .Z(n5642) );
  NAND U6834 ( .A(o[9]), .B(\stack[1][26] ), .Z(n5643) );
  XNOR U6835 ( .A(n5644), .B(n5643), .Z(n5650) );
  AND U6836 ( .A(o[10]), .B(\stack[1][25] ), .Z(n5648) );
  NAND U6837 ( .A(n5476), .B(n5475), .Z(n5480) );
  NAND U6838 ( .A(n5478), .B(n5477), .Z(n5479) );
  NAND U6839 ( .A(n5480), .B(n5479), .Z(n5647) );
  XOR U6840 ( .A(n5648), .B(n5647), .Z(n5649) );
  AND U6841 ( .A(o[11]), .B(\stack[1][24] ), .Z(n5592) );
  AND U6842 ( .A(o[12]), .B(\stack[1][23] ), .Z(n5583) );
  NAND U6843 ( .A(n5482), .B(n5481), .Z(n5486) );
  NAND U6844 ( .A(n5484), .B(n5483), .Z(n5485) );
  AND U6845 ( .A(n5486), .B(n5485), .Z(n5584) );
  XNOR U6846 ( .A(n5586), .B(n5585), .Z(n5577) );
  NAND U6847 ( .A(o[13]), .B(\stack[1][22] ), .Z(n5579) );
  XNOR U6848 ( .A(n5580), .B(n5579), .Z(n5656) );
  AND U6849 ( .A(o[14]), .B(\stack[1][21] ), .Z(n5653) );
  NAND U6850 ( .A(n5488), .B(n5487), .Z(n5492) );
  NAND U6851 ( .A(n5490), .B(n5489), .Z(n5491) );
  NAND U6852 ( .A(n5492), .B(n5491), .Z(n5654) );
  AND U6853 ( .A(o[15]), .B(\stack[1][20] ), .Z(n5574) );
  AND U6854 ( .A(o[16]), .B(\stack[1][19] ), .Z(n5659) );
  NAND U6855 ( .A(n5494), .B(n5493), .Z(n5498) );
  NAND U6856 ( .A(n5496), .B(n5495), .Z(n5497) );
  NAND U6857 ( .A(n5498), .B(n5497), .Z(n5660) );
  XOR U6858 ( .A(n5662), .B(n5661), .Z(n5565) );
  AND U6859 ( .A(\stack[1][18] ), .B(o[17]), .Z(n5568) );
  AND U6860 ( .A(\stack[1][17] ), .B(o[18]), .Z(n5665) );
  NAND U6861 ( .A(n5500), .B(n5499), .Z(n5504) );
  NAND U6862 ( .A(n5502), .B(n5501), .Z(n5503) );
  NAND U6863 ( .A(n5504), .B(n5503), .Z(n5666) );
  XOR U6864 ( .A(n5668), .B(n5667), .Z(n5559) );
  AND U6865 ( .A(\stack[1][16] ), .B(o[19]), .Z(n5562) );
  AND U6866 ( .A(\stack[1][15] ), .B(o[20]), .Z(n5671) );
  NAND U6867 ( .A(n5506), .B(n5505), .Z(n5510) );
  NAND U6868 ( .A(n5508), .B(n5507), .Z(n5509) );
  NAND U6869 ( .A(n5510), .B(n5509), .Z(n5672) );
  XOR U6870 ( .A(n5674), .B(n5673), .Z(n5677) );
  AND U6871 ( .A(\stack[1][14] ), .B(o[21]), .Z(n5680) );
  AND U6872 ( .A(\stack[1][13] ), .B(o[22]), .Z(n5683) );
  NAND U6873 ( .A(n5512), .B(n5511), .Z(n5516) );
  NAND U6874 ( .A(n5514), .B(n5513), .Z(n5515) );
  NAND U6875 ( .A(n5516), .B(n5515), .Z(n5684) );
  XOR U6876 ( .A(n5686), .B(n5685), .Z(n5553) );
  AND U6877 ( .A(\stack[1][12] ), .B(o[23]), .Z(n5556) );
  AND U6878 ( .A(\stack[1][11] ), .B(o[24]), .Z(n5689) );
  NAND U6879 ( .A(n5518), .B(n5517), .Z(n5522) );
  NAND U6880 ( .A(n5520), .B(n5519), .Z(n5521) );
  NAND U6881 ( .A(n5522), .B(n5521), .Z(n5690) );
  XOR U6882 ( .A(n5692), .B(n5691), .Z(n5547) );
  XOR U6883 ( .A(n5550), .B(n5549), .Z(n5698) );
  AND U6884 ( .A(\stack[1][9] ), .B(o[26]), .Z(n5695) );
  NAND U6885 ( .A(n5524), .B(n5523), .Z(n5528) );
  NAND U6886 ( .A(n5526), .B(n5525), .Z(n5527) );
  NAND U6887 ( .A(n5528), .B(n5527), .Z(n5696) );
  XOR U6888 ( .A(n5698), .B(n5697), .Z(n5541) );
  AND U6889 ( .A(\stack[1][8] ), .B(o[27]), .Z(n5544) );
  AND U6890 ( .A(\stack[1][7] ), .B(o[28]), .Z(n5701) );
  NAND U6891 ( .A(n5530), .B(n5529), .Z(n5534) );
  NAND U6892 ( .A(n5532), .B(n5531), .Z(n5533) );
  NAND U6893 ( .A(n5534), .B(n5533), .Z(n5702) );
  XOR U6894 ( .A(n5704), .B(n5703), .Z(n5536) );
  NAND U6895 ( .A(n5535), .B(n5536), .Z(n5538) );
  AND U6896 ( .A(\stack[1][6] ), .B(o[29]), .Z(n12397) );
  NAND U6897 ( .A(n12397), .B(n12396), .Z(n5537) );
  NAND U6898 ( .A(n5538), .B(n5537), .Z(n5539) );
  AND U6899 ( .A(\stack[1][6] ), .B(o[30]), .Z(n5540) );
  NAND U6900 ( .A(n5539), .B(n5540), .Z(n5708) );
  NAND U6901 ( .A(n5542), .B(n5541), .Z(n5546) );
  NAND U6902 ( .A(n5544), .B(n5543), .Z(n5545) );
  NAND U6903 ( .A(n5546), .B(n5545), .Z(n5710) );
  AND U6904 ( .A(\stack[1][8] ), .B(o[28]), .Z(n5709) );
  NAND U6905 ( .A(n5548), .B(n5547), .Z(n5552) );
  NAND U6906 ( .A(n5550), .B(n5549), .Z(n5551) );
  NAND U6907 ( .A(n5552), .B(n5551), .Z(n5716) );
  AND U6908 ( .A(\stack[1][10] ), .B(o[26]), .Z(n5715) );
  NAND U6909 ( .A(n5554), .B(n5553), .Z(n5558) );
  NAND U6910 ( .A(n5556), .B(n5555), .Z(n5557) );
  NAND U6911 ( .A(n5558), .B(n5557), .Z(n5722) );
  AND U6912 ( .A(\stack[1][12] ), .B(o[24]), .Z(n5721) );
  NAND U6913 ( .A(n5560), .B(n5559), .Z(n5564) );
  NAND U6914 ( .A(n5562), .B(n5561), .Z(n5563) );
  NAND U6915 ( .A(n5564), .B(n5563), .Z(n5734) );
  AND U6916 ( .A(\stack[1][16] ), .B(o[20]), .Z(n5733) );
  AND U6917 ( .A(\stack[1][18] ), .B(o[18]), .Z(n16637) );
  NAND U6918 ( .A(n5566), .B(n5565), .Z(n5570) );
  NAND U6919 ( .A(n5568), .B(n5567), .Z(n5569) );
  NAND U6920 ( .A(n5570), .B(n5569), .Z(n5739) );
  NAND U6921 ( .A(n5572), .B(n5571), .Z(n5576) );
  NAND U6922 ( .A(n5574), .B(n5573), .Z(n5575) );
  NAND U6923 ( .A(n5576), .B(n5575), .Z(n5745) );
  AND U6924 ( .A(o[16]), .B(\stack[1][20] ), .Z(n5744) );
  NAND U6925 ( .A(n5578), .B(n5577), .Z(n5582) );
  NAND U6926 ( .A(n5580), .B(n5579), .Z(n5581) );
  AND U6927 ( .A(n5582), .B(n5581), .Z(n5750) );
  AND U6928 ( .A(o[14]), .B(\stack[1][22] ), .Z(n5751) );
  NAND U6929 ( .A(n5584), .B(n5583), .Z(n5588) );
  NAND U6930 ( .A(n5586), .B(n5585), .Z(n5587) );
  NAND U6931 ( .A(n5588), .B(n5587), .Z(n5827) );
  NAND U6932 ( .A(n5590), .B(n5589), .Z(n5594) );
  NAND U6933 ( .A(n5592), .B(n5591), .Z(n5593) );
  AND U6934 ( .A(n5594), .B(n5593), .Z(n5756) );
  NAND U6935 ( .A(o[12]), .B(\stack[1][24] ), .Z(n5757) );
  AND U6936 ( .A(o[6]), .B(\stack[1][30] ), .Z(n5777) );
  AND U6937 ( .A(o[5]), .B(\stack[1][31] ), .Z(n5804) );
  NAND U6938 ( .A(n5596), .B(n5595), .Z(n5600) );
  NAND U6939 ( .A(n5598), .B(n5597), .Z(n5599) );
  NAND U6940 ( .A(n5600), .B(n5599), .Z(n5802) );
  AND U6941 ( .A(o[0]), .B(\stack[1][33] ), .Z(n5602) );
  AND U6942 ( .A(n5602), .B(n5601), .Z(n5603) );
  NAND U6943 ( .A(o[2]), .B(n5603), .Z(n5607) );
  NAND U6944 ( .A(n5605), .B(n5604), .Z(n5606) );
  NAND U6945 ( .A(n5607), .B(n5606), .Z(n5780) );
  AND U6946 ( .A(o[1]), .B(\stack[1][35] ), .Z(n5789) );
  NAND U6947 ( .A(\stack[1][36] ), .B(o[0]), .Z(n5608) );
  XNOR U6948 ( .A(n5789), .B(n5608), .Z(n5793) );
  NAND U6949 ( .A(n5789), .B(o[0]), .Z(n5609) );
  XNOR U6950 ( .A(o[2]), .B(n5609), .Z(n5610) );
  AND U6951 ( .A(\stack[1][34] ), .B(n5610), .Z(n5792) );
  XOR U6952 ( .A(n5793), .B(n5792), .Z(n5781) );
  XOR U6953 ( .A(n5780), .B(n5781), .Z(n5783) );
  AND U6954 ( .A(o[3]), .B(\stack[1][33] ), .Z(n5782) );
  XOR U6955 ( .A(n5783), .B(n5782), .Z(n5799) );
  AND U6956 ( .A(o[4]), .B(\stack[1][32] ), .Z(n5797) );
  NAND U6957 ( .A(n5612), .B(n5611), .Z(n5616) );
  NAND U6958 ( .A(n5614), .B(n5613), .Z(n5615) );
  NAND U6959 ( .A(n5616), .B(n5615), .Z(n5796) );
  XOR U6960 ( .A(n5797), .B(n5796), .Z(n5798) );
  XOR U6961 ( .A(n5799), .B(n5798), .Z(n5803) );
  XOR U6962 ( .A(n5802), .B(n5803), .Z(n5805) );
  NAND U6963 ( .A(n5618), .B(n5617), .Z(n5622) );
  NAND U6964 ( .A(n5620), .B(n5619), .Z(n5621) );
  NAND U6965 ( .A(n5622), .B(n5621), .Z(n5774) );
  XOR U6966 ( .A(n5775), .B(n5774), .Z(n5776) );
  XOR U6967 ( .A(n5777), .B(n5776), .Z(n5809) );
  NAND U6968 ( .A(n5624), .B(n5623), .Z(n5628) );
  NAND U6969 ( .A(n5626), .B(n5625), .Z(n5627) );
  NAND U6970 ( .A(n5628), .B(n5627), .Z(n5808) );
  XOR U6971 ( .A(n5809), .B(n5808), .Z(n5811) );
  AND U6972 ( .A(o[7]), .B(\stack[1][29] ), .Z(n5810) );
  XOR U6973 ( .A(n5811), .B(n5810), .Z(n5770) );
  NAND U6974 ( .A(n5630), .B(n5629), .Z(n5634) );
  NAND U6975 ( .A(n5632), .B(n5631), .Z(n5633) );
  NAND U6976 ( .A(n5634), .B(n5633), .Z(n5768) );
  AND U6977 ( .A(o[8]), .B(\stack[1][28] ), .Z(n5769) );
  XOR U6978 ( .A(n5768), .B(n5769), .Z(n5771) );
  NAND U6979 ( .A(n5636), .B(n5635), .Z(n5640) );
  NAND U6980 ( .A(n5638), .B(n5637), .Z(n5639) );
  NAND U6981 ( .A(n5640), .B(n5639), .Z(n5814) );
  XOR U6982 ( .A(n5815), .B(n5814), .Z(n5817) );
  AND U6983 ( .A(o[9]), .B(\stack[1][27] ), .Z(n5816) );
  XOR U6984 ( .A(n5817), .B(n5816), .Z(n5765) );
  AND U6985 ( .A(o[10]), .B(\stack[1][26] ), .Z(n5763) );
  NAND U6986 ( .A(n5642), .B(n5641), .Z(n5646) );
  NAND U6987 ( .A(n5644), .B(n5643), .Z(n5645) );
  AND U6988 ( .A(n5646), .B(n5645), .Z(n5762) );
  XOR U6989 ( .A(n5763), .B(n5762), .Z(n5764) );
  XNOR U6990 ( .A(n5765), .B(n5764), .Z(n5821) );
  NAND U6991 ( .A(n5648), .B(n5647), .Z(n5652) );
  NAND U6992 ( .A(n5650), .B(n5649), .Z(n5651) );
  AND U6993 ( .A(n5652), .B(n5651), .Z(n5820) );
  NAND U6994 ( .A(o[11]), .B(\stack[1][25] ), .Z(n5822) );
  XOR U6995 ( .A(n5823), .B(n5822), .Z(n5758) );
  XNOR U6996 ( .A(n5759), .B(n5758), .Z(n5826) );
  AND U6997 ( .A(o[13]), .B(\stack[1][23] ), .Z(n5829) );
  XOR U6998 ( .A(n5753), .B(n5752), .Z(n5832) );
  NAND U6999 ( .A(n5654), .B(n5653), .Z(n5658) );
  NAND U7000 ( .A(n5656), .B(n5655), .Z(n5657) );
  NAND U7001 ( .A(n5658), .B(n5657), .Z(n5833) );
  AND U7002 ( .A(o[15]), .B(\stack[1][21] ), .Z(n5835) );
  XOR U7003 ( .A(n5747), .B(n5746), .Z(n5838) );
  NAND U7004 ( .A(n5660), .B(n5659), .Z(n5664) );
  NAND U7005 ( .A(n5662), .B(n5661), .Z(n5663) );
  NAND U7006 ( .A(n5664), .B(n5663), .Z(n5839) );
  AND U7007 ( .A(\stack[1][19] ), .B(o[17]), .Z(n5841) );
  XOR U7008 ( .A(n5741), .B(n5740), .Z(n5844) );
  NAND U7009 ( .A(n5666), .B(n5665), .Z(n5670) );
  NAND U7010 ( .A(n5668), .B(n5667), .Z(n5669) );
  NAND U7011 ( .A(n5670), .B(n5669), .Z(n5845) );
  AND U7012 ( .A(\stack[1][17] ), .B(o[19]), .Z(n5847) );
  XOR U7013 ( .A(n5736), .B(n5735), .Z(n5850) );
  NAND U7014 ( .A(n5672), .B(n5671), .Z(n5676) );
  NAND U7015 ( .A(n5674), .B(n5673), .Z(n5675) );
  NAND U7016 ( .A(n5676), .B(n5675), .Z(n5851) );
  AND U7017 ( .A(\stack[1][15] ), .B(o[21]), .Z(n5852) );
  XNOR U7018 ( .A(n5853), .B(n5852), .Z(n5730) );
  NAND U7019 ( .A(n5678), .B(n5677), .Z(n5682) );
  NAND U7020 ( .A(n5680), .B(n5679), .Z(n5681) );
  AND U7021 ( .A(n5682), .B(n5681), .Z(n5727) );
  NAND U7022 ( .A(\stack[1][14] ), .B(o[22]), .Z(n5728) );
  NAND U7023 ( .A(n5684), .B(n5683), .Z(n5688) );
  NAND U7024 ( .A(n5686), .B(n5685), .Z(n5687) );
  NAND U7025 ( .A(n5688), .B(n5687), .Z(n5856) );
  XOR U7026 ( .A(n5857), .B(n5856), .Z(n5858) );
  AND U7027 ( .A(\stack[1][13] ), .B(o[23]), .Z(n5859) );
  XOR U7028 ( .A(n5724), .B(n5723), .Z(n5862) );
  NAND U7029 ( .A(n5690), .B(n5689), .Z(n5694) );
  NAND U7030 ( .A(n5692), .B(n5691), .Z(n5693) );
  NAND U7031 ( .A(n5694), .B(n5693), .Z(n5863) );
  AND U7032 ( .A(\stack[1][11] ), .B(o[25]), .Z(n5865) );
  XOR U7033 ( .A(n5718), .B(n5717), .Z(n5868) );
  NAND U7034 ( .A(n5696), .B(n5695), .Z(n5700) );
  NAND U7035 ( .A(n5698), .B(n5697), .Z(n5699) );
  NAND U7036 ( .A(n5700), .B(n5699), .Z(n5869) );
  AND U7037 ( .A(\stack[1][9] ), .B(o[27]), .Z(n5871) );
  XOR U7038 ( .A(n5712), .B(n5711), .Z(n5874) );
  NAND U7039 ( .A(n5702), .B(n5701), .Z(n5706) );
  NAND U7040 ( .A(n5704), .B(n5703), .Z(n5705) );
  NAND U7041 ( .A(n5706), .B(n5705), .Z(n5875) );
  AND U7042 ( .A(\stack[1][7] ), .B(o[29]), .Z(n5877) );
  NAND U7043 ( .A(n12403), .B(n12402), .Z(n5707) );
  NAND U7044 ( .A(n5708), .B(n5707), .Z(n5880) );
  NAND U7045 ( .A(n5710), .B(n5709), .Z(n5714) );
  NAND U7046 ( .A(n5712), .B(n5711), .Z(n5713) );
  NAND U7047 ( .A(n5714), .B(n5713), .Z(n6053) );
  AND U7048 ( .A(\stack[1][10] ), .B(o[27]), .Z(n5889) );
  NAND U7049 ( .A(n5716), .B(n5715), .Z(n5720) );
  NAND U7050 ( .A(n5718), .B(n5717), .Z(n5719) );
  NAND U7051 ( .A(n5720), .B(n5719), .Z(n5887) );
  NAND U7052 ( .A(n5722), .B(n5721), .Z(n5726) );
  NAND U7053 ( .A(n5724), .B(n5723), .Z(n5725) );
  NAND U7054 ( .A(n5726), .B(n5725), .Z(n5893) );
  AND U7055 ( .A(\stack[1][14] ), .B(o[23]), .Z(n5901) );
  NAND U7056 ( .A(n5728), .B(n5727), .Z(n5732) );
  NAND U7057 ( .A(n5730), .B(n5729), .Z(n5731) );
  AND U7058 ( .A(n5732), .B(n5731), .Z(n5899) );
  NAND U7059 ( .A(n5734), .B(n5733), .Z(n5738) );
  NAND U7060 ( .A(n5736), .B(n5735), .Z(n5737) );
  NAND U7061 ( .A(n5738), .B(n5737), .Z(n5905) );
  AND U7062 ( .A(\stack[1][18] ), .B(o[19]), .Z(n6019) );
  NAND U7063 ( .A(n5739), .B(n16637), .Z(n5743) );
  NAND U7064 ( .A(n5741), .B(n5740), .Z(n5742) );
  NAND U7065 ( .A(n5743), .B(n5742), .Z(n6017) );
  AND U7066 ( .A(o[17]), .B(\stack[1][20] ), .Z(n5919) );
  NAND U7067 ( .A(n5745), .B(n5744), .Z(n5749) );
  NAND U7068 ( .A(n5747), .B(n5746), .Z(n5748) );
  NAND U7069 ( .A(n5749), .B(n5748), .Z(n5917) );
  NAND U7070 ( .A(n5751), .B(n5750), .Z(n5755) );
  NAND U7071 ( .A(n5753), .B(n5752), .Z(n5754) );
  NAND U7072 ( .A(n5755), .B(n5754), .Z(n5929) );
  NAND U7073 ( .A(n5757), .B(n5756), .Z(n5761) );
  NAND U7074 ( .A(n5759), .B(n5758), .Z(n5760) );
  AND U7075 ( .A(n5761), .B(n5760), .Z(n6005) );
  AND U7076 ( .A(o[11]), .B(\stack[1][26] ), .Z(n5936) );
  NAND U7077 ( .A(n5763), .B(n5762), .Z(n5767) );
  NAND U7078 ( .A(n5765), .B(n5764), .Z(n5766) );
  NAND U7079 ( .A(n5767), .B(n5766), .Z(n5934) );
  NAND U7080 ( .A(n5769), .B(n5768), .Z(n5773) );
  NAND U7081 ( .A(n5771), .B(n5770), .Z(n5772) );
  AND U7082 ( .A(n5773), .B(n5772), .Z(n5986) );
  AND U7083 ( .A(o[7]), .B(\stack[1][30] ), .Z(n5942) );
  NAND U7084 ( .A(n5775), .B(n5774), .Z(n5779) );
  NAND U7085 ( .A(n5777), .B(n5776), .Z(n5778) );
  NAND U7086 ( .A(n5779), .B(n5778), .Z(n5940) );
  AND U7087 ( .A(o[6]), .B(\stack[1][31] ), .Z(n5977) );
  NAND U7088 ( .A(n5781), .B(n5780), .Z(n5785) );
  NAND U7089 ( .A(n5783), .B(n5782), .Z(n5784) );
  NAND U7090 ( .A(n5785), .B(n5784), .Z(n5946) );
  AND U7091 ( .A(o[4]), .B(\stack[1][33] ), .Z(n5947) );
  XOR U7092 ( .A(n5946), .B(n5947), .Z(n5949) );
  AND U7093 ( .A(o[1]), .B(\stack[1][36] ), .Z(n5958) );
  NAND U7094 ( .A(\stack[1][37] ), .B(o[0]), .Z(n5786) );
  XNOR U7095 ( .A(n5958), .B(n5786), .Z(n5962) );
  NAND U7096 ( .A(n5958), .B(o[0]), .Z(n5787) );
  XNOR U7097 ( .A(o[2]), .B(n5787), .Z(n5788) );
  AND U7098 ( .A(\stack[1][35] ), .B(n5788), .Z(n5961) );
  XOR U7099 ( .A(n5962), .B(n5961), .Z(n5953) );
  AND U7100 ( .A(o[0]), .B(\stack[1][34] ), .Z(n5790) );
  AND U7101 ( .A(n5790), .B(n5789), .Z(n5791) );
  NAND U7102 ( .A(o[2]), .B(n5791), .Z(n5795) );
  NAND U7103 ( .A(n5793), .B(n5792), .Z(n5794) );
  NAND U7104 ( .A(n5795), .B(n5794), .Z(n5952) );
  XOR U7105 ( .A(n5953), .B(n5952), .Z(n5955) );
  AND U7106 ( .A(o[3]), .B(\stack[1][34] ), .Z(n5954) );
  XOR U7107 ( .A(n5955), .B(n5954), .Z(n5948) );
  XOR U7108 ( .A(n5949), .B(n5948), .Z(n5969) );
  AND U7109 ( .A(o[5]), .B(\stack[1][32] ), .Z(n5968) );
  XOR U7110 ( .A(n5969), .B(n5968), .Z(n5971) );
  NAND U7111 ( .A(n5797), .B(n5796), .Z(n5801) );
  NAND U7112 ( .A(n5799), .B(n5798), .Z(n5800) );
  NAND U7113 ( .A(n5801), .B(n5800), .Z(n5970) );
  XOR U7114 ( .A(n5971), .B(n5970), .Z(n5975) );
  NAND U7115 ( .A(n5803), .B(n5802), .Z(n5807) );
  NAND U7116 ( .A(n5805), .B(n5804), .Z(n5806) );
  NAND U7117 ( .A(n5807), .B(n5806), .Z(n5974) );
  XOR U7118 ( .A(n5975), .B(n5974), .Z(n5976) );
  XOR U7119 ( .A(n5977), .B(n5976), .Z(n5941) );
  XOR U7120 ( .A(n5940), .B(n5941), .Z(n5943) );
  AND U7121 ( .A(o[8]), .B(\stack[1][29] ), .Z(n5981) );
  NAND U7122 ( .A(n5809), .B(n5808), .Z(n5813) );
  NAND U7123 ( .A(n5811), .B(n5810), .Z(n5812) );
  NAND U7124 ( .A(n5813), .B(n5812), .Z(n5980) );
  XOR U7125 ( .A(n5981), .B(n5980), .Z(n5982) );
  XNOR U7126 ( .A(n5983), .B(n5982), .Z(n5987) );
  NAND U7127 ( .A(o[9]), .B(\stack[1][28] ), .Z(n5988) );
  XNOR U7128 ( .A(n5989), .B(n5988), .Z(n5995) );
  AND U7129 ( .A(o[10]), .B(\stack[1][27] ), .Z(n5993) );
  NAND U7130 ( .A(n5815), .B(n5814), .Z(n5819) );
  NAND U7131 ( .A(n5817), .B(n5816), .Z(n5818) );
  NAND U7132 ( .A(n5819), .B(n5818), .Z(n5992) );
  XOR U7133 ( .A(n5993), .B(n5992), .Z(n5994) );
  XOR U7134 ( .A(n5934), .B(n5935), .Z(n5937) );
  XNOR U7135 ( .A(n5936), .B(n5937), .Z(n6001) );
  AND U7136 ( .A(o[12]), .B(\stack[1][25] ), .Z(n5999) );
  NAND U7137 ( .A(n5821), .B(n5820), .Z(n5825) );
  NAND U7138 ( .A(n5823), .B(n5822), .Z(n5824) );
  AND U7139 ( .A(n5825), .B(n5824), .Z(n5998) );
  XOR U7140 ( .A(n5999), .B(n5998), .Z(n6000) );
  XOR U7141 ( .A(n6001), .B(n6000), .Z(n6004) );
  XOR U7142 ( .A(n6005), .B(n6004), .Z(n6007) );
  AND U7143 ( .A(o[13]), .B(\stack[1][24] ), .Z(n6006) );
  XOR U7144 ( .A(n6007), .B(n6006), .Z(n6013) );
  AND U7145 ( .A(o[14]), .B(\stack[1][23] ), .Z(n6011) );
  NAND U7146 ( .A(n5827), .B(n5826), .Z(n5831) );
  NAND U7147 ( .A(n5829), .B(n5828), .Z(n5830) );
  NAND U7148 ( .A(n5831), .B(n5830), .Z(n6010) );
  XOR U7149 ( .A(n6011), .B(n6010), .Z(n6012) );
  XOR U7150 ( .A(n6013), .B(n6012), .Z(n5928) );
  AND U7151 ( .A(o[15]), .B(\stack[1][22] ), .Z(n5931) );
  AND U7152 ( .A(o[16]), .B(\stack[1][21] ), .Z(n5922) );
  NAND U7153 ( .A(n5833), .B(n5832), .Z(n5837) );
  NAND U7154 ( .A(n5835), .B(n5834), .Z(n5836) );
  NAND U7155 ( .A(n5837), .B(n5836), .Z(n5923) );
  XOR U7156 ( .A(n5925), .B(n5924), .Z(n5916) );
  XOR U7157 ( .A(n5919), .B(n5918), .Z(n5913) );
  AND U7158 ( .A(\stack[1][19] ), .B(o[18]), .Z(n5910) );
  NAND U7159 ( .A(n5839), .B(n5838), .Z(n5843) );
  NAND U7160 ( .A(n5841), .B(n5840), .Z(n5842) );
  NAND U7161 ( .A(n5843), .B(n5842), .Z(n5911) );
  XOR U7162 ( .A(n5913), .B(n5912), .Z(n6016) );
  XOR U7163 ( .A(n6019), .B(n6018), .Z(n6025) );
  AND U7164 ( .A(\stack[1][17] ), .B(o[20]), .Z(n6022) );
  NAND U7165 ( .A(n5845), .B(n5844), .Z(n5849) );
  NAND U7166 ( .A(n5847), .B(n5846), .Z(n5848) );
  NAND U7167 ( .A(n5849), .B(n5848), .Z(n6023) );
  XOR U7168 ( .A(n6025), .B(n6024), .Z(n5904) );
  AND U7169 ( .A(\stack[1][16] ), .B(o[21]), .Z(n5907) );
  AND U7170 ( .A(\stack[1][15] ), .B(o[22]), .Z(n6028) );
  NAND U7171 ( .A(n5851), .B(n5850), .Z(n5855) );
  NAND U7172 ( .A(n5853), .B(n5852), .Z(n5854) );
  NAND U7173 ( .A(n5855), .B(n5854), .Z(n6029) );
  XOR U7174 ( .A(n6031), .B(n6030), .Z(n5898) );
  XOR U7175 ( .A(n5899), .B(n5898), .Z(n5900) );
  XOR U7176 ( .A(n5901), .B(n5900), .Z(n6037) );
  AND U7177 ( .A(\stack[1][13] ), .B(o[24]), .Z(n6034) );
  NAND U7178 ( .A(n5857), .B(n5856), .Z(n5861) );
  NAND U7179 ( .A(n5859), .B(n5858), .Z(n5860) );
  NAND U7180 ( .A(n5861), .B(n5860), .Z(n6035) );
  XOR U7181 ( .A(n6037), .B(n6036), .Z(n5892) );
  AND U7182 ( .A(\stack[1][12] ), .B(o[25]), .Z(n5895) );
  AND U7183 ( .A(\stack[1][11] ), .B(o[26]), .Z(n6040) );
  NAND U7184 ( .A(n5863), .B(n5862), .Z(n5867) );
  NAND U7185 ( .A(n5865), .B(n5864), .Z(n5866) );
  NAND U7186 ( .A(n5867), .B(n5866), .Z(n6041) );
  XOR U7187 ( .A(n6043), .B(n6042), .Z(n5886) );
  XOR U7188 ( .A(n5889), .B(n5888), .Z(n6049) );
  AND U7189 ( .A(\stack[1][9] ), .B(o[28]), .Z(n6046) );
  NAND U7190 ( .A(n5869), .B(n5868), .Z(n5873) );
  NAND U7191 ( .A(n5871), .B(n5870), .Z(n5872) );
  NAND U7192 ( .A(n5873), .B(n5872), .Z(n6047) );
  XOR U7193 ( .A(n6049), .B(n6048), .Z(n6052) );
  AND U7194 ( .A(\stack[1][8] ), .B(o[29]), .Z(n6055) );
  AND U7195 ( .A(\stack[1][7] ), .B(o[30]), .Z(n6058) );
  NAND U7196 ( .A(n5875), .B(n5874), .Z(n5879) );
  NAND U7197 ( .A(n5877), .B(n5876), .Z(n5878) );
  NAND U7198 ( .A(n5879), .B(n5878), .Z(n6059) );
  XOR U7199 ( .A(n6061), .B(n6060), .Z(n5881) );
  NAND U7200 ( .A(n5880), .B(n5881), .Z(n5883) );
  AND U7201 ( .A(\stack[1][6] ), .B(o[31]), .Z(n12408) );
  NAND U7202 ( .A(n12408), .B(n12409), .Z(n5882) );
  AND U7203 ( .A(n5883), .B(n5882), .Z(n5885) );
  NAND U7204 ( .A(n5884), .B(n5885), .Z(n6065) );
  NAND U7205 ( .A(n5887), .B(n5886), .Z(n5891) );
  NAND U7206 ( .A(n5889), .B(n5888), .Z(n5890) );
  AND U7207 ( .A(n5891), .B(n5890), .Z(n6072) );
  NAND U7208 ( .A(\stack[1][10] ), .B(o[28]), .Z(n6073) );
  NAND U7209 ( .A(n5893), .B(n5892), .Z(n5897) );
  NAND U7210 ( .A(n5895), .B(n5894), .Z(n5896) );
  NAND U7211 ( .A(n5897), .B(n5896), .Z(n6079) );
  AND U7212 ( .A(\stack[1][12] ), .B(o[26]), .Z(n6078) );
  NAND U7213 ( .A(n5899), .B(n5898), .Z(n5903) );
  NAND U7214 ( .A(n5901), .B(n5900), .Z(n5902) );
  NAND U7215 ( .A(n5903), .B(n5902), .Z(n6085) );
  AND U7216 ( .A(\stack[1][14] ), .B(o[24]), .Z(n6084) );
  NAND U7217 ( .A(n5905), .B(n5904), .Z(n5909) );
  NAND U7218 ( .A(n5907), .B(n5906), .Z(n5908) );
  NAND U7219 ( .A(n5909), .B(n5908), .Z(n6091) );
  AND U7220 ( .A(\stack[1][16] ), .B(o[22]), .Z(n6090) );
  AND U7221 ( .A(\stack[1][19] ), .B(o[19]), .Z(n6211) );
  NAND U7222 ( .A(n5911), .B(n5910), .Z(n5915) );
  NAND U7223 ( .A(n5913), .B(n5912), .Z(n5914) );
  NAND U7224 ( .A(n5915), .B(n5914), .Z(n6209) );
  NAND U7225 ( .A(n5917), .B(n5916), .Z(n5921) );
  NAND U7226 ( .A(n5919), .B(n5918), .Z(n5920) );
  AND U7227 ( .A(n5921), .B(n5920), .Z(n6102) );
  NAND U7228 ( .A(o[18]), .B(\stack[1][20] ), .Z(n6103) );
  NAND U7229 ( .A(n5923), .B(n5922), .Z(n5927) );
  NAND U7230 ( .A(n5925), .B(n5924), .Z(n5926) );
  NAND U7231 ( .A(n5927), .B(n5926), .Z(n6203) );
  NAND U7232 ( .A(n5929), .B(n5928), .Z(n5933) );
  NAND U7233 ( .A(n5931), .B(n5930), .Z(n5932) );
  AND U7234 ( .A(n5933), .B(n5932), .Z(n6108) );
  NAND U7235 ( .A(o[16]), .B(\stack[1][22] ), .Z(n6109) );
  NANDN U7236 ( .A(n5935), .B(n5934), .Z(n5939) );
  NANDN U7237 ( .A(n5937), .B(n5936), .Z(n5938) );
  AND U7238 ( .A(n5939), .B(n5938), .Z(n6121) );
  NAND U7239 ( .A(o[12]), .B(\stack[1][26] ), .Z(n6120) );
  XOR U7240 ( .A(n6121), .B(n6120), .Z(n6123) );
  NAND U7241 ( .A(n5941), .B(n5940), .Z(n5945) );
  NAND U7242 ( .A(n5943), .B(n5942), .Z(n5944) );
  NAND U7243 ( .A(n5945), .B(n5944), .Z(n6132) );
  AND U7244 ( .A(o[8]), .B(\stack[1][30] ), .Z(n6133) );
  XOR U7245 ( .A(n6132), .B(n6133), .Z(n6135) );
  AND U7246 ( .A(o[5]), .B(\stack[1][33] ), .Z(n6168) );
  NAND U7247 ( .A(n5947), .B(n5946), .Z(n5951) );
  NAND U7248 ( .A(n5949), .B(n5948), .Z(n5950) );
  NAND U7249 ( .A(n5951), .B(n5950), .Z(n6166) );
  AND U7250 ( .A(o[4]), .B(\stack[1][34] ), .Z(n6145) );
  NAND U7251 ( .A(n5953), .B(n5952), .Z(n5957) );
  NAND U7252 ( .A(n5955), .B(n5954), .Z(n5956) );
  NAND U7253 ( .A(n5957), .B(n5956), .Z(n6144) );
  XOR U7254 ( .A(n6145), .B(n6144), .Z(n6147) );
  AND U7255 ( .A(o[0]), .B(\stack[1][35] ), .Z(n5959) );
  AND U7256 ( .A(n5959), .B(n5958), .Z(n5960) );
  NAND U7257 ( .A(o[2]), .B(n5960), .Z(n5964) );
  NAND U7258 ( .A(n5962), .B(n5961), .Z(n5963) );
  NAND U7259 ( .A(n5964), .B(n5963), .Z(n6160) );
  AND U7260 ( .A(o[3]), .B(\stack[1][35] ), .Z(n6161) );
  XOR U7261 ( .A(n6160), .B(n6161), .Z(n6163) );
  AND U7262 ( .A(o[1]), .B(\stack[1][37] ), .Z(n6150) );
  NAND U7263 ( .A(\stack[1][38] ), .B(o[0]), .Z(n5965) );
  XNOR U7264 ( .A(n6150), .B(n5965), .Z(n6154) );
  NAND U7265 ( .A(n6150), .B(o[0]), .Z(n5966) );
  XNOR U7266 ( .A(o[2]), .B(n5966), .Z(n5967) );
  AND U7267 ( .A(\stack[1][36] ), .B(n5967), .Z(n6153) );
  XOR U7268 ( .A(n6154), .B(n6153), .Z(n6162) );
  XOR U7269 ( .A(n6163), .B(n6162), .Z(n6146) );
  XOR U7270 ( .A(n6147), .B(n6146), .Z(n6167) );
  XOR U7271 ( .A(n6166), .B(n6167), .Z(n6169) );
  NAND U7272 ( .A(n5969), .B(n5968), .Z(n5973) );
  NAND U7273 ( .A(n5971), .B(n5970), .Z(n5972) );
  NAND U7274 ( .A(n5973), .B(n5972), .Z(n6138) );
  XOR U7275 ( .A(n6139), .B(n6138), .Z(n6141) );
  AND U7276 ( .A(o[6]), .B(\stack[1][32] ), .Z(n6140) );
  XOR U7277 ( .A(n6141), .B(n6140), .Z(n6173) );
  NAND U7278 ( .A(n5975), .B(n5974), .Z(n5979) );
  NAND U7279 ( .A(n5977), .B(n5976), .Z(n5978) );
  NAND U7280 ( .A(n5979), .B(n5978), .Z(n6172) );
  XOR U7281 ( .A(n6173), .B(n6172), .Z(n6175) );
  AND U7282 ( .A(o[7]), .B(\stack[1][31] ), .Z(n6174) );
  XOR U7283 ( .A(n6175), .B(n6174), .Z(n6134) );
  XOR U7284 ( .A(n6135), .B(n6134), .Z(n6179) );
  NAND U7285 ( .A(n5981), .B(n5980), .Z(n5985) );
  NAND U7286 ( .A(n5983), .B(n5982), .Z(n5984) );
  NAND U7287 ( .A(n5985), .B(n5984), .Z(n6178) );
  XOR U7288 ( .A(n6179), .B(n6178), .Z(n6181) );
  AND U7289 ( .A(o[9]), .B(\stack[1][29] ), .Z(n6180) );
  XOR U7290 ( .A(n6181), .B(n6180), .Z(n6129) );
  AND U7291 ( .A(o[10]), .B(\stack[1][28] ), .Z(n6127) );
  NAND U7292 ( .A(n5987), .B(n5986), .Z(n5991) );
  NAND U7293 ( .A(n5989), .B(n5988), .Z(n5990) );
  AND U7294 ( .A(n5991), .B(n5990), .Z(n6126) );
  XOR U7295 ( .A(n6127), .B(n6126), .Z(n6128) );
  XNOR U7296 ( .A(n6129), .B(n6128), .Z(n6185) );
  NAND U7297 ( .A(n5993), .B(n5992), .Z(n5997) );
  NAND U7298 ( .A(n5995), .B(n5994), .Z(n5996) );
  AND U7299 ( .A(n5997), .B(n5996), .Z(n6184) );
  NAND U7300 ( .A(o[11]), .B(\stack[1][27] ), .Z(n6186) );
  XOR U7301 ( .A(n6187), .B(n6186), .Z(n6122) );
  XNOR U7302 ( .A(n6123), .B(n6122), .Z(n6191) );
  NAND U7303 ( .A(n5999), .B(n5998), .Z(n6003) );
  NAND U7304 ( .A(n6001), .B(n6000), .Z(n6002) );
  NAND U7305 ( .A(n6003), .B(n6002), .Z(n6190) );
  AND U7306 ( .A(o[13]), .B(\stack[1][25] ), .Z(n6192) );
  XOR U7307 ( .A(n6193), .B(n6192), .Z(n6116) );
  NAND U7308 ( .A(n6005), .B(n6004), .Z(n6009) );
  NAND U7309 ( .A(n6007), .B(n6006), .Z(n6008) );
  NAND U7310 ( .A(n6009), .B(n6008), .Z(n6114) );
  AND U7311 ( .A(o[14]), .B(\stack[1][24] ), .Z(n6115) );
  XOR U7312 ( .A(n6114), .B(n6115), .Z(n6117) );
  NAND U7313 ( .A(n6011), .B(n6010), .Z(n6015) );
  NAND U7314 ( .A(n6013), .B(n6012), .Z(n6014) );
  NAND U7315 ( .A(n6015), .B(n6014), .Z(n6196) );
  XOR U7316 ( .A(n6197), .B(n6196), .Z(n6199) );
  AND U7317 ( .A(o[15]), .B(\stack[1][23] ), .Z(n6198) );
  XNOR U7318 ( .A(n6199), .B(n6198), .Z(n6110) );
  XNOR U7319 ( .A(n6111), .B(n6110), .Z(n6202) );
  AND U7320 ( .A(o[17]), .B(\stack[1][21] ), .Z(n6204) );
  XNOR U7321 ( .A(n6205), .B(n6204), .Z(n6104) );
  XNOR U7322 ( .A(n6105), .B(n6104), .Z(n6208) );
  XNOR U7323 ( .A(n6211), .B(n6210), .Z(n6099) );
  NAND U7324 ( .A(n6017), .B(n6016), .Z(n6021) );
  NAND U7325 ( .A(n6019), .B(n6018), .Z(n6020) );
  AND U7326 ( .A(n6021), .B(n6020), .Z(n6096) );
  NAND U7327 ( .A(\stack[1][18] ), .B(o[20]), .Z(n6097) );
  NAND U7328 ( .A(n6023), .B(n6022), .Z(n6027) );
  NAND U7329 ( .A(n6025), .B(n6024), .Z(n6026) );
  NAND U7330 ( .A(n6027), .B(n6026), .Z(n6214) );
  XOR U7331 ( .A(n6215), .B(n6214), .Z(n6216) );
  AND U7332 ( .A(\stack[1][17] ), .B(o[21]), .Z(n6217) );
  XOR U7333 ( .A(n6093), .B(n6092), .Z(n6220) );
  NAND U7334 ( .A(n6029), .B(n6028), .Z(n6033) );
  NAND U7335 ( .A(n6031), .B(n6030), .Z(n6032) );
  NAND U7336 ( .A(n6033), .B(n6032), .Z(n6221) );
  AND U7337 ( .A(\stack[1][15] ), .B(o[23]), .Z(n6223) );
  XOR U7338 ( .A(n6087), .B(n6086), .Z(n6226) );
  NAND U7339 ( .A(n6035), .B(n6034), .Z(n6039) );
  NAND U7340 ( .A(n6037), .B(n6036), .Z(n6038) );
  NAND U7341 ( .A(n6039), .B(n6038), .Z(n6227) );
  AND U7342 ( .A(\stack[1][13] ), .B(o[25]), .Z(n6229) );
  XOR U7343 ( .A(n6081), .B(n6080), .Z(n6232) );
  NAND U7344 ( .A(n6041), .B(n6040), .Z(n6045) );
  NAND U7345 ( .A(n6043), .B(n6042), .Z(n6044) );
  NAND U7346 ( .A(n6045), .B(n6044), .Z(n6233) );
  AND U7347 ( .A(\stack[1][11] ), .B(o[27]), .Z(n6234) );
  XNOR U7348 ( .A(n6235), .B(n6234), .Z(n6074) );
  XNOR U7349 ( .A(n6075), .B(n6074), .Z(n6239) );
  NAND U7350 ( .A(n6047), .B(n6046), .Z(n6051) );
  NAND U7351 ( .A(n6049), .B(n6048), .Z(n6050) );
  NAND U7352 ( .A(n6051), .B(n6050), .Z(n6238) );
  AND U7353 ( .A(\stack[1][9] ), .B(o[29]), .Z(n6240) );
  XNOR U7354 ( .A(n6241), .B(n6240), .Z(n6069) );
  NAND U7355 ( .A(n6053), .B(n6052), .Z(n6057) );
  NAND U7356 ( .A(n6055), .B(n6054), .Z(n6056) );
  AND U7357 ( .A(n6057), .B(n6056), .Z(n6066) );
  NAND U7358 ( .A(\stack[1][8] ), .B(o[30]), .Z(n6067) );
  NAND U7359 ( .A(n6059), .B(n6058), .Z(n6063) );
  NAND U7360 ( .A(n6061), .B(n6060), .Z(n6062) );
  NAND U7361 ( .A(n6063), .B(n6062), .Z(n6244) );
  XOR U7362 ( .A(n6245), .B(n6244), .Z(n6247) );
  AND U7363 ( .A(\stack[1][7] ), .B(o[31]), .Z(n6246) );
  XNOR U7364 ( .A(n6247), .B(n6246), .Z(n12225) );
  NAND U7365 ( .A(n12226), .B(n12225), .Z(n6064) );
  AND U7366 ( .A(n6065), .B(n6064), .Z(n6251) );
  AND U7367 ( .A(\stack[1][8] ), .B(o[31]), .Z(n6259) );
  NAND U7368 ( .A(n6067), .B(n6066), .Z(n6071) );
  NAND U7369 ( .A(n6069), .B(n6068), .Z(n6070) );
  AND U7370 ( .A(n6071), .B(n6070), .Z(n6257) );
  NAND U7371 ( .A(n6073), .B(n6072), .Z(n6077) );
  NAND U7372 ( .A(n6075), .B(n6074), .Z(n6076) );
  AND U7373 ( .A(n6077), .B(n6076), .Z(n6263) );
  NAND U7374 ( .A(n6079), .B(n6078), .Z(n6083) );
  NAND U7375 ( .A(n6081), .B(n6080), .Z(n6082) );
  NAND U7376 ( .A(n6083), .B(n6082), .Z(n6425) );
  NAND U7377 ( .A(n6085), .B(n6084), .Z(n6089) );
  NAND U7378 ( .A(n6087), .B(n6086), .Z(n6088) );
  NAND U7379 ( .A(n6089), .B(n6088), .Z(n6275) );
  AND U7380 ( .A(\stack[1][16] ), .B(o[23]), .Z(n6289) );
  NAND U7381 ( .A(n6091), .B(n6090), .Z(n6095) );
  NAND U7382 ( .A(n6093), .B(n6092), .Z(n6094) );
  NAND U7383 ( .A(n6095), .B(n6094), .Z(n6287) );
  AND U7384 ( .A(\stack[1][18] ), .B(o[21]), .Z(n6301) );
  NAND U7385 ( .A(n6097), .B(n6096), .Z(n6101) );
  NAND U7386 ( .A(n6099), .B(n6098), .Z(n6100) );
  AND U7387 ( .A(n6101), .B(n6100), .Z(n6299) );
  NAND U7388 ( .A(n6103), .B(n6102), .Z(n6107) );
  NAND U7389 ( .A(n6105), .B(n6104), .Z(n6106) );
  AND U7390 ( .A(n6107), .B(n6106), .Z(n6413) );
  NAND U7391 ( .A(n6109), .B(n6108), .Z(n6113) );
  NAND U7392 ( .A(n6111), .B(n6110), .Z(n6112) );
  AND U7393 ( .A(n6113), .B(n6112), .Z(n6305) );
  AND U7394 ( .A(o[15]), .B(\stack[1][24] ), .Z(n6312) );
  NAND U7395 ( .A(n6115), .B(n6114), .Z(n6119) );
  NAND U7396 ( .A(n6117), .B(n6116), .Z(n6118) );
  NAND U7397 ( .A(n6119), .B(n6118), .Z(n6310) );
  NAND U7398 ( .A(n6121), .B(n6120), .Z(n6125) );
  NAND U7399 ( .A(n6123), .B(n6122), .Z(n6124) );
  NAND U7400 ( .A(n6125), .B(n6124), .Z(n6317) );
  AND U7401 ( .A(o[11]), .B(\stack[1][28] ), .Z(n6324) );
  NAND U7402 ( .A(n6127), .B(n6126), .Z(n6131) );
  NAND U7403 ( .A(n6129), .B(n6128), .Z(n6130) );
  NAND U7404 ( .A(n6131), .B(n6130), .Z(n6322) );
  NAND U7405 ( .A(n6133), .B(n6132), .Z(n6137) );
  NAND U7406 ( .A(n6135), .B(n6134), .Z(n6136) );
  AND U7407 ( .A(n6137), .B(n6136), .Z(n6334) );
  NAND U7408 ( .A(n6139), .B(n6138), .Z(n6143) );
  NAND U7409 ( .A(n6141), .B(n6140), .Z(n6142) );
  AND U7410 ( .A(n6143), .B(n6142), .Z(n6376) );
  AND U7411 ( .A(o[5]), .B(\stack[1][34] ), .Z(n6342) );
  NAND U7412 ( .A(n6145), .B(n6144), .Z(n6149) );
  NAND U7413 ( .A(n6147), .B(n6146), .Z(n6148) );
  NAND U7414 ( .A(n6149), .B(n6148), .Z(n6340) );
  AND U7415 ( .A(o[4]), .B(\stack[1][35] ), .Z(n6349) );
  AND U7416 ( .A(o[0]), .B(\stack[1][36] ), .Z(n6151) );
  AND U7417 ( .A(n6151), .B(n6150), .Z(n6152) );
  NAND U7418 ( .A(o[2]), .B(n6152), .Z(n6156) );
  NAND U7419 ( .A(n6154), .B(n6153), .Z(n6155) );
  NAND U7420 ( .A(n6156), .B(n6155), .Z(n6364) );
  AND U7421 ( .A(o[1]), .B(\stack[1][38] ), .Z(n6352) );
  NAND U7422 ( .A(\stack[1][39] ), .B(o[0]), .Z(n6157) );
  XNOR U7423 ( .A(n6352), .B(n6157), .Z(n6356) );
  NAND U7424 ( .A(n6352), .B(o[0]), .Z(n6158) );
  XNOR U7425 ( .A(o[2]), .B(n6158), .Z(n6159) );
  AND U7426 ( .A(\stack[1][37] ), .B(n6159), .Z(n6355) );
  XOR U7427 ( .A(n6356), .B(n6355), .Z(n6365) );
  XOR U7428 ( .A(n6364), .B(n6365), .Z(n6367) );
  AND U7429 ( .A(o[3]), .B(\stack[1][36] ), .Z(n6366) );
  XOR U7430 ( .A(n6367), .B(n6366), .Z(n6347) );
  NAND U7431 ( .A(n6161), .B(n6160), .Z(n6165) );
  NAND U7432 ( .A(n6163), .B(n6162), .Z(n6164) );
  NAND U7433 ( .A(n6165), .B(n6164), .Z(n6346) );
  XOR U7434 ( .A(n6347), .B(n6346), .Z(n6348) );
  XOR U7435 ( .A(n6349), .B(n6348), .Z(n6341) );
  XOR U7436 ( .A(n6340), .B(n6341), .Z(n6343) );
  AND U7437 ( .A(o[6]), .B(\stack[1][33] ), .Z(n6371) );
  NAND U7438 ( .A(n6167), .B(n6166), .Z(n6171) );
  NAND U7439 ( .A(n6169), .B(n6168), .Z(n6170) );
  NAND U7440 ( .A(n6171), .B(n6170), .Z(n6370) );
  XOR U7441 ( .A(n6371), .B(n6370), .Z(n6372) );
  XNOR U7442 ( .A(n6373), .B(n6372), .Z(n6377) );
  NAND U7443 ( .A(o[7]), .B(\stack[1][32] ), .Z(n6378) );
  XNOR U7444 ( .A(n6379), .B(n6378), .Z(n6385) );
  AND U7445 ( .A(o[8]), .B(\stack[1][31] ), .Z(n6383) );
  NAND U7446 ( .A(n6173), .B(n6172), .Z(n6177) );
  NAND U7447 ( .A(n6175), .B(n6174), .Z(n6176) );
  NAND U7448 ( .A(n6177), .B(n6176), .Z(n6382) );
  XOR U7449 ( .A(n6383), .B(n6382), .Z(n6384) );
  NAND U7450 ( .A(o[9]), .B(\stack[1][30] ), .Z(n6336) );
  XNOR U7451 ( .A(n6337), .B(n6336), .Z(n6331) );
  AND U7452 ( .A(o[10]), .B(\stack[1][29] ), .Z(n6329) );
  NAND U7453 ( .A(n6179), .B(n6178), .Z(n6183) );
  NAND U7454 ( .A(n6181), .B(n6180), .Z(n6182) );
  NAND U7455 ( .A(n6183), .B(n6182), .Z(n6328) );
  XOR U7456 ( .A(n6329), .B(n6328), .Z(n6330) );
  XOR U7457 ( .A(n6322), .B(n6323), .Z(n6325) );
  XNOR U7458 ( .A(n6324), .B(n6325), .Z(n6391) );
  AND U7459 ( .A(o[12]), .B(\stack[1][27] ), .Z(n6389) );
  NAND U7460 ( .A(n6185), .B(n6184), .Z(n6189) );
  NAND U7461 ( .A(n6187), .B(n6186), .Z(n6188) );
  AND U7462 ( .A(n6189), .B(n6188), .Z(n6388) );
  XOR U7463 ( .A(n6389), .B(n6388), .Z(n6390) );
  XNOR U7464 ( .A(n6391), .B(n6390), .Z(n6316) );
  XOR U7465 ( .A(n6317), .B(n6316), .Z(n6319) );
  NAND U7466 ( .A(o[13]), .B(\stack[1][26] ), .Z(n6318) );
  XNOR U7467 ( .A(n6319), .B(n6318), .Z(n6397) );
  AND U7468 ( .A(o[14]), .B(\stack[1][25] ), .Z(n6395) );
  NAND U7469 ( .A(n6191), .B(n6190), .Z(n6195) );
  NAND U7470 ( .A(n6193), .B(n6192), .Z(n6194) );
  NAND U7471 ( .A(n6195), .B(n6194), .Z(n6394) );
  XOR U7472 ( .A(n6395), .B(n6394), .Z(n6396) );
  XOR U7473 ( .A(n6310), .B(n6311), .Z(n6313) );
  XNOR U7474 ( .A(n6312), .B(n6313), .Z(n6403) );
  AND U7475 ( .A(o[16]), .B(\stack[1][23] ), .Z(n6401) );
  NAND U7476 ( .A(n6197), .B(n6196), .Z(n6201) );
  NAND U7477 ( .A(n6199), .B(n6198), .Z(n6200) );
  NAND U7478 ( .A(n6201), .B(n6200), .Z(n6400) );
  XOR U7479 ( .A(n6401), .B(n6400), .Z(n6402) );
  XOR U7480 ( .A(n6403), .B(n6402), .Z(n6304) );
  XOR U7481 ( .A(n6305), .B(n6304), .Z(n6306) );
  AND U7482 ( .A(o[17]), .B(\stack[1][22] ), .Z(n6307) );
  AND U7483 ( .A(o[18]), .B(\stack[1][21] ), .Z(n6406) );
  NAND U7484 ( .A(n6203), .B(n6202), .Z(n6207) );
  NAND U7485 ( .A(n6205), .B(n6204), .Z(n6206) );
  NAND U7486 ( .A(n6207), .B(n6206), .Z(n6407) );
  XOR U7487 ( .A(n6409), .B(n6408), .Z(n6412) );
  XOR U7488 ( .A(n6413), .B(n6412), .Z(n6414) );
  AND U7489 ( .A(\stack[1][20] ), .B(o[19]), .Z(n6415) );
  AND U7490 ( .A(\stack[1][19] ), .B(o[20]), .Z(n6418) );
  NAND U7491 ( .A(n6209), .B(n6208), .Z(n6213) );
  NAND U7492 ( .A(n6211), .B(n6210), .Z(n6212) );
  NAND U7493 ( .A(n6213), .B(n6212), .Z(n6419) );
  XOR U7494 ( .A(n6421), .B(n6420), .Z(n6298) );
  XOR U7495 ( .A(n6299), .B(n6298), .Z(n6300) );
  XOR U7496 ( .A(n6301), .B(n6300), .Z(n6295) );
  AND U7497 ( .A(\stack[1][17] ), .B(o[22]), .Z(n6292) );
  NAND U7498 ( .A(n6215), .B(n6214), .Z(n6219) );
  NAND U7499 ( .A(n6217), .B(n6216), .Z(n6218) );
  NAND U7500 ( .A(n6219), .B(n6218), .Z(n6293) );
  XOR U7501 ( .A(n6295), .B(n6294), .Z(n6286) );
  XOR U7502 ( .A(n6289), .B(n6288), .Z(n6283) );
  AND U7503 ( .A(\stack[1][15] ), .B(o[24]), .Z(n6280) );
  NAND U7504 ( .A(n6221), .B(n6220), .Z(n6225) );
  NAND U7505 ( .A(n6223), .B(n6222), .Z(n6224) );
  NAND U7506 ( .A(n6225), .B(n6224), .Z(n6281) );
  XOR U7507 ( .A(n6283), .B(n6282), .Z(n6274) );
  AND U7508 ( .A(\stack[1][14] ), .B(o[25]), .Z(n6277) );
  AND U7509 ( .A(\stack[1][13] ), .B(o[26]), .Z(n6268) );
  NAND U7510 ( .A(n6227), .B(n6226), .Z(n6231) );
  NAND U7511 ( .A(n6229), .B(n6228), .Z(n6230) );
  NAND U7512 ( .A(n6231), .B(n6230), .Z(n6269) );
  XOR U7513 ( .A(n6271), .B(n6270), .Z(n6424) );
  AND U7514 ( .A(\stack[1][12] ), .B(o[27]), .Z(n6427) );
  AND U7515 ( .A(\stack[1][11] ), .B(o[28]), .Z(n6430) );
  NAND U7516 ( .A(n6233), .B(n6232), .Z(n6237) );
  NAND U7517 ( .A(n6235), .B(n6234), .Z(n6236) );
  NAND U7518 ( .A(n6237), .B(n6236), .Z(n6431) );
  XOR U7519 ( .A(n6433), .B(n6432), .Z(n6262) );
  XOR U7520 ( .A(n6263), .B(n6262), .Z(n6264) );
  AND U7521 ( .A(\stack[1][10] ), .B(o[29]), .Z(n6265) );
  AND U7522 ( .A(\stack[1][9] ), .B(o[30]), .Z(n6436) );
  NAND U7523 ( .A(n6239), .B(n6238), .Z(n6243) );
  NAND U7524 ( .A(n6241), .B(n6240), .Z(n6242) );
  NAND U7525 ( .A(n6243), .B(n6242), .Z(n6437) );
  XOR U7526 ( .A(n6439), .B(n6438), .Z(n6256) );
  XOR U7527 ( .A(n6257), .B(n6256), .Z(n6258) );
  XOR U7528 ( .A(n6259), .B(n6258), .Z(n6445) );
  AND U7529 ( .A(\stack[1][7] ), .B(o[32]), .Z(n6442) );
  NAND U7530 ( .A(n6245), .B(n6244), .Z(n6249) );
  NAND U7531 ( .A(n6247), .B(n6246), .Z(n6248) );
  NAND U7532 ( .A(n6249), .B(n6248), .Z(n6443) );
  XOR U7533 ( .A(n6445), .B(n6444), .Z(n6250) );
  NAND U7534 ( .A(n6251), .B(n6250), .Z(n6253) );
  AND U7535 ( .A(\stack[1][6] ), .B(o[33]), .Z(n12418) );
  XOR U7536 ( .A(n6251), .B(n6250), .Z(n12419) );
  NAND U7537 ( .A(n12418), .B(n12419), .Z(n6252) );
  NAND U7538 ( .A(n6253), .B(n6252), .Z(n6254) );
  AND U7539 ( .A(\stack[1][6] ), .B(o[34]), .Z(n6255) );
  NAND U7540 ( .A(n6254), .B(n6255), .Z(n6449) );
  NAND U7541 ( .A(n6257), .B(n6256), .Z(n6261) );
  NAND U7542 ( .A(n6259), .B(n6258), .Z(n6260) );
  NAND U7543 ( .A(n6261), .B(n6260), .Z(n6451) );
  AND U7544 ( .A(\stack[1][8] ), .B(o[32]), .Z(n6450) );
  NAND U7545 ( .A(n6263), .B(n6262), .Z(n6267) );
  NAND U7546 ( .A(n6265), .B(n6264), .Z(n6266) );
  NAND U7547 ( .A(n6267), .B(n6266), .Z(n6457) );
  AND U7548 ( .A(\stack[1][10] ), .B(o[30]), .Z(n6456) );
  NAND U7549 ( .A(n6269), .B(n6268), .Z(n6273) );
  NAND U7550 ( .A(n6271), .B(n6270), .Z(n6272) );
  NAND U7551 ( .A(n6273), .B(n6272), .Z(n6618) );
  NAND U7552 ( .A(n6275), .B(n6274), .Z(n6279) );
  NAND U7553 ( .A(n6277), .B(n6276), .Z(n6278) );
  AND U7554 ( .A(n6279), .B(n6278), .Z(n6468) );
  NAND U7555 ( .A(\stack[1][14] ), .B(o[26]), .Z(n6469) );
  NAND U7556 ( .A(n6281), .B(n6280), .Z(n6285) );
  NAND U7557 ( .A(n6283), .B(n6282), .Z(n6284) );
  NAND U7558 ( .A(n6285), .B(n6284), .Z(n6612) );
  NAND U7559 ( .A(n6287), .B(n6286), .Z(n6291) );
  NAND U7560 ( .A(n6289), .B(n6288), .Z(n6290) );
  AND U7561 ( .A(n6291), .B(n6290), .Z(n6474) );
  NAND U7562 ( .A(\stack[1][16] ), .B(o[24]), .Z(n6475) );
  NAND U7563 ( .A(n6293), .B(n6292), .Z(n6297) );
  NAND U7564 ( .A(n6295), .B(n6294), .Z(n6296) );
  NAND U7565 ( .A(n6297), .B(n6296), .Z(n6606) );
  NAND U7566 ( .A(n6299), .B(n6298), .Z(n6303) );
  NAND U7567 ( .A(n6301), .B(n6300), .Z(n6302) );
  AND U7568 ( .A(n6303), .B(n6302), .Z(n6480) );
  NAND U7569 ( .A(\stack[1][18] ), .B(o[22]), .Z(n6481) );
  NAND U7570 ( .A(n6305), .B(n6304), .Z(n6309) );
  NAND U7571 ( .A(n6307), .B(n6306), .Z(n6308) );
  NAND U7572 ( .A(n6309), .B(n6308), .Z(n6492) );
  AND U7573 ( .A(o[18]), .B(\stack[1][22] ), .Z(n6491) );
  NANDN U7574 ( .A(n6311), .B(n6310), .Z(n6315) );
  NANDN U7575 ( .A(n6313), .B(n6312), .Z(n6314) );
  NAND U7576 ( .A(n6315), .B(n6314), .Z(n6497) );
  AND U7577 ( .A(o[16]), .B(\stack[1][24] ), .Z(n6498) );
  XOR U7578 ( .A(n6497), .B(n6498), .Z(n6500) );
  NAND U7579 ( .A(n6317), .B(n6316), .Z(n6321) );
  NAND U7580 ( .A(n6319), .B(n6318), .Z(n6320) );
  AND U7581 ( .A(n6321), .B(n6320), .Z(n6504) );
  AND U7582 ( .A(o[14]), .B(\stack[1][26] ), .Z(n6503) );
  XOR U7583 ( .A(n6504), .B(n6503), .Z(n6506) );
  NANDN U7584 ( .A(n6323), .B(n6322), .Z(n6327) );
  NANDN U7585 ( .A(n6325), .B(n6324), .Z(n6326) );
  AND U7586 ( .A(n6327), .B(n6326), .Z(n6510) );
  NAND U7587 ( .A(o[12]), .B(\stack[1][28] ), .Z(n6509) );
  XOR U7588 ( .A(n6510), .B(n6509), .Z(n6512) );
  NAND U7589 ( .A(n6329), .B(n6328), .Z(n6333) );
  NAND U7590 ( .A(n6331), .B(n6330), .Z(n6332) );
  AND U7591 ( .A(n6333), .B(n6332), .Z(n6570) );
  NAND U7592 ( .A(n6335), .B(n6334), .Z(n6339) );
  NAND U7593 ( .A(n6337), .B(n6336), .Z(n6338) );
  NAND U7594 ( .A(n6339), .B(n6338), .Z(n6516) );
  NAND U7595 ( .A(o[10]), .B(\stack[1][30] ), .Z(n6515) );
  XOR U7596 ( .A(n6516), .B(n6515), .Z(n6518) );
  NAND U7597 ( .A(n6341), .B(n6340), .Z(n6345) );
  NAND U7598 ( .A(n6343), .B(n6342), .Z(n6344) );
  NAND U7599 ( .A(n6345), .B(n6344), .Z(n6533) );
  AND U7600 ( .A(o[6]), .B(\stack[1][34] ), .Z(n6534) );
  XOR U7601 ( .A(n6533), .B(n6534), .Z(n6536) );
  NAND U7602 ( .A(n6347), .B(n6346), .Z(n6351) );
  NAND U7603 ( .A(n6349), .B(n6348), .Z(n6350) );
  NAND U7604 ( .A(n6351), .B(n6350), .Z(n6558) );
  AND U7605 ( .A(o[3]), .B(\stack[1][37] ), .Z(n6547) );
  AND U7606 ( .A(o[0]), .B(\stack[1][37] ), .Z(n6353) );
  AND U7607 ( .A(n6353), .B(n6352), .Z(n6354) );
  NAND U7608 ( .A(o[2]), .B(n6354), .Z(n6358) );
  NAND U7609 ( .A(n6356), .B(n6355), .Z(n6357) );
  NAND U7610 ( .A(n6358), .B(n6357), .Z(n6545) );
  AND U7611 ( .A(o[2]), .B(\stack[1][38] ), .Z(n6555) );
  AND U7612 ( .A(o[0]), .B(\stack[1][38] ), .Z(n6359) );
  AND U7613 ( .A(o[1]), .B(\stack[1][39] ), .Z(n6361) );
  AND U7614 ( .A(n6359), .B(n6361), .Z(n6554) );
  AND U7615 ( .A(o[0]), .B(\stack[1][39] ), .Z(n6360) );
  AND U7616 ( .A(o[1]), .B(\stack[1][40] ), .Z(n6551) );
  AND U7617 ( .A(n6360), .B(n6551), .Z(n6724) );
  XNOR U7618 ( .A(n6554), .B(n6724), .Z(n6363) );
  AND U7619 ( .A(o[0]), .B(\stack[1][40] ), .Z(n6719) );
  OR U7620 ( .A(n6361), .B(n6719), .Z(n6362) );
  NAND U7621 ( .A(n6363), .B(n6362), .Z(n6556) );
  XNOR U7622 ( .A(n6555), .B(n6556), .Z(n6546) );
  XNOR U7623 ( .A(n6547), .B(n6548), .Z(n6542) );
  NAND U7624 ( .A(n6365), .B(n6364), .Z(n6369) );
  NAND U7625 ( .A(n6367), .B(n6366), .Z(n6368) );
  AND U7626 ( .A(n6369), .B(n6368), .Z(n6540) );
  NAND U7627 ( .A(o[4]), .B(\stack[1][36] ), .Z(n6539) );
  XOR U7628 ( .A(n6540), .B(n6539), .Z(n6541) );
  XOR U7629 ( .A(n6542), .B(n6541), .Z(n6557) );
  XOR U7630 ( .A(n6558), .B(n6557), .Z(n6560) );
  AND U7631 ( .A(o[5]), .B(\stack[1][35] ), .Z(n6559) );
  XOR U7632 ( .A(n6560), .B(n6559), .Z(n6535) );
  XOR U7633 ( .A(n6536), .B(n6535), .Z(n6528) );
  NAND U7634 ( .A(n6371), .B(n6370), .Z(n6375) );
  NAND U7635 ( .A(n6373), .B(n6372), .Z(n6374) );
  NAND U7636 ( .A(n6375), .B(n6374), .Z(n6527) );
  XOR U7637 ( .A(n6528), .B(n6527), .Z(n6530) );
  AND U7638 ( .A(o[7]), .B(\stack[1][33] ), .Z(n6529) );
  XOR U7639 ( .A(n6530), .B(n6529), .Z(n6524) );
  AND U7640 ( .A(o[8]), .B(\stack[1][32] ), .Z(n6522) );
  NAND U7641 ( .A(n6377), .B(n6376), .Z(n6381) );
  NAND U7642 ( .A(n6379), .B(n6378), .Z(n6380) );
  AND U7643 ( .A(n6381), .B(n6380), .Z(n6521) );
  XOR U7644 ( .A(n6522), .B(n6521), .Z(n6523) );
  XOR U7645 ( .A(n6524), .B(n6523), .Z(n6564) );
  NAND U7646 ( .A(n6383), .B(n6382), .Z(n6387) );
  NAND U7647 ( .A(n6385), .B(n6384), .Z(n6386) );
  NAND U7648 ( .A(n6387), .B(n6386), .Z(n6563) );
  XOR U7649 ( .A(n6564), .B(n6563), .Z(n6566) );
  AND U7650 ( .A(o[9]), .B(\stack[1][31] ), .Z(n6565) );
  XNOR U7651 ( .A(n6566), .B(n6565), .Z(n6517) );
  XOR U7652 ( .A(n6518), .B(n6517), .Z(n6569) );
  XOR U7653 ( .A(n6570), .B(n6569), .Z(n6572) );
  NAND U7654 ( .A(o[11]), .B(\stack[1][29] ), .Z(n6571) );
  XOR U7655 ( .A(n6572), .B(n6571), .Z(n6511) );
  XNOR U7656 ( .A(n6512), .B(n6511), .Z(n6576) );
  NAND U7657 ( .A(n6389), .B(n6388), .Z(n6393) );
  NAND U7658 ( .A(n6391), .B(n6390), .Z(n6392) );
  NAND U7659 ( .A(n6393), .B(n6392), .Z(n6575) );
  AND U7660 ( .A(o[13]), .B(\stack[1][27] ), .Z(n6577) );
  XOR U7661 ( .A(n6578), .B(n6577), .Z(n6505) );
  XOR U7662 ( .A(n6506), .B(n6505), .Z(n6582) );
  NAND U7663 ( .A(n6395), .B(n6394), .Z(n6399) );
  NAND U7664 ( .A(n6397), .B(n6396), .Z(n6398) );
  NAND U7665 ( .A(n6399), .B(n6398), .Z(n6581) );
  XOR U7666 ( .A(n6582), .B(n6581), .Z(n6584) );
  AND U7667 ( .A(o[15]), .B(\stack[1][25] ), .Z(n6583) );
  XOR U7668 ( .A(n6584), .B(n6583), .Z(n6499) );
  XOR U7669 ( .A(n6500), .B(n6499), .Z(n6588) );
  NAND U7670 ( .A(n6401), .B(n6400), .Z(n6405) );
  NAND U7671 ( .A(n6403), .B(n6402), .Z(n6404) );
  NAND U7672 ( .A(n6405), .B(n6404), .Z(n6587) );
  XOR U7673 ( .A(n6588), .B(n6587), .Z(n6590) );
  AND U7674 ( .A(o[17]), .B(\stack[1][23] ), .Z(n6589) );
  XOR U7675 ( .A(n6590), .B(n6589), .Z(n6493) );
  XOR U7676 ( .A(n6494), .B(n6493), .Z(n6593) );
  NAND U7677 ( .A(n6407), .B(n6406), .Z(n6411) );
  NAND U7678 ( .A(n6409), .B(n6408), .Z(n6410) );
  NAND U7679 ( .A(n6411), .B(n6410), .Z(n6594) );
  AND U7680 ( .A(\stack[1][21] ), .B(o[19]), .Z(n6596) );
  AND U7681 ( .A(\stack[1][20] ), .B(o[20]), .Z(n16560) );
  NAND U7682 ( .A(n6413), .B(n6412), .Z(n6417) );
  NAND U7683 ( .A(n6415), .B(n6414), .Z(n6416) );
  NAND U7684 ( .A(n6417), .B(n6416), .Z(n6486) );
  XOR U7685 ( .A(n6488), .B(n6487), .Z(n6599) );
  NAND U7686 ( .A(n6419), .B(n6418), .Z(n6423) );
  NAND U7687 ( .A(n6421), .B(n6420), .Z(n6422) );
  NAND U7688 ( .A(n6423), .B(n6422), .Z(n6600) );
  AND U7689 ( .A(\stack[1][19] ), .B(o[21]), .Z(n6601) );
  XNOR U7690 ( .A(n6602), .B(n6601), .Z(n6482) );
  XNOR U7691 ( .A(n6483), .B(n6482), .Z(n6605) );
  AND U7692 ( .A(\stack[1][17] ), .B(o[23]), .Z(n6607) );
  XNOR U7693 ( .A(n6608), .B(n6607), .Z(n6476) );
  XNOR U7694 ( .A(n6477), .B(n6476), .Z(n6611) );
  AND U7695 ( .A(\stack[1][15] ), .B(o[25]), .Z(n6613) );
  XNOR U7696 ( .A(n6614), .B(n6613), .Z(n6470) );
  XNOR U7697 ( .A(n6471), .B(n6470), .Z(n6617) );
  AND U7698 ( .A(\stack[1][13] ), .B(o[27]), .Z(n6619) );
  XNOR U7699 ( .A(n6620), .B(n6619), .Z(n6465) );
  NAND U7700 ( .A(n6425), .B(n6424), .Z(n6429) );
  NAND U7701 ( .A(n6427), .B(n6426), .Z(n6428) );
  AND U7702 ( .A(n6429), .B(n6428), .Z(n6462) );
  NAND U7703 ( .A(\stack[1][12] ), .B(o[28]), .Z(n6463) );
  NAND U7704 ( .A(n6431), .B(n6430), .Z(n6435) );
  NAND U7705 ( .A(n6433), .B(n6432), .Z(n6434) );
  NAND U7706 ( .A(n6435), .B(n6434), .Z(n6623) );
  XOR U7707 ( .A(n6624), .B(n6623), .Z(n6625) );
  AND U7708 ( .A(\stack[1][11] ), .B(o[29]), .Z(n6626) );
  XOR U7709 ( .A(n6459), .B(n6458), .Z(n6629) );
  NAND U7710 ( .A(n6437), .B(n6436), .Z(n6441) );
  NAND U7711 ( .A(n6439), .B(n6438), .Z(n6440) );
  NAND U7712 ( .A(n6441), .B(n6440), .Z(n6630) );
  AND U7713 ( .A(\stack[1][9] ), .B(o[31]), .Z(n6632) );
  XOR U7714 ( .A(n6453), .B(n6452), .Z(n6635) );
  NAND U7715 ( .A(n6443), .B(n6442), .Z(n6447) );
  NAND U7716 ( .A(n6445), .B(n6444), .Z(n6446) );
  NAND U7717 ( .A(n6447), .B(n6446), .Z(n6636) );
  AND U7718 ( .A(\stack[1][7] ), .B(o[33]), .Z(n6638) );
  NAND U7719 ( .A(n12425), .B(n12424), .Z(n6448) );
  NAND U7720 ( .A(n6449), .B(n6448), .Z(n6641) );
  AND U7721 ( .A(\stack[1][8] ), .B(o[33]), .Z(n6650) );
  NAND U7722 ( .A(n6451), .B(n6450), .Z(n6455) );
  NAND U7723 ( .A(n6453), .B(n6452), .Z(n6454) );
  NAND U7724 ( .A(n6455), .B(n6454), .Z(n6648) );
  NAND U7725 ( .A(n6457), .B(n6456), .Z(n6461) );
  NAND U7726 ( .A(n6459), .B(n6458), .Z(n6460) );
  NAND U7727 ( .A(n6461), .B(n6460), .Z(n6832) );
  NAND U7728 ( .A(n6463), .B(n6462), .Z(n6467) );
  NAND U7729 ( .A(n6465), .B(n6464), .Z(n6466) );
  AND U7730 ( .A(n6467), .B(n6466), .Z(n6660) );
  AND U7731 ( .A(\stack[1][14] ), .B(o[27]), .Z(n6822) );
  NAND U7732 ( .A(n6469), .B(n6468), .Z(n6473) );
  NAND U7733 ( .A(n6471), .B(n6470), .Z(n6472) );
  AND U7734 ( .A(n6473), .B(n6472), .Z(n6820) );
  NAND U7735 ( .A(n6475), .B(n6474), .Z(n6479) );
  NAND U7736 ( .A(n6477), .B(n6476), .Z(n6478) );
  AND U7737 ( .A(n6479), .B(n6478), .Z(n6808) );
  AND U7738 ( .A(\stack[1][18] ), .B(o[23]), .Z(n6798) );
  NAND U7739 ( .A(n6481), .B(n6480), .Z(n6485) );
  NAND U7740 ( .A(n6483), .B(n6482), .Z(n6484) );
  AND U7741 ( .A(n6485), .B(n6484), .Z(n6796) );
  NAND U7742 ( .A(n6486), .B(n16560), .Z(n6490) );
  NAND U7743 ( .A(n6488), .B(n6487), .Z(n6489) );
  NAND U7744 ( .A(n6490), .B(n6489), .Z(n6666) );
  NAND U7745 ( .A(n6492), .B(n6491), .Z(n6496) );
  NAND U7746 ( .A(n6494), .B(n6493), .Z(n6495) );
  NAND U7747 ( .A(n6496), .B(n6495), .Z(n6777) );
  NAND U7748 ( .A(n6498), .B(n6497), .Z(n6502) );
  NAND U7749 ( .A(n6500), .B(n6499), .Z(n6501) );
  NAND U7750 ( .A(n6502), .B(n6501), .Z(n6671) );
  AND U7751 ( .A(o[15]), .B(\stack[1][26] ), .Z(n6685) );
  NAND U7752 ( .A(n6504), .B(n6503), .Z(n6508) );
  NAND U7753 ( .A(n6506), .B(n6505), .Z(n6507) );
  NAND U7754 ( .A(n6508), .B(n6507), .Z(n6683) );
  NAND U7755 ( .A(n6510), .B(n6509), .Z(n6514) );
  NAND U7756 ( .A(n6512), .B(n6511), .Z(n6513) );
  NAND U7757 ( .A(n6514), .B(n6513), .Z(n6760) );
  NAND U7758 ( .A(n6516), .B(n6515), .Z(n6520) );
  NAND U7759 ( .A(n6518), .B(n6517), .Z(n6519) );
  AND U7760 ( .A(n6520), .B(n6519), .Z(n6690) );
  NAND U7761 ( .A(n6522), .B(n6521), .Z(n6526) );
  NAND U7762 ( .A(n6524), .B(n6523), .Z(n6525) );
  NAND U7763 ( .A(n6526), .B(n6525), .Z(n6695) );
  AND U7764 ( .A(o[8]), .B(\stack[1][33] ), .Z(n6702) );
  NAND U7765 ( .A(n6528), .B(n6527), .Z(n6532) );
  NAND U7766 ( .A(n6530), .B(n6529), .Z(n6531) );
  NAND U7767 ( .A(n6532), .B(n6531), .Z(n6701) );
  XOR U7768 ( .A(n6702), .B(n6701), .Z(n6704) );
  AND U7769 ( .A(o[7]), .B(\stack[1][34] ), .Z(n6710) );
  NAND U7770 ( .A(n6534), .B(n6533), .Z(n6538) );
  NAND U7771 ( .A(n6536), .B(n6535), .Z(n6537) );
  NAND U7772 ( .A(n6538), .B(n6537), .Z(n6707) );
  AND U7773 ( .A(o[6]), .B(\stack[1][35] ), .Z(n6744) );
  NAND U7774 ( .A(n6540), .B(n6539), .Z(n6544) );
  NANDN U7775 ( .A(n6542), .B(n6541), .Z(n6543) );
  AND U7776 ( .A(n6544), .B(n6543), .Z(n6714) );
  NAND U7777 ( .A(n6546), .B(n6545), .Z(n6550) );
  NANDN U7778 ( .A(n6548), .B(n6547), .Z(n6549) );
  NAND U7779 ( .A(n6550), .B(n6549), .Z(n6735) );
  AND U7780 ( .A(o[4]), .B(\stack[1][37] ), .Z(n6736) );
  XOR U7781 ( .A(n6735), .B(n6736), .Z(n6738) );
  AND U7782 ( .A(o[3]), .B(\stack[1][38] ), .Z(n6732) );
  AND U7783 ( .A(o[2]), .B(\stack[1][39] ), .Z(n6725) );
  AND U7784 ( .A(o[1]), .B(\stack[1][41] ), .Z(n6721) );
  NAND U7785 ( .A(n6719), .B(n6721), .Z(n6947) );
  XOR U7786 ( .A(n6724), .B(n6947), .Z(n6553) );
  AND U7787 ( .A(o[0]), .B(\stack[1][41] ), .Z(n6952) );
  OR U7788 ( .A(n6551), .B(n6952), .Z(n6552) );
  NAND U7789 ( .A(n6553), .B(n6552), .Z(n6726) );
  XNOR U7790 ( .A(n6725), .B(n6726), .Z(n6730) );
  XOR U7791 ( .A(n6730), .B(n6729), .Z(n6731) );
  XOR U7792 ( .A(n6732), .B(n6731), .Z(n6737) );
  XOR U7793 ( .A(n6738), .B(n6737), .Z(n6713) );
  XOR U7794 ( .A(n6714), .B(n6713), .Z(n6716) );
  AND U7795 ( .A(o[5]), .B(\stack[1][36] ), .Z(n6715) );
  XOR U7796 ( .A(n6716), .B(n6715), .Z(n6742) );
  NAND U7797 ( .A(n6558), .B(n6557), .Z(n6562) );
  NAND U7798 ( .A(n6560), .B(n6559), .Z(n6561) );
  NAND U7799 ( .A(n6562), .B(n6561), .Z(n6741) );
  XOR U7800 ( .A(n6742), .B(n6741), .Z(n6743) );
  XOR U7801 ( .A(n6744), .B(n6743), .Z(n6708) );
  XOR U7802 ( .A(n6707), .B(n6708), .Z(n6709) );
  XOR U7803 ( .A(n6710), .B(n6709), .Z(n6703) );
  XOR U7804 ( .A(n6704), .B(n6703), .Z(n6696) );
  XOR U7805 ( .A(n6695), .B(n6696), .Z(n6698) );
  AND U7806 ( .A(o[9]), .B(\stack[1][32] ), .Z(n6697) );
  XOR U7807 ( .A(n6698), .B(n6697), .Z(n6750) );
  AND U7808 ( .A(o[10]), .B(\stack[1][31] ), .Z(n6748) );
  NAND U7809 ( .A(n6564), .B(n6563), .Z(n6568) );
  NAND U7810 ( .A(n6566), .B(n6565), .Z(n6567) );
  NAND U7811 ( .A(n6568), .B(n6567), .Z(n6747) );
  XOR U7812 ( .A(n6748), .B(n6747), .Z(n6749) );
  XOR U7813 ( .A(n6750), .B(n6749), .Z(n6689) );
  XOR U7814 ( .A(n6690), .B(n6689), .Z(n6692) );
  AND U7815 ( .A(o[11]), .B(\stack[1][30] ), .Z(n6691) );
  XOR U7816 ( .A(n6692), .B(n6691), .Z(n6756) );
  AND U7817 ( .A(o[12]), .B(\stack[1][29] ), .Z(n6754) );
  NAND U7818 ( .A(n6570), .B(n6569), .Z(n6574) );
  NAND U7819 ( .A(n6572), .B(n6571), .Z(n6573) );
  AND U7820 ( .A(n6574), .B(n6573), .Z(n6753) );
  XOR U7821 ( .A(n6754), .B(n6753), .Z(n6755) );
  XNOR U7822 ( .A(n6756), .B(n6755), .Z(n6759) );
  XOR U7823 ( .A(n6760), .B(n6759), .Z(n6762) );
  NAND U7824 ( .A(o[13]), .B(\stack[1][28] ), .Z(n6761) );
  XNOR U7825 ( .A(n6762), .B(n6761), .Z(n6768) );
  AND U7826 ( .A(o[14]), .B(\stack[1][27] ), .Z(n6766) );
  NAND U7827 ( .A(n6576), .B(n6575), .Z(n6580) );
  NAND U7828 ( .A(n6578), .B(n6577), .Z(n6579) );
  NAND U7829 ( .A(n6580), .B(n6579), .Z(n6765) );
  XOR U7830 ( .A(n6766), .B(n6765), .Z(n6767) );
  XOR U7831 ( .A(n6683), .B(n6684), .Z(n6686) );
  XNOR U7832 ( .A(n6685), .B(n6686), .Z(n6680) );
  AND U7833 ( .A(o[16]), .B(\stack[1][25] ), .Z(n6678) );
  NAND U7834 ( .A(n6582), .B(n6581), .Z(n6586) );
  NAND U7835 ( .A(n6584), .B(n6583), .Z(n6585) );
  NAND U7836 ( .A(n6586), .B(n6585), .Z(n6677) );
  XOR U7837 ( .A(n6678), .B(n6677), .Z(n6679) );
  XOR U7838 ( .A(n6680), .B(n6679), .Z(n6672) );
  XOR U7839 ( .A(n6671), .B(n6672), .Z(n6674) );
  AND U7840 ( .A(o[17]), .B(\stack[1][24] ), .Z(n6673) );
  XOR U7841 ( .A(n6674), .B(n6673), .Z(n6774) );
  AND U7842 ( .A(o[18]), .B(\stack[1][23] ), .Z(n6772) );
  NAND U7843 ( .A(n6588), .B(n6587), .Z(n6592) );
  NAND U7844 ( .A(n6590), .B(n6589), .Z(n6591) );
  NAND U7845 ( .A(n6592), .B(n6591), .Z(n6771) );
  XOR U7846 ( .A(n6772), .B(n6771), .Z(n6773) );
  XOR U7847 ( .A(n6774), .B(n6773), .Z(n6778) );
  XOR U7848 ( .A(n6777), .B(n6778), .Z(n6780) );
  AND U7849 ( .A(o[19]), .B(\stack[1][22] ), .Z(n6779) );
  XOR U7850 ( .A(n6780), .B(n6779), .Z(n6786) );
  AND U7851 ( .A(\stack[1][21] ), .B(o[20]), .Z(n6784) );
  NAND U7852 ( .A(n6594), .B(n6593), .Z(n6598) );
  NAND U7853 ( .A(n6596), .B(n6595), .Z(n6597) );
  NAND U7854 ( .A(n6598), .B(n6597), .Z(n6783) );
  XOR U7855 ( .A(n6784), .B(n6783), .Z(n6785) );
  XOR U7856 ( .A(n6786), .B(n6785), .Z(n6665) );
  AND U7857 ( .A(\stack[1][20] ), .B(o[21]), .Z(n6668) );
  AND U7858 ( .A(\stack[1][19] ), .B(o[22]), .Z(n6789) );
  NAND U7859 ( .A(n6600), .B(n6599), .Z(n6604) );
  NAND U7860 ( .A(n6602), .B(n6601), .Z(n6603) );
  NAND U7861 ( .A(n6604), .B(n6603), .Z(n6790) );
  XOR U7862 ( .A(n6792), .B(n6791), .Z(n6795) );
  XOR U7863 ( .A(n6796), .B(n6795), .Z(n6797) );
  XOR U7864 ( .A(n6798), .B(n6797), .Z(n6804) );
  AND U7865 ( .A(\stack[1][17] ), .B(o[24]), .Z(n6801) );
  NAND U7866 ( .A(n6606), .B(n6605), .Z(n6610) );
  NAND U7867 ( .A(n6608), .B(n6607), .Z(n6609) );
  NAND U7868 ( .A(n6610), .B(n6609), .Z(n6802) );
  XOR U7869 ( .A(n6804), .B(n6803), .Z(n6807) );
  XOR U7870 ( .A(n6808), .B(n6807), .Z(n6809) );
  AND U7871 ( .A(\stack[1][16] ), .B(o[25]), .Z(n6810) );
  AND U7872 ( .A(\stack[1][15] ), .B(o[26]), .Z(n6813) );
  NAND U7873 ( .A(n6612), .B(n6611), .Z(n6616) );
  NAND U7874 ( .A(n6614), .B(n6613), .Z(n6615) );
  NAND U7875 ( .A(n6616), .B(n6615), .Z(n6814) );
  XOR U7876 ( .A(n6816), .B(n6815), .Z(n6819) );
  XOR U7877 ( .A(n6820), .B(n6819), .Z(n6821) );
  XOR U7878 ( .A(n6822), .B(n6821), .Z(n6828) );
  AND U7879 ( .A(\stack[1][13] ), .B(o[28]), .Z(n6825) );
  NAND U7880 ( .A(n6618), .B(n6617), .Z(n6622) );
  NAND U7881 ( .A(n6620), .B(n6619), .Z(n6621) );
  NAND U7882 ( .A(n6622), .B(n6621), .Z(n6826) );
  XOR U7883 ( .A(n6828), .B(n6827), .Z(n6659) );
  XOR U7884 ( .A(n6660), .B(n6659), .Z(n6661) );
  AND U7885 ( .A(\stack[1][12] ), .B(o[29]), .Z(n6662) );
  AND U7886 ( .A(\stack[1][11] ), .B(o[30]), .Z(n6653) );
  NAND U7887 ( .A(n6624), .B(n6623), .Z(n6628) );
  NAND U7888 ( .A(n6626), .B(n6625), .Z(n6627) );
  NAND U7889 ( .A(n6628), .B(n6627), .Z(n6654) );
  XOR U7890 ( .A(n6656), .B(n6655), .Z(n6831) );
  AND U7891 ( .A(\stack[1][10] ), .B(o[31]), .Z(n6834) );
  AND U7892 ( .A(\stack[1][9] ), .B(o[32]), .Z(n6837) );
  NAND U7893 ( .A(n6630), .B(n6629), .Z(n6634) );
  NAND U7894 ( .A(n6632), .B(n6631), .Z(n6633) );
  NAND U7895 ( .A(n6634), .B(n6633), .Z(n6838) );
  XOR U7896 ( .A(n6840), .B(n6839), .Z(n6647) );
  XOR U7897 ( .A(n6650), .B(n6649), .Z(n6846) );
  AND U7898 ( .A(\stack[1][7] ), .B(o[34]), .Z(n6843) );
  NAND U7899 ( .A(n6636), .B(n6635), .Z(n6640) );
  NAND U7900 ( .A(n6638), .B(n6637), .Z(n6639) );
  NAND U7901 ( .A(n6640), .B(n6639), .Z(n6844) );
  XOR U7902 ( .A(n6846), .B(n6845), .Z(n6642) );
  NAND U7903 ( .A(n6641), .B(n6642), .Z(n6644) );
  AND U7904 ( .A(\stack[1][6] ), .B(o[35]), .Z(n12431) );
  NAND U7905 ( .A(n12431), .B(n12430), .Z(n6643) );
  NAND U7906 ( .A(n6644), .B(n6643), .Z(n6645) );
  AND U7907 ( .A(\stack[1][6] ), .B(o[36]), .Z(n6646) );
  NAND U7908 ( .A(n6645), .B(n6646), .Z(n6850) );
  NAND U7909 ( .A(n6648), .B(n6647), .Z(n6652) );
  NAND U7910 ( .A(n6650), .B(n6649), .Z(n6651) );
  NAND U7911 ( .A(n6652), .B(n6651), .Z(n6852) );
  AND U7912 ( .A(\stack[1][8] ), .B(o[34]), .Z(n6851) );
  NAND U7913 ( .A(n6654), .B(n6653), .Z(n6658) );
  NAND U7914 ( .A(n6656), .B(n6655), .Z(n6657) );
  NAND U7915 ( .A(n6658), .B(n6657), .Z(n7041) );
  NAND U7916 ( .A(n6660), .B(n6659), .Z(n6664) );
  NAND U7917 ( .A(n6662), .B(n6661), .Z(n6663) );
  AND U7918 ( .A(n6664), .B(n6663), .Z(n6863) );
  NAND U7919 ( .A(\stack[1][12] ), .B(o[30]), .Z(n6864) );
  NAND U7920 ( .A(n6666), .B(n6665), .Z(n6670) );
  NAND U7921 ( .A(n6668), .B(n6667), .Z(n6669) );
  AND U7922 ( .A(n6670), .B(n6669), .Z(n6887) );
  NAND U7923 ( .A(\stack[1][20] ), .B(o[22]), .Z(n6888) );
  AND U7924 ( .A(\stack[1][21] ), .B(o[21]), .Z(n16521) );
  NAND U7925 ( .A(n6672), .B(n6671), .Z(n6676) );
  NAND U7926 ( .A(n6674), .B(n6673), .Z(n6675) );
  AND U7927 ( .A(n6676), .B(n6675), .Z(n6900) );
  NAND U7928 ( .A(o[18]), .B(\stack[1][24] ), .Z(n6899) );
  XOR U7929 ( .A(n6900), .B(n6899), .Z(n6901) );
  NAND U7930 ( .A(n6678), .B(n6677), .Z(n6682) );
  NAND U7931 ( .A(n6680), .B(n6679), .Z(n6681) );
  NAND U7932 ( .A(n6682), .B(n6681), .Z(n7000) );
  NANDN U7933 ( .A(n6684), .B(n6683), .Z(n6688) );
  NANDN U7934 ( .A(n6686), .B(n6685), .Z(n6687) );
  AND U7935 ( .A(n6688), .B(n6687), .Z(n6906) );
  NAND U7936 ( .A(o[16]), .B(\stack[1][26] ), .Z(n6905) );
  XOR U7937 ( .A(n6906), .B(n6905), .Z(n6908) );
  NAND U7938 ( .A(n6690), .B(n6689), .Z(n6694) );
  NAND U7939 ( .A(n6692), .B(n6691), .Z(n6693) );
  NAND U7940 ( .A(n6694), .B(n6693), .Z(n6923) );
  AND U7941 ( .A(o[12]), .B(\stack[1][30] ), .Z(n6924) );
  XOR U7942 ( .A(n6923), .B(n6924), .Z(n6926) );
  NAND U7943 ( .A(n6696), .B(n6695), .Z(n6700) );
  NAND U7944 ( .A(n6698), .B(n6697), .Z(n6699) );
  NAND U7945 ( .A(n6700), .B(n6699), .Z(n6929) );
  AND U7946 ( .A(o[10]), .B(\stack[1][32] ), .Z(n6930) );
  XOR U7947 ( .A(n6929), .B(n6930), .Z(n6932) );
  NAND U7948 ( .A(n6702), .B(n6701), .Z(n6706) );
  NAND U7949 ( .A(n6704), .B(n6703), .Z(n6705) );
  NAND U7950 ( .A(n6706), .B(n6705), .Z(n6982) );
  NAND U7951 ( .A(n6708), .B(n6707), .Z(n6712) );
  NAND U7952 ( .A(n6710), .B(n6709), .Z(n6711) );
  AND U7953 ( .A(n6712), .B(n6711), .Z(n6936) );
  NAND U7954 ( .A(o[8]), .B(\stack[1][34] ), .Z(n6935) );
  XOR U7955 ( .A(n6936), .B(n6935), .Z(n6938) );
  NAND U7956 ( .A(n6714), .B(n6713), .Z(n6718) );
  NAND U7957 ( .A(n6716), .B(n6715), .Z(n6717) );
  NAND U7958 ( .A(n6718), .B(n6717), .Z(n6941) );
  AND U7959 ( .A(o[6]), .B(\stack[1][36] ), .Z(n6942) );
  XOR U7960 ( .A(n6941), .B(n6942), .Z(n6944) );
  AND U7961 ( .A(o[5]), .B(\stack[1][37] ), .Z(n6972) );
  AND U7962 ( .A(o[2]), .B(\stack[1][40] ), .Z(n6948) );
  AND U7963 ( .A(n6719), .B(n6721), .Z(n6720) );
  AND U7964 ( .A(o[1]), .B(\stack[1][42] ), .Z(n6954) );
  NAND U7965 ( .A(n6952), .B(n6954), .Z(n7178) );
  XOR U7966 ( .A(n6720), .B(n7178), .Z(n6723) );
  AND U7967 ( .A(o[0]), .B(\stack[1][42] ), .Z(n7183) );
  OR U7968 ( .A(n6721), .B(n7183), .Z(n6722) );
  NAND U7969 ( .A(n6723), .B(n6722), .Z(n6949) );
  XNOR U7970 ( .A(n6948), .B(n6949), .Z(n6958) );
  NAND U7971 ( .A(n6724), .B(n6947), .Z(n6728) );
  NANDN U7972 ( .A(n6726), .B(n6725), .Z(n6727) );
  NAND U7973 ( .A(n6728), .B(n6727), .Z(n6957) );
  XOR U7974 ( .A(n6958), .B(n6957), .Z(n6960) );
  AND U7975 ( .A(o[3]), .B(\stack[1][39] ), .Z(n6959) );
  XNOR U7976 ( .A(n6960), .B(n6959), .Z(n6964) );
  NAND U7977 ( .A(n6730), .B(n6729), .Z(n6734) );
  NAND U7978 ( .A(n6732), .B(n6731), .Z(n6733) );
  AND U7979 ( .A(n6734), .B(n6733), .Z(n6963) );
  NAND U7980 ( .A(o[4]), .B(\stack[1][38] ), .Z(n6965) );
  XNOR U7981 ( .A(n6966), .B(n6965), .Z(n6970) );
  NAND U7982 ( .A(n6736), .B(n6735), .Z(n6740) );
  NAND U7983 ( .A(n6738), .B(n6737), .Z(n6739) );
  NAND U7984 ( .A(n6740), .B(n6739), .Z(n6969) );
  XOR U7985 ( .A(n6972), .B(n6971), .Z(n6943) );
  XOR U7986 ( .A(n6944), .B(n6943), .Z(n6976) );
  NAND U7987 ( .A(n6742), .B(n6741), .Z(n6746) );
  NAND U7988 ( .A(n6744), .B(n6743), .Z(n6745) );
  NAND U7989 ( .A(n6746), .B(n6745), .Z(n6975) );
  XOR U7990 ( .A(n6976), .B(n6975), .Z(n6978) );
  AND U7991 ( .A(o[7]), .B(\stack[1][35] ), .Z(n6977) );
  XNOR U7992 ( .A(n6978), .B(n6977), .Z(n6937) );
  XNOR U7993 ( .A(n6938), .B(n6937), .Z(n6981) );
  XOR U7994 ( .A(n6982), .B(n6981), .Z(n6984) );
  AND U7995 ( .A(o[9]), .B(\stack[1][33] ), .Z(n6983) );
  XOR U7996 ( .A(n6984), .B(n6983), .Z(n6931) );
  XOR U7997 ( .A(n6932), .B(n6931), .Z(n6988) );
  NAND U7998 ( .A(n6748), .B(n6747), .Z(n6752) );
  NAND U7999 ( .A(n6750), .B(n6749), .Z(n6751) );
  NAND U8000 ( .A(n6752), .B(n6751), .Z(n6987) );
  XOR U8001 ( .A(n6988), .B(n6987), .Z(n6990) );
  AND U8002 ( .A(o[11]), .B(\stack[1][31] ), .Z(n6989) );
  XOR U8003 ( .A(n6990), .B(n6989), .Z(n6925) );
  XOR U8004 ( .A(n6926), .B(n6925), .Z(n6918) );
  NAND U8005 ( .A(n6754), .B(n6753), .Z(n6758) );
  NAND U8006 ( .A(n6756), .B(n6755), .Z(n6757) );
  NAND U8007 ( .A(n6758), .B(n6757), .Z(n6917) );
  XOR U8008 ( .A(n6918), .B(n6917), .Z(n6920) );
  AND U8009 ( .A(o[13]), .B(\stack[1][29] ), .Z(n6919) );
  XOR U8010 ( .A(n6920), .B(n6919), .Z(n6914) );
  NAND U8011 ( .A(n6760), .B(n6759), .Z(n6764) );
  NAND U8012 ( .A(n6762), .B(n6761), .Z(n6763) );
  AND U8013 ( .A(n6764), .B(n6763), .Z(n6912) );
  AND U8014 ( .A(o[14]), .B(\stack[1][28] ), .Z(n6911) );
  XOR U8015 ( .A(n6912), .B(n6911), .Z(n6913) );
  XOR U8016 ( .A(n6914), .B(n6913), .Z(n6994) );
  NAND U8017 ( .A(n6766), .B(n6765), .Z(n6770) );
  NAND U8018 ( .A(n6768), .B(n6767), .Z(n6769) );
  NAND U8019 ( .A(n6770), .B(n6769), .Z(n6993) );
  XOR U8020 ( .A(n6994), .B(n6993), .Z(n6996) );
  AND U8021 ( .A(o[15]), .B(\stack[1][27] ), .Z(n6995) );
  XNOR U8022 ( .A(n6996), .B(n6995), .Z(n6907) );
  XNOR U8023 ( .A(n6908), .B(n6907), .Z(n6999) );
  XOR U8024 ( .A(n7000), .B(n6999), .Z(n7002) );
  AND U8025 ( .A(o[17]), .B(\stack[1][25] ), .Z(n7001) );
  XNOR U8026 ( .A(n7002), .B(n7001), .Z(n6902) );
  NAND U8027 ( .A(n6772), .B(n6771), .Z(n6776) );
  NAND U8028 ( .A(n6774), .B(n6773), .Z(n6775) );
  NAND U8029 ( .A(n6776), .B(n6775), .Z(n7005) );
  AND U8030 ( .A(o[19]), .B(\stack[1][23] ), .Z(n7007) );
  XNOR U8031 ( .A(n7008), .B(n7007), .Z(n6896) );
  NAND U8032 ( .A(n6778), .B(n6777), .Z(n6782) );
  NAND U8033 ( .A(n6780), .B(n6779), .Z(n6781) );
  AND U8034 ( .A(n6782), .B(n6781), .Z(n6894) );
  NAND U8035 ( .A(o[20]), .B(\stack[1][22] ), .Z(n6893) );
  XOR U8036 ( .A(n6894), .B(n6893), .Z(n6895) );
  NAND U8037 ( .A(n6784), .B(n6783), .Z(n6788) );
  NAND U8038 ( .A(n6786), .B(n6785), .Z(n6787) );
  NAND U8039 ( .A(n6788), .B(n6787), .Z(n7011) );
  XNOR U8040 ( .A(n16521), .B(n7013), .Z(n6889) );
  XNOR U8041 ( .A(n6890), .B(n6889), .Z(n7017) );
  NAND U8042 ( .A(n6790), .B(n6789), .Z(n6794) );
  NAND U8043 ( .A(n6792), .B(n6791), .Z(n6793) );
  NAND U8044 ( .A(n6794), .B(n6793), .Z(n7016) );
  AND U8045 ( .A(\stack[1][19] ), .B(o[23]), .Z(n7019) );
  NAND U8046 ( .A(n6796), .B(n6795), .Z(n6800) );
  NAND U8047 ( .A(n6798), .B(n6797), .Z(n6799) );
  NAND U8048 ( .A(n6800), .B(n6799), .Z(n6882) );
  AND U8049 ( .A(\stack[1][18] ), .B(o[24]), .Z(n6881) );
  XOR U8050 ( .A(n6884), .B(n6883), .Z(n7022) );
  NAND U8051 ( .A(n6802), .B(n6801), .Z(n6806) );
  NAND U8052 ( .A(n6804), .B(n6803), .Z(n6805) );
  NAND U8053 ( .A(n6806), .B(n6805), .Z(n7023) );
  AND U8054 ( .A(\stack[1][17] ), .B(o[25]), .Z(n7025) );
  NAND U8055 ( .A(n6808), .B(n6807), .Z(n6812) );
  NAND U8056 ( .A(n6810), .B(n6809), .Z(n6811) );
  NAND U8057 ( .A(n6812), .B(n6811), .Z(n6876) );
  AND U8058 ( .A(\stack[1][16] ), .B(o[26]), .Z(n6875) );
  XOR U8059 ( .A(n6878), .B(n6877), .Z(n7028) );
  NAND U8060 ( .A(n6814), .B(n6813), .Z(n6818) );
  NAND U8061 ( .A(n6816), .B(n6815), .Z(n6817) );
  NAND U8062 ( .A(n6818), .B(n6817), .Z(n7029) );
  AND U8063 ( .A(\stack[1][15] ), .B(o[27]), .Z(n7031) );
  NAND U8064 ( .A(n6820), .B(n6819), .Z(n6824) );
  NAND U8065 ( .A(n6822), .B(n6821), .Z(n6823) );
  NAND U8066 ( .A(n6824), .B(n6823), .Z(n6870) );
  AND U8067 ( .A(\stack[1][14] ), .B(o[28]), .Z(n6869) );
  XOR U8068 ( .A(n6872), .B(n6871), .Z(n7034) );
  NAND U8069 ( .A(n6826), .B(n6825), .Z(n6830) );
  NAND U8070 ( .A(n6828), .B(n6827), .Z(n6829) );
  NAND U8071 ( .A(n6830), .B(n6829), .Z(n7035) );
  AND U8072 ( .A(\stack[1][13] ), .B(o[29]), .Z(n7036) );
  XNOR U8073 ( .A(n7037), .B(n7036), .Z(n6865) );
  XNOR U8074 ( .A(n6866), .B(n6865), .Z(n7040) );
  AND U8075 ( .A(\stack[1][11] ), .B(o[31]), .Z(n7042) );
  XNOR U8076 ( .A(n7043), .B(n7042), .Z(n6860) );
  NAND U8077 ( .A(n6832), .B(n6831), .Z(n6836) );
  NAND U8078 ( .A(n6834), .B(n6833), .Z(n6835) );
  AND U8079 ( .A(n6836), .B(n6835), .Z(n6857) );
  NAND U8080 ( .A(\stack[1][10] ), .B(o[32]), .Z(n6858) );
  NAND U8081 ( .A(n6838), .B(n6837), .Z(n6842) );
  NAND U8082 ( .A(n6840), .B(n6839), .Z(n6841) );
  NAND U8083 ( .A(n6842), .B(n6841), .Z(n7046) );
  XOR U8084 ( .A(n7047), .B(n7046), .Z(n7048) );
  AND U8085 ( .A(\stack[1][9] ), .B(o[33]), .Z(n7049) );
  XOR U8086 ( .A(n6854), .B(n6853), .Z(n7052) );
  NAND U8087 ( .A(n6844), .B(n6843), .Z(n6848) );
  NAND U8088 ( .A(n6846), .B(n6845), .Z(n6847) );
  NAND U8089 ( .A(n6848), .B(n6847), .Z(n7053) );
  AND U8090 ( .A(\stack[1][7] ), .B(o[35]), .Z(n7055) );
  NAND U8091 ( .A(n12437), .B(n12436), .Z(n6849) );
  NAND U8092 ( .A(n6850), .B(n6849), .Z(n7058) );
  AND U8093 ( .A(\stack[1][8] ), .B(o[35]), .Z(n7067) );
  NAND U8094 ( .A(n6852), .B(n6851), .Z(n6856) );
  NAND U8095 ( .A(n6854), .B(n6853), .Z(n6855) );
  NAND U8096 ( .A(n6856), .B(n6855), .Z(n7065) );
  NAND U8097 ( .A(n6858), .B(n6857), .Z(n6862) );
  NAND U8098 ( .A(n6860), .B(n6859), .Z(n6861) );
  AND U8099 ( .A(n6862), .B(n6861), .Z(n7071) );
  AND U8100 ( .A(\stack[1][12] ), .B(o[31]), .Z(n7079) );
  NAND U8101 ( .A(n6864), .B(n6863), .Z(n6868) );
  NAND U8102 ( .A(n6866), .B(n6865), .Z(n6867) );
  AND U8103 ( .A(n6868), .B(n6867), .Z(n7077) );
  AND U8104 ( .A(\stack[1][14] ), .B(o[29]), .Z(n7085) );
  NAND U8105 ( .A(n6870), .B(n6869), .Z(n6874) );
  NAND U8106 ( .A(n6872), .B(n6871), .Z(n6873) );
  NAND U8107 ( .A(n6874), .B(n6873), .Z(n7083) );
  AND U8108 ( .A(\stack[1][16] ), .B(o[27]), .Z(n7091) );
  NAND U8109 ( .A(n6876), .B(n6875), .Z(n6880) );
  NAND U8110 ( .A(n6878), .B(n6877), .Z(n6879) );
  NAND U8111 ( .A(n6880), .B(n6879), .Z(n7089) );
  NAND U8112 ( .A(n6882), .B(n6881), .Z(n6886) );
  NAND U8113 ( .A(n6884), .B(n6883), .Z(n6885) );
  NAND U8114 ( .A(n6886), .B(n6885), .Z(n7237) );
  NAND U8115 ( .A(n6888), .B(n6887), .Z(n6892) );
  NAND U8116 ( .A(n6890), .B(n6889), .Z(n6891) );
  AND U8117 ( .A(n6892), .B(n6891), .Z(n7101) );
  NAND U8118 ( .A(n6894), .B(n6893), .Z(n6898) );
  NAND U8119 ( .A(n6896), .B(n6895), .Z(n6897) );
  AND U8120 ( .A(n6898), .B(n6897), .Z(n7113) );
  NAND U8121 ( .A(n6900), .B(n6899), .Z(n6904) );
  NAND U8122 ( .A(n6902), .B(n6901), .Z(n6903) );
  AND U8123 ( .A(n6904), .B(n6903), .Z(n7119) );
  NAND U8124 ( .A(n6906), .B(n6905), .Z(n6910) );
  NAND U8125 ( .A(n6908), .B(n6907), .Z(n6909) );
  AND U8126 ( .A(n6910), .B(n6909), .Z(n7125) );
  AND U8127 ( .A(o[15]), .B(\stack[1][28] ), .Z(n7132) );
  NAND U8128 ( .A(n6912), .B(n6911), .Z(n6916) );
  NAND U8129 ( .A(n6914), .B(n6913), .Z(n6915) );
  NAND U8130 ( .A(n6916), .B(n6915), .Z(n7130) );
  AND U8131 ( .A(o[14]), .B(\stack[1][29] ), .Z(n7137) );
  NAND U8132 ( .A(n6918), .B(n6917), .Z(n6922) );
  NAND U8133 ( .A(n6920), .B(n6919), .Z(n6921) );
  NAND U8134 ( .A(n6922), .B(n6921), .Z(n7136) );
  XOR U8135 ( .A(n7137), .B(n7136), .Z(n7139) );
  NAND U8136 ( .A(n6924), .B(n6923), .Z(n6928) );
  NAND U8137 ( .A(n6926), .B(n6925), .Z(n6927) );
  NAND U8138 ( .A(n6928), .B(n6927), .Z(n7212) );
  NAND U8139 ( .A(n6930), .B(n6929), .Z(n6934) );
  NAND U8140 ( .A(n6932), .B(n6931), .Z(n6933) );
  NAND U8141 ( .A(n6934), .B(n6933), .Z(n7148) );
  NAND U8142 ( .A(n6936), .B(n6935), .Z(n6940) );
  NAND U8143 ( .A(n6938), .B(n6937), .Z(n6939) );
  NAND U8144 ( .A(n6940), .B(n6939), .Z(n7155) );
  NAND U8145 ( .A(n6942), .B(n6941), .Z(n6946) );
  NAND U8146 ( .A(n6944), .B(n6943), .Z(n6945) );
  AND U8147 ( .A(n6946), .B(n6945), .Z(n7200) );
  NAND U8148 ( .A(o[5]), .B(\stack[1][38] ), .Z(n7196) );
  AND U8149 ( .A(o[4]), .B(\stack[1][39] ), .Z(n7175) );
  AND U8150 ( .A(o[3]), .B(\stack[1][40] ), .Z(n7190) );
  NANDN U8151 ( .A(n6947), .B(n7178), .Z(n6951) );
  NANDN U8152 ( .A(n6949), .B(n6948), .Z(n6950) );
  NAND U8153 ( .A(n6951), .B(n6950), .Z(n7188) );
  AND U8154 ( .A(o[2]), .B(\stack[1][41] ), .Z(n7179) );
  AND U8155 ( .A(n6952), .B(n6954), .Z(n6953) );
  AND U8156 ( .A(o[1]), .B(\stack[1][43] ), .Z(n7185) );
  NAND U8157 ( .A(n7183), .B(n7185), .Z(n7370) );
  XOR U8158 ( .A(n6953), .B(n7370), .Z(n6956) );
  AND U8159 ( .A(o[0]), .B(\stack[1][43] ), .Z(n7375) );
  OR U8160 ( .A(n6954), .B(n7375), .Z(n6955) );
  NAND U8161 ( .A(n6956), .B(n6955), .Z(n7180) );
  XNOR U8162 ( .A(n7179), .B(n7180), .Z(n7189) );
  XNOR U8163 ( .A(n7190), .B(n7191), .Z(n7173) );
  NAND U8164 ( .A(n6958), .B(n6957), .Z(n6962) );
  NAND U8165 ( .A(n6960), .B(n6959), .Z(n6961) );
  NAND U8166 ( .A(n6962), .B(n6961), .Z(n7172) );
  XOR U8167 ( .A(n7173), .B(n7172), .Z(n7174) );
  XNOR U8168 ( .A(n7175), .B(n7174), .Z(n7195) );
  NAND U8169 ( .A(n6964), .B(n6963), .Z(n6968) );
  NAND U8170 ( .A(n6966), .B(n6965), .Z(n6967) );
  NAND U8171 ( .A(n6968), .B(n6967), .Z(n7194) );
  XNOR U8172 ( .A(n7196), .B(n7197), .Z(n7169) );
  AND U8173 ( .A(o[6]), .B(\stack[1][37] ), .Z(n7167) );
  NAND U8174 ( .A(n6970), .B(n6969), .Z(n6974) );
  NAND U8175 ( .A(n6972), .B(n6971), .Z(n6973) );
  NAND U8176 ( .A(n6974), .B(n6973), .Z(n7166) );
  XOR U8177 ( .A(n7167), .B(n7166), .Z(n7168) );
  NAND U8178 ( .A(o[7]), .B(\stack[1][36] ), .Z(n7202) );
  XNOR U8179 ( .A(n7203), .B(n7202), .Z(n7162) );
  NAND U8180 ( .A(n6976), .B(n6975), .Z(n6980) );
  NAND U8181 ( .A(n6978), .B(n6977), .Z(n6979) );
  NAND U8182 ( .A(n6980), .B(n6979), .Z(n7160) );
  AND U8183 ( .A(o[8]), .B(\stack[1][35] ), .Z(n7161) );
  XNOR U8184 ( .A(n7160), .B(n7161), .Z(n7163) );
  XOR U8185 ( .A(n7162), .B(n7163), .Z(n7154) );
  XOR U8186 ( .A(n7155), .B(n7154), .Z(n7157) );
  NAND U8187 ( .A(o[9]), .B(\stack[1][34] ), .Z(n7156) );
  XNOR U8188 ( .A(n7157), .B(n7156), .Z(n7209) );
  AND U8189 ( .A(o[10]), .B(\stack[1][33] ), .Z(n7207) );
  NAND U8190 ( .A(n6982), .B(n6981), .Z(n6986) );
  NAND U8191 ( .A(n6984), .B(n6983), .Z(n6985) );
  NAND U8192 ( .A(n6986), .B(n6985), .Z(n7206) );
  XOR U8193 ( .A(n7207), .B(n7206), .Z(n7208) );
  XOR U8194 ( .A(n7148), .B(n7149), .Z(n7151) );
  AND U8195 ( .A(o[11]), .B(\stack[1][32] ), .Z(n7150) );
  XOR U8196 ( .A(n7151), .B(n7150), .Z(n7145) );
  AND U8197 ( .A(o[12]), .B(\stack[1][31] ), .Z(n7143) );
  NAND U8198 ( .A(n6988), .B(n6987), .Z(n6992) );
  NAND U8199 ( .A(n6990), .B(n6989), .Z(n6991) );
  NAND U8200 ( .A(n6992), .B(n6991), .Z(n7142) );
  XOR U8201 ( .A(n7143), .B(n7142), .Z(n7144) );
  XOR U8202 ( .A(n7145), .B(n7144), .Z(n7213) );
  XOR U8203 ( .A(n7212), .B(n7213), .Z(n7215) );
  AND U8204 ( .A(o[13]), .B(\stack[1][30] ), .Z(n7214) );
  XOR U8205 ( .A(n7215), .B(n7214), .Z(n7138) );
  XOR U8206 ( .A(n7139), .B(n7138), .Z(n7131) );
  XOR U8207 ( .A(n7130), .B(n7131), .Z(n7133) );
  AND U8208 ( .A(o[16]), .B(\stack[1][27] ), .Z(n7219) );
  NAND U8209 ( .A(n6994), .B(n6993), .Z(n6998) );
  NAND U8210 ( .A(n6996), .B(n6995), .Z(n6997) );
  NAND U8211 ( .A(n6998), .B(n6997), .Z(n7218) );
  XOR U8212 ( .A(n7219), .B(n7218), .Z(n7220) );
  XOR U8213 ( .A(n7221), .B(n7220), .Z(n7124) );
  XOR U8214 ( .A(n7125), .B(n7124), .Z(n7127) );
  AND U8215 ( .A(o[17]), .B(\stack[1][26] ), .Z(n7126) );
  XOR U8216 ( .A(n7127), .B(n7126), .Z(n7227) );
  AND U8217 ( .A(o[18]), .B(\stack[1][25] ), .Z(n7225) );
  NAND U8218 ( .A(n7000), .B(n6999), .Z(n7004) );
  NAND U8219 ( .A(n7002), .B(n7001), .Z(n7003) );
  NAND U8220 ( .A(n7004), .B(n7003), .Z(n7224) );
  XOR U8221 ( .A(n7225), .B(n7224), .Z(n7226) );
  XOR U8222 ( .A(n7227), .B(n7226), .Z(n7118) );
  XOR U8223 ( .A(n7119), .B(n7118), .Z(n7121) );
  AND U8224 ( .A(o[19]), .B(\stack[1][24] ), .Z(n7120) );
  XOR U8225 ( .A(n7121), .B(n7120), .Z(n7233) );
  AND U8226 ( .A(o[20]), .B(\stack[1][23] ), .Z(n7231) );
  NAND U8227 ( .A(n7006), .B(n7005), .Z(n7010) );
  NAND U8228 ( .A(n7008), .B(n7007), .Z(n7009) );
  NAND U8229 ( .A(n7010), .B(n7009), .Z(n7230) );
  XOR U8230 ( .A(n7231), .B(n7230), .Z(n7232) );
  XOR U8231 ( .A(n7233), .B(n7232), .Z(n7112) );
  XOR U8232 ( .A(n7113), .B(n7112), .Z(n7115) );
  AND U8233 ( .A(\stack[1][22] ), .B(o[21]), .Z(n7114) );
  XOR U8234 ( .A(n7115), .B(n7114), .Z(n7109) );
  AND U8235 ( .A(\stack[1][21] ), .B(o[22]), .Z(n7107) );
  NAND U8236 ( .A(n7012), .B(n7011), .Z(n7015) );
  NAND U8237 ( .A(n16521), .B(n7013), .Z(n7014) );
  NAND U8238 ( .A(n7015), .B(n7014), .Z(n7106) );
  XOR U8239 ( .A(n7107), .B(n7106), .Z(n7108) );
  XOR U8240 ( .A(n7109), .B(n7108), .Z(n7100) );
  XOR U8241 ( .A(n7101), .B(n7100), .Z(n7102) );
  AND U8242 ( .A(\stack[1][20] ), .B(o[23]), .Z(n7103) );
  AND U8243 ( .A(\stack[1][19] ), .B(o[24]), .Z(n7094) );
  NAND U8244 ( .A(n7017), .B(n7016), .Z(n7021) );
  NAND U8245 ( .A(n7019), .B(n7018), .Z(n7020) );
  NAND U8246 ( .A(n7021), .B(n7020), .Z(n7095) );
  XOR U8247 ( .A(n7097), .B(n7096), .Z(n7236) );
  AND U8248 ( .A(\stack[1][18] ), .B(o[25]), .Z(n7239) );
  AND U8249 ( .A(\stack[1][17] ), .B(o[26]), .Z(n7242) );
  NAND U8250 ( .A(n7023), .B(n7022), .Z(n7027) );
  NAND U8251 ( .A(n7025), .B(n7024), .Z(n7026) );
  NAND U8252 ( .A(n7027), .B(n7026), .Z(n7243) );
  XOR U8253 ( .A(n7245), .B(n7244), .Z(n7088) );
  XOR U8254 ( .A(n7091), .B(n7090), .Z(n7251) );
  AND U8255 ( .A(\stack[1][15] ), .B(o[28]), .Z(n7248) );
  NAND U8256 ( .A(n7029), .B(n7028), .Z(n7033) );
  NAND U8257 ( .A(n7031), .B(n7030), .Z(n7032) );
  NAND U8258 ( .A(n7033), .B(n7032), .Z(n7249) );
  XOR U8259 ( .A(n7251), .B(n7250), .Z(n7082) );
  XOR U8260 ( .A(n7085), .B(n7084), .Z(n7257) );
  AND U8261 ( .A(\stack[1][13] ), .B(o[30]), .Z(n7254) );
  NAND U8262 ( .A(n7035), .B(n7034), .Z(n7039) );
  NAND U8263 ( .A(n7037), .B(n7036), .Z(n7038) );
  NAND U8264 ( .A(n7039), .B(n7038), .Z(n7255) );
  XOR U8265 ( .A(n7257), .B(n7256), .Z(n7076) );
  XOR U8266 ( .A(n7077), .B(n7076), .Z(n7078) );
  XOR U8267 ( .A(n7079), .B(n7078), .Z(n7263) );
  AND U8268 ( .A(\stack[1][11] ), .B(o[32]), .Z(n7260) );
  NAND U8269 ( .A(n7041), .B(n7040), .Z(n7045) );
  NAND U8270 ( .A(n7043), .B(n7042), .Z(n7044) );
  NAND U8271 ( .A(n7045), .B(n7044), .Z(n7261) );
  XOR U8272 ( .A(n7263), .B(n7262), .Z(n7070) );
  XOR U8273 ( .A(n7071), .B(n7070), .Z(n7072) );
  AND U8274 ( .A(\stack[1][10] ), .B(o[33]), .Z(n7073) );
  AND U8275 ( .A(\stack[1][9] ), .B(o[34]), .Z(n7266) );
  NAND U8276 ( .A(n7047), .B(n7046), .Z(n7051) );
  NAND U8277 ( .A(n7049), .B(n7048), .Z(n7050) );
  NAND U8278 ( .A(n7051), .B(n7050), .Z(n7267) );
  XOR U8279 ( .A(n7269), .B(n7268), .Z(n7064) );
  XOR U8280 ( .A(n7067), .B(n7066), .Z(n7275) );
  AND U8281 ( .A(\stack[1][7] ), .B(o[36]), .Z(n7272) );
  NAND U8282 ( .A(n7053), .B(n7052), .Z(n7057) );
  NAND U8283 ( .A(n7055), .B(n7054), .Z(n7056) );
  NAND U8284 ( .A(n7057), .B(n7056), .Z(n7273) );
  XOR U8285 ( .A(n7275), .B(n7274), .Z(n7059) );
  NAND U8286 ( .A(n7058), .B(n7059), .Z(n7061) );
  AND U8287 ( .A(\stack[1][6] ), .B(o[37]), .Z(n12443) );
  NAND U8288 ( .A(n12443), .B(n12442), .Z(n7060) );
  AND U8289 ( .A(n7061), .B(n7060), .Z(n7063) );
  NAND U8290 ( .A(n7062), .B(n7063), .Z(n7279) );
  NAND U8291 ( .A(n7065), .B(n7064), .Z(n7069) );
  NAND U8292 ( .A(n7067), .B(n7066), .Z(n7068) );
  NAND U8293 ( .A(n7069), .B(n7068), .Z(n7281) );
  AND U8294 ( .A(\stack[1][8] ), .B(o[36]), .Z(n7280) );
  NAND U8295 ( .A(n7071), .B(n7070), .Z(n7075) );
  NAND U8296 ( .A(n7073), .B(n7072), .Z(n7074) );
  NAND U8297 ( .A(n7075), .B(n7074), .Z(n7287) );
  AND U8298 ( .A(\stack[1][10] ), .B(o[34]), .Z(n7286) );
  NAND U8299 ( .A(n7077), .B(n7076), .Z(n7081) );
  NAND U8300 ( .A(n7079), .B(n7078), .Z(n7080) );
  NAND U8301 ( .A(n7081), .B(n7080), .Z(n7293) );
  AND U8302 ( .A(\stack[1][12] ), .B(o[32]), .Z(n7292) );
  NAND U8303 ( .A(n7083), .B(n7082), .Z(n7087) );
  NAND U8304 ( .A(n7085), .B(n7084), .Z(n7086) );
  NAND U8305 ( .A(n7087), .B(n7086), .Z(n7299) );
  AND U8306 ( .A(\stack[1][14] ), .B(o[30]), .Z(n7298) );
  NAND U8307 ( .A(n7089), .B(n7088), .Z(n7093) );
  NAND U8308 ( .A(n7091), .B(n7090), .Z(n7092) );
  NAND U8309 ( .A(n7093), .B(n7092), .Z(n7305) );
  AND U8310 ( .A(\stack[1][16] ), .B(o[28]), .Z(n7304) );
  NAND U8311 ( .A(n7095), .B(n7094), .Z(n7099) );
  NAND U8312 ( .A(n7097), .B(n7096), .Z(n7098) );
  NAND U8313 ( .A(n7099), .B(n7098), .Z(n7459) );
  NAND U8314 ( .A(n7101), .B(n7100), .Z(n7105) );
  NAND U8315 ( .A(n7103), .B(n7102), .Z(n7104) );
  AND U8316 ( .A(n7105), .B(n7104), .Z(n7316) );
  NAND U8317 ( .A(\stack[1][20] ), .B(o[24]), .Z(n7317) );
  NAND U8318 ( .A(n7107), .B(n7106), .Z(n7111) );
  NAND U8319 ( .A(n7109), .B(n7108), .Z(n7110) );
  NAND U8320 ( .A(n7111), .B(n7110), .Z(n7453) );
  NAND U8321 ( .A(n7113), .B(n7112), .Z(n7117) );
  NAND U8322 ( .A(n7115), .B(n7114), .Z(n7116) );
  AND U8323 ( .A(n7117), .B(n7116), .Z(n7323) );
  NAND U8324 ( .A(\stack[1][22] ), .B(o[22]), .Z(n7322) );
  XOR U8325 ( .A(n7323), .B(n7322), .Z(n7325) );
  NAND U8326 ( .A(n7119), .B(n7118), .Z(n7123) );
  NAND U8327 ( .A(n7121), .B(n7120), .Z(n7122) );
  NAND U8328 ( .A(n7123), .B(n7122), .Z(n7328) );
  AND U8329 ( .A(o[20]), .B(\stack[1][24] ), .Z(n7329) );
  XOR U8330 ( .A(n7328), .B(n7329), .Z(n7331) );
  NAND U8331 ( .A(n7125), .B(n7124), .Z(n7129) );
  NAND U8332 ( .A(n7127), .B(n7126), .Z(n7128) );
  NAND U8333 ( .A(n7129), .B(n7128), .Z(n7334) );
  AND U8334 ( .A(o[18]), .B(\stack[1][26] ), .Z(n7335) );
  XOR U8335 ( .A(n7334), .B(n7335), .Z(n7337) );
  NAND U8336 ( .A(n7131), .B(n7130), .Z(n7135) );
  NAND U8337 ( .A(n7133), .B(n7132), .Z(n7134) );
  NAND U8338 ( .A(n7135), .B(n7134), .Z(n7340) );
  AND U8339 ( .A(o[16]), .B(\stack[1][28] ), .Z(n7341) );
  XOR U8340 ( .A(n7340), .B(n7341), .Z(n7343) );
  NAND U8341 ( .A(n7137), .B(n7136), .Z(n7141) );
  NAND U8342 ( .A(n7139), .B(n7138), .Z(n7140) );
  NAND U8343 ( .A(n7141), .B(n7140), .Z(n7429) );
  NAND U8344 ( .A(n7143), .B(n7142), .Z(n7147) );
  NAND U8345 ( .A(n7145), .B(n7144), .Z(n7146) );
  NAND U8346 ( .A(n7147), .B(n7146), .Z(n7423) );
  NAND U8347 ( .A(n7149), .B(n7148), .Z(n7153) );
  NAND U8348 ( .A(n7151), .B(n7150), .Z(n7152) );
  AND U8349 ( .A(n7153), .B(n7152), .Z(n7353) );
  NAND U8350 ( .A(o[12]), .B(\stack[1][32] ), .Z(n7352) );
  XOR U8351 ( .A(n7353), .B(n7352), .Z(n7355) );
  AND U8352 ( .A(o[10]), .B(\stack[1][34] ), .Z(n7359) );
  NAND U8353 ( .A(n7155), .B(n7154), .Z(n7159) );
  NAND U8354 ( .A(n7157), .B(n7156), .Z(n7158) );
  AND U8355 ( .A(n7159), .B(n7158), .Z(n7358) );
  XOR U8356 ( .A(n7359), .B(n7358), .Z(n7361) );
  AND U8357 ( .A(o[9]), .B(\stack[1][35] ), .Z(n7413) );
  NAND U8358 ( .A(n7161), .B(n7160), .Z(n7165) );
  NANDN U8359 ( .A(n7163), .B(n7162), .Z(n7164) );
  NAND U8360 ( .A(n7165), .B(n7164), .Z(n7410) );
  AND U8361 ( .A(o[8]), .B(\stack[1][36] ), .Z(n7367) );
  NAND U8362 ( .A(n7167), .B(n7166), .Z(n7171) );
  NAND U8363 ( .A(n7169), .B(n7168), .Z(n7170) );
  NAND U8364 ( .A(n7171), .B(n7170), .Z(n7405) );
  NAND U8365 ( .A(o[6]), .B(\stack[1][38] ), .Z(n7400) );
  NAND U8366 ( .A(n7173), .B(n7172), .Z(n7177) );
  NAND U8367 ( .A(n7175), .B(n7174), .Z(n7176) );
  NAND U8368 ( .A(n7177), .B(n7176), .Z(n7393) );
  NANDN U8369 ( .A(n7178), .B(n7370), .Z(n7182) );
  NANDN U8370 ( .A(n7180), .B(n7179), .Z(n7181) );
  NAND U8371 ( .A(n7182), .B(n7181), .Z(n7380) );
  AND U8372 ( .A(o[3]), .B(\stack[1][41] ), .Z(n7381) );
  XOR U8373 ( .A(n7380), .B(n7381), .Z(n7382) );
  AND U8374 ( .A(o[2]), .B(\stack[1][42] ), .Z(n7371) );
  AND U8375 ( .A(n7183), .B(n7185), .Z(n7184) );
  AND U8376 ( .A(o[1]), .B(\stack[1][44] ), .Z(n7377) );
  NAND U8377 ( .A(n7375), .B(n7377), .Z(n7625) );
  XOR U8378 ( .A(n7184), .B(n7625), .Z(n7187) );
  AND U8379 ( .A(o[0]), .B(\stack[1][44] ), .Z(n7620) );
  OR U8380 ( .A(n7185), .B(n7620), .Z(n7186) );
  NAND U8381 ( .A(n7187), .B(n7186), .Z(n7372) );
  XNOR U8382 ( .A(n7371), .B(n7372), .Z(n7383) );
  NAND U8383 ( .A(n7189), .B(n7188), .Z(n7193) );
  NANDN U8384 ( .A(n7191), .B(n7190), .Z(n7192) );
  AND U8385 ( .A(n7193), .B(n7192), .Z(n7386) );
  NAND U8386 ( .A(o[4]), .B(\stack[1][40] ), .Z(n7388) );
  XNOR U8387 ( .A(n7389), .B(n7388), .Z(n7392) );
  XOR U8388 ( .A(n7393), .B(n7392), .Z(n7395) );
  AND U8389 ( .A(o[5]), .B(\stack[1][39] ), .Z(n7394) );
  XNOR U8390 ( .A(n7395), .B(n7394), .Z(n7399) );
  NAND U8391 ( .A(n7195), .B(n7194), .Z(n7199) );
  NAND U8392 ( .A(n7197), .B(n7196), .Z(n7198) );
  NAND U8393 ( .A(n7199), .B(n7198), .Z(n7398) );
  XOR U8394 ( .A(n7400), .B(n7401), .Z(n7404) );
  XOR U8395 ( .A(n7405), .B(n7404), .Z(n7407) );
  AND U8396 ( .A(o[7]), .B(\stack[1][37] ), .Z(n7406) );
  XOR U8397 ( .A(n7407), .B(n7406), .Z(n7365) );
  NAND U8398 ( .A(n7201), .B(n7200), .Z(n7205) );
  NAND U8399 ( .A(n7203), .B(n7202), .Z(n7204) );
  AND U8400 ( .A(n7205), .B(n7204), .Z(n7364) );
  XOR U8401 ( .A(n7365), .B(n7364), .Z(n7366) );
  XOR U8402 ( .A(n7367), .B(n7366), .Z(n7411) );
  XOR U8403 ( .A(n7410), .B(n7411), .Z(n7412) );
  XOR U8404 ( .A(n7413), .B(n7412), .Z(n7360) );
  XOR U8405 ( .A(n7361), .B(n7360), .Z(n7417) );
  NAND U8406 ( .A(n7207), .B(n7206), .Z(n7211) );
  NAND U8407 ( .A(n7209), .B(n7208), .Z(n7210) );
  NAND U8408 ( .A(n7211), .B(n7210), .Z(n7416) );
  XOR U8409 ( .A(n7417), .B(n7416), .Z(n7419) );
  AND U8410 ( .A(o[11]), .B(\stack[1][33] ), .Z(n7418) );
  XNOR U8411 ( .A(n7419), .B(n7418), .Z(n7354) );
  XNOR U8412 ( .A(n7355), .B(n7354), .Z(n7422) );
  XOR U8413 ( .A(n7423), .B(n7422), .Z(n7425) );
  AND U8414 ( .A(o[13]), .B(\stack[1][31] ), .Z(n7424) );
  XOR U8415 ( .A(n7425), .B(n7424), .Z(n7349) );
  NAND U8416 ( .A(n7213), .B(n7212), .Z(n7217) );
  NAND U8417 ( .A(n7215), .B(n7214), .Z(n7216) );
  AND U8418 ( .A(n7217), .B(n7216), .Z(n7347) );
  NAND U8419 ( .A(o[14]), .B(\stack[1][30] ), .Z(n7346) );
  XOR U8420 ( .A(n7347), .B(n7346), .Z(n7348) );
  XOR U8421 ( .A(n7349), .B(n7348), .Z(n7428) );
  XOR U8422 ( .A(n7429), .B(n7428), .Z(n7431) );
  AND U8423 ( .A(o[15]), .B(\stack[1][29] ), .Z(n7430) );
  XOR U8424 ( .A(n7431), .B(n7430), .Z(n7342) );
  XOR U8425 ( .A(n7343), .B(n7342), .Z(n7435) );
  NAND U8426 ( .A(n7219), .B(n7218), .Z(n7223) );
  NAND U8427 ( .A(n7221), .B(n7220), .Z(n7222) );
  NAND U8428 ( .A(n7223), .B(n7222), .Z(n7434) );
  XOR U8429 ( .A(n7435), .B(n7434), .Z(n7437) );
  AND U8430 ( .A(o[17]), .B(\stack[1][27] ), .Z(n7436) );
  XOR U8431 ( .A(n7437), .B(n7436), .Z(n7336) );
  XOR U8432 ( .A(n7337), .B(n7336), .Z(n7441) );
  NAND U8433 ( .A(n7225), .B(n7224), .Z(n7229) );
  NAND U8434 ( .A(n7227), .B(n7226), .Z(n7228) );
  NAND U8435 ( .A(n7229), .B(n7228), .Z(n7440) );
  XOR U8436 ( .A(n7441), .B(n7440), .Z(n7443) );
  AND U8437 ( .A(o[19]), .B(\stack[1][25] ), .Z(n7442) );
  XOR U8438 ( .A(n7443), .B(n7442), .Z(n7330) );
  XOR U8439 ( .A(n7331), .B(n7330), .Z(n7447) );
  NAND U8440 ( .A(n7231), .B(n7230), .Z(n7235) );
  NAND U8441 ( .A(n7233), .B(n7232), .Z(n7234) );
  NAND U8442 ( .A(n7235), .B(n7234), .Z(n7446) );
  XOR U8443 ( .A(n7447), .B(n7446), .Z(n7449) );
  AND U8444 ( .A(\stack[1][23] ), .B(o[21]), .Z(n7448) );
  XNOR U8445 ( .A(n7449), .B(n7448), .Z(n7324) );
  XNOR U8446 ( .A(n7325), .B(n7324), .Z(n7452) );
  XOR U8447 ( .A(n7453), .B(n7452), .Z(n7455) );
  AND U8448 ( .A(\stack[1][21] ), .B(o[23]), .Z(n7454) );
  XNOR U8449 ( .A(n7455), .B(n7454), .Z(n7318) );
  XNOR U8450 ( .A(n7319), .B(n7318), .Z(n7458) );
  AND U8451 ( .A(\stack[1][19] ), .B(o[25]), .Z(n7460) );
  XNOR U8452 ( .A(n7461), .B(n7460), .Z(n7313) );
  NAND U8453 ( .A(n7237), .B(n7236), .Z(n7241) );
  NAND U8454 ( .A(n7239), .B(n7238), .Z(n7240) );
  AND U8455 ( .A(n7241), .B(n7240), .Z(n7310) );
  NAND U8456 ( .A(\stack[1][18] ), .B(o[26]), .Z(n7311) );
  NAND U8457 ( .A(n7243), .B(n7242), .Z(n7247) );
  NAND U8458 ( .A(n7245), .B(n7244), .Z(n7246) );
  NAND U8459 ( .A(n7247), .B(n7246), .Z(n7464) );
  XOR U8460 ( .A(n7465), .B(n7464), .Z(n7466) );
  AND U8461 ( .A(\stack[1][17] ), .B(o[27]), .Z(n7467) );
  XOR U8462 ( .A(n7307), .B(n7306), .Z(n7470) );
  NAND U8463 ( .A(n7249), .B(n7248), .Z(n7253) );
  NAND U8464 ( .A(n7251), .B(n7250), .Z(n7252) );
  NAND U8465 ( .A(n7253), .B(n7252), .Z(n7471) );
  AND U8466 ( .A(\stack[1][15] ), .B(o[29]), .Z(n7473) );
  XOR U8467 ( .A(n7301), .B(n7300), .Z(n7476) );
  NAND U8468 ( .A(n7255), .B(n7254), .Z(n7259) );
  NAND U8469 ( .A(n7257), .B(n7256), .Z(n7258) );
  NAND U8470 ( .A(n7259), .B(n7258), .Z(n7477) );
  AND U8471 ( .A(\stack[1][13] ), .B(o[31]), .Z(n7479) );
  XOR U8472 ( .A(n7295), .B(n7294), .Z(n7482) );
  NAND U8473 ( .A(n7261), .B(n7260), .Z(n7265) );
  NAND U8474 ( .A(n7263), .B(n7262), .Z(n7264) );
  NAND U8475 ( .A(n7265), .B(n7264), .Z(n7483) );
  AND U8476 ( .A(\stack[1][11] ), .B(o[33]), .Z(n7485) );
  XOR U8477 ( .A(n7289), .B(n7288), .Z(n7488) );
  NAND U8478 ( .A(n7267), .B(n7266), .Z(n7271) );
  NAND U8479 ( .A(n7269), .B(n7268), .Z(n7270) );
  NAND U8480 ( .A(n7271), .B(n7270), .Z(n7489) );
  AND U8481 ( .A(\stack[1][9] ), .B(o[35]), .Z(n7491) );
  XOR U8482 ( .A(n7283), .B(n7282), .Z(n7494) );
  NAND U8483 ( .A(n7273), .B(n7272), .Z(n7277) );
  NAND U8484 ( .A(n7275), .B(n7274), .Z(n7276) );
  NAND U8485 ( .A(n7277), .B(n7276), .Z(n7495) );
  AND U8486 ( .A(\stack[1][7] ), .B(o[37]), .Z(n7496) );
  XNOR U8487 ( .A(n7497), .B(n7496), .Z(n12448) );
  NAND U8488 ( .A(n12449), .B(n12448), .Z(n7278) );
  AND U8489 ( .A(n7279), .B(n7278), .Z(n7501) );
  NAND U8490 ( .A(n7281), .B(n7280), .Z(n7285) );
  NAND U8491 ( .A(n7283), .B(n7282), .Z(n7284) );
  NAND U8492 ( .A(n7285), .B(n7284), .Z(n7507) );
  NAND U8493 ( .A(n7287), .B(n7286), .Z(n7291) );
  NAND U8494 ( .A(n7289), .B(n7288), .Z(n7290) );
  NAND U8495 ( .A(n7291), .B(n7290), .Z(n7513) );
  NAND U8496 ( .A(n7293), .B(n7292), .Z(n7297) );
  NAND U8497 ( .A(n7295), .B(n7294), .Z(n7296) );
  NAND U8498 ( .A(n7297), .B(n7296), .Z(n7519) );
  NAND U8499 ( .A(n7299), .B(n7298), .Z(n7303) );
  NAND U8500 ( .A(n7301), .B(n7300), .Z(n7302) );
  NAND U8501 ( .A(n7303), .B(n7302), .Z(n7525) );
  NAND U8502 ( .A(n7305), .B(n7304), .Z(n7309) );
  NAND U8503 ( .A(n7307), .B(n7306), .Z(n7308) );
  NAND U8504 ( .A(n7309), .B(n7308), .Z(n7537) );
  NAND U8505 ( .A(n7311), .B(n7310), .Z(n7315) );
  NAND U8506 ( .A(n7313), .B(n7312), .Z(n7314) );
  AND U8507 ( .A(n7315), .B(n7314), .Z(n7543) );
  NAND U8508 ( .A(n7317), .B(n7316), .Z(n7321) );
  NAND U8509 ( .A(n7319), .B(n7318), .Z(n7320) );
  AND U8510 ( .A(n7321), .B(n7320), .Z(n7549) );
  AND U8511 ( .A(\stack[1][22] ), .B(o[23]), .Z(n7557) );
  NAND U8512 ( .A(n7323), .B(n7322), .Z(n7327) );
  NAND U8513 ( .A(n7325), .B(n7324), .Z(n7326) );
  AND U8514 ( .A(n7327), .B(n7326), .Z(n7555) );
  AND U8515 ( .A(o[21]), .B(\stack[1][24] ), .Z(n7562) );
  NAND U8516 ( .A(n7329), .B(n7328), .Z(n7333) );
  NAND U8517 ( .A(n7331), .B(n7330), .Z(n7332) );
  NAND U8518 ( .A(n7333), .B(n7332), .Z(n7560) );
  NAND U8519 ( .A(n7335), .B(n7334), .Z(n7339) );
  NAND U8520 ( .A(n7337), .B(n7336), .Z(n7338) );
  NAND U8521 ( .A(n7339), .B(n7338), .Z(n7566) );
  NAND U8522 ( .A(n7341), .B(n7340), .Z(n7345) );
  NAND U8523 ( .A(n7343), .B(n7342), .Z(n7344) );
  NAND U8524 ( .A(n7345), .B(n7344), .Z(n7572) );
  AND U8525 ( .A(o[15]), .B(\stack[1][30] ), .Z(n7587) );
  NAND U8526 ( .A(n7347), .B(n7346), .Z(n7351) );
  NANDN U8527 ( .A(n7349), .B(n7348), .Z(n7350) );
  AND U8528 ( .A(n7351), .B(n7350), .Z(n7585) );
  AND U8529 ( .A(o[13]), .B(\stack[1][32] ), .Z(n7593) );
  NAND U8530 ( .A(n7353), .B(n7352), .Z(n7357) );
  NAND U8531 ( .A(n7355), .B(n7354), .Z(n7356) );
  AND U8532 ( .A(n7357), .B(n7356), .Z(n7591) );
  AND U8533 ( .A(o[11]), .B(\stack[1][34] ), .Z(n7598) );
  NAND U8534 ( .A(n7359), .B(n7358), .Z(n7363) );
  NAND U8535 ( .A(n7361), .B(n7360), .Z(n7362) );
  NAND U8536 ( .A(n7363), .B(n7362), .Z(n7596) );
  AND U8537 ( .A(o[10]), .B(\stack[1][35] ), .Z(n7605) );
  NAND U8538 ( .A(n7365), .B(n7364), .Z(n7369) );
  NAND U8539 ( .A(n7367), .B(n7366), .Z(n7368) );
  NAND U8540 ( .A(n7369), .B(n7368), .Z(n7654) );
  NAND U8541 ( .A(o[7]), .B(\stack[1][38] ), .Z(n7650) );
  AND U8542 ( .A(o[6]), .B(\stack[1][39] ), .Z(n7617) );
  AND U8543 ( .A(o[4]), .B(\stack[1][41] ), .Z(n7639) );
  NANDN U8544 ( .A(n7370), .B(n7625), .Z(n7374) );
  NANDN U8545 ( .A(n7372), .B(n7371), .Z(n7373) );
  NAND U8546 ( .A(n7374), .B(n7373), .Z(n7630) );
  AND U8547 ( .A(o[3]), .B(\stack[1][42] ), .Z(n7631) );
  XOR U8548 ( .A(n7630), .B(n7631), .Z(n7632) );
  AND U8549 ( .A(o[2]), .B(\stack[1][43] ), .Z(n7626) );
  AND U8550 ( .A(n7375), .B(n7377), .Z(n7376) );
  AND U8551 ( .A(o[1]), .B(\stack[1][45] ), .Z(n7622) );
  NAND U8552 ( .A(n7620), .B(n7622), .Z(n7853) );
  XOR U8553 ( .A(n7376), .B(n7853), .Z(n7379) );
  AND U8554 ( .A(o[0]), .B(\stack[1][45] ), .Z(n7848) );
  OR U8555 ( .A(n7377), .B(n7848), .Z(n7378) );
  NAND U8556 ( .A(n7379), .B(n7378), .Z(n7627) );
  XNOR U8557 ( .A(n7626), .B(n7627), .Z(n7633) );
  NAND U8558 ( .A(n7381), .B(n7380), .Z(n7385) );
  NAND U8559 ( .A(n7383), .B(n7382), .Z(n7384) );
  NAND U8560 ( .A(n7385), .B(n7384), .Z(n7636) );
  XOR U8561 ( .A(n7637), .B(n7636), .Z(n7638) );
  XOR U8562 ( .A(n7639), .B(n7638), .Z(n7643) );
  NAND U8563 ( .A(n7387), .B(n7386), .Z(n7391) );
  NAND U8564 ( .A(n7389), .B(n7388), .Z(n7390) );
  AND U8565 ( .A(n7391), .B(n7390), .Z(n7642) );
  XOR U8566 ( .A(n7643), .B(n7642), .Z(n7645) );
  AND U8567 ( .A(o[5]), .B(\stack[1][40] ), .Z(n7644) );
  XOR U8568 ( .A(n7645), .B(n7644), .Z(n7615) );
  NAND U8569 ( .A(n7393), .B(n7392), .Z(n7397) );
  NAND U8570 ( .A(n7395), .B(n7394), .Z(n7396) );
  NAND U8571 ( .A(n7397), .B(n7396), .Z(n7614) );
  XOR U8572 ( .A(n7615), .B(n7614), .Z(n7616) );
  XNOR U8573 ( .A(n7617), .B(n7616), .Z(n7649) );
  NAND U8574 ( .A(n7399), .B(n7398), .Z(n7403) );
  NANDN U8575 ( .A(n7401), .B(n7400), .Z(n7402) );
  NAND U8576 ( .A(n7403), .B(n7402), .Z(n7648) );
  XNOR U8577 ( .A(n7650), .B(n7651), .Z(n7611) );
  AND U8578 ( .A(o[8]), .B(\stack[1][37] ), .Z(n7609) );
  NAND U8579 ( .A(n7405), .B(n7404), .Z(n7409) );
  NAND U8580 ( .A(n7407), .B(n7406), .Z(n7408) );
  NAND U8581 ( .A(n7409), .B(n7408), .Z(n7608) );
  XOR U8582 ( .A(n7609), .B(n7608), .Z(n7610) );
  XOR U8583 ( .A(n7654), .B(n7655), .Z(n7657) );
  AND U8584 ( .A(o[9]), .B(\stack[1][36] ), .Z(n7656) );
  XOR U8585 ( .A(n7657), .B(n7656), .Z(n7603) );
  NAND U8586 ( .A(n7411), .B(n7410), .Z(n7415) );
  NAND U8587 ( .A(n7413), .B(n7412), .Z(n7414) );
  NAND U8588 ( .A(n7415), .B(n7414), .Z(n7602) );
  XOR U8589 ( .A(n7603), .B(n7602), .Z(n7604) );
  XOR U8590 ( .A(n7605), .B(n7604), .Z(n7597) );
  XOR U8591 ( .A(n7596), .B(n7597), .Z(n7599) );
  AND U8592 ( .A(o[12]), .B(\stack[1][33] ), .Z(n7661) );
  NAND U8593 ( .A(n7417), .B(n7416), .Z(n7421) );
  NAND U8594 ( .A(n7419), .B(n7418), .Z(n7420) );
  NAND U8595 ( .A(n7421), .B(n7420), .Z(n7660) );
  XOR U8596 ( .A(n7661), .B(n7660), .Z(n7662) );
  XOR U8597 ( .A(n7663), .B(n7662), .Z(n7590) );
  XOR U8598 ( .A(n7591), .B(n7590), .Z(n7592) );
  XOR U8599 ( .A(n7593), .B(n7592), .Z(n7669) );
  AND U8600 ( .A(o[14]), .B(\stack[1][31] ), .Z(n7667) );
  NAND U8601 ( .A(n7423), .B(n7422), .Z(n7427) );
  NAND U8602 ( .A(n7425), .B(n7424), .Z(n7426) );
  NAND U8603 ( .A(n7427), .B(n7426), .Z(n7666) );
  XOR U8604 ( .A(n7667), .B(n7666), .Z(n7668) );
  XOR U8605 ( .A(n7669), .B(n7668), .Z(n7584) );
  XOR U8606 ( .A(n7585), .B(n7584), .Z(n7586) );
  XOR U8607 ( .A(n7587), .B(n7586), .Z(n7581) );
  AND U8608 ( .A(o[16]), .B(\stack[1][29] ), .Z(n7579) );
  NAND U8609 ( .A(n7429), .B(n7428), .Z(n7433) );
  NAND U8610 ( .A(n7431), .B(n7430), .Z(n7432) );
  NAND U8611 ( .A(n7433), .B(n7432), .Z(n7578) );
  XOR U8612 ( .A(n7579), .B(n7578), .Z(n7580) );
  XOR U8613 ( .A(n7581), .B(n7580), .Z(n7573) );
  XOR U8614 ( .A(n7572), .B(n7573), .Z(n7575) );
  AND U8615 ( .A(o[17]), .B(\stack[1][28] ), .Z(n7574) );
  XOR U8616 ( .A(n7575), .B(n7574), .Z(n7675) );
  AND U8617 ( .A(o[18]), .B(\stack[1][27] ), .Z(n7673) );
  NAND U8618 ( .A(n7435), .B(n7434), .Z(n7439) );
  NAND U8619 ( .A(n7437), .B(n7436), .Z(n7438) );
  NAND U8620 ( .A(n7439), .B(n7438), .Z(n7672) );
  XOR U8621 ( .A(n7673), .B(n7672), .Z(n7674) );
  XOR U8622 ( .A(n7675), .B(n7674), .Z(n7567) );
  XOR U8623 ( .A(n7566), .B(n7567), .Z(n7569) );
  AND U8624 ( .A(o[19]), .B(\stack[1][26] ), .Z(n7568) );
  XOR U8625 ( .A(n7569), .B(n7568), .Z(n7681) );
  AND U8626 ( .A(o[20]), .B(\stack[1][25] ), .Z(n7679) );
  NAND U8627 ( .A(n7441), .B(n7440), .Z(n7445) );
  NAND U8628 ( .A(n7443), .B(n7442), .Z(n7444) );
  NAND U8629 ( .A(n7445), .B(n7444), .Z(n7678) );
  XOR U8630 ( .A(n7679), .B(n7678), .Z(n7680) );
  XOR U8631 ( .A(n7681), .B(n7680), .Z(n7561) );
  XOR U8632 ( .A(n7560), .B(n7561), .Z(n7563) );
  AND U8633 ( .A(\stack[1][23] ), .B(o[22]), .Z(n7685) );
  NAND U8634 ( .A(n7447), .B(n7446), .Z(n7451) );
  NAND U8635 ( .A(n7449), .B(n7448), .Z(n7450) );
  NAND U8636 ( .A(n7451), .B(n7450), .Z(n7684) );
  XOR U8637 ( .A(n7685), .B(n7684), .Z(n7686) );
  XOR U8638 ( .A(n7687), .B(n7686), .Z(n7554) );
  XOR U8639 ( .A(n7555), .B(n7554), .Z(n7556) );
  XOR U8640 ( .A(n7557), .B(n7556), .Z(n7693) );
  AND U8641 ( .A(\stack[1][21] ), .B(o[24]), .Z(n7691) );
  NAND U8642 ( .A(n7453), .B(n7452), .Z(n7457) );
  NAND U8643 ( .A(n7455), .B(n7454), .Z(n7456) );
  NAND U8644 ( .A(n7457), .B(n7456), .Z(n7690) );
  XOR U8645 ( .A(n7691), .B(n7690), .Z(n7692) );
  XOR U8646 ( .A(n7693), .B(n7692), .Z(n7548) );
  XOR U8647 ( .A(n7549), .B(n7548), .Z(n7550) );
  AND U8648 ( .A(\stack[1][20] ), .B(o[25]), .Z(n7551) );
  AND U8649 ( .A(\stack[1][19] ), .B(o[26]), .Z(n7696) );
  NAND U8650 ( .A(n7459), .B(n7458), .Z(n7463) );
  NAND U8651 ( .A(n7461), .B(n7460), .Z(n7462) );
  NAND U8652 ( .A(n7463), .B(n7462), .Z(n7697) );
  XOR U8653 ( .A(n7699), .B(n7698), .Z(n7542) );
  XOR U8654 ( .A(n7543), .B(n7542), .Z(n7544) );
  AND U8655 ( .A(\stack[1][18] ), .B(o[27]), .Z(n7545) );
  AND U8656 ( .A(\stack[1][17] ), .B(o[28]), .Z(n7702) );
  NAND U8657 ( .A(n7465), .B(n7464), .Z(n7469) );
  NAND U8658 ( .A(n7467), .B(n7466), .Z(n7468) );
  NAND U8659 ( .A(n7469), .B(n7468), .Z(n7703) );
  XOR U8660 ( .A(n7705), .B(n7704), .Z(n7536) );
  AND U8661 ( .A(\stack[1][16] ), .B(o[29]), .Z(n7539) );
  AND U8662 ( .A(\stack[1][15] ), .B(o[30]), .Z(n7530) );
  NAND U8663 ( .A(n7471), .B(n7470), .Z(n7475) );
  NAND U8664 ( .A(n7473), .B(n7472), .Z(n7474) );
  NAND U8665 ( .A(n7475), .B(n7474), .Z(n7531) );
  XOR U8666 ( .A(n7533), .B(n7532), .Z(n7524) );
  AND U8667 ( .A(\stack[1][14] ), .B(o[31]), .Z(n7527) );
  AND U8668 ( .A(\stack[1][13] ), .B(o[32]), .Z(n7708) );
  NAND U8669 ( .A(n7477), .B(n7476), .Z(n7481) );
  NAND U8670 ( .A(n7479), .B(n7478), .Z(n7480) );
  NAND U8671 ( .A(n7481), .B(n7480), .Z(n7709) );
  XOR U8672 ( .A(n7711), .B(n7710), .Z(n7518) );
  AND U8673 ( .A(\stack[1][12] ), .B(o[33]), .Z(n7521) );
  AND U8674 ( .A(\stack[1][11] ), .B(o[34]), .Z(n7714) );
  NAND U8675 ( .A(n7483), .B(n7482), .Z(n7487) );
  NAND U8676 ( .A(n7485), .B(n7484), .Z(n7486) );
  NAND U8677 ( .A(n7487), .B(n7486), .Z(n7715) );
  XOR U8678 ( .A(n7717), .B(n7716), .Z(n7512) );
  AND U8679 ( .A(\stack[1][10] ), .B(o[35]), .Z(n7515) );
  AND U8680 ( .A(\stack[1][9] ), .B(o[36]), .Z(n7720) );
  NAND U8681 ( .A(n7489), .B(n7488), .Z(n7493) );
  NAND U8682 ( .A(n7491), .B(n7490), .Z(n7492) );
  NAND U8683 ( .A(n7493), .B(n7492), .Z(n7721) );
  XOR U8684 ( .A(n7723), .B(n7722), .Z(n7506) );
  AND U8685 ( .A(\stack[1][8] ), .B(o[37]), .Z(n7509) );
  AND U8686 ( .A(\stack[1][7] ), .B(o[38]), .Z(n7726) );
  NAND U8687 ( .A(n7495), .B(n7494), .Z(n7499) );
  NAND U8688 ( .A(n7497), .B(n7496), .Z(n7498) );
  NAND U8689 ( .A(n7499), .B(n7498), .Z(n7727) );
  XOR U8690 ( .A(n7729), .B(n7728), .Z(n7500) );
  NAND U8691 ( .A(n7501), .B(n7500), .Z(n7503) );
  AND U8692 ( .A(\stack[1][6] ), .B(o[39]), .Z(n12454) );
  XOR U8693 ( .A(n7501), .B(n7500), .Z(n12455) );
  NAND U8694 ( .A(n12454), .B(n12455), .Z(n7502) );
  NAND U8695 ( .A(n7503), .B(n7502), .Z(n7504) );
  AND U8696 ( .A(\stack[1][6] ), .B(o[40]), .Z(n7505) );
  NAND U8697 ( .A(n7504), .B(n7505), .Z(n7733) );
  NAND U8698 ( .A(n7507), .B(n7506), .Z(n7511) );
  NAND U8699 ( .A(n7509), .B(n7508), .Z(n7510) );
  NAND U8700 ( .A(n7511), .B(n7510), .Z(n7735) );
  AND U8701 ( .A(\stack[1][8] ), .B(o[38]), .Z(n7734) );
  NAND U8702 ( .A(n7513), .B(n7512), .Z(n7517) );
  NAND U8703 ( .A(n7515), .B(n7514), .Z(n7516) );
  NAND U8704 ( .A(n7517), .B(n7516), .Z(n7741) );
  AND U8705 ( .A(\stack[1][10] ), .B(o[36]), .Z(n7740) );
  NAND U8706 ( .A(n7519), .B(n7518), .Z(n7523) );
  NAND U8707 ( .A(n7521), .B(n7520), .Z(n7522) );
  NAND U8708 ( .A(n7523), .B(n7522), .Z(n7747) );
  AND U8709 ( .A(\stack[1][12] ), .B(o[34]), .Z(n7746) );
  NAND U8710 ( .A(n7525), .B(n7524), .Z(n7529) );
  NAND U8711 ( .A(n7527), .B(n7526), .Z(n7528) );
  AND U8712 ( .A(n7529), .B(n7528), .Z(n7752) );
  NAND U8713 ( .A(\stack[1][14] ), .B(o[32]), .Z(n7753) );
  NAND U8714 ( .A(n7531), .B(n7530), .Z(n7535) );
  NAND U8715 ( .A(n7533), .B(n7532), .Z(n7534) );
  NAND U8716 ( .A(n7535), .B(n7534), .Z(n7937) );
  NAND U8717 ( .A(n7537), .B(n7536), .Z(n7541) );
  NAND U8718 ( .A(n7539), .B(n7538), .Z(n7540) );
  AND U8719 ( .A(n7541), .B(n7540), .Z(n7758) );
  NAND U8720 ( .A(\stack[1][16] ), .B(o[30]), .Z(n7759) );
  NAND U8721 ( .A(n7543), .B(n7542), .Z(n7547) );
  NAND U8722 ( .A(n7545), .B(n7544), .Z(n7546) );
  NAND U8723 ( .A(n7547), .B(n7546), .Z(n7765) );
  AND U8724 ( .A(\stack[1][18] ), .B(o[28]), .Z(n7764) );
  NAND U8725 ( .A(n7549), .B(n7548), .Z(n7553) );
  NAND U8726 ( .A(n7551), .B(n7550), .Z(n7552) );
  NAND U8727 ( .A(n7553), .B(n7552), .Z(n7771) );
  AND U8728 ( .A(\stack[1][20] ), .B(o[26]), .Z(n7770) );
  NAND U8729 ( .A(n7555), .B(n7554), .Z(n7559) );
  NAND U8730 ( .A(n7557), .B(n7556), .Z(n7558) );
  NAND U8731 ( .A(n7559), .B(n7558), .Z(n7776) );
  AND U8732 ( .A(\stack[1][22] ), .B(o[24]), .Z(n7777) );
  XOR U8733 ( .A(n7776), .B(n7777), .Z(n7779) );
  AND U8734 ( .A(\stack[1][23] ), .B(o[23]), .Z(n7915) );
  NAND U8735 ( .A(n7561), .B(n7560), .Z(n7565) );
  NAND U8736 ( .A(n7563), .B(n7562), .Z(n7564) );
  NAND U8737 ( .A(n7565), .B(n7564), .Z(n7782) );
  AND U8738 ( .A(o[22]), .B(\stack[1][24] ), .Z(n7783) );
  XOR U8739 ( .A(n7782), .B(n7783), .Z(n7785) );
  NAND U8740 ( .A(n7567), .B(n7566), .Z(n7571) );
  NAND U8741 ( .A(n7569), .B(n7568), .Z(n7570) );
  AND U8742 ( .A(n7571), .B(n7570), .Z(n7789) );
  NAND U8743 ( .A(o[20]), .B(\stack[1][26] ), .Z(n7788) );
  XOR U8744 ( .A(n7789), .B(n7788), .Z(n7790) );
  NAND U8745 ( .A(n7573), .B(n7572), .Z(n7577) );
  NAND U8746 ( .A(n7575), .B(n7574), .Z(n7576) );
  NAND U8747 ( .A(n7577), .B(n7576), .Z(n7794) );
  AND U8748 ( .A(o[18]), .B(\stack[1][28] ), .Z(n7795) );
  XOR U8749 ( .A(n7794), .B(n7795), .Z(n7797) );
  NAND U8750 ( .A(n7579), .B(n7578), .Z(n7583) );
  NAND U8751 ( .A(n7581), .B(n7580), .Z(n7582) );
  NAND U8752 ( .A(n7583), .B(n7582), .Z(n7801) );
  NAND U8753 ( .A(n7585), .B(n7584), .Z(n7589) );
  NAND U8754 ( .A(n7587), .B(n7586), .Z(n7588) );
  AND U8755 ( .A(n7589), .B(n7588), .Z(n7807) );
  NAND U8756 ( .A(o[16]), .B(\stack[1][30] ), .Z(n7806) );
  XOR U8757 ( .A(n7807), .B(n7806), .Z(n7809) );
  NAND U8758 ( .A(n7591), .B(n7590), .Z(n7595) );
  NAND U8759 ( .A(n7593), .B(n7592), .Z(n7594) );
  NAND U8760 ( .A(n7595), .B(n7594), .Z(n7812) );
  AND U8761 ( .A(o[14]), .B(\stack[1][32] ), .Z(n7813) );
  XOR U8762 ( .A(n7812), .B(n7813), .Z(n7815) );
  AND U8763 ( .A(o[13]), .B(\stack[1][33] ), .Z(n7891) );
  AND U8764 ( .A(o[12]), .B(\stack[1][34] ), .Z(n7819) );
  NAND U8765 ( .A(n7597), .B(n7596), .Z(n7601) );
  NAND U8766 ( .A(n7599), .B(n7598), .Z(n7600) );
  NAND U8767 ( .A(n7601), .B(n7600), .Z(n7818) );
  XOR U8768 ( .A(n7819), .B(n7818), .Z(n7821) );
  AND U8769 ( .A(o[11]), .B(\stack[1][35] ), .Z(n7885) );
  NAND U8770 ( .A(n7603), .B(n7602), .Z(n7607) );
  NAND U8771 ( .A(n7605), .B(n7604), .Z(n7606) );
  NAND U8772 ( .A(n7607), .B(n7606), .Z(n7882) );
  AND U8773 ( .A(o[10]), .B(\stack[1][36] ), .Z(n7827) );
  NAND U8774 ( .A(n7609), .B(n7608), .Z(n7613) );
  NAND U8775 ( .A(n7611), .B(n7610), .Z(n7612) );
  NAND U8776 ( .A(n7613), .B(n7612), .Z(n7877) );
  NAND U8777 ( .A(o[8]), .B(\stack[1][38] ), .Z(n7872) );
  NAND U8778 ( .A(n7615), .B(n7614), .Z(n7619) );
  NAND U8779 ( .A(n7617), .B(n7616), .Z(n7618) );
  NAND U8780 ( .A(n7619), .B(n7618), .Z(n7832) );
  AND U8781 ( .A(o[7]), .B(\stack[1][39] ), .Z(n7831) );
  AND U8782 ( .A(o[6]), .B(\stack[1][40] ), .Z(n7839) );
  AND U8783 ( .A(o[4]), .B(\stack[1][42] ), .Z(n7845) );
  AND U8784 ( .A(o[2]), .B(\stack[1][44] ), .Z(n7854) );
  AND U8785 ( .A(n7620), .B(n7622), .Z(n7621) );
  AND U8786 ( .A(o[1]), .B(\stack[1][46] ), .Z(n7850) );
  NAND U8787 ( .A(n7848), .B(n7850), .Z(n8055) );
  XOR U8788 ( .A(n7621), .B(n8055), .Z(n7624) );
  AND U8789 ( .A(o[0]), .B(\stack[1][46] ), .Z(n8050) );
  OR U8790 ( .A(n7622), .B(n8050), .Z(n7623) );
  NAND U8791 ( .A(n7624), .B(n7623), .Z(n7855) );
  XNOR U8792 ( .A(n7854), .B(n7855), .Z(n7860) );
  NANDN U8793 ( .A(n7625), .B(n7853), .Z(n7629) );
  NANDN U8794 ( .A(n7627), .B(n7626), .Z(n7628) );
  NAND U8795 ( .A(n7629), .B(n7628), .Z(n7858) );
  AND U8796 ( .A(o[3]), .B(\stack[1][43] ), .Z(n7859) );
  XOR U8797 ( .A(n7858), .B(n7859), .Z(n7861) );
  NAND U8798 ( .A(n7631), .B(n7630), .Z(n7635) );
  NAND U8799 ( .A(n7633), .B(n7632), .Z(n7634) );
  NAND U8800 ( .A(n7635), .B(n7634), .Z(n7842) );
  XOR U8801 ( .A(n7843), .B(n7842), .Z(n7844) );
  XOR U8802 ( .A(n7845), .B(n7844), .Z(n7865) );
  NAND U8803 ( .A(n7637), .B(n7636), .Z(n7641) );
  NAND U8804 ( .A(n7639), .B(n7638), .Z(n7640) );
  NAND U8805 ( .A(n7641), .B(n7640), .Z(n7864) );
  XOR U8806 ( .A(n7865), .B(n7864), .Z(n7867) );
  AND U8807 ( .A(o[5]), .B(\stack[1][41] ), .Z(n7866) );
  XOR U8808 ( .A(n7867), .B(n7866), .Z(n7837) );
  NAND U8809 ( .A(n7643), .B(n7642), .Z(n7647) );
  NAND U8810 ( .A(n7645), .B(n7644), .Z(n7646) );
  NAND U8811 ( .A(n7647), .B(n7646), .Z(n7836) );
  XOR U8812 ( .A(n7837), .B(n7836), .Z(n7838) );
  XOR U8813 ( .A(n7839), .B(n7838), .Z(n7830) );
  XOR U8814 ( .A(n7831), .B(n7830), .Z(n7833) );
  XNOR U8815 ( .A(n7832), .B(n7833), .Z(n7871) );
  NAND U8816 ( .A(n7649), .B(n7648), .Z(n7653) );
  NAND U8817 ( .A(n7651), .B(n7650), .Z(n7652) );
  NAND U8818 ( .A(n7653), .B(n7652), .Z(n7870) );
  XOR U8819 ( .A(n7872), .B(n7873), .Z(n7876) );
  XOR U8820 ( .A(n7877), .B(n7876), .Z(n7879) );
  AND U8821 ( .A(o[9]), .B(\stack[1][37] ), .Z(n7878) );
  XOR U8822 ( .A(n7879), .B(n7878), .Z(n7825) );
  NAND U8823 ( .A(n7655), .B(n7654), .Z(n7659) );
  NAND U8824 ( .A(n7657), .B(n7656), .Z(n7658) );
  NAND U8825 ( .A(n7659), .B(n7658), .Z(n7824) );
  XOR U8826 ( .A(n7825), .B(n7824), .Z(n7826) );
  XOR U8827 ( .A(n7827), .B(n7826), .Z(n7883) );
  XOR U8828 ( .A(n7882), .B(n7883), .Z(n7884) );
  XOR U8829 ( .A(n7885), .B(n7884), .Z(n7820) );
  XOR U8830 ( .A(n7821), .B(n7820), .Z(n7889) );
  NAND U8831 ( .A(n7661), .B(n7660), .Z(n7665) );
  NAND U8832 ( .A(n7663), .B(n7662), .Z(n7664) );
  NAND U8833 ( .A(n7665), .B(n7664), .Z(n7888) );
  XOR U8834 ( .A(n7889), .B(n7888), .Z(n7890) );
  XOR U8835 ( .A(n7891), .B(n7890), .Z(n7814) );
  XOR U8836 ( .A(n7815), .B(n7814), .Z(n7895) );
  NAND U8837 ( .A(n7667), .B(n7666), .Z(n7671) );
  NAND U8838 ( .A(n7669), .B(n7668), .Z(n7670) );
  NAND U8839 ( .A(n7671), .B(n7670), .Z(n7894) );
  XOR U8840 ( .A(n7895), .B(n7894), .Z(n7897) );
  AND U8841 ( .A(o[15]), .B(\stack[1][31] ), .Z(n7896) );
  XNOR U8842 ( .A(n7897), .B(n7896), .Z(n7808) );
  XNOR U8843 ( .A(n7809), .B(n7808), .Z(n7800) );
  XOR U8844 ( .A(n7801), .B(n7800), .Z(n7803) );
  AND U8845 ( .A(o[17]), .B(\stack[1][29] ), .Z(n7802) );
  XOR U8846 ( .A(n7803), .B(n7802), .Z(n7796) );
  XOR U8847 ( .A(n7797), .B(n7796), .Z(n7901) );
  NAND U8848 ( .A(n7673), .B(n7672), .Z(n7677) );
  NAND U8849 ( .A(n7675), .B(n7674), .Z(n7676) );
  NAND U8850 ( .A(n7677), .B(n7676), .Z(n7900) );
  XOR U8851 ( .A(n7901), .B(n7900), .Z(n7903) );
  AND U8852 ( .A(o[19]), .B(\stack[1][27] ), .Z(n7902) );
  XNOR U8853 ( .A(n7903), .B(n7902), .Z(n7791) );
  NAND U8854 ( .A(n7679), .B(n7678), .Z(n7683) );
  NAND U8855 ( .A(n7681), .B(n7680), .Z(n7682) );
  NAND U8856 ( .A(n7683), .B(n7682), .Z(n7906) );
  AND U8857 ( .A(o[21]), .B(\stack[1][25] ), .Z(n7908) );
  XOR U8858 ( .A(n7909), .B(n7908), .Z(n7784) );
  XOR U8859 ( .A(n7785), .B(n7784), .Z(n7913) );
  NAND U8860 ( .A(n7685), .B(n7684), .Z(n7689) );
  NAND U8861 ( .A(n7687), .B(n7686), .Z(n7688) );
  NAND U8862 ( .A(n7689), .B(n7688), .Z(n7912) );
  XOR U8863 ( .A(n7913), .B(n7912), .Z(n7914) );
  XOR U8864 ( .A(n7915), .B(n7914), .Z(n7778) );
  XOR U8865 ( .A(n7779), .B(n7778), .Z(n7919) );
  NAND U8866 ( .A(n7691), .B(n7690), .Z(n7695) );
  NAND U8867 ( .A(n7693), .B(n7692), .Z(n7694) );
  NAND U8868 ( .A(n7695), .B(n7694), .Z(n7918) );
  XOR U8869 ( .A(n7919), .B(n7918), .Z(n7921) );
  AND U8870 ( .A(\stack[1][21] ), .B(o[25]), .Z(n7920) );
  XOR U8871 ( .A(n7921), .B(n7920), .Z(n7772) );
  XOR U8872 ( .A(n7773), .B(n7772), .Z(n7924) );
  NAND U8873 ( .A(n7697), .B(n7696), .Z(n7701) );
  NAND U8874 ( .A(n7699), .B(n7698), .Z(n7700) );
  NAND U8875 ( .A(n7701), .B(n7700), .Z(n7925) );
  AND U8876 ( .A(\stack[1][19] ), .B(o[27]), .Z(n7927) );
  XOR U8877 ( .A(n7767), .B(n7766), .Z(n7930) );
  NAND U8878 ( .A(n7703), .B(n7702), .Z(n7707) );
  NAND U8879 ( .A(n7705), .B(n7704), .Z(n7706) );
  NAND U8880 ( .A(n7707), .B(n7706), .Z(n7931) );
  AND U8881 ( .A(\stack[1][17] ), .B(o[29]), .Z(n7932) );
  XNOR U8882 ( .A(n7933), .B(n7932), .Z(n7760) );
  XNOR U8883 ( .A(n7761), .B(n7760), .Z(n7936) );
  AND U8884 ( .A(\stack[1][15] ), .B(o[31]), .Z(n7938) );
  XNOR U8885 ( .A(n7939), .B(n7938), .Z(n7754) );
  XNOR U8886 ( .A(n7755), .B(n7754), .Z(n7943) );
  NAND U8887 ( .A(n7709), .B(n7708), .Z(n7713) );
  NAND U8888 ( .A(n7711), .B(n7710), .Z(n7712) );
  NAND U8889 ( .A(n7713), .B(n7712), .Z(n7942) );
  AND U8890 ( .A(\stack[1][13] ), .B(o[33]), .Z(n7945) );
  XOR U8891 ( .A(n7749), .B(n7748), .Z(n7948) );
  NAND U8892 ( .A(n7715), .B(n7714), .Z(n7719) );
  NAND U8893 ( .A(n7717), .B(n7716), .Z(n7718) );
  NAND U8894 ( .A(n7719), .B(n7718), .Z(n7949) );
  AND U8895 ( .A(\stack[1][11] ), .B(o[35]), .Z(n7951) );
  XOR U8896 ( .A(n7743), .B(n7742), .Z(n7954) );
  NAND U8897 ( .A(n7721), .B(n7720), .Z(n7725) );
  NAND U8898 ( .A(n7723), .B(n7722), .Z(n7724) );
  NAND U8899 ( .A(n7725), .B(n7724), .Z(n7955) );
  AND U8900 ( .A(\stack[1][9] ), .B(o[37]), .Z(n7957) );
  XOR U8901 ( .A(n7737), .B(n7736), .Z(n7960) );
  NAND U8902 ( .A(n7727), .B(n7726), .Z(n7731) );
  NAND U8903 ( .A(n7729), .B(n7728), .Z(n7730) );
  NAND U8904 ( .A(n7731), .B(n7730), .Z(n7961) );
  AND U8905 ( .A(\stack[1][7] ), .B(o[39]), .Z(n7963) );
  NAND U8906 ( .A(n12461), .B(n12460), .Z(n7732) );
  NAND U8907 ( .A(n7733), .B(n7732), .Z(n7966) );
  AND U8908 ( .A(\stack[1][8] ), .B(o[39]), .Z(n7975) );
  NAND U8909 ( .A(n7735), .B(n7734), .Z(n7739) );
  NAND U8910 ( .A(n7737), .B(n7736), .Z(n7738) );
  NAND U8911 ( .A(n7739), .B(n7738), .Z(n7973) );
  AND U8912 ( .A(\stack[1][10] ), .B(o[37]), .Z(n7981) );
  NAND U8913 ( .A(n7741), .B(n7740), .Z(n7745) );
  NAND U8914 ( .A(n7743), .B(n7742), .Z(n7744) );
  NAND U8915 ( .A(n7745), .B(n7744), .Z(n7979) );
  AND U8916 ( .A(\stack[1][12] ), .B(o[35]), .Z(n8189) );
  NAND U8917 ( .A(n7747), .B(n7746), .Z(n7751) );
  NAND U8918 ( .A(n7749), .B(n7748), .Z(n7750) );
  NAND U8919 ( .A(n7751), .B(n7750), .Z(n8187) );
  NAND U8920 ( .A(n7753), .B(n7752), .Z(n7757) );
  NAND U8921 ( .A(n7755), .B(n7754), .Z(n7756) );
  AND U8922 ( .A(n7757), .B(n7756), .Z(n7991) );
  NAND U8923 ( .A(n7759), .B(n7758), .Z(n7763) );
  NAND U8924 ( .A(n7761), .B(n7760), .Z(n7762) );
  AND U8925 ( .A(n7763), .B(n7762), .Z(n8175) );
  NAND U8926 ( .A(n7765), .B(n7764), .Z(n7769) );
  NAND U8927 ( .A(n7767), .B(n7766), .Z(n7768) );
  NAND U8928 ( .A(n7769), .B(n7768), .Z(n7997) );
  NAND U8929 ( .A(n7771), .B(n7770), .Z(n7775) );
  NAND U8930 ( .A(n7773), .B(n7772), .Z(n7774) );
  NAND U8931 ( .A(n7775), .B(n7774), .Z(n8002) );
  AND U8932 ( .A(\stack[1][22] ), .B(o[25]), .Z(n8152) );
  NAND U8933 ( .A(n7777), .B(n7776), .Z(n7781) );
  NAND U8934 ( .A(n7779), .B(n7778), .Z(n7780) );
  NAND U8935 ( .A(n7781), .B(n7780), .Z(n8150) );
  NAND U8936 ( .A(n7783), .B(n7782), .Z(n7787) );
  NAND U8937 ( .A(n7785), .B(n7784), .Z(n7786) );
  NAND U8938 ( .A(n7787), .B(n7786), .Z(n8138) );
  AND U8939 ( .A(o[21]), .B(\stack[1][26] ), .Z(n8017) );
  NAND U8940 ( .A(n7789), .B(n7788), .Z(n7793) );
  NAND U8941 ( .A(n7791), .B(n7790), .Z(n7792) );
  AND U8942 ( .A(n7793), .B(n7792), .Z(n8015) );
  AND U8943 ( .A(o[19]), .B(\stack[1][28] ), .Z(n8128) );
  NAND U8944 ( .A(n7795), .B(n7794), .Z(n7799) );
  NAND U8945 ( .A(n7797), .B(n7796), .Z(n7798) );
  NAND U8946 ( .A(n7799), .B(n7798), .Z(n8126) );
  AND U8947 ( .A(o[18]), .B(\stack[1][29] ), .Z(n8121) );
  NAND U8948 ( .A(n7801), .B(n7800), .Z(n7805) );
  NAND U8949 ( .A(n7803), .B(n7802), .Z(n7804) );
  NAND U8950 ( .A(n7805), .B(n7804), .Z(n8120) );
  XOR U8951 ( .A(n8121), .B(n8120), .Z(n8123) );
  NAND U8952 ( .A(n7807), .B(n7806), .Z(n7811) );
  NAND U8953 ( .A(n7809), .B(n7808), .Z(n7810) );
  AND U8954 ( .A(n7811), .B(n7810), .Z(n8021) );
  AND U8955 ( .A(o[15]), .B(\stack[1][32] ), .Z(n8028) );
  NAND U8956 ( .A(n7813), .B(n7812), .Z(n7817) );
  NAND U8957 ( .A(n7815), .B(n7814), .Z(n7816) );
  NAND U8958 ( .A(n7817), .B(n7816), .Z(n8026) );
  NAND U8959 ( .A(n7819), .B(n7818), .Z(n7823) );
  NAND U8960 ( .A(n7821), .B(n7820), .Z(n7822) );
  AND U8961 ( .A(n7823), .B(n7822), .Z(n8102) );
  NAND U8962 ( .A(n7825), .B(n7824), .Z(n7829) );
  NAND U8963 ( .A(n7827), .B(n7826), .Z(n7828) );
  AND U8964 ( .A(n7829), .B(n7828), .Z(n8096) );
  AND U8965 ( .A(o[10]), .B(\stack[1][37] ), .Z(n8090) );
  NAND U8966 ( .A(o[9]), .B(\stack[1][38] ), .Z(n8040) );
  NAND U8967 ( .A(n7831), .B(n7830), .Z(n7835) );
  NAND U8968 ( .A(n7833), .B(n7832), .Z(n7834) );
  NAND U8969 ( .A(n7835), .B(n7834), .Z(n8086) );
  NAND U8970 ( .A(n7837), .B(n7836), .Z(n7841) );
  NAND U8971 ( .A(n7839), .B(n7838), .Z(n7840) );
  NAND U8972 ( .A(n7841), .B(n7840), .Z(n8080) );
  AND U8973 ( .A(o[7]), .B(\stack[1][40] ), .Z(n8079) );
  AND U8974 ( .A(o[6]), .B(\stack[1][41] ), .Z(n8047) );
  AND U8975 ( .A(o[5]), .B(\stack[1][42] ), .Z(n8074) );
  NAND U8976 ( .A(n7843), .B(n7842), .Z(n7847) );
  NAND U8977 ( .A(n7845), .B(n7844), .Z(n7846) );
  NAND U8978 ( .A(n7847), .B(n7846), .Z(n8072) );
  AND U8979 ( .A(o[2]), .B(\stack[1][45] ), .Z(n8056) );
  AND U8980 ( .A(n7848), .B(n7850), .Z(n7849) );
  AND U8981 ( .A(o[1]), .B(\stack[1][47] ), .Z(n8052) );
  NAND U8982 ( .A(n8050), .B(n8052), .Z(n8326) );
  XOR U8983 ( .A(n7849), .B(n8326), .Z(n7852) );
  AND U8984 ( .A(o[0]), .B(\stack[1][47] ), .Z(n8331) );
  OR U8985 ( .A(n7850), .B(n8331), .Z(n7851) );
  NAND U8986 ( .A(n7852), .B(n7851), .Z(n8057) );
  XNOR U8987 ( .A(n8056), .B(n8057), .Z(n8061) );
  NANDN U8988 ( .A(n7853), .B(n8055), .Z(n7857) );
  NANDN U8989 ( .A(n7855), .B(n7854), .Z(n7856) );
  NAND U8990 ( .A(n7857), .B(n7856), .Z(n8060) );
  XOR U8991 ( .A(n8061), .B(n8060), .Z(n8063) );
  AND U8992 ( .A(o[3]), .B(\stack[1][44] ), .Z(n8062) );
  XOR U8993 ( .A(n8063), .B(n8062), .Z(n8067) );
  NAND U8994 ( .A(n7859), .B(n7858), .Z(n7863) );
  NAND U8995 ( .A(n7861), .B(n7860), .Z(n7862) );
  NAND U8996 ( .A(n7863), .B(n7862), .Z(n8066) );
  XOR U8997 ( .A(n8067), .B(n8066), .Z(n8069) );
  AND U8998 ( .A(o[4]), .B(\stack[1][43] ), .Z(n8068) );
  XOR U8999 ( .A(n8069), .B(n8068), .Z(n8073) );
  XOR U9000 ( .A(n8072), .B(n8073), .Z(n8075) );
  NAND U9001 ( .A(n7865), .B(n7864), .Z(n7869) );
  NAND U9002 ( .A(n7867), .B(n7866), .Z(n7868) );
  NAND U9003 ( .A(n7869), .B(n7868), .Z(n8044) );
  XOR U9004 ( .A(n8045), .B(n8044), .Z(n8046) );
  XOR U9005 ( .A(n8047), .B(n8046), .Z(n8078) );
  XOR U9006 ( .A(n8079), .B(n8078), .Z(n8081) );
  XOR U9007 ( .A(n8080), .B(n8081), .Z(n8085) );
  AND U9008 ( .A(o[8]), .B(\stack[1][39] ), .Z(n8084) );
  XOR U9009 ( .A(n8085), .B(n8084), .Z(n8087) );
  XNOR U9010 ( .A(n8086), .B(n8087), .Z(n8039) );
  NAND U9011 ( .A(n7871), .B(n7870), .Z(n7875) );
  NANDN U9012 ( .A(n7873), .B(n7872), .Z(n7874) );
  NAND U9013 ( .A(n7875), .B(n7874), .Z(n8038) );
  XNOR U9014 ( .A(n8040), .B(n8041), .Z(n8091) );
  NAND U9015 ( .A(n7877), .B(n7876), .Z(n7881) );
  NAND U9016 ( .A(n7879), .B(n7878), .Z(n7880) );
  NAND U9017 ( .A(n7881), .B(n7880), .Z(n8092) );
  XNOR U9018 ( .A(n8093), .B(n8092), .Z(n8097) );
  NAND U9019 ( .A(o[11]), .B(\stack[1][36] ), .Z(n8098) );
  XNOR U9020 ( .A(n8099), .B(n8098), .Z(n8035) );
  NAND U9021 ( .A(n7883), .B(n7882), .Z(n7887) );
  NAND U9022 ( .A(n7885), .B(n7884), .Z(n7886) );
  NAND U9023 ( .A(n7887), .B(n7886), .Z(n8032) );
  AND U9024 ( .A(o[12]), .B(\stack[1][35] ), .Z(n8033) );
  XOR U9025 ( .A(n8032), .B(n8033), .Z(n8034) );
  NAND U9026 ( .A(o[13]), .B(\stack[1][34] ), .Z(n8104) );
  XNOR U9027 ( .A(n8105), .B(n8104), .Z(n8111) );
  AND U9028 ( .A(o[14]), .B(\stack[1][33] ), .Z(n8109) );
  NAND U9029 ( .A(n7889), .B(n7888), .Z(n7893) );
  NAND U9030 ( .A(n7891), .B(n7890), .Z(n7892) );
  NAND U9031 ( .A(n7893), .B(n7892), .Z(n8108) );
  XOR U9032 ( .A(n8109), .B(n8108), .Z(n8110) );
  XOR U9033 ( .A(n8026), .B(n8027), .Z(n8029) );
  XNOR U9034 ( .A(n8028), .B(n8029), .Z(n8117) );
  AND U9035 ( .A(o[16]), .B(\stack[1][31] ), .Z(n8115) );
  NAND U9036 ( .A(n7895), .B(n7894), .Z(n7899) );
  NAND U9037 ( .A(n7897), .B(n7896), .Z(n7898) );
  NAND U9038 ( .A(n7899), .B(n7898), .Z(n8114) );
  XOR U9039 ( .A(n8115), .B(n8114), .Z(n8116) );
  XOR U9040 ( .A(n8117), .B(n8116), .Z(n8020) );
  XOR U9041 ( .A(n8021), .B(n8020), .Z(n8023) );
  AND U9042 ( .A(o[17]), .B(\stack[1][30] ), .Z(n8022) );
  XOR U9043 ( .A(n8023), .B(n8022), .Z(n8122) );
  XOR U9044 ( .A(n8123), .B(n8122), .Z(n8127) );
  XOR U9045 ( .A(n8126), .B(n8127), .Z(n8129) );
  AND U9046 ( .A(o[20]), .B(\stack[1][27] ), .Z(n8133) );
  NAND U9047 ( .A(n7901), .B(n7900), .Z(n7905) );
  NAND U9048 ( .A(n7903), .B(n7902), .Z(n7904) );
  NAND U9049 ( .A(n7905), .B(n7904), .Z(n8132) );
  XOR U9050 ( .A(n8133), .B(n8132), .Z(n8134) );
  XOR U9051 ( .A(n8135), .B(n8134), .Z(n8014) );
  XOR U9052 ( .A(n8015), .B(n8014), .Z(n8016) );
  XOR U9053 ( .A(n8017), .B(n8016), .Z(n8011) );
  AND U9054 ( .A(o[22]), .B(\stack[1][25] ), .Z(n8009) );
  NAND U9055 ( .A(n7907), .B(n7906), .Z(n7911) );
  NAND U9056 ( .A(n7909), .B(n7908), .Z(n7910) );
  NAND U9057 ( .A(n7911), .B(n7910), .Z(n8008) );
  XOR U9058 ( .A(n8009), .B(n8008), .Z(n8010) );
  XOR U9059 ( .A(n8011), .B(n8010), .Z(n8139) );
  XOR U9060 ( .A(n8138), .B(n8139), .Z(n8141) );
  AND U9061 ( .A(\stack[1][24] ), .B(o[23]), .Z(n8140) );
  XOR U9062 ( .A(n8141), .B(n8140), .Z(n8147) );
  AND U9063 ( .A(\stack[1][23] ), .B(o[24]), .Z(n8145) );
  NAND U9064 ( .A(n7913), .B(n7912), .Z(n7917) );
  NAND U9065 ( .A(n7915), .B(n7914), .Z(n7916) );
  NAND U9066 ( .A(n7917), .B(n7916), .Z(n8144) );
  XOR U9067 ( .A(n8145), .B(n8144), .Z(n8146) );
  XOR U9068 ( .A(n8147), .B(n8146), .Z(n8151) );
  XOR U9069 ( .A(n8150), .B(n8151), .Z(n8153) );
  AND U9070 ( .A(\stack[1][21] ), .B(o[26]), .Z(n8157) );
  NAND U9071 ( .A(n7919), .B(n7918), .Z(n7923) );
  NAND U9072 ( .A(n7921), .B(n7920), .Z(n7922) );
  NAND U9073 ( .A(n7923), .B(n7922), .Z(n8156) );
  XOR U9074 ( .A(n8157), .B(n8156), .Z(n8158) );
  XOR U9075 ( .A(n8159), .B(n8158), .Z(n8003) );
  XOR U9076 ( .A(n8002), .B(n8003), .Z(n8005) );
  AND U9077 ( .A(\stack[1][20] ), .B(o[27]), .Z(n8004) );
  XOR U9078 ( .A(n8005), .B(n8004), .Z(n8165) );
  AND U9079 ( .A(\stack[1][19] ), .B(o[28]), .Z(n8163) );
  NAND U9080 ( .A(n7925), .B(n7924), .Z(n7929) );
  NAND U9081 ( .A(n7927), .B(n7926), .Z(n7928) );
  NAND U9082 ( .A(n7929), .B(n7928), .Z(n8162) );
  XOR U9083 ( .A(n8163), .B(n8162), .Z(n8164) );
  XOR U9084 ( .A(n8165), .B(n8164), .Z(n7996) );
  AND U9085 ( .A(\stack[1][18] ), .B(o[29]), .Z(n7999) );
  AND U9086 ( .A(\stack[1][17] ), .B(o[30]), .Z(n8168) );
  NAND U9087 ( .A(n7931), .B(n7930), .Z(n7935) );
  NAND U9088 ( .A(n7933), .B(n7932), .Z(n7934) );
  NAND U9089 ( .A(n7935), .B(n7934), .Z(n8169) );
  XOR U9090 ( .A(n8171), .B(n8170), .Z(n8174) );
  XOR U9091 ( .A(n8175), .B(n8174), .Z(n8176) );
  AND U9092 ( .A(\stack[1][16] ), .B(o[31]), .Z(n8177) );
  AND U9093 ( .A(\stack[1][15] ), .B(o[32]), .Z(n8180) );
  NAND U9094 ( .A(n7937), .B(n7936), .Z(n7941) );
  NAND U9095 ( .A(n7939), .B(n7938), .Z(n7940) );
  NAND U9096 ( .A(n7941), .B(n7940), .Z(n8181) );
  XOR U9097 ( .A(n8183), .B(n8182), .Z(n7990) );
  XOR U9098 ( .A(n7991), .B(n7990), .Z(n7992) );
  AND U9099 ( .A(\stack[1][14] ), .B(o[33]), .Z(n7993) );
  AND U9100 ( .A(\stack[1][13] ), .B(o[34]), .Z(n7984) );
  NAND U9101 ( .A(n7943), .B(n7942), .Z(n7947) );
  NAND U9102 ( .A(n7945), .B(n7944), .Z(n7946) );
  NAND U9103 ( .A(n7947), .B(n7946), .Z(n7985) );
  XOR U9104 ( .A(n7987), .B(n7986), .Z(n8186) );
  XOR U9105 ( .A(n8189), .B(n8188), .Z(n8195) );
  AND U9106 ( .A(\stack[1][11] ), .B(o[36]), .Z(n8192) );
  NAND U9107 ( .A(n7949), .B(n7948), .Z(n7953) );
  NAND U9108 ( .A(n7951), .B(n7950), .Z(n7952) );
  NAND U9109 ( .A(n7953), .B(n7952), .Z(n8193) );
  XOR U9110 ( .A(n8195), .B(n8194), .Z(n7978) );
  XOR U9111 ( .A(n7981), .B(n7980), .Z(n8201) );
  AND U9112 ( .A(\stack[1][9] ), .B(o[38]), .Z(n8198) );
  NAND U9113 ( .A(n7955), .B(n7954), .Z(n7959) );
  NAND U9114 ( .A(n7957), .B(n7956), .Z(n7958) );
  NAND U9115 ( .A(n7959), .B(n7958), .Z(n8199) );
  XOR U9116 ( .A(n8201), .B(n8200), .Z(n7972) );
  XOR U9117 ( .A(n7975), .B(n7974), .Z(n8207) );
  AND U9118 ( .A(\stack[1][7] ), .B(o[40]), .Z(n8204) );
  NAND U9119 ( .A(n7961), .B(n7960), .Z(n7965) );
  NAND U9120 ( .A(n7963), .B(n7962), .Z(n7964) );
  NAND U9121 ( .A(n7965), .B(n7964), .Z(n8205) );
  XOR U9122 ( .A(n8207), .B(n8206), .Z(n7967) );
  NAND U9123 ( .A(n7966), .B(n7967), .Z(n7969) );
  AND U9124 ( .A(\stack[1][6] ), .B(o[41]), .Z(n12466) );
  NAND U9125 ( .A(n12466), .B(n12467), .Z(n7968) );
  NAND U9126 ( .A(n7969), .B(n7968), .Z(n7970) );
  AND U9127 ( .A(\stack[1][6] ), .B(o[42]), .Z(n7971) );
  NAND U9128 ( .A(n7970), .B(n7971), .Z(n8211) );
  NAND U9129 ( .A(n7973), .B(n7972), .Z(n7977) );
  NAND U9130 ( .A(n7975), .B(n7974), .Z(n7976) );
  NAND U9131 ( .A(n7977), .B(n7976), .Z(n8213) );
  AND U9132 ( .A(\stack[1][8] ), .B(o[40]), .Z(n8212) );
  NAND U9133 ( .A(n7979), .B(n7978), .Z(n7983) );
  NAND U9134 ( .A(n7981), .B(n7980), .Z(n7982) );
  NAND U9135 ( .A(n7983), .B(n7982), .Z(n8219) );
  AND U9136 ( .A(\stack[1][10] ), .B(o[38]), .Z(n8218) );
  NAND U9137 ( .A(n7985), .B(n7984), .Z(n7989) );
  NAND U9138 ( .A(n7987), .B(n7986), .Z(n7988) );
  NAND U9139 ( .A(n7989), .B(n7988), .Z(n8433) );
  NAND U9140 ( .A(n7991), .B(n7990), .Z(n7995) );
  NAND U9141 ( .A(n7993), .B(n7992), .Z(n7994) );
  AND U9142 ( .A(n7995), .B(n7994), .Z(n8230) );
  NAND U9143 ( .A(\stack[1][14] ), .B(o[34]), .Z(n8231) );
  NAND U9144 ( .A(n7997), .B(n7996), .Z(n8001) );
  NAND U9145 ( .A(n7999), .B(n7998), .Z(n8000) );
  NAND U9146 ( .A(n8001), .B(n8000), .Z(n8243) );
  AND U9147 ( .A(\stack[1][18] ), .B(o[30]), .Z(n8242) );
  NAND U9148 ( .A(n8003), .B(n8002), .Z(n8007) );
  NAND U9149 ( .A(n8005), .B(n8004), .Z(n8006) );
  NAND U9150 ( .A(n8007), .B(n8006), .Z(n8248) );
  AND U9151 ( .A(\stack[1][20] ), .B(o[28]), .Z(n8249) );
  XOR U9152 ( .A(n8248), .B(n8249), .Z(n8251) );
  NAND U9153 ( .A(n8009), .B(n8008), .Z(n8013) );
  NAND U9154 ( .A(n8011), .B(n8010), .Z(n8012) );
  NAND U9155 ( .A(n8013), .B(n8012), .Z(n8397) );
  NAND U9156 ( .A(n8015), .B(n8014), .Z(n8019) );
  NAND U9157 ( .A(n8017), .B(n8016), .Z(n8018) );
  AND U9158 ( .A(n8019), .B(n8018), .Z(n8267) );
  NAND U9159 ( .A(o[22]), .B(\stack[1][26] ), .Z(n8266) );
  XOR U9160 ( .A(n8267), .B(n8266), .Z(n8269) );
  NAND U9161 ( .A(n8021), .B(n8020), .Z(n8025) );
  NAND U9162 ( .A(n8023), .B(n8022), .Z(n8024) );
  NAND U9163 ( .A(n8025), .B(n8024), .Z(n8278) );
  AND U9164 ( .A(o[18]), .B(\stack[1][30] ), .Z(n8279) );
  XOR U9165 ( .A(n8278), .B(n8279), .Z(n8281) );
  NANDN U9166 ( .A(n8027), .B(n8026), .Z(n8031) );
  NANDN U9167 ( .A(n8029), .B(n8028), .Z(n8030) );
  NAND U9168 ( .A(n8031), .B(n8030), .Z(n8290) );
  AND U9169 ( .A(o[16]), .B(\stack[1][32] ), .Z(n8291) );
  XOR U9170 ( .A(n8290), .B(n8291), .Z(n8293) );
  NAND U9171 ( .A(n8033), .B(n8032), .Z(n8037) );
  NAND U9172 ( .A(n8035), .B(n8034), .Z(n8036) );
  NAND U9173 ( .A(n8037), .B(n8036), .Z(n8372) );
  NAND U9174 ( .A(o[10]), .B(\stack[1][38] ), .Z(n8368) );
  NAND U9175 ( .A(n8039), .B(n8038), .Z(n8043) );
  NAND U9176 ( .A(n8041), .B(n8040), .Z(n8042) );
  NAND U9177 ( .A(n8043), .B(n8042), .Z(n8366) );
  NAND U9178 ( .A(o[9]), .B(\stack[1][39] ), .Z(n8316) );
  NAND U9179 ( .A(n8045), .B(n8044), .Z(n8049) );
  NAND U9180 ( .A(n8047), .B(n8046), .Z(n8048) );
  NAND U9181 ( .A(n8049), .B(n8048), .Z(n8356) );
  AND U9182 ( .A(o[6]), .B(\stack[1][42] ), .Z(n8323) );
  AND U9183 ( .A(o[5]), .B(\stack[1][43] ), .Z(n8351) );
  AND U9184 ( .A(o[4]), .B(\stack[1][44] ), .Z(n8345) );
  AND U9185 ( .A(o[2]), .B(\stack[1][46] ), .Z(n8327) );
  AND U9186 ( .A(n8050), .B(n8052), .Z(n8051) );
  AND U9187 ( .A(o[1]), .B(\stack[1][48] ), .Z(n8333) );
  NAND U9188 ( .A(n8331), .B(n8333), .Z(n8568) );
  XOR U9189 ( .A(n8051), .B(n8568), .Z(n8054) );
  AND U9190 ( .A(o[0]), .B(\stack[1][48] ), .Z(n8573) );
  OR U9191 ( .A(n8052), .B(n8573), .Z(n8053) );
  NAND U9192 ( .A(n8054), .B(n8053), .Z(n8328) );
  XNOR U9193 ( .A(n8327), .B(n8328), .Z(n8337) );
  NANDN U9194 ( .A(n8055), .B(n8326), .Z(n8059) );
  NANDN U9195 ( .A(n8057), .B(n8056), .Z(n8058) );
  NAND U9196 ( .A(n8059), .B(n8058), .Z(n8336) );
  XOR U9197 ( .A(n8337), .B(n8336), .Z(n8339) );
  AND U9198 ( .A(o[3]), .B(\stack[1][45] ), .Z(n8338) );
  XOR U9199 ( .A(n8339), .B(n8338), .Z(n8343) );
  NAND U9200 ( .A(n8061), .B(n8060), .Z(n8065) );
  NAND U9201 ( .A(n8063), .B(n8062), .Z(n8064) );
  NAND U9202 ( .A(n8065), .B(n8064), .Z(n8342) );
  XOR U9203 ( .A(n8343), .B(n8342), .Z(n8344) );
  XOR U9204 ( .A(n8345), .B(n8344), .Z(n8349) );
  NAND U9205 ( .A(n8067), .B(n8066), .Z(n8071) );
  NAND U9206 ( .A(n8069), .B(n8068), .Z(n8070) );
  NAND U9207 ( .A(n8071), .B(n8070), .Z(n8348) );
  XOR U9208 ( .A(n8349), .B(n8348), .Z(n8350) );
  XOR U9209 ( .A(n8351), .B(n8350), .Z(n8321) );
  NAND U9210 ( .A(n8073), .B(n8072), .Z(n8077) );
  NAND U9211 ( .A(n8075), .B(n8074), .Z(n8076) );
  NAND U9212 ( .A(n8077), .B(n8076), .Z(n8320) );
  XOR U9213 ( .A(n8321), .B(n8320), .Z(n8322) );
  XOR U9214 ( .A(n8323), .B(n8322), .Z(n8355) );
  AND U9215 ( .A(o[7]), .B(\stack[1][41] ), .Z(n8354) );
  XOR U9216 ( .A(n8355), .B(n8354), .Z(n8357) );
  XNOR U9217 ( .A(n8356), .B(n8357), .Z(n8363) );
  NAND U9218 ( .A(o[8]), .B(\stack[1][40] ), .Z(n8360) );
  NAND U9219 ( .A(n8079), .B(n8078), .Z(n8083) );
  NAND U9220 ( .A(n8081), .B(n8080), .Z(n8082) );
  AND U9221 ( .A(n8083), .B(n8082), .Z(n8361) );
  XOR U9222 ( .A(n8360), .B(n8361), .Z(n8362) );
  NAND U9223 ( .A(n8085), .B(n8084), .Z(n8089) );
  NAND U9224 ( .A(n8087), .B(n8086), .Z(n8088) );
  AND U9225 ( .A(n8089), .B(n8088), .Z(n8314) );
  XOR U9226 ( .A(n8315), .B(n8314), .Z(n8317) );
  XOR U9227 ( .A(n8316), .B(n8317), .Z(n8367) );
  XOR U9228 ( .A(n8366), .B(n8367), .Z(n8369) );
  XNOR U9229 ( .A(n8368), .B(n8369), .Z(n8311) );
  AND U9230 ( .A(o[11]), .B(\stack[1][37] ), .Z(n8309) );
  NAND U9231 ( .A(n8091), .B(n8090), .Z(n8095) );
  NAND U9232 ( .A(n8093), .B(n8092), .Z(n8094) );
  NAND U9233 ( .A(n8095), .B(n8094), .Z(n8308) );
  XOR U9234 ( .A(n8309), .B(n8308), .Z(n8310) );
  AND U9235 ( .A(o[12]), .B(\stack[1][36] ), .Z(n8303) );
  NAND U9236 ( .A(n8097), .B(n8096), .Z(n8101) );
  NAND U9237 ( .A(n8099), .B(n8098), .Z(n8100) );
  AND U9238 ( .A(n8101), .B(n8100), .Z(n8302) );
  XOR U9239 ( .A(n8303), .B(n8302), .Z(n8304) );
  XOR U9240 ( .A(n8305), .B(n8304), .Z(n8373) );
  XOR U9241 ( .A(n8372), .B(n8373), .Z(n8375) );
  AND U9242 ( .A(o[13]), .B(\stack[1][35] ), .Z(n8374) );
  XOR U9243 ( .A(n8375), .B(n8374), .Z(n8299) );
  AND U9244 ( .A(o[14]), .B(\stack[1][34] ), .Z(n8297) );
  NAND U9245 ( .A(n8103), .B(n8102), .Z(n8107) );
  NAND U9246 ( .A(n8105), .B(n8104), .Z(n8106) );
  AND U9247 ( .A(n8107), .B(n8106), .Z(n8296) );
  XOR U9248 ( .A(n8297), .B(n8296), .Z(n8298) );
  XOR U9249 ( .A(n8299), .B(n8298), .Z(n8379) );
  NAND U9250 ( .A(n8109), .B(n8108), .Z(n8113) );
  NAND U9251 ( .A(n8111), .B(n8110), .Z(n8112) );
  NAND U9252 ( .A(n8113), .B(n8112), .Z(n8378) );
  XOR U9253 ( .A(n8379), .B(n8378), .Z(n8381) );
  AND U9254 ( .A(o[15]), .B(\stack[1][33] ), .Z(n8380) );
  XOR U9255 ( .A(n8381), .B(n8380), .Z(n8292) );
  XOR U9256 ( .A(n8293), .B(n8292), .Z(n8285) );
  NAND U9257 ( .A(n8115), .B(n8114), .Z(n8119) );
  NAND U9258 ( .A(n8117), .B(n8116), .Z(n8118) );
  NAND U9259 ( .A(n8119), .B(n8118), .Z(n8284) );
  XOR U9260 ( .A(n8285), .B(n8284), .Z(n8287) );
  AND U9261 ( .A(o[17]), .B(\stack[1][31] ), .Z(n8286) );
  XOR U9262 ( .A(n8287), .B(n8286), .Z(n8280) );
  XOR U9263 ( .A(n8281), .B(n8280), .Z(n8385) );
  NAND U9264 ( .A(n8121), .B(n8120), .Z(n8125) );
  NAND U9265 ( .A(n8123), .B(n8122), .Z(n8124) );
  NAND U9266 ( .A(n8125), .B(n8124), .Z(n8384) );
  XOR U9267 ( .A(n8385), .B(n8384), .Z(n8387) );
  AND U9268 ( .A(o[19]), .B(\stack[1][29] ), .Z(n8386) );
  XOR U9269 ( .A(n8387), .B(n8386), .Z(n8274) );
  NAND U9270 ( .A(n8127), .B(n8126), .Z(n8131) );
  NAND U9271 ( .A(n8129), .B(n8128), .Z(n8130) );
  NAND U9272 ( .A(n8131), .B(n8130), .Z(n8272) );
  AND U9273 ( .A(o[20]), .B(\stack[1][28] ), .Z(n8273) );
  XOR U9274 ( .A(n8272), .B(n8273), .Z(n8275) );
  NAND U9275 ( .A(n8133), .B(n8132), .Z(n8137) );
  NAND U9276 ( .A(n8135), .B(n8134), .Z(n8136) );
  NAND U9277 ( .A(n8137), .B(n8136), .Z(n8390) );
  XOR U9278 ( .A(n8391), .B(n8390), .Z(n8393) );
  AND U9279 ( .A(o[21]), .B(\stack[1][27] ), .Z(n8392) );
  XNOR U9280 ( .A(n8393), .B(n8392), .Z(n8268) );
  XNOR U9281 ( .A(n8269), .B(n8268), .Z(n8396) );
  XOR U9282 ( .A(n8397), .B(n8396), .Z(n8399) );
  AND U9283 ( .A(\stack[1][25] ), .B(o[23]), .Z(n8398) );
  XNOR U9284 ( .A(n8399), .B(n8398), .Z(n8263) );
  NAND U9285 ( .A(\stack[1][24] ), .B(o[24]), .Z(n8260) );
  NAND U9286 ( .A(n8139), .B(n8138), .Z(n8143) );
  NAND U9287 ( .A(n8141), .B(n8140), .Z(n8142) );
  AND U9288 ( .A(n8143), .B(n8142), .Z(n8261) );
  XOR U9289 ( .A(n8260), .B(n8261), .Z(n8262) );
  NAND U9290 ( .A(n8145), .B(n8144), .Z(n8149) );
  NAND U9291 ( .A(n8147), .B(n8146), .Z(n8148) );
  NAND U9292 ( .A(n8149), .B(n8148), .Z(n8402) );
  AND U9293 ( .A(\stack[1][23] ), .B(o[25]), .Z(n8404) );
  XNOR U9294 ( .A(n8405), .B(n8404), .Z(n8257) );
  NAND U9295 ( .A(\stack[1][22] ), .B(o[26]), .Z(n8254) );
  NAND U9296 ( .A(n8151), .B(n8150), .Z(n8155) );
  NAND U9297 ( .A(n8153), .B(n8152), .Z(n8154) );
  AND U9298 ( .A(n8155), .B(n8154), .Z(n8255) );
  XOR U9299 ( .A(n8254), .B(n8255), .Z(n8256) );
  NAND U9300 ( .A(n8157), .B(n8156), .Z(n8161) );
  NAND U9301 ( .A(n8159), .B(n8158), .Z(n8160) );
  NAND U9302 ( .A(n8161), .B(n8160), .Z(n8408) );
  AND U9303 ( .A(\stack[1][21] ), .B(o[27]), .Z(n8410) );
  XOR U9304 ( .A(n8411), .B(n8410), .Z(n8250) );
  XOR U9305 ( .A(n8251), .B(n8250), .Z(n8415) );
  NAND U9306 ( .A(n8163), .B(n8162), .Z(n8167) );
  NAND U9307 ( .A(n8165), .B(n8164), .Z(n8166) );
  NAND U9308 ( .A(n8167), .B(n8166), .Z(n8414) );
  XOR U9309 ( .A(n8415), .B(n8414), .Z(n8417) );
  AND U9310 ( .A(\stack[1][19] ), .B(o[29]), .Z(n8416) );
  XOR U9311 ( .A(n8417), .B(n8416), .Z(n8244) );
  XOR U9312 ( .A(n8245), .B(n8244), .Z(n8420) );
  NAND U9313 ( .A(n8169), .B(n8168), .Z(n8173) );
  NAND U9314 ( .A(n8171), .B(n8170), .Z(n8172) );
  NAND U9315 ( .A(n8173), .B(n8172), .Z(n8421) );
  AND U9316 ( .A(\stack[1][17] ), .B(o[31]), .Z(n8423) );
  NAND U9317 ( .A(n8175), .B(n8174), .Z(n8179) );
  NAND U9318 ( .A(n8177), .B(n8176), .Z(n8178) );
  NAND U9319 ( .A(n8179), .B(n8178), .Z(n8237) );
  AND U9320 ( .A(\stack[1][16] ), .B(o[32]), .Z(n8236) );
  XOR U9321 ( .A(n8239), .B(n8238), .Z(n8426) );
  NAND U9322 ( .A(n8181), .B(n8180), .Z(n8185) );
  NAND U9323 ( .A(n8183), .B(n8182), .Z(n8184) );
  NAND U9324 ( .A(n8185), .B(n8184), .Z(n8427) );
  AND U9325 ( .A(\stack[1][15] ), .B(o[33]), .Z(n8428) );
  XNOR U9326 ( .A(n8429), .B(n8428), .Z(n8232) );
  XNOR U9327 ( .A(n8233), .B(n8232), .Z(n8432) );
  AND U9328 ( .A(\stack[1][13] ), .B(o[35]), .Z(n8434) );
  XNOR U9329 ( .A(n8435), .B(n8434), .Z(n8227) );
  NAND U9330 ( .A(n8187), .B(n8186), .Z(n8191) );
  NAND U9331 ( .A(n8189), .B(n8188), .Z(n8190) );
  AND U9332 ( .A(n8191), .B(n8190), .Z(n8224) );
  NAND U9333 ( .A(\stack[1][12] ), .B(o[36]), .Z(n8225) );
  NAND U9334 ( .A(n8193), .B(n8192), .Z(n8197) );
  NAND U9335 ( .A(n8195), .B(n8194), .Z(n8196) );
  NAND U9336 ( .A(n8197), .B(n8196), .Z(n8438) );
  XOR U9337 ( .A(n8439), .B(n8438), .Z(n8440) );
  AND U9338 ( .A(\stack[1][11] ), .B(o[37]), .Z(n8441) );
  XOR U9339 ( .A(n8221), .B(n8220), .Z(n8444) );
  NAND U9340 ( .A(n8199), .B(n8198), .Z(n8203) );
  NAND U9341 ( .A(n8201), .B(n8200), .Z(n8202) );
  NAND U9342 ( .A(n8203), .B(n8202), .Z(n8445) );
  AND U9343 ( .A(\stack[1][9] ), .B(o[39]), .Z(n8447) );
  XOR U9344 ( .A(n8215), .B(n8214), .Z(n8450) );
  NAND U9345 ( .A(n8205), .B(n8204), .Z(n8209) );
  NAND U9346 ( .A(n8207), .B(n8206), .Z(n8208) );
  NAND U9347 ( .A(n8209), .B(n8208), .Z(n8451) );
  AND U9348 ( .A(\stack[1][7] ), .B(o[41]), .Z(n8453) );
  NAND U9349 ( .A(n12473), .B(n12472), .Z(n8210) );
  NAND U9350 ( .A(n8211), .B(n8210), .Z(n8456) );
  AND U9351 ( .A(\stack[1][8] ), .B(o[41]), .Z(n8463) );
  NAND U9352 ( .A(n8213), .B(n8212), .Z(n8217) );
  NAND U9353 ( .A(n8215), .B(n8214), .Z(n8216) );
  NAND U9354 ( .A(n8217), .B(n8216), .Z(n8461) );
  AND U9355 ( .A(\stack[1][10] ), .B(o[39]), .Z(n8469) );
  NAND U9356 ( .A(n8219), .B(n8218), .Z(n8223) );
  NAND U9357 ( .A(n8221), .B(n8220), .Z(n8222) );
  NAND U9358 ( .A(n8223), .B(n8222), .Z(n8467) );
  NAND U9359 ( .A(n8225), .B(n8224), .Z(n8229) );
  NAND U9360 ( .A(n8227), .B(n8226), .Z(n8228) );
  AND U9361 ( .A(n8229), .B(n8228), .Z(n8473) );
  AND U9362 ( .A(\stack[1][14] ), .B(o[35]), .Z(n8481) );
  NAND U9363 ( .A(n8231), .B(n8230), .Z(n8235) );
  NAND U9364 ( .A(n8233), .B(n8232), .Z(n8234) );
  AND U9365 ( .A(n8235), .B(n8234), .Z(n8479) );
  NAND U9366 ( .A(n8237), .B(n8236), .Z(n8241) );
  NAND U9367 ( .A(n8239), .B(n8238), .Z(n8240) );
  NAND U9368 ( .A(n8241), .B(n8240), .Z(n8485) );
  AND U9369 ( .A(\stack[1][18] ), .B(o[31]), .Z(n8492) );
  NAND U9370 ( .A(n8243), .B(n8242), .Z(n8247) );
  NAND U9371 ( .A(n8245), .B(n8244), .Z(n8246) );
  NAND U9372 ( .A(n8247), .B(n8246), .Z(n8490) );
  AND U9373 ( .A(\stack[1][20] ), .B(o[29]), .Z(n8498) );
  NAND U9374 ( .A(n8249), .B(n8248), .Z(n8253) );
  NAND U9375 ( .A(n8251), .B(n8250), .Z(n8252) );
  NAND U9376 ( .A(n8253), .B(n8252), .Z(n8496) );
  AND U9377 ( .A(\stack[1][22] ), .B(o[27]), .Z(n8505) );
  NAND U9378 ( .A(n8255), .B(n8254), .Z(n8259) );
  NAND U9379 ( .A(n8257), .B(n8256), .Z(n8258) );
  AND U9380 ( .A(n8259), .B(n8258), .Z(n8503) );
  AND U9381 ( .A(\stack[1][24] ), .B(o[25]), .Z(n8511) );
  NAND U9382 ( .A(n8261), .B(n8260), .Z(n8265) );
  NAND U9383 ( .A(n8263), .B(n8262), .Z(n8264) );
  AND U9384 ( .A(n8265), .B(n8264), .Z(n8509) );
  NAND U9385 ( .A(n8267), .B(n8266), .Z(n8271) );
  NAND U9386 ( .A(n8269), .B(n8268), .Z(n8270) );
  AND U9387 ( .A(n8271), .B(n8270), .Z(n8515) );
  AND U9388 ( .A(o[21]), .B(\stack[1][28] ), .Z(n8522) );
  NAND U9389 ( .A(n8273), .B(n8272), .Z(n8277) );
  NAND U9390 ( .A(n8275), .B(n8274), .Z(n8276) );
  NAND U9391 ( .A(n8277), .B(n8276), .Z(n8520) );
  AND U9392 ( .A(o[19]), .B(\stack[1][30] ), .Z(n8528) );
  NAND U9393 ( .A(n8279), .B(n8278), .Z(n8283) );
  NAND U9394 ( .A(n8281), .B(n8280), .Z(n8282) );
  NAND U9395 ( .A(n8283), .B(n8282), .Z(n8526) );
  AND U9396 ( .A(o[18]), .B(\stack[1][31] ), .Z(n8633) );
  NAND U9397 ( .A(n8285), .B(n8284), .Z(n8289) );
  NAND U9398 ( .A(n8287), .B(n8286), .Z(n8288) );
  NAND U9399 ( .A(n8289), .B(n8288), .Z(n8632) );
  XOR U9400 ( .A(n8633), .B(n8632), .Z(n8635) );
  NAND U9401 ( .A(n8291), .B(n8290), .Z(n8295) );
  NAND U9402 ( .A(n8293), .B(n8292), .Z(n8294) );
  NAND U9403 ( .A(n8295), .B(n8294), .Z(n8532) );
  AND U9404 ( .A(o[15]), .B(\stack[1][34] ), .Z(n8540) );
  NAND U9405 ( .A(n8297), .B(n8296), .Z(n8301) );
  NAND U9406 ( .A(n8299), .B(n8298), .Z(n8300) );
  NAND U9407 ( .A(n8301), .B(n8300), .Z(n8538) );
  AND U9408 ( .A(o[13]), .B(\stack[1][36] ), .Z(n8622) );
  NAND U9409 ( .A(n8303), .B(n8302), .Z(n8307) );
  NAND U9410 ( .A(n8305), .B(n8304), .Z(n8306) );
  NAND U9411 ( .A(n8307), .B(n8306), .Z(n8620) );
  NAND U9412 ( .A(n8309), .B(n8308), .Z(n8313) );
  NAND U9413 ( .A(n8311), .B(n8310), .Z(n8312) );
  NAND U9414 ( .A(n8313), .B(n8312), .Z(n8616) );
  AND U9415 ( .A(o[12]), .B(\stack[1][37] ), .Z(n8615) );
  NAND U9416 ( .A(o[11]), .B(\stack[1][38] ), .Z(n8610) );
  AND U9417 ( .A(o[10]), .B(\stack[1][39] ), .Z(n8605) );
  NAND U9418 ( .A(n8315), .B(n8314), .Z(n8319) );
  NAND U9419 ( .A(n8317), .B(n8316), .Z(n8318) );
  AND U9420 ( .A(n8319), .B(n8318), .Z(n8603) );
  NAND U9421 ( .A(o[9]), .B(\stack[1][40] ), .Z(n8552) );
  NAND U9422 ( .A(n8321), .B(n8320), .Z(n8325) );
  NAND U9423 ( .A(n8323), .B(n8322), .Z(n8324) );
  NAND U9424 ( .A(n8325), .B(n8324), .Z(n8592) );
  AND U9425 ( .A(o[6]), .B(\stack[1][43] ), .Z(n8559) );
  AND U9426 ( .A(o[5]), .B(\stack[1][44] ), .Z(n8587) );
  NANDN U9427 ( .A(n8326), .B(n8568), .Z(n8330) );
  NANDN U9428 ( .A(n8328), .B(n8327), .Z(n8329) );
  NAND U9429 ( .A(n8330), .B(n8329), .Z(n8578) );
  AND U9430 ( .A(o[3]), .B(\stack[1][46] ), .Z(n8579) );
  XOR U9431 ( .A(n8578), .B(n8579), .Z(n8580) );
  AND U9432 ( .A(o[2]), .B(\stack[1][47] ), .Z(n8569) );
  AND U9433 ( .A(n8331), .B(n8333), .Z(n8332) );
  AND U9434 ( .A(o[1]), .B(\stack[1][49] ), .Z(n8575) );
  NAND U9435 ( .A(n8573), .B(n8575), .Z(n8846) );
  XOR U9436 ( .A(n8332), .B(n8846), .Z(n8335) );
  AND U9437 ( .A(o[0]), .B(\stack[1][49] ), .Z(n8851) );
  OR U9438 ( .A(n8333), .B(n8851), .Z(n8334) );
  NAND U9439 ( .A(n8335), .B(n8334), .Z(n8570) );
  XNOR U9440 ( .A(n8569), .B(n8570), .Z(n8581) );
  NAND U9441 ( .A(n8337), .B(n8336), .Z(n8341) );
  NAND U9442 ( .A(n8339), .B(n8338), .Z(n8340) );
  NAND U9443 ( .A(n8341), .B(n8340), .Z(n8562) );
  XOR U9444 ( .A(n8563), .B(n8562), .Z(n8565) );
  AND U9445 ( .A(o[4]), .B(\stack[1][45] ), .Z(n8564) );
  XOR U9446 ( .A(n8565), .B(n8564), .Z(n8585) );
  NAND U9447 ( .A(n8343), .B(n8342), .Z(n8347) );
  NAND U9448 ( .A(n8345), .B(n8344), .Z(n8346) );
  NAND U9449 ( .A(n8347), .B(n8346), .Z(n8584) );
  XOR U9450 ( .A(n8585), .B(n8584), .Z(n8586) );
  XOR U9451 ( .A(n8587), .B(n8586), .Z(n8557) );
  NAND U9452 ( .A(n8349), .B(n8348), .Z(n8353) );
  NAND U9453 ( .A(n8351), .B(n8350), .Z(n8352) );
  NAND U9454 ( .A(n8353), .B(n8352), .Z(n8556) );
  XOR U9455 ( .A(n8557), .B(n8556), .Z(n8558) );
  XOR U9456 ( .A(n8559), .B(n8558), .Z(n8591) );
  AND U9457 ( .A(o[7]), .B(\stack[1][42] ), .Z(n8590) );
  XOR U9458 ( .A(n8591), .B(n8590), .Z(n8593) );
  XOR U9459 ( .A(n8592), .B(n8593), .Z(n8599) );
  AND U9460 ( .A(o[8]), .B(\stack[1][41] ), .Z(n8597) );
  NAND U9461 ( .A(n8355), .B(n8354), .Z(n8359) );
  NAND U9462 ( .A(n8357), .B(n8356), .Z(n8358) );
  NAND U9463 ( .A(n8359), .B(n8358), .Z(n8596) );
  XOR U9464 ( .A(n8597), .B(n8596), .Z(n8598) );
  XNOR U9465 ( .A(n8599), .B(n8598), .Z(n8551) );
  NAND U9466 ( .A(n8361), .B(n8360), .Z(n8365) );
  NAND U9467 ( .A(n8363), .B(n8362), .Z(n8364) );
  NAND U9468 ( .A(n8365), .B(n8364), .Z(n8550) );
  XOR U9469 ( .A(n8552), .B(n8553), .Z(n8602) );
  XOR U9470 ( .A(n8603), .B(n8602), .Z(n8604) );
  XNOR U9471 ( .A(n8605), .B(n8604), .Z(n8609) );
  NAND U9472 ( .A(n8367), .B(n8366), .Z(n8371) );
  NAND U9473 ( .A(n8369), .B(n8368), .Z(n8370) );
  NAND U9474 ( .A(n8371), .B(n8370), .Z(n8608) );
  XOR U9475 ( .A(n8610), .B(n8611), .Z(n8614) );
  XOR U9476 ( .A(n8615), .B(n8614), .Z(n8617) );
  XOR U9477 ( .A(n8616), .B(n8617), .Z(n8621) );
  XNOR U9478 ( .A(n8622), .B(n8623), .Z(n8547) );
  NAND U9479 ( .A(n8373), .B(n8372), .Z(n8377) );
  NAND U9480 ( .A(n8375), .B(n8374), .Z(n8376) );
  NAND U9481 ( .A(n8377), .B(n8376), .Z(n8544) );
  AND U9482 ( .A(o[14]), .B(\stack[1][35] ), .Z(n8545) );
  XOR U9483 ( .A(n8544), .B(n8545), .Z(n8546) );
  XOR U9484 ( .A(n8547), .B(n8546), .Z(n8539) );
  XOR U9485 ( .A(n8538), .B(n8539), .Z(n8541) );
  AND U9486 ( .A(o[16]), .B(\stack[1][33] ), .Z(n8627) );
  NAND U9487 ( .A(n8379), .B(n8378), .Z(n8383) );
  NAND U9488 ( .A(n8381), .B(n8380), .Z(n8382) );
  NAND U9489 ( .A(n8383), .B(n8382), .Z(n8626) );
  XOR U9490 ( .A(n8627), .B(n8626), .Z(n8628) );
  XOR U9491 ( .A(n8629), .B(n8628), .Z(n8533) );
  XOR U9492 ( .A(n8532), .B(n8533), .Z(n8535) );
  AND U9493 ( .A(o[17]), .B(\stack[1][32] ), .Z(n8534) );
  XOR U9494 ( .A(n8535), .B(n8534), .Z(n8634) );
  XOR U9495 ( .A(n8635), .B(n8634), .Z(n8527) );
  XOR U9496 ( .A(n8526), .B(n8527), .Z(n8529) );
  AND U9497 ( .A(o[20]), .B(\stack[1][29] ), .Z(n8639) );
  NAND U9498 ( .A(n8385), .B(n8384), .Z(n8389) );
  NAND U9499 ( .A(n8387), .B(n8386), .Z(n8388) );
  NAND U9500 ( .A(n8389), .B(n8388), .Z(n8638) );
  XOR U9501 ( .A(n8639), .B(n8638), .Z(n8640) );
  XOR U9502 ( .A(n8641), .B(n8640), .Z(n8521) );
  XOR U9503 ( .A(n8520), .B(n8521), .Z(n8523) );
  AND U9504 ( .A(o[22]), .B(\stack[1][27] ), .Z(n8645) );
  NAND U9505 ( .A(n8391), .B(n8390), .Z(n8395) );
  NAND U9506 ( .A(n8393), .B(n8392), .Z(n8394) );
  NAND U9507 ( .A(n8395), .B(n8394), .Z(n8644) );
  XOR U9508 ( .A(n8645), .B(n8644), .Z(n8646) );
  XOR U9509 ( .A(n8647), .B(n8646), .Z(n8514) );
  XOR U9510 ( .A(n8515), .B(n8514), .Z(n8517) );
  AND U9511 ( .A(o[23]), .B(\stack[1][26] ), .Z(n8516) );
  XOR U9512 ( .A(n8517), .B(n8516), .Z(n8653) );
  AND U9513 ( .A(\stack[1][25] ), .B(o[24]), .Z(n8651) );
  NAND U9514 ( .A(n8397), .B(n8396), .Z(n8401) );
  NAND U9515 ( .A(n8399), .B(n8398), .Z(n8400) );
  NAND U9516 ( .A(n8401), .B(n8400), .Z(n8650) );
  XOR U9517 ( .A(n8651), .B(n8650), .Z(n8652) );
  XOR U9518 ( .A(n8653), .B(n8652), .Z(n8508) );
  XOR U9519 ( .A(n8509), .B(n8508), .Z(n8510) );
  XOR U9520 ( .A(n8511), .B(n8510), .Z(n8659) );
  AND U9521 ( .A(\stack[1][23] ), .B(o[26]), .Z(n8657) );
  NAND U9522 ( .A(n8403), .B(n8402), .Z(n8407) );
  NAND U9523 ( .A(n8405), .B(n8404), .Z(n8406) );
  NAND U9524 ( .A(n8407), .B(n8406), .Z(n8656) );
  XOR U9525 ( .A(n8657), .B(n8656), .Z(n8658) );
  XOR U9526 ( .A(n8659), .B(n8658), .Z(n8502) );
  XOR U9527 ( .A(n8503), .B(n8502), .Z(n8504) );
  XOR U9528 ( .A(n8505), .B(n8504), .Z(n8665) );
  AND U9529 ( .A(\stack[1][21] ), .B(o[28]), .Z(n8663) );
  NAND U9530 ( .A(n8409), .B(n8408), .Z(n8413) );
  NAND U9531 ( .A(n8411), .B(n8410), .Z(n8412) );
  NAND U9532 ( .A(n8413), .B(n8412), .Z(n8662) );
  XOR U9533 ( .A(n8663), .B(n8662), .Z(n8664) );
  XOR U9534 ( .A(n8665), .B(n8664), .Z(n8497) );
  XOR U9535 ( .A(n8496), .B(n8497), .Z(n8499) );
  AND U9536 ( .A(\stack[1][19] ), .B(o[30]), .Z(n8669) );
  NAND U9537 ( .A(n8415), .B(n8414), .Z(n8419) );
  NAND U9538 ( .A(n8417), .B(n8416), .Z(n8418) );
  NAND U9539 ( .A(n8419), .B(n8418), .Z(n8668) );
  XOR U9540 ( .A(n8669), .B(n8668), .Z(n8670) );
  XOR U9541 ( .A(n8671), .B(n8670), .Z(n8491) );
  XOR U9542 ( .A(n8490), .B(n8491), .Z(n8493) );
  AND U9543 ( .A(\stack[1][17] ), .B(o[32]), .Z(n8675) );
  NAND U9544 ( .A(n8421), .B(n8420), .Z(n8425) );
  NAND U9545 ( .A(n8423), .B(n8422), .Z(n8424) );
  NAND U9546 ( .A(n8425), .B(n8424), .Z(n8674) );
  XOR U9547 ( .A(n8675), .B(n8674), .Z(n8676) );
  XOR U9548 ( .A(n8677), .B(n8676), .Z(n8484) );
  AND U9549 ( .A(\stack[1][16] ), .B(o[33]), .Z(n8487) );
  AND U9550 ( .A(\stack[1][15] ), .B(o[34]), .Z(n8680) );
  NAND U9551 ( .A(n8427), .B(n8426), .Z(n8431) );
  NAND U9552 ( .A(n8429), .B(n8428), .Z(n8430) );
  NAND U9553 ( .A(n8431), .B(n8430), .Z(n8681) );
  XOR U9554 ( .A(n8683), .B(n8682), .Z(n8478) );
  XOR U9555 ( .A(n8479), .B(n8478), .Z(n8480) );
  XOR U9556 ( .A(n8481), .B(n8480), .Z(n8689) );
  AND U9557 ( .A(\stack[1][13] ), .B(o[36]), .Z(n8686) );
  NAND U9558 ( .A(n8433), .B(n8432), .Z(n8437) );
  NAND U9559 ( .A(n8435), .B(n8434), .Z(n8436) );
  NAND U9560 ( .A(n8437), .B(n8436), .Z(n8687) );
  XOR U9561 ( .A(n8689), .B(n8688), .Z(n8472) );
  XOR U9562 ( .A(n8473), .B(n8472), .Z(n8474) );
  AND U9563 ( .A(\stack[1][12] ), .B(o[37]), .Z(n8475) );
  AND U9564 ( .A(\stack[1][11] ), .B(o[38]), .Z(n8692) );
  NAND U9565 ( .A(n8439), .B(n8438), .Z(n8443) );
  NAND U9566 ( .A(n8441), .B(n8440), .Z(n8442) );
  NAND U9567 ( .A(n8443), .B(n8442), .Z(n8693) );
  XOR U9568 ( .A(n8695), .B(n8694), .Z(n8466) );
  XOR U9569 ( .A(n8469), .B(n8468), .Z(n8701) );
  AND U9570 ( .A(\stack[1][9] ), .B(o[40]), .Z(n8698) );
  NAND U9571 ( .A(n8445), .B(n8444), .Z(n8449) );
  NAND U9572 ( .A(n8447), .B(n8446), .Z(n8448) );
  NAND U9573 ( .A(n8449), .B(n8448), .Z(n8699) );
  XOR U9574 ( .A(n8701), .B(n8700), .Z(n8460) );
  XOR U9575 ( .A(n8463), .B(n8462), .Z(n8707) );
  AND U9576 ( .A(\stack[1][7] ), .B(o[42]), .Z(n8704) );
  NAND U9577 ( .A(n8451), .B(n8450), .Z(n8455) );
  NAND U9578 ( .A(n8453), .B(n8452), .Z(n8454) );
  NAND U9579 ( .A(n8455), .B(n8454), .Z(n8705) );
  XOR U9580 ( .A(n8707), .B(n8706), .Z(n8457) );
  NAND U9581 ( .A(n8456), .B(n8457), .Z(n8459) );
  AND U9582 ( .A(\stack[1][6] ), .B(o[43]), .Z(n12479) );
  NAND U9583 ( .A(n12479), .B(n12478), .Z(n8458) );
  AND U9584 ( .A(n8459), .B(n8458), .Z(n8711) );
  NAND U9585 ( .A(n8710), .B(n8711), .Z(n8713) );
  NAND U9586 ( .A(n8461), .B(n8460), .Z(n8465) );
  NAND U9587 ( .A(n8463), .B(n8462), .Z(n8464) );
  AND U9588 ( .A(n8465), .B(n8464), .Z(n8714) );
  NAND U9589 ( .A(\stack[1][8] ), .B(o[42]), .Z(n8715) );
  NAND U9590 ( .A(n8467), .B(n8466), .Z(n8471) );
  NAND U9591 ( .A(n8469), .B(n8468), .Z(n8470) );
  NAND U9592 ( .A(n8471), .B(n8470), .Z(n8721) );
  AND U9593 ( .A(\stack[1][10] ), .B(o[40]), .Z(n8720) );
  NAND U9594 ( .A(n8473), .B(n8472), .Z(n8477) );
  NAND U9595 ( .A(n8475), .B(n8474), .Z(n8476) );
  NAND U9596 ( .A(n8477), .B(n8476), .Z(n8727) );
  AND U9597 ( .A(\stack[1][12] ), .B(o[38]), .Z(n8726) );
  NAND U9598 ( .A(n8479), .B(n8478), .Z(n8483) );
  NAND U9599 ( .A(n8481), .B(n8480), .Z(n8482) );
  NAND U9600 ( .A(n8483), .B(n8482), .Z(n8733) );
  AND U9601 ( .A(\stack[1][14] ), .B(o[36]), .Z(n8732) );
  NAND U9602 ( .A(n8485), .B(n8484), .Z(n8489) );
  NAND U9603 ( .A(n8487), .B(n8486), .Z(n8488) );
  NAND U9604 ( .A(n8489), .B(n8488), .Z(n8739) );
  AND U9605 ( .A(\stack[1][16] ), .B(o[34]), .Z(n8738) );
  NAND U9606 ( .A(n8491), .B(n8490), .Z(n8495) );
  NAND U9607 ( .A(n8493), .B(n8492), .Z(n8494) );
  AND U9608 ( .A(n8495), .B(n8494), .Z(n8745) );
  NAND U9609 ( .A(\stack[1][18] ), .B(o[32]), .Z(n8744) );
  XOR U9610 ( .A(n8745), .B(n8744), .Z(n8746) );
  NAND U9611 ( .A(n8497), .B(n8496), .Z(n8501) );
  NAND U9612 ( .A(n8499), .B(n8498), .Z(n8500) );
  NAND U9613 ( .A(n8501), .B(n8500), .Z(n8750) );
  AND U9614 ( .A(\stack[1][20] ), .B(o[30]), .Z(n8751) );
  XOR U9615 ( .A(n8750), .B(n8751), .Z(n8753) );
  NAND U9616 ( .A(n8503), .B(n8502), .Z(n8507) );
  NAND U9617 ( .A(n8505), .B(n8504), .Z(n8506) );
  NAND U9618 ( .A(n8507), .B(n8506), .Z(n8756) );
  AND U9619 ( .A(\stack[1][22] ), .B(o[28]), .Z(n8757) );
  XOR U9620 ( .A(n8756), .B(n8757), .Z(n8759) );
  NAND U9621 ( .A(n8509), .B(n8508), .Z(n8513) );
  NAND U9622 ( .A(n8511), .B(n8510), .Z(n8512) );
  NAND U9623 ( .A(n8513), .B(n8512), .Z(n8762) );
  AND U9624 ( .A(\stack[1][24] ), .B(o[26]), .Z(n8763) );
  XOR U9625 ( .A(n8762), .B(n8763), .Z(n8765) );
  AND U9626 ( .A(\stack[1][25] ), .B(o[25]), .Z(n16368) );
  NAND U9627 ( .A(n8515), .B(n8514), .Z(n8519) );
  NAND U9628 ( .A(n8517), .B(n8516), .Z(n8518) );
  NAND U9629 ( .A(n8519), .B(n8518), .Z(n8768) );
  AND U9630 ( .A(o[24]), .B(\stack[1][26] ), .Z(n8769) );
  XOR U9631 ( .A(n8768), .B(n8769), .Z(n8771) );
  NAND U9632 ( .A(n8521), .B(n8520), .Z(n8525) );
  NAND U9633 ( .A(n8523), .B(n8522), .Z(n8524) );
  NAND U9634 ( .A(n8525), .B(n8524), .Z(n8774) );
  AND U9635 ( .A(o[22]), .B(\stack[1][28] ), .Z(n8775) );
  XOR U9636 ( .A(n8774), .B(n8775), .Z(n8777) );
  NAND U9637 ( .A(n8527), .B(n8526), .Z(n8531) );
  NAND U9638 ( .A(n8529), .B(n8528), .Z(n8530) );
  NAND U9639 ( .A(n8531), .B(n8530), .Z(n8786) );
  AND U9640 ( .A(o[20]), .B(\stack[1][30] ), .Z(n8787) );
  XOR U9641 ( .A(n8786), .B(n8787), .Z(n8789) );
  NAND U9642 ( .A(n8533), .B(n8532), .Z(n8537) );
  NAND U9643 ( .A(n8535), .B(n8534), .Z(n8536) );
  NAND U9644 ( .A(n8537), .B(n8536), .Z(n8792) );
  AND U9645 ( .A(o[18]), .B(\stack[1][32] ), .Z(n8793) );
  XOR U9646 ( .A(n8792), .B(n8793), .Z(n8795) );
  NAND U9647 ( .A(n8539), .B(n8538), .Z(n8543) );
  NAND U9648 ( .A(n8541), .B(n8540), .Z(n8542) );
  NAND U9649 ( .A(n8543), .B(n8542), .Z(n8804) );
  AND U9650 ( .A(o[16]), .B(\stack[1][34] ), .Z(n8805) );
  XOR U9651 ( .A(n8804), .B(n8805), .Z(n8807) );
  NAND U9652 ( .A(n8545), .B(n8544), .Z(n8549) );
  NAND U9653 ( .A(n8547), .B(n8546), .Z(n8548) );
  NAND U9654 ( .A(n8549), .B(n8548), .Z(n8892) );
  AND U9655 ( .A(o[14]), .B(\stack[1][36] ), .Z(n8886) );
  NAND U9656 ( .A(o[12]), .B(\stack[1][38] ), .Z(n8882) );
  NAND U9657 ( .A(n8551), .B(n8550), .Z(n8555) );
  NANDN U9658 ( .A(n8553), .B(n8552), .Z(n8554) );
  AND U9659 ( .A(n8555), .B(n8554), .Z(n8822) );
  NAND U9660 ( .A(o[9]), .B(\stack[1][41] ), .Z(n8830) );
  NAND U9661 ( .A(n8557), .B(n8556), .Z(n8561) );
  NAND U9662 ( .A(n8559), .B(n8558), .Z(n8560) );
  NAND U9663 ( .A(n8561), .B(n8560), .Z(n8870) );
  NAND U9664 ( .A(o[6]), .B(\stack[1][44] ), .Z(n8836) );
  NAND U9665 ( .A(n8563), .B(n8562), .Z(n8567) );
  NAND U9666 ( .A(n8565), .B(n8564), .Z(n8566) );
  NAND U9667 ( .A(n8567), .B(n8566), .Z(n8862) );
  AND U9668 ( .A(o[4]), .B(\stack[1][46] ), .Z(n8843) );
  NANDN U9669 ( .A(n8568), .B(n8846), .Z(n8572) );
  NANDN U9670 ( .A(n8570), .B(n8569), .Z(n8571) );
  NAND U9671 ( .A(n8572), .B(n8571), .Z(n8856) );
  AND U9672 ( .A(o[3]), .B(\stack[1][47] ), .Z(n8857) );
  XOR U9673 ( .A(n8856), .B(n8857), .Z(n8858) );
  AND U9674 ( .A(o[2]), .B(\stack[1][48] ), .Z(n8847) );
  AND U9675 ( .A(n8573), .B(n8575), .Z(n8574) );
  AND U9676 ( .A(o[1]), .B(\stack[1][50] ), .Z(n8853) );
  NAND U9677 ( .A(n8851), .B(n8853), .Z(n9089) );
  XOR U9678 ( .A(n8574), .B(n9089), .Z(n8577) );
  AND U9679 ( .A(o[0]), .B(\stack[1][50] ), .Z(n9094) );
  OR U9680 ( .A(n8575), .B(n9094), .Z(n8576) );
  NAND U9681 ( .A(n8577), .B(n8576), .Z(n8848) );
  XNOR U9682 ( .A(n8847), .B(n8848), .Z(n8859) );
  NAND U9683 ( .A(n8579), .B(n8578), .Z(n8583) );
  NAND U9684 ( .A(n8581), .B(n8580), .Z(n8582) );
  NAND U9685 ( .A(n8583), .B(n8582), .Z(n8840) );
  XOR U9686 ( .A(n8841), .B(n8840), .Z(n8842) );
  XOR U9687 ( .A(n8843), .B(n8842), .Z(n8863) );
  XOR U9688 ( .A(n8862), .B(n8863), .Z(n8865) );
  AND U9689 ( .A(o[5]), .B(\stack[1][45] ), .Z(n8864) );
  XNOR U9690 ( .A(n8865), .B(n8864), .Z(n8835) );
  NAND U9691 ( .A(n8585), .B(n8584), .Z(n8589) );
  NAND U9692 ( .A(n8587), .B(n8586), .Z(n8588) );
  AND U9693 ( .A(n8589), .B(n8588), .Z(n8834) );
  XNOR U9694 ( .A(n8836), .B(n8837), .Z(n8869) );
  AND U9695 ( .A(o[7]), .B(\stack[1][43] ), .Z(n8868) );
  XOR U9696 ( .A(n8870), .B(n8871), .Z(n8877) );
  AND U9697 ( .A(o[8]), .B(\stack[1][42] ), .Z(n8875) );
  NAND U9698 ( .A(n8591), .B(n8590), .Z(n8595) );
  NAND U9699 ( .A(n8593), .B(n8592), .Z(n8594) );
  NAND U9700 ( .A(n8595), .B(n8594), .Z(n8874) );
  XOR U9701 ( .A(n8875), .B(n8874), .Z(n8876) );
  XNOR U9702 ( .A(n8877), .B(n8876), .Z(n8829) );
  NAND U9703 ( .A(n8597), .B(n8596), .Z(n8601) );
  NAND U9704 ( .A(n8599), .B(n8598), .Z(n8600) );
  AND U9705 ( .A(n8601), .B(n8600), .Z(n8828) );
  XNOR U9706 ( .A(n8830), .B(n8831), .Z(n8823) );
  AND U9707 ( .A(o[10]), .B(\stack[1][40] ), .Z(n8824) );
  XOR U9708 ( .A(n8825), .B(n8824), .Z(n8819) );
  AND U9709 ( .A(o[11]), .B(\stack[1][39] ), .Z(n8817) );
  NAND U9710 ( .A(n8603), .B(n8602), .Z(n8607) );
  NAND U9711 ( .A(n8605), .B(n8604), .Z(n8606) );
  NAND U9712 ( .A(n8607), .B(n8606), .Z(n8816) );
  XOR U9713 ( .A(n8817), .B(n8816), .Z(n8818) );
  XNOR U9714 ( .A(n8819), .B(n8818), .Z(n8881) );
  NAND U9715 ( .A(n8609), .B(n8608), .Z(n8613) );
  NANDN U9716 ( .A(n8611), .B(n8610), .Z(n8612) );
  NAND U9717 ( .A(n8613), .B(n8612), .Z(n8880) );
  XNOR U9718 ( .A(n8882), .B(n8883), .Z(n8813) );
  AND U9719 ( .A(o[13]), .B(\stack[1][37] ), .Z(n8811) );
  NAND U9720 ( .A(n8615), .B(n8614), .Z(n8619) );
  NAND U9721 ( .A(n8617), .B(n8616), .Z(n8618) );
  NAND U9722 ( .A(n8619), .B(n8618), .Z(n8810) );
  XOR U9723 ( .A(n8811), .B(n8810), .Z(n8812) );
  XNOR U9724 ( .A(n8886), .B(n8887), .Z(n8889) );
  NAND U9725 ( .A(n8621), .B(n8620), .Z(n8625) );
  NANDN U9726 ( .A(n8623), .B(n8622), .Z(n8624) );
  NAND U9727 ( .A(n8625), .B(n8624), .Z(n8888) );
  XOR U9728 ( .A(n8889), .B(n8888), .Z(n8893) );
  XOR U9729 ( .A(n8892), .B(n8893), .Z(n8895) );
  AND U9730 ( .A(o[15]), .B(\stack[1][35] ), .Z(n8894) );
  XOR U9731 ( .A(n8895), .B(n8894), .Z(n8806) );
  XOR U9732 ( .A(n8807), .B(n8806), .Z(n8799) );
  NAND U9733 ( .A(n8627), .B(n8626), .Z(n8631) );
  NAND U9734 ( .A(n8629), .B(n8628), .Z(n8630) );
  NAND U9735 ( .A(n8631), .B(n8630), .Z(n8798) );
  XOR U9736 ( .A(n8799), .B(n8798), .Z(n8801) );
  AND U9737 ( .A(o[17]), .B(\stack[1][33] ), .Z(n8800) );
  XOR U9738 ( .A(n8801), .B(n8800), .Z(n8794) );
  XOR U9739 ( .A(n8795), .B(n8794), .Z(n8899) );
  NAND U9740 ( .A(n8633), .B(n8632), .Z(n8637) );
  NAND U9741 ( .A(n8635), .B(n8634), .Z(n8636) );
  NAND U9742 ( .A(n8637), .B(n8636), .Z(n8898) );
  XOR U9743 ( .A(n8899), .B(n8898), .Z(n8901) );
  AND U9744 ( .A(o[19]), .B(\stack[1][31] ), .Z(n8900) );
  XOR U9745 ( .A(n8901), .B(n8900), .Z(n8788) );
  XOR U9746 ( .A(n8789), .B(n8788), .Z(n8781) );
  NAND U9747 ( .A(n8639), .B(n8638), .Z(n8643) );
  NAND U9748 ( .A(n8641), .B(n8640), .Z(n8642) );
  NAND U9749 ( .A(n8643), .B(n8642), .Z(n8780) );
  XOR U9750 ( .A(n8781), .B(n8780), .Z(n8783) );
  AND U9751 ( .A(o[21]), .B(\stack[1][29] ), .Z(n8782) );
  XOR U9752 ( .A(n8783), .B(n8782), .Z(n8776) );
  XOR U9753 ( .A(n8777), .B(n8776), .Z(n8905) );
  NAND U9754 ( .A(n8645), .B(n8644), .Z(n8649) );
  NAND U9755 ( .A(n8647), .B(n8646), .Z(n8648) );
  NAND U9756 ( .A(n8649), .B(n8648), .Z(n8904) );
  XOR U9757 ( .A(n8905), .B(n8904), .Z(n8907) );
  AND U9758 ( .A(o[23]), .B(\stack[1][27] ), .Z(n8906) );
  XOR U9759 ( .A(n8907), .B(n8906), .Z(n8770) );
  XOR U9760 ( .A(n8771), .B(n8770), .Z(n8911) );
  NAND U9761 ( .A(n8651), .B(n8650), .Z(n8655) );
  NAND U9762 ( .A(n8653), .B(n8652), .Z(n8654) );
  NAND U9763 ( .A(n8655), .B(n8654), .Z(n8910) );
  XOR U9764 ( .A(n8911), .B(n8910), .Z(n8912) );
  XOR U9765 ( .A(n16368), .B(n8912), .Z(n8764) );
  XOR U9766 ( .A(n8765), .B(n8764), .Z(n8916) );
  NAND U9767 ( .A(n8657), .B(n8656), .Z(n8661) );
  NAND U9768 ( .A(n8659), .B(n8658), .Z(n8660) );
  NAND U9769 ( .A(n8661), .B(n8660), .Z(n8915) );
  XOR U9770 ( .A(n8916), .B(n8915), .Z(n8918) );
  AND U9771 ( .A(\stack[1][23] ), .B(o[27]), .Z(n8917) );
  XOR U9772 ( .A(n8918), .B(n8917), .Z(n8758) );
  XOR U9773 ( .A(n8759), .B(n8758), .Z(n8922) );
  NAND U9774 ( .A(n8663), .B(n8662), .Z(n8667) );
  NAND U9775 ( .A(n8665), .B(n8664), .Z(n8666) );
  NAND U9776 ( .A(n8667), .B(n8666), .Z(n8921) );
  XOR U9777 ( .A(n8922), .B(n8921), .Z(n8924) );
  AND U9778 ( .A(\stack[1][21] ), .B(o[29]), .Z(n8923) );
  XOR U9779 ( .A(n8924), .B(n8923), .Z(n8752) );
  XOR U9780 ( .A(n8753), .B(n8752), .Z(n8928) );
  NAND U9781 ( .A(n8669), .B(n8668), .Z(n8673) );
  NAND U9782 ( .A(n8671), .B(n8670), .Z(n8672) );
  NAND U9783 ( .A(n8673), .B(n8672), .Z(n8927) );
  XOR U9784 ( .A(n8928), .B(n8927), .Z(n8930) );
  AND U9785 ( .A(\stack[1][19] ), .B(o[31]), .Z(n8929) );
  XNOR U9786 ( .A(n8930), .B(n8929), .Z(n8747) );
  NAND U9787 ( .A(n8675), .B(n8674), .Z(n8679) );
  NAND U9788 ( .A(n8677), .B(n8676), .Z(n8678) );
  NAND U9789 ( .A(n8679), .B(n8678), .Z(n8933) );
  AND U9790 ( .A(\stack[1][17] ), .B(o[33]), .Z(n8935) );
  XOR U9791 ( .A(n8936), .B(n8935), .Z(n8740) );
  XOR U9792 ( .A(n8741), .B(n8740), .Z(n8939) );
  NAND U9793 ( .A(n8681), .B(n8680), .Z(n8685) );
  NAND U9794 ( .A(n8683), .B(n8682), .Z(n8684) );
  NAND U9795 ( .A(n8685), .B(n8684), .Z(n8940) );
  AND U9796 ( .A(\stack[1][15] ), .B(o[35]), .Z(n8942) );
  XOR U9797 ( .A(n8735), .B(n8734), .Z(n8945) );
  NAND U9798 ( .A(n8687), .B(n8686), .Z(n8691) );
  NAND U9799 ( .A(n8689), .B(n8688), .Z(n8690) );
  NAND U9800 ( .A(n8691), .B(n8690), .Z(n8946) );
  AND U9801 ( .A(\stack[1][13] ), .B(o[37]), .Z(n8948) );
  XOR U9802 ( .A(n8729), .B(n8728), .Z(n8951) );
  NAND U9803 ( .A(n8693), .B(n8692), .Z(n8697) );
  NAND U9804 ( .A(n8695), .B(n8694), .Z(n8696) );
  NAND U9805 ( .A(n8697), .B(n8696), .Z(n8952) );
  AND U9806 ( .A(\stack[1][11] ), .B(o[39]), .Z(n8954) );
  XOR U9807 ( .A(n8723), .B(n8722), .Z(n8957) );
  NAND U9808 ( .A(n8699), .B(n8698), .Z(n8703) );
  NAND U9809 ( .A(n8701), .B(n8700), .Z(n8702) );
  NAND U9810 ( .A(n8703), .B(n8702), .Z(n8958) );
  AND U9811 ( .A(\stack[1][9] ), .B(o[41]), .Z(n8959) );
  XNOR U9812 ( .A(n8960), .B(n8959), .Z(n8716) );
  XNOR U9813 ( .A(n8717), .B(n8716), .Z(n8964) );
  NAND U9814 ( .A(n8705), .B(n8704), .Z(n8709) );
  NAND U9815 ( .A(n8707), .B(n8706), .Z(n8708) );
  NAND U9816 ( .A(n8709), .B(n8708), .Z(n8963) );
  AND U9817 ( .A(\stack[1][7] ), .B(o[43]), .Z(n8965) );
  XNOR U9818 ( .A(n8966), .B(n8965), .Z(n12223) );
  NAND U9819 ( .A(n12223), .B(n12224), .Z(n8712) );
  AND U9820 ( .A(n8713), .B(n8712), .Z(n8970) );
  AND U9821 ( .A(\stack[1][8] ), .B(o[43]), .Z(n8984) );
  NAND U9822 ( .A(n8715), .B(n8714), .Z(n8719) );
  NAND U9823 ( .A(n8717), .B(n8716), .Z(n8718) );
  AND U9824 ( .A(n8719), .B(n8718), .Z(n8982) );
  NAND U9825 ( .A(n8721), .B(n8720), .Z(n8725) );
  NAND U9826 ( .A(n8723), .B(n8722), .Z(n8724) );
  NAND U9827 ( .A(n8725), .B(n8724), .Z(n9226) );
  NAND U9828 ( .A(n8727), .B(n8726), .Z(n8731) );
  NAND U9829 ( .A(n8729), .B(n8728), .Z(n8730) );
  NAND U9830 ( .A(n8731), .B(n8730), .Z(n8988) );
  NAND U9831 ( .A(n8733), .B(n8732), .Z(n8737) );
  NAND U9832 ( .A(n8735), .B(n8734), .Z(n8736) );
  NAND U9833 ( .A(n8737), .B(n8736), .Z(n9208) );
  AND U9834 ( .A(\stack[1][16] ), .B(o[35]), .Z(n9197) );
  NAND U9835 ( .A(n8739), .B(n8738), .Z(n8743) );
  NAND U9836 ( .A(n8741), .B(n8740), .Z(n8742) );
  NAND U9837 ( .A(n8743), .B(n8742), .Z(n9195) );
  NAND U9838 ( .A(n8745), .B(n8744), .Z(n8749) );
  NAND U9839 ( .A(n8747), .B(n8746), .Z(n8748) );
  AND U9840 ( .A(n8749), .B(n8748), .Z(n9000) );
  AND U9841 ( .A(\stack[1][20] ), .B(o[31]), .Z(n9185) );
  NAND U9842 ( .A(n8751), .B(n8750), .Z(n8755) );
  NAND U9843 ( .A(n8753), .B(n8752), .Z(n8754) );
  NAND U9844 ( .A(n8755), .B(n8754), .Z(n9183) );
  AND U9845 ( .A(\stack[1][22] ), .B(o[29]), .Z(n9007) );
  NAND U9846 ( .A(n8757), .B(n8756), .Z(n8761) );
  NAND U9847 ( .A(n8759), .B(n8758), .Z(n8760) );
  NAND U9848 ( .A(n8761), .B(n8760), .Z(n9005) );
  NAND U9849 ( .A(n8763), .B(n8762), .Z(n8767) );
  NAND U9850 ( .A(n8765), .B(n8764), .Z(n8766) );
  NAND U9851 ( .A(n8767), .B(n8766), .Z(n9165) );
  AND U9852 ( .A(\stack[1][26] ), .B(o[25]), .Z(n9013) );
  NAND U9853 ( .A(n8769), .B(n8768), .Z(n8773) );
  NAND U9854 ( .A(n8771), .B(n8770), .Z(n8772) );
  NAND U9855 ( .A(n8773), .B(n8772), .Z(n9011) );
  AND U9856 ( .A(o[23]), .B(\stack[1][28] ), .Z(n9019) );
  NAND U9857 ( .A(n8775), .B(n8774), .Z(n8779) );
  NAND U9858 ( .A(n8777), .B(n8776), .Z(n8778) );
  NAND U9859 ( .A(n8779), .B(n8778), .Z(n9017) );
  AND U9860 ( .A(o[22]), .B(\stack[1][29] ), .Z(n9148) );
  NAND U9861 ( .A(n8781), .B(n8780), .Z(n8785) );
  NAND U9862 ( .A(n8783), .B(n8782), .Z(n8784) );
  NAND U9863 ( .A(n8785), .B(n8784), .Z(n9147) );
  XOR U9864 ( .A(n9148), .B(n9147), .Z(n9150) );
  AND U9865 ( .A(o[21]), .B(\stack[1][30] ), .Z(n9025) );
  NAND U9866 ( .A(n8787), .B(n8786), .Z(n8791) );
  NAND U9867 ( .A(n8789), .B(n8788), .Z(n8790) );
  NAND U9868 ( .A(n8791), .B(n8790), .Z(n9023) );
  AND U9869 ( .A(o[19]), .B(\stack[1][32] ), .Z(n9037) );
  NAND U9870 ( .A(n8793), .B(n8792), .Z(n8797) );
  NAND U9871 ( .A(n8795), .B(n8794), .Z(n8796) );
  NAND U9872 ( .A(n8797), .B(n8796), .Z(n9035) );
  AND U9873 ( .A(o[18]), .B(\stack[1][33] ), .Z(n9142) );
  NAND U9874 ( .A(n8799), .B(n8798), .Z(n8803) );
  NAND U9875 ( .A(n8801), .B(n8800), .Z(n8802) );
  NAND U9876 ( .A(n8803), .B(n8802), .Z(n9141) );
  XOR U9877 ( .A(n9142), .B(n9141), .Z(n9144) );
  AND U9878 ( .A(o[17]), .B(\stack[1][34] ), .Z(n9043) );
  NAND U9879 ( .A(n8805), .B(n8804), .Z(n8809) );
  NAND U9880 ( .A(n8807), .B(n8806), .Z(n8808) );
  NAND U9881 ( .A(n8809), .B(n8808), .Z(n9041) );
  AND U9882 ( .A(o[16]), .B(\stack[1][35] ), .Z(n9138) );
  NAND U9883 ( .A(n8811), .B(n8810), .Z(n8815) );
  NAND U9884 ( .A(n8813), .B(n8812), .Z(n8814) );
  NAND U9885 ( .A(n8815), .B(n8814), .Z(n9055) );
  AND U9886 ( .A(o[13]), .B(\stack[1][38] ), .Z(n9132) );
  AND U9887 ( .A(o[12]), .B(\stack[1][39] ), .Z(n9061) );
  NAND U9888 ( .A(n8817), .B(n8816), .Z(n8821) );
  NAND U9889 ( .A(n8819), .B(n8818), .Z(n8820) );
  NAND U9890 ( .A(n8821), .B(n8820), .Z(n9059) );
  NAND U9891 ( .A(n8823), .B(n8822), .Z(n8827) );
  NAND U9892 ( .A(n8825), .B(n8824), .Z(n8826) );
  AND U9893 ( .A(n8827), .B(n8826), .Z(n9065) );
  NAND U9894 ( .A(n8829), .B(n8828), .Z(n8833) );
  NAND U9895 ( .A(n8831), .B(n8830), .Z(n8832) );
  AND U9896 ( .A(n8833), .B(n8832), .Z(n9123) );
  NAND U9897 ( .A(o[9]), .B(\stack[1][42] ), .Z(n9073) );
  NAND U9898 ( .A(n8835), .B(n8834), .Z(n8839) );
  NAND U9899 ( .A(n8837), .B(n8836), .Z(n8838) );
  AND U9900 ( .A(n8839), .B(n8838), .Z(n9114) );
  AND U9901 ( .A(o[6]), .B(\stack[1][45] ), .Z(n9080) );
  NAND U9902 ( .A(n8841), .B(n8840), .Z(n8845) );
  NAND U9903 ( .A(n8843), .B(n8842), .Z(n8844) );
  NAND U9904 ( .A(n8845), .B(n8844), .Z(n9105) );
  NANDN U9905 ( .A(n8846), .B(n9089), .Z(n8850) );
  NANDN U9906 ( .A(n8848), .B(n8847), .Z(n8849) );
  NAND U9907 ( .A(n8850), .B(n8849), .Z(n9099) );
  AND U9908 ( .A(o[2]), .B(\stack[1][49] ), .Z(n9090) );
  AND U9909 ( .A(n8851), .B(n8853), .Z(n8852) );
  AND U9910 ( .A(o[1]), .B(\stack[1][51] ), .Z(n9096) );
  NAND U9911 ( .A(n9094), .B(n9096), .Z(n9364) );
  XOR U9912 ( .A(n8852), .B(n9364), .Z(n8855) );
  AND U9913 ( .A(o[0]), .B(\stack[1][51] ), .Z(n9369) );
  OR U9914 ( .A(n8853), .B(n9369), .Z(n8854) );
  NAND U9915 ( .A(n8855), .B(n8854), .Z(n9091) );
  XNOR U9916 ( .A(n9090), .B(n9091), .Z(n9100) );
  XOR U9917 ( .A(n9099), .B(n9100), .Z(n9102) );
  AND U9918 ( .A(o[3]), .B(\stack[1][48] ), .Z(n9101) );
  XOR U9919 ( .A(n9102), .B(n9101), .Z(n9084) );
  NAND U9920 ( .A(n8857), .B(n8856), .Z(n8861) );
  NAND U9921 ( .A(n8859), .B(n8858), .Z(n8860) );
  NAND U9922 ( .A(n8861), .B(n8860), .Z(n9083) );
  XOR U9923 ( .A(n9084), .B(n9083), .Z(n9086) );
  AND U9924 ( .A(o[4]), .B(\stack[1][47] ), .Z(n9085) );
  XOR U9925 ( .A(n9086), .B(n9085), .Z(n9106) );
  XOR U9926 ( .A(n9105), .B(n9106), .Z(n9108) );
  AND U9927 ( .A(o[5]), .B(\stack[1][46] ), .Z(n9107) );
  XOR U9928 ( .A(n9108), .B(n9107), .Z(n9078) );
  NAND U9929 ( .A(n8863), .B(n8862), .Z(n8867) );
  NAND U9930 ( .A(n8865), .B(n8864), .Z(n8866) );
  NAND U9931 ( .A(n8867), .B(n8866), .Z(n9077) );
  XOR U9932 ( .A(n9078), .B(n9077), .Z(n9079) );
  XOR U9933 ( .A(n9080), .B(n9079), .Z(n9112) );
  AND U9934 ( .A(o[7]), .B(\stack[1][44] ), .Z(n9111) );
  XOR U9935 ( .A(n9112), .B(n9111), .Z(n9113) );
  XOR U9936 ( .A(n9114), .B(n9113), .Z(n9120) );
  AND U9937 ( .A(o[8]), .B(\stack[1][43] ), .Z(n9118) );
  NAND U9938 ( .A(n8869), .B(n8868), .Z(n8873) );
  NAND U9939 ( .A(n8871), .B(n8870), .Z(n8872) );
  NAND U9940 ( .A(n8873), .B(n8872), .Z(n9117) );
  XOR U9941 ( .A(n9118), .B(n9117), .Z(n9119) );
  XNOR U9942 ( .A(n9120), .B(n9119), .Z(n9072) );
  NAND U9943 ( .A(n8875), .B(n8874), .Z(n8879) );
  NAND U9944 ( .A(n8877), .B(n8876), .Z(n8878) );
  AND U9945 ( .A(n8879), .B(n8878), .Z(n9071) );
  XNOR U9946 ( .A(n9073), .B(n9074), .Z(n9124) );
  AND U9947 ( .A(o[10]), .B(\stack[1][41] ), .Z(n9125) );
  XNOR U9948 ( .A(n9126), .B(n9125), .Z(n9066) );
  NAND U9949 ( .A(o[11]), .B(\stack[1][40] ), .Z(n9067) );
  XNOR U9950 ( .A(n9068), .B(n9067), .Z(n9060) );
  XNOR U9951 ( .A(n9061), .B(n9062), .Z(n9130) );
  NAND U9952 ( .A(n8881), .B(n8880), .Z(n8885) );
  NAND U9953 ( .A(n8883), .B(n8882), .Z(n8884) );
  AND U9954 ( .A(n8885), .B(n8884), .Z(n9129) );
  XOR U9955 ( .A(n9130), .B(n9129), .Z(n9131) );
  XOR U9956 ( .A(n9132), .B(n9131), .Z(n9054) );
  AND U9957 ( .A(o[14]), .B(\stack[1][37] ), .Z(n9053) );
  XOR U9958 ( .A(n9054), .B(n9053), .Z(n9056) );
  XOR U9959 ( .A(n9055), .B(n9056), .Z(n9049) );
  NANDN U9960 ( .A(n8887), .B(n8886), .Z(n8891) );
  NAND U9961 ( .A(n8889), .B(n8888), .Z(n8890) );
  NAND U9962 ( .A(n8891), .B(n8890), .Z(n9047) );
  AND U9963 ( .A(o[15]), .B(\stack[1][36] ), .Z(n9048) );
  XOR U9964 ( .A(n9047), .B(n9048), .Z(n9050) );
  NAND U9965 ( .A(n8893), .B(n8892), .Z(n8897) );
  NAND U9966 ( .A(n8895), .B(n8894), .Z(n8896) );
  NAND U9967 ( .A(n8897), .B(n8896), .Z(n9135) );
  XOR U9968 ( .A(n9136), .B(n9135), .Z(n9137) );
  XOR U9969 ( .A(n9138), .B(n9137), .Z(n9042) );
  XOR U9970 ( .A(n9041), .B(n9042), .Z(n9044) );
  XOR U9971 ( .A(n9144), .B(n9143), .Z(n9036) );
  XOR U9972 ( .A(n9035), .B(n9036), .Z(n9038) );
  AND U9973 ( .A(o[20]), .B(\stack[1][31] ), .Z(n9030) );
  NAND U9974 ( .A(n8899), .B(n8898), .Z(n8903) );
  NAND U9975 ( .A(n8901), .B(n8900), .Z(n8902) );
  NAND U9976 ( .A(n8903), .B(n8902), .Z(n9029) );
  XOR U9977 ( .A(n9030), .B(n9029), .Z(n9031) );
  XOR U9978 ( .A(n9032), .B(n9031), .Z(n9024) );
  XOR U9979 ( .A(n9023), .B(n9024), .Z(n9026) );
  XOR U9980 ( .A(n9150), .B(n9149), .Z(n9018) );
  XOR U9981 ( .A(n9017), .B(n9018), .Z(n9020) );
  AND U9982 ( .A(o[24]), .B(\stack[1][27] ), .Z(n9154) );
  NAND U9983 ( .A(n8905), .B(n8904), .Z(n8909) );
  NAND U9984 ( .A(n8907), .B(n8906), .Z(n8908) );
  NAND U9985 ( .A(n8909), .B(n8908), .Z(n9153) );
  XOR U9986 ( .A(n9154), .B(n9153), .Z(n9155) );
  XOR U9987 ( .A(n9156), .B(n9155), .Z(n9012) );
  XOR U9988 ( .A(n9011), .B(n9012), .Z(n9014) );
  AND U9989 ( .A(\stack[1][25] ), .B(o[26]), .Z(n9160) );
  NAND U9990 ( .A(n8911), .B(n8910), .Z(n8914) );
  NAND U9991 ( .A(n16368), .B(n8912), .Z(n8913) );
  NAND U9992 ( .A(n8914), .B(n8913), .Z(n9159) );
  XOR U9993 ( .A(n9160), .B(n9159), .Z(n9161) );
  XOR U9994 ( .A(n9162), .B(n9161), .Z(n9166) );
  XOR U9995 ( .A(n9165), .B(n9166), .Z(n9168) );
  AND U9996 ( .A(\stack[1][24] ), .B(o[27]), .Z(n9167) );
  XOR U9997 ( .A(n9168), .B(n9167), .Z(n9174) );
  AND U9998 ( .A(\stack[1][23] ), .B(o[28]), .Z(n9172) );
  NAND U9999 ( .A(n8916), .B(n8915), .Z(n8920) );
  NAND U10000 ( .A(n8918), .B(n8917), .Z(n8919) );
  NAND U10001 ( .A(n8920), .B(n8919), .Z(n9171) );
  XOR U10002 ( .A(n9172), .B(n9171), .Z(n9173) );
  XOR U10003 ( .A(n9174), .B(n9173), .Z(n9006) );
  XOR U10004 ( .A(n9005), .B(n9006), .Z(n9008) );
  AND U10005 ( .A(\stack[1][21] ), .B(o[30]), .Z(n9178) );
  NAND U10006 ( .A(n8922), .B(n8921), .Z(n8926) );
  NAND U10007 ( .A(n8924), .B(n8923), .Z(n8925) );
  NAND U10008 ( .A(n8926), .B(n8925), .Z(n9177) );
  XOR U10009 ( .A(n9178), .B(n9177), .Z(n9179) );
  XOR U10010 ( .A(n9180), .B(n9179), .Z(n9184) );
  XOR U10011 ( .A(n9183), .B(n9184), .Z(n9186) );
  AND U10012 ( .A(\stack[1][19] ), .B(o[32]), .Z(n9190) );
  NAND U10013 ( .A(n8928), .B(n8927), .Z(n8932) );
  NAND U10014 ( .A(n8930), .B(n8929), .Z(n8931) );
  NAND U10015 ( .A(n8932), .B(n8931), .Z(n9189) );
  XOR U10016 ( .A(n9190), .B(n9189), .Z(n9191) );
  XOR U10017 ( .A(n9192), .B(n9191), .Z(n8999) );
  XOR U10018 ( .A(n9000), .B(n8999), .Z(n9002) );
  AND U10019 ( .A(\stack[1][18] ), .B(o[33]), .Z(n9001) );
  XOR U10020 ( .A(n9002), .B(n9001), .Z(n8996) );
  AND U10021 ( .A(\stack[1][17] ), .B(o[34]), .Z(n8994) );
  NAND U10022 ( .A(n8934), .B(n8933), .Z(n8938) );
  NAND U10023 ( .A(n8936), .B(n8935), .Z(n8937) );
  NAND U10024 ( .A(n8938), .B(n8937), .Z(n8993) );
  XOR U10025 ( .A(n8994), .B(n8993), .Z(n8995) );
  XOR U10026 ( .A(n8996), .B(n8995), .Z(n9196) );
  XOR U10027 ( .A(n9195), .B(n9196), .Z(n9198) );
  AND U10028 ( .A(\stack[1][15] ), .B(o[36]), .Z(n9202) );
  NAND U10029 ( .A(n8940), .B(n8939), .Z(n8944) );
  NAND U10030 ( .A(n8942), .B(n8941), .Z(n8943) );
  NAND U10031 ( .A(n8944), .B(n8943), .Z(n9201) );
  XOR U10032 ( .A(n9202), .B(n9201), .Z(n9203) );
  XOR U10033 ( .A(n9204), .B(n9203), .Z(n9207) );
  AND U10034 ( .A(\stack[1][14] ), .B(o[37]), .Z(n9210) );
  AND U10035 ( .A(\stack[1][13] ), .B(o[38]), .Z(n9213) );
  NAND U10036 ( .A(n8946), .B(n8945), .Z(n8950) );
  NAND U10037 ( .A(n8948), .B(n8947), .Z(n8949) );
  NAND U10038 ( .A(n8950), .B(n8949), .Z(n9214) );
  XOR U10039 ( .A(n9216), .B(n9215), .Z(n8987) );
  AND U10040 ( .A(\stack[1][12] ), .B(o[39]), .Z(n8990) );
  AND U10041 ( .A(\stack[1][11] ), .B(o[40]), .Z(n9219) );
  NAND U10042 ( .A(n8952), .B(n8951), .Z(n8956) );
  NAND U10043 ( .A(n8954), .B(n8953), .Z(n8955) );
  NAND U10044 ( .A(n8956), .B(n8955), .Z(n9220) );
  XOR U10045 ( .A(n9222), .B(n9221), .Z(n9225) );
  AND U10046 ( .A(\stack[1][10] ), .B(o[41]), .Z(n9228) );
  AND U10047 ( .A(\stack[1][9] ), .B(o[42]), .Z(n9231) );
  NAND U10048 ( .A(n8958), .B(n8957), .Z(n8962) );
  NAND U10049 ( .A(n8960), .B(n8959), .Z(n8961) );
  NAND U10050 ( .A(n8962), .B(n8961), .Z(n9232) );
  XOR U10051 ( .A(n9234), .B(n9233), .Z(n8981) );
  XOR U10052 ( .A(n8982), .B(n8981), .Z(n8983) );
  XOR U10053 ( .A(n8984), .B(n8983), .Z(n8978) );
  AND U10054 ( .A(\stack[1][7] ), .B(o[44]), .Z(n8975) );
  NAND U10055 ( .A(n8964), .B(n8963), .Z(n8968) );
  NAND U10056 ( .A(n8966), .B(n8965), .Z(n8967) );
  NAND U10057 ( .A(n8968), .B(n8967), .Z(n8976) );
  XOR U10058 ( .A(n8978), .B(n8977), .Z(n8969) );
  NAND U10059 ( .A(n8970), .B(n8969), .Z(n8972) );
  AND U10060 ( .A(\stack[1][6] ), .B(o[45]), .Z(n12488) );
  XOR U10061 ( .A(n8970), .B(n8969), .Z(n12489) );
  NAND U10062 ( .A(n12488), .B(n12489), .Z(n8971) );
  AND U10063 ( .A(n8972), .B(n8971), .Z(n8974) );
  NAND U10064 ( .A(n8973), .B(n8974), .Z(n9238) );
  NAND U10065 ( .A(n8976), .B(n8975), .Z(n8980) );
  NAND U10066 ( .A(n8978), .B(n8977), .Z(n8979) );
  NAND U10067 ( .A(n8980), .B(n8979), .Z(n9501) );
  NAND U10068 ( .A(n8982), .B(n8981), .Z(n8986) );
  NAND U10069 ( .A(n8984), .B(n8983), .Z(n8985) );
  AND U10070 ( .A(n8986), .B(n8985), .Z(n9239) );
  NAND U10071 ( .A(\stack[1][8] ), .B(o[44]), .Z(n9240) );
  NAND U10072 ( .A(n8988), .B(n8987), .Z(n8992) );
  NAND U10073 ( .A(n8990), .B(n8989), .Z(n8991) );
  AND U10074 ( .A(n8992), .B(n8991), .Z(n9251) );
  NAND U10075 ( .A(\stack[1][12] ), .B(o[40]), .Z(n9252) );
  NAND U10076 ( .A(n8994), .B(n8993), .Z(n8998) );
  NAND U10077 ( .A(n8996), .B(n8995), .Z(n8997) );
  NAND U10078 ( .A(n8998), .B(n8997), .Z(n9471) );
  NAND U10079 ( .A(n9000), .B(n8999), .Z(n9004) );
  NAND U10080 ( .A(n9002), .B(n9001), .Z(n9003) );
  AND U10081 ( .A(n9004), .B(n9003), .Z(n9270) );
  NAND U10082 ( .A(\stack[1][18] ), .B(o[34]), .Z(n9269) );
  XOR U10083 ( .A(n9270), .B(n9269), .Z(n9272) );
  NAND U10084 ( .A(n9006), .B(n9005), .Z(n9010) );
  NAND U10085 ( .A(n9008), .B(n9007), .Z(n9009) );
  NAND U10086 ( .A(n9010), .B(n9009), .Z(n9281) );
  AND U10087 ( .A(\stack[1][22] ), .B(o[30]), .Z(n9282) );
  XOR U10088 ( .A(n9281), .B(n9282), .Z(n9284) );
  AND U10089 ( .A(\stack[1][26] ), .B(o[26]), .Z(n16327) );
  NAND U10090 ( .A(n9012), .B(n9011), .Z(n9016) );
  NAND U10091 ( .A(n9014), .B(n9013), .Z(n9015) );
  NAND U10092 ( .A(n9016), .B(n9015), .Z(n9293) );
  XOR U10093 ( .A(n16327), .B(n9293), .Z(n9295) );
  NAND U10094 ( .A(n9018), .B(n9017), .Z(n9022) );
  NAND U10095 ( .A(n9020), .B(n9019), .Z(n9021) );
  NAND U10096 ( .A(n9022), .B(n9021), .Z(n9298) );
  AND U10097 ( .A(o[24]), .B(\stack[1][28] ), .Z(n9299) );
  XOR U10098 ( .A(n9298), .B(n9299), .Z(n9301) );
  NAND U10099 ( .A(n9024), .B(n9023), .Z(n9028) );
  NAND U10100 ( .A(n9026), .B(n9025), .Z(n9027) );
  NAND U10101 ( .A(n9028), .B(n9027), .Z(n9428) );
  AND U10102 ( .A(o[22]), .B(\stack[1][30] ), .Z(n9429) );
  XOR U10103 ( .A(n9428), .B(n9429), .Z(n9431) );
  NAND U10104 ( .A(n9030), .B(n9029), .Z(n9034) );
  NAND U10105 ( .A(n9032), .B(n9031), .Z(n9033) );
  NAND U10106 ( .A(n9034), .B(n9033), .Z(n9423) );
  NAND U10107 ( .A(n9036), .B(n9035), .Z(n9040) );
  NAND U10108 ( .A(n9038), .B(n9037), .Z(n9039) );
  AND U10109 ( .A(n9040), .B(n9039), .Z(n9305) );
  NAND U10110 ( .A(o[20]), .B(\stack[1][32] ), .Z(n9304) );
  XOR U10111 ( .A(n9305), .B(n9304), .Z(n9307) );
  NAND U10112 ( .A(n9042), .B(n9041), .Z(n9046) );
  NAND U10113 ( .A(n9044), .B(n9043), .Z(n9045) );
  NAND U10114 ( .A(n9046), .B(n9045), .Z(n9310) );
  AND U10115 ( .A(o[18]), .B(\stack[1][34] ), .Z(n9311) );
  XOR U10116 ( .A(n9310), .B(n9311), .Z(n9313) );
  AND U10117 ( .A(o[17]), .B(\stack[1][35] ), .Z(n9413) );
  NAND U10118 ( .A(n9048), .B(n9047), .Z(n9052) );
  NAND U10119 ( .A(n9050), .B(n9049), .Z(n9051) );
  NAND U10120 ( .A(n9052), .B(n9051), .Z(n9316) );
  AND U10121 ( .A(o[16]), .B(\stack[1][36] ), .Z(n9317) );
  XOR U10122 ( .A(n9316), .B(n9317), .Z(n9319) );
  AND U10123 ( .A(o[15]), .B(\stack[1][37] ), .Z(n9407) );
  NAND U10124 ( .A(n9054), .B(n9053), .Z(n9058) );
  NAND U10125 ( .A(n9056), .B(n9055), .Z(n9057) );
  NAND U10126 ( .A(n9058), .B(n9057), .Z(n9404) );
  AND U10127 ( .A(o[14]), .B(\stack[1][38] ), .Z(n9401) );
  NAND U10128 ( .A(n9060), .B(n9059), .Z(n9064) );
  NANDN U10129 ( .A(n9062), .B(n9061), .Z(n9063) );
  NAND U10130 ( .A(n9064), .B(n9063), .Z(n9323) );
  NAND U10131 ( .A(n9066), .B(n9065), .Z(n9070) );
  NAND U10132 ( .A(n9068), .B(n9067), .Z(n9069) );
  NAND U10133 ( .A(n9070), .B(n9069), .Z(n9328) );
  NAND U10134 ( .A(o[11]), .B(\stack[1][41] ), .Z(n9336) );
  NAND U10135 ( .A(n9072), .B(n9071), .Z(n9076) );
  NAND U10136 ( .A(n9074), .B(n9073), .Z(n9075) );
  NAND U10137 ( .A(n9076), .B(n9075), .Z(n9392) );
  NAND U10138 ( .A(o[9]), .B(\stack[1][43] ), .Z(n9342) );
  NAND U10139 ( .A(n9078), .B(n9077), .Z(n9082) );
  NAND U10140 ( .A(n9080), .B(n9079), .Z(n9081) );
  NAND U10141 ( .A(n9082), .B(n9081), .Z(n9348) );
  AND U10142 ( .A(o[6]), .B(\stack[1][46] ), .Z(n9355) );
  NAND U10143 ( .A(n9084), .B(n9083), .Z(n9088) );
  NAND U10144 ( .A(n9086), .B(n9085), .Z(n9087) );
  NAND U10145 ( .A(n9088), .B(n9087), .Z(n9381) );
  NANDN U10146 ( .A(n9089), .B(n9364), .Z(n9093) );
  NANDN U10147 ( .A(n9091), .B(n9090), .Z(n9092) );
  NAND U10148 ( .A(n9093), .B(n9092), .Z(n9374) );
  AND U10149 ( .A(o[2]), .B(\stack[1][50] ), .Z(n9365) );
  AND U10150 ( .A(n9094), .B(n9096), .Z(n9095) );
  AND U10151 ( .A(o[1]), .B(\stack[1][52] ), .Z(n9371) );
  NAND U10152 ( .A(n9369), .B(n9371), .Z(n9614) );
  XOR U10153 ( .A(n9095), .B(n9614), .Z(n9098) );
  AND U10154 ( .A(o[0]), .B(\stack[1][52] ), .Z(n9619) );
  OR U10155 ( .A(n9096), .B(n9619), .Z(n9097) );
  NAND U10156 ( .A(n9098), .B(n9097), .Z(n9366) );
  XNOR U10157 ( .A(n9365), .B(n9366), .Z(n9375) );
  XOR U10158 ( .A(n9374), .B(n9375), .Z(n9377) );
  AND U10159 ( .A(o[3]), .B(\stack[1][49] ), .Z(n9376) );
  XNOR U10160 ( .A(n9377), .B(n9376), .Z(n9359) );
  NAND U10161 ( .A(n9100), .B(n9099), .Z(n9104) );
  NAND U10162 ( .A(n9102), .B(n9101), .Z(n9103) );
  AND U10163 ( .A(n9104), .B(n9103), .Z(n9358) );
  NAND U10164 ( .A(o[4]), .B(\stack[1][48] ), .Z(n9360) );
  XNOR U10165 ( .A(n9361), .B(n9360), .Z(n9380) );
  XOR U10166 ( .A(n9381), .B(n9380), .Z(n9383) );
  AND U10167 ( .A(o[5]), .B(\stack[1][47] ), .Z(n9382) );
  XOR U10168 ( .A(n9383), .B(n9382), .Z(n9353) );
  NAND U10169 ( .A(n9106), .B(n9105), .Z(n9110) );
  NAND U10170 ( .A(n9108), .B(n9107), .Z(n9109) );
  NAND U10171 ( .A(n9110), .B(n9109), .Z(n9352) );
  XOR U10172 ( .A(n9353), .B(n9352), .Z(n9354) );
  XOR U10173 ( .A(n9355), .B(n9354), .Z(n9347) );
  AND U10174 ( .A(o[7]), .B(\stack[1][45] ), .Z(n9346) );
  XOR U10175 ( .A(n9347), .B(n9346), .Z(n9349) );
  XOR U10176 ( .A(n9348), .B(n9349), .Z(n9387) );
  AND U10177 ( .A(o[8]), .B(\stack[1][44] ), .Z(n9386) );
  XOR U10178 ( .A(n9387), .B(n9386), .Z(n9389) );
  NAND U10179 ( .A(n9112), .B(n9111), .Z(n9116) );
  NAND U10180 ( .A(n9114), .B(n9113), .Z(n9115) );
  NAND U10181 ( .A(n9116), .B(n9115), .Z(n9388) );
  XNOR U10182 ( .A(n9389), .B(n9388), .Z(n9341) );
  NAND U10183 ( .A(n9118), .B(n9117), .Z(n9122) );
  NAND U10184 ( .A(n9120), .B(n9119), .Z(n9121) );
  AND U10185 ( .A(n9122), .B(n9121), .Z(n9340) );
  XOR U10186 ( .A(n9342), .B(n9343), .Z(n9393) );
  XOR U10187 ( .A(n9392), .B(n9393), .Z(n9395) );
  NAND U10188 ( .A(o[10]), .B(\stack[1][42] ), .Z(n9394) );
  XOR U10189 ( .A(n9395), .B(n9394), .Z(n9335) );
  NAND U10190 ( .A(n9124), .B(n9123), .Z(n9128) );
  NAND U10191 ( .A(n9126), .B(n9125), .Z(n9127) );
  AND U10192 ( .A(n9128), .B(n9127), .Z(n9334) );
  XOR U10193 ( .A(n9335), .B(n9334), .Z(n9337) );
  XOR U10194 ( .A(n9336), .B(n9337), .Z(n9329) );
  XOR U10195 ( .A(n9328), .B(n9329), .Z(n9331) );
  NAND U10196 ( .A(o[12]), .B(\stack[1][40] ), .Z(n9330) );
  XNOR U10197 ( .A(n9331), .B(n9330), .Z(n9322) );
  XOR U10198 ( .A(n9323), .B(n9322), .Z(n9325) );
  AND U10199 ( .A(o[13]), .B(\stack[1][39] ), .Z(n9324) );
  XOR U10200 ( .A(n9325), .B(n9324), .Z(n9399) );
  NAND U10201 ( .A(n9130), .B(n9129), .Z(n9134) );
  NAND U10202 ( .A(n9132), .B(n9131), .Z(n9133) );
  NAND U10203 ( .A(n9134), .B(n9133), .Z(n9398) );
  XOR U10204 ( .A(n9399), .B(n9398), .Z(n9400) );
  XOR U10205 ( .A(n9401), .B(n9400), .Z(n9405) );
  XOR U10206 ( .A(n9404), .B(n9405), .Z(n9406) );
  XOR U10207 ( .A(n9407), .B(n9406), .Z(n9318) );
  XOR U10208 ( .A(n9319), .B(n9318), .Z(n9411) );
  NAND U10209 ( .A(n9136), .B(n9135), .Z(n9140) );
  NAND U10210 ( .A(n9138), .B(n9137), .Z(n9139) );
  NAND U10211 ( .A(n9140), .B(n9139), .Z(n9410) );
  XOR U10212 ( .A(n9411), .B(n9410), .Z(n9412) );
  XOR U10213 ( .A(n9413), .B(n9412), .Z(n9312) );
  XOR U10214 ( .A(n9313), .B(n9312), .Z(n9417) );
  NAND U10215 ( .A(n9142), .B(n9141), .Z(n9146) );
  NAND U10216 ( .A(n9144), .B(n9143), .Z(n9145) );
  NAND U10217 ( .A(n9146), .B(n9145), .Z(n9416) );
  XOR U10218 ( .A(n9417), .B(n9416), .Z(n9419) );
  AND U10219 ( .A(o[19]), .B(\stack[1][33] ), .Z(n9418) );
  XNOR U10220 ( .A(n9419), .B(n9418), .Z(n9306) );
  XNOR U10221 ( .A(n9307), .B(n9306), .Z(n9422) );
  XOR U10222 ( .A(n9423), .B(n9422), .Z(n9425) );
  AND U10223 ( .A(o[21]), .B(\stack[1][31] ), .Z(n9424) );
  XOR U10224 ( .A(n9425), .B(n9424), .Z(n9430) );
  XOR U10225 ( .A(n9431), .B(n9430), .Z(n9435) );
  NAND U10226 ( .A(n9148), .B(n9147), .Z(n9152) );
  NAND U10227 ( .A(n9150), .B(n9149), .Z(n9151) );
  NAND U10228 ( .A(n9152), .B(n9151), .Z(n9434) );
  XOR U10229 ( .A(n9435), .B(n9434), .Z(n9437) );
  AND U10230 ( .A(o[23]), .B(\stack[1][29] ), .Z(n9436) );
  XOR U10231 ( .A(n9437), .B(n9436), .Z(n9300) );
  XOR U10232 ( .A(n9301), .B(n9300), .Z(n9441) );
  NAND U10233 ( .A(n9154), .B(n9153), .Z(n9158) );
  NAND U10234 ( .A(n9156), .B(n9155), .Z(n9157) );
  NAND U10235 ( .A(n9158), .B(n9157), .Z(n9440) );
  XOR U10236 ( .A(n9441), .B(n9440), .Z(n9443) );
  AND U10237 ( .A(\stack[1][27] ), .B(o[25]), .Z(n9442) );
  XOR U10238 ( .A(n9443), .B(n9442), .Z(n9294) );
  XOR U10239 ( .A(n9295), .B(n9294), .Z(n9447) );
  NAND U10240 ( .A(n9160), .B(n9159), .Z(n9164) );
  NAND U10241 ( .A(n9162), .B(n9161), .Z(n9163) );
  NAND U10242 ( .A(n9164), .B(n9163), .Z(n9446) );
  XOR U10243 ( .A(n9447), .B(n9446), .Z(n9449) );
  AND U10244 ( .A(\stack[1][25] ), .B(o[27]), .Z(n9448) );
  XOR U10245 ( .A(n9449), .B(n9448), .Z(n9289) );
  NAND U10246 ( .A(n9166), .B(n9165), .Z(n9170) );
  NAND U10247 ( .A(n9168), .B(n9167), .Z(n9169) );
  NAND U10248 ( .A(n9170), .B(n9169), .Z(n9287) );
  AND U10249 ( .A(\stack[1][24] ), .B(o[28]), .Z(n9288) );
  XOR U10250 ( .A(n9287), .B(n9288), .Z(n9290) );
  NAND U10251 ( .A(n9172), .B(n9171), .Z(n9176) );
  NAND U10252 ( .A(n9174), .B(n9173), .Z(n9175) );
  NAND U10253 ( .A(n9176), .B(n9175), .Z(n9452) );
  XOR U10254 ( .A(n9453), .B(n9452), .Z(n9455) );
  AND U10255 ( .A(\stack[1][23] ), .B(o[29]), .Z(n9454) );
  XOR U10256 ( .A(n9455), .B(n9454), .Z(n9283) );
  XOR U10257 ( .A(n9284), .B(n9283), .Z(n9459) );
  NAND U10258 ( .A(n9178), .B(n9177), .Z(n9182) );
  NAND U10259 ( .A(n9180), .B(n9179), .Z(n9181) );
  NAND U10260 ( .A(n9182), .B(n9181), .Z(n9458) );
  XOR U10261 ( .A(n9459), .B(n9458), .Z(n9461) );
  AND U10262 ( .A(\stack[1][21] ), .B(o[31]), .Z(n9460) );
  XOR U10263 ( .A(n9461), .B(n9460), .Z(n9277) );
  NAND U10264 ( .A(n9184), .B(n9183), .Z(n9188) );
  NAND U10265 ( .A(n9186), .B(n9185), .Z(n9187) );
  NAND U10266 ( .A(n9188), .B(n9187), .Z(n9275) );
  AND U10267 ( .A(\stack[1][20] ), .B(o[32]), .Z(n9276) );
  XOR U10268 ( .A(n9275), .B(n9276), .Z(n9278) );
  NAND U10269 ( .A(n9190), .B(n9189), .Z(n9194) );
  NAND U10270 ( .A(n9192), .B(n9191), .Z(n9193) );
  NAND U10271 ( .A(n9194), .B(n9193), .Z(n9464) );
  XOR U10272 ( .A(n9465), .B(n9464), .Z(n9467) );
  AND U10273 ( .A(\stack[1][19] ), .B(o[33]), .Z(n9466) );
  XNOR U10274 ( .A(n9467), .B(n9466), .Z(n9271) );
  XNOR U10275 ( .A(n9272), .B(n9271), .Z(n9470) );
  XOR U10276 ( .A(n9471), .B(n9470), .Z(n9473) );
  AND U10277 ( .A(\stack[1][17] ), .B(o[35]), .Z(n9472) );
  XNOR U10278 ( .A(n9473), .B(n9472), .Z(n9266) );
  NAND U10279 ( .A(n9196), .B(n9195), .Z(n9200) );
  NAND U10280 ( .A(n9198), .B(n9197), .Z(n9199) );
  AND U10281 ( .A(n9200), .B(n9199), .Z(n9264) );
  NAND U10282 ( .A(\stack[1][16] ), .B(o[36]), .Z(n9263) );
  XOR U10283 ( .A(n9264), .B(n9263), .Z(n9265) );
  NAND U10284 ( .A(n9202), .B(n9201), .Z(n9206) );
  NAND U10285 ( .A(n9204), .B(n9203), .Z(n9205) );
  NAND U10286 ( .A(n9206), .B(n9205), .Z(n9476) );
  AND U10287 ( .A(\stack[1][15] ), .B(o[37]), .Z(n9478) );
  XNOR U10288 ( .A(n9479), .B(n9478), .Z(n9260) );
  NAND U10289 ( .A(n9208), .B(n9207), .Z(n9212) );
  NAND U10290 ( .A(n9210), .B(n9209), .Z(n9211) );
  AND U10291 ( .A(n9212), .B(n9211), .Z(n9257) );
  NAND U10292 ( .A(\stack[1][14] ), .B(o[38]), .Z(n9258) );
  NAND U10293 ( .A(n9214), .B(n9213), .Z(n9218) );
  NAND U10294 ( .A(n9216), .B(n9215), .Z(n9217) );
  NAND U10295 ( .A(n9218), .B(n9217), .Z(n9482) );
  XOR U10296 ( .A(n9483), .B(n9482), .Z(n9485) );
  AND U10297 ( .A(\stack[1][13] ), .B(o[39]), .Z(n9484) );
  XNOR U10298 ( .A(n9485), .B(n9484), .Z(n9253) );
  XNOR U10299 ( .A(n9254), .B(n9253), .Z(n9489) );
  NAND U10300 ( .A(n9220), .B(n9219), .Z(n9224) );
  NAND U10301 ( .A(n9222), .B(n9221), .Z(n9223) );
  NAND U10302 ( .A(n9224), .B(n9223), .Z(n9488) );
  AND U10303 ( .A(\stack[1][11] ), .B(o[41]), .Z(n9490) );
  XNOR U10304 ( .A(n9491), .B(n9490), .Z(n9248) );
  NAND U10305 ( .A(n9226), .B(n9225), .Z(n9230) );
  NAND U10306 ( .A(n9228), .B(n9227), .Z(n9229) );
  AND U10307 ( .A(n9230), .B(n9229), .Z(n9245) );
  NAND U10308 ( .A(\stack[1][10] ), .B(o[42]), .Z(n9246) );
  NAND U10309 ( .A(n9232), .B(n9231), .Z(n9236) );
  NAND U10310 ( .A(n9234), .B(n9233), .Z(n9235) );
  NAND U10311 ( .A(n9236), .B(n9235), .Z(n9494) );
  XOR U10312 ( .A(n9495), .B(n9494), .Z(n9497) );
  AND U10313 ( .A(\stack[1][9] ), .B(o[43]), .Z(n9496) );
  XNOR U10314 ( .A(n9497), .B(n9496), .Z(n9241) );
  XNOR U10315 ( .A(n9242), .B(n9241), .Z(n9500) );
  AND U10316 ( .A(\stack[1][7] ), .B(o[45]), .Z(n9502) );
  XNOR U10317 ( .A(n9503), .B(n9502), .Z(n12494) );
  NAND U10318 ( .A(n12495), .B(n12494), .Z(n9237) );
  AND U10319 ( .A(n9238), .B(n9237), .Z(n9507) );
  AND U10320 ( .A(\stack[1][8] ), .B(o[45]), .Z(n9777) );
  NAND U10321 ( .A(n9240), .B(n9239), .Z(n9244) );
  NAND U10322 ( .A(n9242), .B(n9241), .Z(n9243) );
  AND U10323 ( .A(n9244), .B(n9243), .Z(n9775) );
  NAND U10324 ( .A(n9246), .B(n9245), .Z(n9250) );
  NAND U10325 ( .A(n9248), .B(n9247), .Z(n9249) );
  AND U10326 ( .A(n9250), .B(n9249), .Z(n9763) );
  NAND U10327 ( .A(n9252), .B(n9251), .Z(n9256) );
  NAND U10328 ( .A(n9254), .B(n9253), .Z(n9255) );
  AND U10329 ( .A(n9256), .B(n9255), .Z(n9751) );
  AND U10330 ( .A(\stack[1][14] ), .B(o[39]), .Z(n9741) );
  NAND U10331 ( .A(n9258), .B(n9257), .Z(n9262) );
  NAND U10332 ( .A(n9260), .B(n9259), .Z(n9261) );
  AND U10333 ( .A(n9262), .B(n9261), .Z(n9739) );
  AND U10334 ( .A(\stack[1][16] ), .B(o[37]), .Z(n9515) );
  NAND U10335 ( .A(n9264), .B(n9263), .Z(n9268) );
  NAND U10336 ( .A(n9266), .B(n9265), .Z(n9267) );
  AND U10337 ( .A(n9268), .B(n9267), .Z(n9513) );
  NAND U10338 ( .A(n9270), .B(n9269), .Z(n9274) );
  NAND U10339 ( .A(n9272), .B(n9271), .Z(n9273) );
  AND U10340 ( .A(n9274), .B(n9273), .Z(n9721) );
  AND U10341 ( .A(\stack[1][20] ), .B(o[33]), .Z(n9710) );
  NAND U10342 ( .A(n9276), .B(n9275), .Z(n9280) );
  NAND U10343 ( .A(n9278), .B(n9277), .Z(n9279) );
  NAND U10344 ( .A(n9280), .B(n9279), .Z(n9708) );
  NAND U10345 ( .A(n9282), .B(n9281), .Z(n9286) );
  NAND U10346 ( .A(n9284), .B(n9283), .Z(n9285) );
  NAND U10347 ( .A(n9286), .B(n9285), .Z(n9518) );
  AND U10348 ( .A(\stack[1][24] ), .B(o[29]), .Z(n9526) );
  NAND U10349 ( .A(n9288), .B(n9287), .Z(n9292) );
  NAND U10350 ( .A(n9290), .B(n9289), .Z(n9291) );
  NAND U10351 ( .A(n9292), .B(n9291), .Z(n9524) );
  AND U10352 ( .A(\stack[1][26] ), .B(o[27]), .Z(n9532) );
  NAND U10353 ( .A(n16327), .B(n9293), .Z(n9297) );
  NAND U10354 ( .A(n9295), .B(n9294), .Z(n9296) );
  NAND U10355 ( .A(n9297), .B(n9296), .Z(n9530) );
  AND U10356 ( .A(o[25]), .B(\stack[1][28] ), .Z(n9538) );
  NAND U10357 ( .A(n9299), .B(n9298), .Z(n9303) );
  NAND U10358 ( .A(n9301), .B(n9300), .Z(n9302) );
  NAND U10359 ( .A(n9303), .B(n9302), .Z(n9536) );
  AND U10360 ( .A(o[23]), .B(\stack[1][30] ), .Z(n9544) );
  AND U10361 ( .A(o[21]), .B(\stack[1][32] ), .Z(n9551) );
  NAND U10362 ( .A(n9305), .B(n9304), .Z(n9309) );
  NAND U10363 ( .A(n9307), .B(n9306), .Z(n9308) );
  AND U10364 ( .A(n9309), .B(n9308), .Z(n9549) );
  NAND U10365 ( .A(n9311), .B(n9310), .Z(n9315) );
  NAND U10366 ( .A(n9313), .B(n9312), .Z(n9314) );
  NAND U10367 ( .A(n9315), .B(n9314), .Z(n9554) );
  NAND U10368 ( .A(n9317), .B(n9316), .Z(n9321) );
  NAND U10369 ( .A(n9319), .B(n9318), .Z(n9320) );
  AND U10370 ( .A(n9321), .B(n9320), .Z(n9660) );
  NAND U10371 ( .A(o[15]), .B(\stack[1][38] ), .Z(n9656) );
  NAND U10372 ( .A(n9323), .B(n9322), .Z(n9327) );
  NAND U10373 ( .A(n9325), .B(n9324), .Z(n9326) );
  NAND U10374 ( .A(n9327), .B(n9326), .Z(n9574) );
  AND U10375 ( .A(o[14]), .B(\stack[1][39] ), .Z(n9573) );
  NAND U10376 ( .A(n9329), .B(n9328), .Z(n9333) );
  NAND U10377 ( .A(n9331), .B(n9330), .Z(n9332) );
  AND U10378 ( .A(n9333), .B(n9332), .Z(n9579) );
  AND U10379 ( .A(o[12]), .B(\stack[1][41] ), .Z(n9651) );
  NAND U10380 ( .A(n9335), .B(n9334), .Z(n9339) );
  NAND U10381 ( .A(n9337), .B(n9336), .Z(n9338) );
  AND U10382 ( .A(n9339), .B(n9338), .Z(n9648) );
  NAND U10383 ( .A(o[11]), .B(\stack[1][42] ), .Z(n9586) );
  AND U10384 ( .A(o[10]), .B(\stack[1][43] ), .Z(n9593) );
  NAND U10385 ( .A(n9341), .B(n9340), .Z(n9345) );
  NAND U10386 ( .A(n9343), .B(n9342), .Z(n9344) );
  AND U10387 ( .A(n9345), .B(n9344), .Z(n9591) );
  NAND U10388 ( .A(o[9]), .B(\stack[1][44] ), .Z(n9598) );
  NAND U10389 ( .A(n9347), .B(n9346), .Z(n9351) );
  NAND U10390 ( .A(n9349), .B(n9348), .Z(n9350) );
  NAND U10391 ( .A(n9351), .B(n9350), .Z(n9644) );
  NAND U10392 ( .A(n9353), .B(n9352), .Z(n9357) );
  NAND U10393 ( .A(n9355), .B(n9354), .Z(n9356) );
  NAND U10394 ( .A(n9357), .B(n9356), .Z(n9638) );
  AND U10395 ( .A(o[6]), .B(\stack[1][47] ), .Z(n9605) );
  NAND U10396 ( .A(n9359), .B(n9358), .Z(n9363) );
  NAND U10397 ( .A(n9361), .B(n9360), .Z(n9362) );
  AND U10398 ( .A(n9363), .B(n9362), .Z(n9631) );
  NANDN U10399 ( .A(n9364), .B(n9614), .Z(n9368) );
  NANDN U10400 ( .A(n9366), .B(n9365), .Z(n9367) );
  NAND U10401 ( .A(n9368), .B(n9367), .Z(n9624) );
  AND U10402 ( .A(o[2]), .B(\stack[1][51] ), .Z(n9615) );
  AND U10403 ( .A(n9369), .B(n9371), .Z(n9370) );
  AND U10404 ( .A(o[1]), .B(\stack[1][53] ), .Z(n9621) );
  NAND U10405 ( .A(n9619), .B(n9621), .Z(n9944) );
  XOR U10406 ( .A(n9370), .B(n9944), .Z(n9373) );
  AND U10407 ( .A(o[0]), .B(\stack[1][53] ), .Z(n9949) );
  OR U10408 ( .A(n9371), .B(n9949), .Z(n9372) );
  NAND U10409 ( .A(n9373), .B(n9372), .Z(n9616) );
  XNOR U10410 ( .A(n9615), .B(n9616), .Z(n9625) );
  XOR U10411 ( .A(n9624), .B(n9625), .Z(n9627) );
  AND U10412 ( .A(o[3]), .B(\stack[1][50] ), .Z(n9626) );
  XOR U10413 ( .A(n9627), .B(n9626), .Z(n9609) );
  NAND U10414 ( .A(n9375), .B(n9374), .Z(n9379) );
  NAND U10415 ( .A(n9377), .B(n9376), .Z(n9378) );
  NAND U10416 ( .A(n9379), .B(n9378), .Z(n9608) );
  XOR U10417 ( .A(n9609), .B(n9608), .Z(n9611) );
  AND U10418 ( .A(o[4]), .B(\stack[1][49] ), .Z(n9610) );
  XOR U10419 ( .A(n9611), .B(n9610), .Z(n9630) );
  XOR U10420 ( .A(n9631), .B(n9630), .Z(n9633) );
  AND U10421 ( .A(o[5]), .B(\stack[1][48] ), .Z(n9632) );
  XOR U10422 ( .A(n9633), .B(n9632), .Z(n9603) );
  NAND U10423 ( .A(n9381), .B(n9380), .Z(n9385) );
  NAND U10424 ( .A(n9383), .B(n9382), .Z(n9384) );
  NAND U10425 ( .A(n9385), .B(n9384), .Z(n9602) );
  XOR U10426 ( .A(n9603), .B(n9602), .Z(n9604) );
  XOR U10427 ( .A(n9605), .B(n9604), .Z(n9637) );
  AND U10428 ( .A(o[7]), .B(\stack[1][46] ), .Z(n9636) );
  XOR U10429 ( .A(n9637), .B(n9636), .Z(n9639) );
  XOR U10430 ( .A(n9638), .B(n9639), .Z(n9643) );
  AND U10431 ( .A(o[8]), .B(\stack[1][45] ), .Z(n9642) );
  XOR U10432 ( .A(n9643), .B(n9642), .Z(n9645) );
  XNOR U10433 ( .A(n9644), .B(n9645), .Z(n9597) );
  NAND U10434 ( .A(n9387), .B(n9386), .Z(n9391) );
  NAND U10435 ( .A(n9389), .B(n9388), .Z(n9390) );
  AND U10436 ( .A(n9391), .B(n9390), .Z(n9596) );
  XOR U10437 ( .A(n9598), .B(n9599), .Z(n9590) );
  XOR U10438 ( .A(n9591), .B(n9590), .Z(n9592) );
  XNOR U10439 ( .A(n9593), .B(n9592), .Z(n9585) );
  NAND U10440 ( .A(n9393), .B(n9392), .Z(n9397) );
  NAND U10441 ( .A(n9395), .B(n9394), .Z(n9396) );
  NAND U10442 ( .A(n9397), .B(n9396), .Z(n9584) );
  XNOR U10443 ( .A(n9586), .B(n9587), .Z(n9649) );
  XOR U10444 ( .A(n9651), .B(n9650), .Z(n9578) );
  XOR U10445 ( .A(n9579), .B(n9578), .Z(n9581) );
  AND U10446 ( .A(o[13]), .B(\stack[1][40] ), .Z(n9580) );
  XOR U10447 ( .A(n9581), .B(n9580), .Z(n9572) );
  XOR U10448 ( .A(n9573), .B(n9572), .Z(n9575) );
  XNOR U10449 ( .A(n9574), .B(n9575), .Z(n9655) );
  NAND U10450 ( .A(n9399), .B(n9398), .Z(n9403) );
  NAND U10451 ( .A(n9401), .B(n9400), .Z(n9402) );
  AND U10452 ( .A(n9403), .B(n9402), .Z(n9654) );
  XNOR U10453 ( .A(n9656), .B(n9657), .Z(n9569) );
  AND U10454 ( .A(o[16]), .B(\stack[1][37] ), .Z(n9567) );
  NAND U10455 ( .A(n9405), .B(n9404), .Z(n9409) );
  NAND U10456 ( .A(n9407), .B(n9406), .Z(n9408) );
  NAND U10457 ( .A(n9409), .B(n9408), .Z(n9566) );
  XOR U10458 ( .A(n9567), .B(n9566), .Z(n9568) );
  NAND U10459 ( .A(o[17]), .B(\stack[1][36] ), .Z(n9662) );
  XNOR U10460 ( .A(n9663), .B(n9662), .Z(n9563) );
  NAND U10461 ( .A(n9411), .B(n9410), .Z(n9415) );
  NAND U10462 ( .A(n9413), .B(n9412), .Z(n9414) );
  NAND U10463 ( .A(n9415), .B(n9414), .Z(n9560) );
  AND U10464 ( .A(o[18]), .B(\stack[1][35] ), .Z(n9561) );
  XOR U10465 ( .A(n9560), .B(n9561), .Z(n9562) );
  XOR U10466 ( .A(n9554), .B(n9555), .Z(n9557) );
  AND U10467 ( .A(o[19]), .B(\stack[1][34] ), .Z(n9556) );
  XOR U10468 ( .A(n9557), .B(n9556), .Z(n9669) );
  AND U10469 ( .A(o[20]), .B(\stack[1][33] ), .Z(n9667) );
  NAND U10470 ( .A(n9417), .B(n9416), .Z(n9421) );
  NAND U10471 ( .A(n9419), .B(n9418), .Z(n9420) );
  NAND U10472 ( .A(n9421), .B(n9420), .Z(n9666) );
  XOR U10473 ( .A(n9667), .B(n9666), .Z(n9668) );
  XOR U10474 ( .A(n9669), .B(n9668), .Z(n9548) );
  XOR U10475 ( .A(n9549), .B(n9548), .Z(n9550) );
  XNOR U10476 ( .A(n9551), .B(n9550), .Z(n9675) );
  NAND U10477 ( .A(o[22]), .B(\stack[1][31] ), .Z(n9672) );
  NAND U10478 ( .A(n9423), .B(n9422), .Z(n9427) );
  NAND U10479 ( .A(n9425), .B(n9424), .Z(n9426) );
  AND U10480 ( .A(n9427), .B(n9426), .Z(n9673) );
  XOR U10481 ( .A(n9672), .B(n9673), .Z(n9674) );
  NAND U10482 ( .A(n9429), .B(n9428), .Z(n9433) );
  NAND U10483 ( .A(n9431), .B(n9430), .Z(n9432) );
  NAND U10484 ( .A(n9433), .B(n9432), .Z(n9542) );
  XNOR U10485 ( .A(n9544), .B(n9545), .Z(n9681) );
  AND U10486 ( .A(o[24]), .B(\stack[1][29] ), .Z(n9679) );
  NAND U10487 ( .A(n9435), .B(n9434), .Z(n9439) );
  NAND U10488 ( .A(n9437), .B(n9436), .Z(n9438) );
  NAND U10489 ( .A(n9439), .B(n9438), .Z(n9678) );
  XOR U10490 ( .A(n9679), .B(n9678), .Z(n9680) );
  XOR U10491 ( .A(n9681), .B(n9680), .Z(n9537) );
  XOR U10492 ( .A(n9536), .B(n9537), .Z(n9539) );
  AND U10493 ( .A(\stack[1][27] ), .B(o[26]), .Z(n9685) );
  NAND U10494 ( .A(n9441), .B(n9440), .Z(n9445) );
  NAND U10495 ( .A(n9443), .B(n9442), .Z(n9444) );
  NAND U10496 ( .A(n9445), .B(n9444), .Z(n9684) );
  XOR U10497 ( .A(n9685), .B(n9684), .Z(n9686) );
  XOR U10498 ( .A(n9687), .B(n9686), .Z(n9531) );
  XOR U10499 ( .A(n9530), .B(n9531), .Z(n9533) );
  AND U10500 ( .A(\stack[1][25] ), .B(o[28]), .Z(n9691) );
  NAND U10501 ( .A(n9447), .B(n9446), .Z(n9451) );
  NAND U10502 ( .A(n9449), .B(n9448), .Z(n9450) );
  NAND U10503 ( .A(n9451), .B(n9450), .Z(n9690) );
  XOR U10504 ( .A(n9691), .B(n9690), .Z(n9692) );
  XOR U10505 ( .A(n9693), .B(n9692), .Z(n9525) );
  XOR U10506 ( .A(n9524), .B(n9525), .Z(n9527) );
  AND U10507 ( .A(\stack[1][23] ), .B(o[30]), .Z(n9697) );
  NAND U10508 ( .A(n9453), .B(n9452), .Z(n9457) );
  NAND U10509 ( .A(n9455), .B(n9454), .Z(n9456) );
  NAND U10510 ( .A(n9457), .B(n9456), .Z(n9696) );
  XOR U10511 ( .A(n9697), .B(n9696), .Z(n9698) );
  XOR U10512 ( .A(n9699), .B(n9698), .Z(n9519) );
  XOR U10513 ( .A(n9518), .B(n9519), .Z(n9521) );
  AND U10514 ( .A(\stack[1][22] ), .B(o[31]), .Z(n9520) );
  XOR U10515 ( .A(n9521), .B(n9520), .Z(n9705) );
  AND U10516 ( .A(\stack[1][21] ), .B(o[32]), .Z(n9703) );
  NAND U10517 ( .A(n9459), .B(n9458), .Z(n9463) );
  NAND U10518 ( .A(n9461), .B(n9460), .Z(n9462) );
  NAND U10519 ( .A(n9463), .B(n9462), .Z(n9702) );
  XOR U10520 ( .A(n9703), .B(n9702), .Z(n9704) );
  XOR U10521 ( .A(n9705), .B(n9704), .Z(n9709) );
  XOR U10522 ( .A(n9708), .B(n9709), .Z(n9711) );
  AND U10523 ( .A(\stack[1][19] ), .B(o[34]), .Z(n9715) );
  NAND U10524 ( .A(n9465), .B(n9464), .Z(n9469) );
  NAND U10525 ( .A(n9467), .B(n9466), .Z(n9468) );
  NAND U10526 ( .A(n9469), .B(n9468), .Z(n9714) );
  XOR U10527 ( .A(n9715), .B(n9714), .Z(n9716) );
  XOR U10528 ( .A(n9717), .B(n9716), .Z(n9720) );
  XOR U10529 ( .A(n9721), .B(n9720), .Z(n9723) );
  AND U10530 ( .A(\stack[1][18] ), .B(o[35]), .Z(n9722) );
  XOR U10531 ( .A(n9723), .B(n9722), .Z(n9729) );
  AND U10532 ( .A(\stack[1][17] ), .B(o[36]), .Z(n9727) );
  NAND U10533 ( .A(n9471), .B(n9470), .Z(n9475) );
  NAND U10534 ( .A(n9473), .B(n9472), .Z(n9474) );
  NAND U10535 ( .A(n9475), .B(n9474), .Z(n9726) );
  XOR U10536 ( .A(n9727), .B(n9726), .Z(n9728) );
  XOR U10537 ( .A(n9729), .B(n9728), .Z(n9512) );
  XOR U10538 ( .A(n9513), .B(n9512), .Z(n9514) );
  XOR U10539 ( .A(n9515), .B(n9514), .Z(n9735) );
  AND U10540 ( .A(\stack[1][15] ), .B(o[38]), .Z(n9733) );
  NAND U10541 ( .A(n9477), .B(n9476), .Z(n9481) );
  NAND U10542 ( .A(n9479), .B(n9478), .Z(n9480) );
  NAND U10543 ( .A(n9481), .B(n9480), .Z(n9732) );
  XOR U10544 ( .A(n9733), .B(n9732), .Z(n9734) );
  XOR U10545 ( .A(n9735), .B(n9734), .Z(n9738) );
  XOR U10546 ( .A(n9739), .B(n9738), .Z(n9740) );
  XOR U10547 ( .A(n9741), .B(n9740), .Z(n9747) );
  AND U10548 ( .A(\stack[1][13] ), .B(o[40]), .Z(n9744) );
  NAND U10549 ( .A(n9483), .B(n9482), .Z(n9487) );
  NAND U10550 ( .A(n9485), .B(n9484), .Z(n9486) );
  NAND U10551 ( .A(n9487), .B(n9486), .Z(n9745) );
  XOR U10552 ( .A(n9747), .B(n9746), .Z(n9750) );
  XOR U10553 ( .A(n9751), .B(n9750), .Z(n9752) );
  AND U10554 ( .A(\stack[1][12] ), .B(o[41]), .Z(n9753) );
  AND U10555 ( .A(\stack[1][11] ), .B(o[42]), .Z(n9756) );
  NAND U10556 ( .A(n9489), .B(n9488), .Z(n9493) );
  NAND U10557 ( .A(n9491), .B(n9490), .Z(n9492) );
  NAND U10558 ( .A(n9493), .B(n9492), .Z(n9757) );
  XOR U10559 ( .A(n9759), .B(n9758), .Z(n9762) );
  XOR U10560 ( .A(n9763), .B(n9762), .Z(n9764) );
  AND U10561 ( .A(\stack[1][10] ), .B(o[43]), .Z(n9765) );
  AND U10562 ( .A(\stack[1][9] ), .B(o[44]), .Z(n9768) );
  NAND U10563 ( .A(n9495), .B(n9494), .Z(n9499) );
  NAND U10564 ( .A(n9497), .B(n9496), .Z(n9498) );
  NAND U10565 ( .A(n9499), .B(n9498), .Z(n9769) );
  XOR U10566 ( .A(n9771), .B(n9770), .Z(n9774) );
  XOR U10567 ( .A(n9775), .B(n9774), .Z(n9776) );
  XOR U10568 ( .A(n9777), .B(n9776), .Z(n9783) );
  AND U10569 ( .A(\stack[1][7] ), .B(o[46]), .Z(n9780) );
  NAND U10570 ( .A(n9501), .B(n9500), .Z(n9505) );
  NAND U10571 ( .A(n9503), .B(n9502), .Z(n9504) );
  NAND U10572 ( .A(n9505), .B(n9504), .Z(n9781) );
  XOR U10573 ( .A(n9783), .B(n9782), .Z(n9506) );
  NAND U10574 ( .A(n9507), .B(n9506), .Z(n9509) );
  AND U10575 ( .A(\stack[1][6] ), .B(o[47]), .Z(n12501) );
  XOR U10576 ( .A(n9507), .B(n9506), .Z(n12500) );
  NAND U10577 ( .A(n12501), .B(n12500), .Z(n9508) );
  NAND U10578 ( .A(n9509), .B(n9508), .Z(n9510) );
  AND U10579 ( .A(\stack[1][6] ), .B(o[48]), .Z(n9511) );
  NAND U10580 ( .A(n9510), .B(n9511), .Z(n9787) );
  NAND U10581 ( .A(n9513), .B(n9512), .Z(n9517) );
  NAND U10582 ( .A(n9515), .B(n9514), .Z(n9516) );
  NAND U10583 ( .A(n9517), .B(n9516), .Z(n9812) );
  AND U10584 ( .A(\stack[1][16] ), .B(o[38]), .Z(n9813) );
  XOR U10585 ( .A(n9812), .B(n9813), .Z(n9815) );
  NAND U10586 ( .A(n9519), .B(n9518), .Z(n9523) );
  NAND U10587 ( .A(n9521), .B(n9520), .Z(n9522) );
  NAND U10588 ( .A(n9523), .B(n9522), .Z(n9830) );
  AND U10589 ( .A(\stack[1][22] ), .B(o[32]), .Z(n9831) );
  XOR U10590 ( .A(n9830), .B(n9831), .Z(n9833) );
  NAND U10591 ( .A(n9525), .B(n9524), .Z(n9529) );
  NAND U10592 ( .A(n9527), .B(n9526), .Z(n9528) );
  NAND U10593 ( .A(n9529), .B(n9528), .Z(n9836) );
  AND U10594 ( .A(\stack[1][24] ), .B(o[30]), .Z(n9837) );
  XOR U10595 ( .A(n9836), .B(n9837), .Z(n9839) );
  NAND U10596 ( .A(n9531), .B(n9530), .Z(n9535) );
  NAND U10597 ( .A(n9533), .B(n9532), .Z(n9534) );
  NAND U10598 ( .A(n9535), .B(n9534), .Z(n9842) );
  AND U10599 ( .A(\stack[1][26] ), .B(o[28]), .Z(n9843) );
  XOR U10600 ( .A(n9842), .B(n9843), .Z(n9845) );
  AND U10601 ( .A(\stack[1][27] ), .B(o[27]), .Z(n16290) );
  NAND U10602 ( .A(n9537), .B(n9536), .Z(n9541) );
  NAND U10603 ( .A(n9539), .B(n9538), .Z(n9540) );
  NAND U10604 ( .A(n9541), .B(n9540), .Z(n9848) );
  AND U10605 ( .A(o[26]), .B(\stack[1][28] ), .Z(n9849) );
  XOR U10606 ( .A(n9848), .B(n9849), .Z(n9851) );
  NAND U10607 ( .A(n9543), .B(n9542), .Z(n9547) );
  NANDN U10608 ( .A(n9545), .B(n9544), .Z(n9546) );
  NAND U10609 ( .A(n9547), .B(n9546), .Z(n9860) );
  AND U10610 ( .A(o[24]), .B(\stack[1][30] ), .Z(n9861) );
  XOR U10611 ( .A(n9860), .B(n9861), .Z(n9863) );
  NAND U10612 ( .A(n9549), .B(n9548), .Z(n9553) );
  NAND U10613 ( .A(n9551), .B(n9550), .Z(n9552) );
  NAND U10614 ( .A(n9553), .B(n9552), .Z(n9866) );
  AND U10615 ( .A(o[22]), .B(\stack[1][32] ), .Z(n9867) );
  XOR U10616 ( .A(n9866), .B(n9867), .Z(n9869) );
  NAND U10617 ( .A(n9555), .B(n9554), .Z(n9559) );
  NAND U10618 ( .A(n9557), .B(n9556), .Z(n9558) );
  NAND U10619 ( .A(n9559), .B(n9558), .Z(n9878) );
  AND U10620 ( .A(o[20]), .B(\stack[1][34] ), .Z(n9879) );
  XOR U10621 ( .A(n9878), .B(n9879), .Z(n9881) );
  NAND U10622 ( .A(n9561), .B(n9560), .Z(n9565) );
  NAND U10623 ( .A(n9563), .B(n9562), .Z(n9564) );
  NAND U10624 ( .A(n9565), .B(n9564), .Z(n9990) );
  AND U10625 ( .A(o[18]), .B(\stack[1][36] ), .Z(n9887) );
  NAND U10626 ( .A(n9567), .B(n9566), .Z(n9571) );
  NAND U10627 ( .A(n9569), .B(n9568), .Z(n9570) );
  NAND U10628 ( .A(n9571), .B(n9570), .Z(n9985) );
  NAND U10629 ( .A(o[16]), .B(\stack[1][38] ), .Z(n9892) );
  NAND U10630 ( .A(n9573), .B(n9572), .Z(n9577) );
  NAND U10631 ( .A(n9575), .B(n9574), .Z(n9576) );
  NAND U10632 ( .A(n9577), .B(n9576), .Z(n9898) );
  AND U10633 ( .A(o[15]), .B(\stack[1][39] ), .Z(n9896) );
  NAND U10634 ( .A(n9579), .B(n9578), .Z(n9583) );
  NAND U10635 ( .A(n9581), .B(n9580), .Z(n9582) );
  NAND U10636 ( .A(n9583), .B(n9582), .Z(n9904) );
  AND U10637 ( .A(o[12]), .B(\stack[1][42] ), .Z(n9981) );
  NAND U10638 ( .A(n9585), .B(n9584), .Z(n9589) );
  NAND U10639 ( .A(n9587), .B(n9586), .Z(n9588) );
  AND U10640 ( .A(n9589), .B(n9588), .Z(n9979) );
  NAND U10641 ( .A(o[11]), .B(\stack[1][43] ), .Z(n9916) );
  NAND U10642 ( .A(n9591), .B(n9590), .Z(n9595) );
  NAND U10643 ( .A(n9593), .B(n9592), .Z(n9594) );
  AND U10644 ( .A(n9595), .B(n9594), .Z(n9915) );
  AND U10645 ( .A(o[10]), .B(\stack[1][44] ), .Z(n9923) );
  NAND U10646 ( .A(n9597), .B(n9596), .Z(n9601) );
  NANDN U10647 ( .A(n9599), .B(n9598), .Z(n9600) );
  AND U10648 ( .A(n9601), .B(n9600), .Z(n9920) );
  NAND U10649 ( .A(o[9]), .B(\stack[1][45] ), .Z(n9928) );
  NAND U10650 ( .A(n9603), .B(n9602), .Z(n9607) );
  NAND U10651 ( .A(n9605), .B(n9604), .Z(n9606) );
  NAND U10652 ( .A(n9607), .B(n9606), .Z(n9968) );
  AND U10653 ( .A(o[6]), .B(\stack[1][48] ), .Z(n9935) );
  NAND U10654 ( .A(n9609), .B(n9608), .Z(n9613) );
  NAND U10655 ( .A(n9611), .B(n9610), .Z(n9612) );
  NAND U10656 ( .A(n9613), .B(n9612), .Z(n9960) );
  AND U10657 ( .A(o[4]), .B(\stack[1][50] ), .Z(n9941) );
  NANDN U10658 ( .A(n9614), .B(n9944), .Z(n9618) );
  NANDN U10659 ( .A(n9616), .B(n9615), .Z(n9617) );
  NAND U10660 ( .A(n9618), .B(n9617), .Z(n9954) );
  AND U10661 ( .A(o[2]), .B(\stack[1][52] ), .Z(n9945) );
  AND U10662 ( .A(n9619), .B(n9621), .Z(n9620) );
  AND U10663 ( .A(o[1]), .B(\stack[1][54] ), .Z(n9951) );
  NAND U10664 ( .A(n9949), .B(n9951), .Z(n10218) );
  XOR U10665 ( .A(n9620), .B(n10218), .Z(n9623) );
  AND U10666 ( .A(o[0]), .B(\stack[1][54] ), .Z(n10223) );
  OR U10667 ( .A(n9621), .B(n10223), .Z(n9622) );
  NAND U10668 ( .A(n9623), .B(n9622), .Z(n9946) );
  XNOR U10669 ( .A(n9945), .B(n9946), .Z(n9955) );
  XOR U10670 ( .A(n9954), .B(n9955), .Z(n9957) );
  AND U10671 ( .A(o[3]), .B(\stack[1][51] ), .Z(n9956) );
  XOR U10672 ( .A(n9957), .B(n9956), .Z(n9939) );
  NAND U10673 ( .A(n9625), .B(n9624), .Z(n9629) );
  NAND U10674 ( .A(n9627), .B(n9626), .Z(n9628) );
  NAND U10675 ( .A(n9629), .B(n9628), .Z(n9938) );
  XOR U10676 ( .A(n9939), .B(n9938), .Z(n9940) );
  XOR U10677 ( .A(n9941), .B(n9940), .Z(n9961) );
  XOR U10678 ( .A(n9960), .B(n9961), .Z(n9963) );
  AND U10679 ( .A(o[5]), .B(\stack[1][49] ), .Z(n9962) );
  XOR U10680 ( .A(n9963), .B(n9962), .Z(n9933) );
  NAND U10681 ( .A(n9631), .B(n9630), .Z(n9635) );
  NAND U10682 ( .A(n9633), .B(n9632), .Z(n9634) );
  NAND U10683 ( .A(n9635), .B(n9634), .Z(n9932) );
  XOR U10684 ( .A(n9933), .B(n9932), .Z(n9934) );
  XOR U10685 ( .A(n9935), .B(n9934), .Z(n9967) );
  AND U10686 ( .A(o[7]), .B(\stack[1][47] ), .Z(n9966) );
  XOR U10687 ( .A(n9967), .B(n9966), .Z(n9969) );
  XOR U10688 ( .A(n9968), .B(n9969), .Z(n9973) );
  AND U10689 ( .A(o[8]), .B(\stack[1][46] ), .Z(n9972) );
  XOR U10690 ( .A(n9973), .B(n9972), .Z(n9975) );
  NAND U10691 ( .A(n9637), .B(n9636), .Z(n9641) );
  NAND U10692 ( .A(n9639), .B(n9638), .Z(n9640) );
  NAND U10693 ( .A(n9641), .B(n9640), .Z(n9974) );
  XNOR U10694 ( .A(n9975), .B(n9974), .Z(n9927) );
  NAND U10695 ( .A(n9643), .B(n9642), .Z(n9647) );
  NAND U10696 ( .A(n9645), .B(n9644), .Z(n9646) );
  AND U10697 ( .A(n9647), .B(n9646), .Z(n9926) );
  XNOR U10698 ( .A(n9928), .B(n9929), .Z(n9921) );
  XNOR U10699 ( .A(n9923), .B(n9922), .Z(n9914) );
  XOR U10700 ( .A(n9915), .B(n9914), .Z(n9917) );
  XNOR U10701 ( .A(n9916), .B(n9917), .Z(n9978) );
  XOR U10702 ( .A(n9979), .B(n9978), .Z(n9980) );
  XOR U10703 ( .A(n9981), .B(n9980), .Z(n9909) );
  NAND U10704 ( .A(n9649), .B(n9648), .Z(n9653) );
  NAND U10705 ( .A(n9651), .B(n9650), .Z(n9652) );
  NAND U10706 ( .A(n9653), .B(n9652), .Z(n9908) );
  XOR U10707 ( .A(n9909), .B(n9908), .Z(n9911) );
  AND U10708 ( .A(o[13]), .B(\stack[1][41] ), .Z(n9910) );
  XOR U10709 ( .A(n9911), .B(n9910), .Z(n9903) );
  AND U10710 ( .A(o[14]), .B(\stack[1][40] ), .Z(n9902) );
  XOR U10711 ( .A(n9903), .B(n9902), .Z(n9905) );
  XOR U10712 ( .A(n9904), .B(n9905), .Z(n9897) );
  XNOR U10713 ( .A(n9898), .B(n9899), .Z(n9891) );
  NAND U10714 ( .A(n9655), .B(n9654), .Z(n9659) );
  NAND U10715 ( .A(n9657), .B(n9656), .Z(n9658) );
  NAND U10716 ( .A(n9659), .B(n9658), .Z(n9890) );
  XOR U10717 ( .A(n9892), .B(n9893), .Z(n9984) );
  XOR U10718 ( .A(n9985), .B(n9984), .Z(n9987) );
  AND U10719 ( .A(o[17]), .B(\stack[1][37] ), .Z(n9986) );
  XOR U10720 ( .A(n9987), .B(n9986), .Z(n9885) );
  NAND U10721 ( .A(n9661), .B(n9660), .Z(n9665) );
  NAND U10722 ( .A(n9663), .B(n9662), .Z(n9664) );
  AND U10723 ( .A(n9665), .B(n9664), .Z(n9884) );
  XOR U10724 ( .A(n9885), .B(n9884), .Z(n9886) );
  XOR U10725 ( .A(n9887), .B(n9886), .Z(n9991) );
  XOR U10726 ( .A(n9990), .B(n9991), .Z(n9993) );
  AND U10727 ( .A(o[19]), .B(\stack[1][35] ), .Z(n9992) );
  XOR U10728 ( .A(n9993), .B(n9992), .Z(n9880) );
  XOR U10729 ( .A(n9881), .B(n9880), .Z(n9873) );
  NAND U10730 ( .A(n9667), .B(n9666), .Z(n9671) );
  NAND U10731 ( .A(n9669), .B(n9668), .Z(n9670) );
  NAND U10732 ( .A(n9671), .B(n9670), .Z(n9872) );
  XOR U10733 ( .A(n9873), .B(n9872), .Z(n9875) );
  AND U10734 ( .A(o[21]), .B(\stack[1][33] ), .Z(n9874) );
  XOR U10735 ( .A(n9875), .B(n9874), .Z(n9868) );
  XOR U10736 ( .A(n9869), .B(n9868), .Z(n9997) );
  NAND U10737 ( .A(n9673), .B(n9672), .Z(n9677) );
  NAND U10738 ( .A(n9675), .B(n9674), .Z(n9676) );
  AND U10739 ( .A(n9677), .B(n9676), .Z(n9996) );
  XOR U10740 ( .A(n9997), .B(n9996), .Z(n9999) );
  AND U10741 ( .A(o[23]), .B(\stack[1][31] ), .Z(n9998) );
  XOR U10742 ( .A(n9999), .B(n9998), .Z(n9862) );
  XOR U10743 ( .A(n9863), .B(n9862), .Z(n9855) );
  NAND U10744 ( .A(n9679), .B(n9678), .Z(n9683) );
  NAND U10745 ( .A(n9681), .B(n9680), .Z(n9682) );
  NAND U10746 ( .A(n9683), .B(n9682), .Z(n9854) );
  XOR U10747 ( .A(n9855), .B(n9854), .Z(n9857) );
  AND U10748 ( .A(o[25]), .B(\stack[1][29] ), .Z(n9856) );
  XOR U10749 ( .A(n9857), .B(n9856), .Z(n9850) );
  XOR U10750 ( .A(n9851), .B(n9850), .Z(n10003) );
  NAND U10751 ( .A(n9685), .B(n9684), .Z(n9689) );
  NAND U10752 ( .A(n9687), .B(n9686), .Z(n9688) );
  NAND U10753 ( .A(n9689), .B(n9688), .Z(n10002) );
  XOR U10754 ( .A(n10003), .B(n10002), .Z(n10004) );
  XOR U10755 ( .A(n16290), .B(n10004), .Z(n9844) );
  XOR U10756 ( .A(n9845), .B(n9844), .Z(n10008) );
  NAND U10757 ( .A(n9691), .B(n9690), .Z(n9695) );
  NAND U10758 ( .A(n9693), .B(n9692), .Z(n9694) );
  NAND U10759 ( .A(n9695), .B(n9694), .Z(n10007) );
  XOR U10760 ( .A(n10008), .B(n10007), .Z(n10010) );
  AND U10761 ( .A(\stack[1][25] ), .B(o[29]), .Z(n10009) );
  XOR U10762 ( .A(n10010), .B(n10009), .Z(n9838) );
  XOR U10763 ( .A(n9839), .B(n9838), .Z(n10014) );
  NAND U10764 ( .A(n9697), .B(n9696), .Z(n9701) );
  NAND U10765 ( .A(n9699), .B(n9698), .Z(n9700) );
  NAND U10766 ( .A(n9701), .B(n9700), .Z(n10013) );
  XOR U10767 ( .A(n10014), .B(n10013), .Z(n10016) );
  AND U10768 ( .A(\stack[1][23] ), .B(o[31]), .Z(n10015) );
  XOR U10769 ( .A(n10016), .B(n10015), .Z(n9832) );
  XOR U10770 ( .A(n9833), .B(n9832), .Z(n10020) );
  NAND U10771 ( .A(n9703), .B(n9702), .Z(n9707) );
  NAND U10772 ( .A(n9705), .B(n9704), .Z(n9706) );
  NAND U10773 ( .A(n9707), .B(n9706), .Z(n10019) );
  XOR U10774 ( .A(n10020), .B(n10019), .Z(n10022) );
  AND U10775 ( .A(\stack[1][21] ), .B(o[33]), .Z(n10021) );
  XOR U10776 ( .A(n10022), .B(n10021), .Z(n9826) );
  NAND U10777 ( .A(n9709), .B(n9708), .Z(n9713) );
  NAND U10778 ( .A(n9711), .B(n9710), .Z(n9712) );
  NAND U10779 ( .A(n9713), .B(n9712), .Z(n9824) );
  AND U10780 ( .A(\stack[1][20] ), .B(o[34]), .Z(n9825) );
  XOR U10781 ( .A(n9824), .B(n9825), .Z(n9827) );
  NAND U10782 ( .A(n9715), .B(n9714), .Z(n9719) );
  NAND U10783 ( .A(n9717), .B(n9716), .Z(n9718) );
  NAND U10784 ( .A(n9719), .B(n9718), .Z(n10025) );
  XOR U10785 ( .A(n10026), .B(n10025), .Z(n10028) );
  AND U10786 ( .A(\stack[1][19] ), .B(o[35]), .Z(n10027) );
  XOR U10787 ( .A(n10028), .B(n10027), .Z(n9820) );
  NAND U10788 ( .A(n9721), .B(n9720), .Z(n9725) );
  NAND U10789 ( .A(n9723), .B(n9722), .Z(n9724) );
  NAND U10790 ( .A(n9725), .B(n9724), .Z(n9818) );
  AND U10791 ( .A(\stack[1][18] ), .B(o[36]), .Z(n9819) );
  XOR U10792 ( .A(n9818), .B(n9819), .Z(n9821) );
  NAND U10793 ( .A(n9727), .B(n9726), .Z(n9731) );
  NAND U10794 ( .A(n9729), .B(n9728), .Z(n9730) );
  NAND U10795 ( .A(n9731), .B(n9730), .Z(n10031) );
  XOR U10796 ( .A(n10032), .B(n10031), .Z(n10034) );
  AND U10797 ( .A(\stack[1][17] ), .B(o[37]), .Z(n10033) );
  XOR U10798 ( .A(n10034), .B(n10033), .Z(n9814) );
  XOR U10799 ( .A(n9815), .B(n9814), .Z(n10038) );
  NAND U10800 ( .A(n9733), .B(n9732), .Z(n9737) );
  NAND U10801 ( .A(n9735), .B(n9734), .Z(n9736) );
  NAND U10802 ( .A(n9737), .B(n9736), .Z(n10037) );
  XOR U10803 ( .A(n10038), .B(n10037), .Z(n10040) );
  AND U10804 ( .A(\stack[1][15] ), .B(o[39]), .Z(n10039) );
  XOR U10805 ( .A(n10040), .B(n10039), .Z(n9809) );
  NAND U10806 ( .A(n9739), .B(n9738), .Z(n9743) );
  NAND U10807 ( .A(n9741), .B(n9740), .Z(n9742) );
  NAND U10808 ( .A(n9743), .B(n9742), .Z(n9807) );
  AND U10809 ( .A(\stack[1][14] ), .B(o[40]), .Z(n9806) );
  XOR U10810 ( .A(n9809), .B(n9808), .Z(n10043) );
  NAND U10811 ( .A(n9745), .B(n9744), .Z(n9749) );
  NAND U10812 ( .A(n9747), .B(n9746), .Z(n9748) );
  NAND U10813 ( .A(n9749), .B(n9748), .Z(n10044) );
  AND U10814 ( .A(\stack[1][13] ), .B(o[41]), .Z(n10046) );
  NAND U10815 ( .A(n9751), .B(n9750), .Z(n9755) );
  NAND U10816 ( .A(n9753), .B(n9752), .Z(n9754) );
  NAND U10817 ( .A(n9755), .B(n9754), .Z(n9801) );
  AND U10818 ( .A(\stack[1][12] ), .B(o[42]), .Z(n9800) );
  XOR U10819 ( .A(n9803), .B(n9802), .Z(n10049) );
  NAND U10820 ( .A(n9757), .B(n9756), .Z(n9761) );
  NAND U10821 ( .A(n9759), .B(n9758), .Z(n9760) );
  NAND U10822 ( .A(n9761), .B(n9760), .Z(n10050) );
  AND U10823 ( .A(\stack[1][11] ), .B(o[43]), .Z(n10052) );
  NAND U10824 ( .A(n9763), .B(n9762), .Z(n9767) );
  NAND U10825 ( .A(n9765), .B(n9764), .Z(n9766) );
  NAND U10826 ( .A(n9767), .B(n9766), .Z(n9795) );
  AND U10827 ( .A(\stack[1][10] ), .B(o[44]), .Z(n9794) );
  XOR U10828 ( .A(n9797), .B(n9796), .Z(n10055) );
  NAND U10829 ( .A(n9769), .B(n9768), .Z(n9773) );
  NAND U10830 ( .A(n9771), .B(n9770), .Z(n9772) );
  NAND U10831 ( .A(n9773), .B(n9772), .Z(n10056) );
  AND U10832 ( .A(\stack[1][9] ), .B(o[45]), .Z(n10058) );
  NAND U10833 ( .A(n9775), .B(n9774), .Z(n9779) );
  NAND U10834 ( .A(n9777), .B(n9776), .Z(n9778) );
  NAND U10835 ( .A(n9779), .B(n9778), .Z(n9789) );
  AND U10836 ( .A(\stack[1][8] ), .B(o[46]), .Z(n9788) );
  XOR U10837 ( .A(n9791), .B(n9790), .Z(n10061) );
  NAND U10838 ( .A(n9781), .B(n9780), .Z(n9785) );
  NAND U10839 ( .A(n9783), .B(n9782), .Z(n9784) );
  NAND U10840 ( .A(n9785), .B(n9784), .Z(n10062) );
  AND U10841 ( .A(\stack[1][7] ), .B(o[47]), .Z(n10064) );
  NAND U10842 ( .A(n12507), .B(n12506), .Z(n9786) );
  NAND U10843 ( .A(n9787), .B(n9786), .Z(n10067) );
  NAND U10844 ( .A(n9789), .B(n9788), .Z(n9793) );
  NAND U10845 ( .A(n9791), .B(n9790), .Z(n9792) );
  NAND U10846 ( .A(n9793), .B(n9792), .Z(n10349) );
  AND U10847 ( .A(\stack[1][10] ), .B(o[45]), .Z(n10077) );
  NAND U10848 ( .A(n9795), .B(n9794), .Z(n9799) );
  NAND U10849 ( .A(n9797), .B(n9796), .Z(n9798) );
  NAND U10850 ( .A(n9799), .B(n9798), .Z(n10075) );
  NAND U10851 ( .A(n9801), .B(n9800), .Z(n9805) );
  NAND U10852 ( .A(n9803), .B(n9802), .Z(n9804) );
  NAND U10853 ( .A(n9805), .B(n9804), .Z(n10081) );
  AND U10854 ( .A(\stack[1][14] ), .B(o[41]), .Z(n10088) );
  NAND U10855 ( .A(n9807), .B(n9806), .Z(n9811) );
  NAND U10856 ( .A(n9809), .B(n9808), .Z(n9810) );
  NAND U10857 ( .A(n9811), .B(n9810), .Z(n10086) );
  AND U10858 ( .A(\stack[1][16] ), .B(o[39]), .Z(n10320) );
  NAND U10859 ( .A(n9813), .B(n9812), .Z(n9817) );
  NAND U10860 ( .A(n9815), .B(n9814), .Z(n9816) );
  NAND U10861 ( .A(n9817), .B(n9816), .Z(n10318) );
  NAND U10862 ( .A(n9819), .B(n9818), .Z(n9823) );
  NAND U10863 ( .A(n9821), .B(n9820), .Z(n9822) );
  NAND U10864 ( .A(n9823), .B(n9822), .Z(n10306) );
  AND U10865 ( .A(\stack[1][20] ), .B(o[35]), .Z(n10094) );
  NAND U10866 ( .A(n9825), .B(n9824), .Z(n9829) );
  NAND U10867 ( .A(n9827), .B(n9826), .Z(n9828) );
  NAND U10868 ( .A(n9829), .B(n9828), .Z(n10092) );
  NAND U10869 ( .A(n9831), .B(n9830), .Z(n9835) );
  NAND U10870 ( .A(n9833), .B(n9832), .Z(n9834) );
  NAND U10871 ( .A(n9835), .B(n9834), .Z(n10104) );
  NAND U10872 ( .A(n9837), .B(n9836), .Z(n9841) );
  NAND U10873 ( .A(n9839), .B(n9838), .Z(n9840) );
  NAND U10874 ( .A(n9841), .B(n9840), .Z(n10116) );
  NAND U10875 ( .A(n9843), .B(n9842), .Z(n9847) );
  NAND U10876 ( .A(n9845), .B(n9844), .Z(n9846) );
  NAND U10877 ( .A(n9847), .B(n9846), .Z(n10288) );
  AND U10878 ( .A(\stack[1][28] ), .B(o[27]), .Z(n10124) );
  NAND U10879 ( .A(n9849), .B(n9848), .Z(n9853) );
  NAND U10880 ( .A(n9851), .B(n9850), .Z(n9852) );
  NAND U10881 ( .A(n9853), .B(n9852), .Z(n10122) );
  AND U10882 ( .A(o[26]), .B(\stack[1][29] ), .Z(n10129) );
  NAND U10883 ( .A(n9855), .B(n9854), .Z(n9859) );
  NAND U10884 ( .A(n9857), .B(n9856), .Z(n9858) );
  NAND U10885 ( .A(n9859), .B(n9858), .Z(n10128) );
  XOR U10886 ( .A(n10129), .B(n10128), .Z(n10131) );
  AND U10887 ( .A(o[25]), .B(\stack[1][30] ), .Z(n10136) );
  NAND U10888 ( .A(n9861), .B(n9860), .Z(n9865) );
  NAND U10889 ( .A(n9863), .B(n9862), .Z(n9864) );
  NAND U10890 ( .A(n9865), .B(n9864), .Z(n10134) );
  AND U10891 ( .A(o[23]), .B(\stack[1][32] ), .Z(n10142) );
  NAND U10892 ( .A(n9867), .B(n9866), .Z(n9871) );
  NAND U10893 ( .A(n9869), .B(n9868), .Z(n9870) );
  NAND U10894 ( .A(n9871), .B(n9870), .Z(n10140) );
  AND U10895 ( .A(o[22]), .B(\stack[1][33] ), .Z(n10271) );
  NAND U10896 ( .A(n9873), .B(n9872), .Z(n9877) );
  NAND U10897 ( .A(n9875), .B(n9874), .Z(n9876) );
  NAND U10898 ( .A(n9877), .B(n9876), .Z(n10270) );
  XOR U10899 ( .A(n10271), .B(n10270), .Z(n10273) );
  AND U10900 ( .A(o[21]), .B(\stack[1][34] ), .Z(n10148) );
  NAND U10901 ( .A(n9879), .B(n9878), .Z(n9883) );
  NAND U10902 ( .A(n9881), .B(n9880), .Z(n9882) );
  NAND U10903 ( .A(n9883), .B(n9882), .Z(n10146) );
  NAND U10904 ( .A(n9885), .B(n9884), .Z(n9889) );
  NAND U10905 ( .A(n9887), .B(n9886), .Z(n9888) );
  NAND U10906 ( .A(n9889), .B(n9888), .Z(n10152) );
  AND U10907 ( .A(o[19]), .B(\stack[1][36] ), .Z(n10153) );
  XOR U10908 ( .A(n10152), .B(n10153), .Z(n10154) );
  NAND U10909 ( .A(o[17]), .B(\stack[1][38] ), .Z(n10166) );
  NAND U10910 ( .A(n9891), .B(n9890), .Z(n9895) );
  NANDN U10911 ( .A(n9893), .B(n9892), .Z(n9894) );
  NAND U10912 ( .A(n9895), .B(n9894), .Z(n10165) );
  NAND U10913 ( .A(n9897), .B(n9896), .Z(n9901) );
  NAND U10914 ( .A(n9899), .B(n9898), .Z(n9900) );
  NAND U10915 ( .A(n9901), .B(n9900), .Z(n10260) );
  NAND U10916 ( .A(n9903), .B(n9902), .Z(n9907) );
  NAND U10917 ( .A(n9905), .B(n9904), .Z(n9906) );
  NAND U10918 ( .A(n9907), .B(n9906), .Z(n10254) );
  NAND U10919 ( .A(n9909), .B(n9908), .Z(n9913) );
  NAND U10920 ( .A(n9911), .B(n9910), .Z(n9912) );
  NAND U10921 ( .A(n9913), .B(n9912), .Z(n10172) );
  AND U10922 ( .A(o[12]), .B(\stack[1][43] ), .Z(n10185) );
  NAND U10923 ( .A(n9915), .B(n9914), .Z(n9919) );
  NAND U10924 ( .A(n9917), .B(n9916), .Z(n9918) );
  AND U10925 ( .A(n9919), .B(n9918), .Z(n10183) );
  NAND U10926 ( .A(o[11]), .B(\stack[1][44] ), .Z(n10190) );
  NAND U10927 ( .A(n9921), .B(n9920), .Z(n9925) );
  NAND U10928 ( .A(n9923), .B(n9922), .Z(n9924) );
  AND U10929 ( .A(n9925), .B(n9924), .Z(n10189) );
  AND U10930 ( .A(o[10]), .B(\stack[1][45] ), .Z(n10197) );
  NAND U10931 ( .A(n9927), .B(n9926), .Z(n9931) );
  NAND U10932 ( .A(n9929), .B(n9928), .Z(n9930) );
  AND U10933 ( .A(n9931), .B(n9930), .Z(n10194) );
  NAND U10934 ( .A(o[9]), .B(\stack[1][46] ), .Z(n10202) );
  NAND U10935 ( .A(n9933), .B(n9932), .Z(n9937) );
  NAND U10936 ( .A(n9935), .B(n9934), .Z(n9936) );
  NAND U10937 ( .A(n9937), .B(n9936), .Z(n10242) );
  AND U10938 ( .A(o[6]), .B(\stack[1][49] ), .Z(n10209) );
  NAND U10939 ( .A(n9939), .B(n9938), .Z(n9943) );
  NAND U10940 ( .A(n9941), .B(n9940), .Z(n9942) );
  NAND U10941 ( .A(n9943), .B(n9942), .Z(n10234) );
  AND U10942 ( .A(o[4]), .B(\stack[1][51] ), .Z(n10215) );
  NANDN U10943 ( .A(n9944), .B(n10218), .Z(n9948) );
  NANDN U10944 ( .A(n9946), .B(n9945), .Z(n9947) );
  NAND U10945 ( .A(n9948), .B(n9947), .Z(n10228) );
  AND U10946 ( .A(o[2]), .B(\stack[1][53] ), .Z(n10219) );
  AND U10947 ( .A(n9949), .B(n9951), .Z(n9950) );
  AND U10948 ( .A(o[1]), .B(\stack[1][55] ), .Z(n10225) );
  NAND U10949 ( .A(n10223), .B(n10225), .Z(n10511) );
  XOR U10950 ( .A(n9950), .B(n10511), .Z(n9953) );
  AND U10951 ( .A(o[0]), .B(\stack[1][55] ), .Z(n10516) );
  OR U10952 ( .A(n9951), .B(n10516), .Z(n9952) );
  NAND U10953 ( .A(n9953), .B(n9952), .Z(n10220) );
  XNOR U10954 ( .A(n10219), .B(n10220), .Z(n10229) );
  XOR U10955 ( .A(n10228), .B(n10229), .Z(n10231) );
  AND U10956 ( .A(o[3]), .B(\stack[1][52] ), .Z(n10230) );
  XOR U10957 ( .A(n10231), .B(n10230), .Z(n10213) );
  NAND U10958 ( .A(n9955), .B(n9954), .Z(n9959) );
  NAND U10959 ( .A(n9957), .B(n9956), .Z(n9958) );
  NAND U10960 ( .A(n9959), .B(n9958), .Z(n10212) );
  XOR U10961 ( .A(n10213), .B(n10212), .Z(n10214) );
  XOR U10962 ( .A(n10215), .B(n10214), .Z(n10235) );
  XOR U10963 ( .A(n10234), .B(n10235), .Z(n10237) );
  AND U10964 ( .A(o[5]), .B(\stack[1][50] ), .Z(n10236) );
  XOR U10965 ( .A(n10237), .B(n10236), .Z(n10207) );
  NAND U10966 ( .A(n9961), .B(n9960), .Z(n9965) );
  NAND U10967 ( .A(n9963), .B(n9962), .Z(n9964) );
  NAND U10968 ( .A(n9965), .B(n9964), .Z(n10206) );
  XOR U10969 ( .A(n10207), .B(n10206), .Z(n10208) );
  XOR U10970 ( .A(n10209), .B(n10208), .Z(n10241) );
  AND U10971 ( .A(o[7]), .B(\stack[1][48] ), .Z(n10240) );
  XOR U10972 ( .A(n10241), .B(n10240), .Z(n10243) );
  XOR U10973 ( .A(n10242), .B(n10243), .Z(n10247) );
  AND U10974 ( .A(o[8]), .B(\stack[1][47] ), .Z(n10246) );
  XOR U10975 ( .A(n10247), .B(n10246), .Z(n10249) );
  NAND U10976 ( .A(n9967), .B(n9966), .Z(n9971) );
  NAND U10977 ( .A(n9969), .B(n9968), .Z(n9970) );
  NAND U10978 ( .A(n9971), .B(n9970), .Z(n10248) );
  XNOR U10979 ( .A(n10249), .B(n10248), .Z(n10201) );
  NAND U10980 ( .A(n9973), .B(n9972), .Z(n9977) );
  NAND U10981 ( .A(n9975), .B(n9974), .Z(n9976) );
  AND U10982 ( .A(n9977), .B(n9976), .Z(n10200) );
  XNOR U10983 ( .A(n10202), .B(n10203), .Z(n10195) );
  XNOR U10984 ( .A(n10197), .B(n10196), .Z(n10188) );
  XOR U10985 ( .A(n10189), .B(n10188), .Z(n10191) );
  XNOR U10986 ( .A(n10190), .B(n10191), .Z(n10182) );
  XOR U10987 ( .A(n10183), .B(n10182), .Z(n10184) );
  XOR U10988 ( .A(n10185), .B(n10184), .Z(n10177) );
  NAND U10989 ( .A(n9979), .B(n9978), .Z(n9983) );
  NAND U10990 ( .A(n9981), .B(n9980), .Z(n9982) );
  NAND U10991 ( .A(n9983), .B(n9982), .Z(n10176) );
  XOR U10992 ( .A(n10177), .B(n10176), .Z(n10179) );
  AND U10993 ( .A(o[13]), .B(\stack[1][42] ), .Z(n10178) );
  XOR U10994 ( .A(n10179), .B(n10178), .Z(n10171) );
  AND U10995 ( .A(o[14]), .B(\stack[1][41] ), .Z(n10170) );
  XOR U10996 ( .A(n10171), .B(n10170), .Z(n10173) );
  XOR U10997 ( .A(n10172), .B(n10173), .Z(n10253) );
  AND U10998 ( .A(o[15]), .B(\stack[1][40] ), .Z(n10252) );
  XOR U10999 ( .A(n10253), .B(n10252), .Z(n10255) );
  XOR U11000 ( .A(n10254), .B(n10255), .Z(n10259) );
  AND U11001 ( .A(o[16]), .B(\stack[1][39] ), .Z(n10258) );
  XOR U11002 ( .A(n10259), .B(n10258), .Z(n10261) );
  XNOR U11003 ( .A(n10260), .B(n10261), .Z(n10164) );
  XOR U11004 ( .A(n10165), .B(n10164), .Z(n10167) );
  XNOR U11005 ( .A(n10166), .B(n10167), .Z(n10161) );
  AND U11006 ( .A(o[18]), .B(\stack[1][37] ), .Z(n10159) );
  NAND U11007 ( .A(n9985), .B(n9984), .Z(n9989) );
  NAND U11008 ( .A(n9987), .B(n9986), .Z(n9988) );
  NAND U11009 ( .A(n9989), .B(n9988), .Z(n10158) );
  XOR U11010 ( .A(n10159), .B(n10158), .Z(n10160) );
  XNOR U11011 ( .A(n10154), .B(n10155), .Z(n10267) );
  AND U11012 ( .A(o[20]), .B(\stack[1][35] ), .Z(n10265) );
  NAND U11013 ( .A(n9991), .B(n9990), .Z(n9995) );
  NAND U11014 ( .A(n9993), .B(n9992), .Z(n9994) );
  NAND U11015 ( .A(n9995), .B(n9994), .Z(n10264) );
  XOR U11016 ( .A(n10265), .B(n10264), .Z(n10266) );
  XOR U11017 ( .A(n10267), .B(n10266), .Z(n10147) );
  XOR U11018 ( .A(n10146), .B(n10147), .Z(n10149) );
  XOR U11019 ( .A(n10273), .B(n10272), .Z(n10141) );
  XOR U11020 ( .A(n10140), .B(n10141), .Z(n10143) );
  AND U11021 ( .A(o[24]), .B(\stack[1][31] ), .Z(n10277) );
  NAND U11022 ( .A(n9997), .B(n9996), .Z(n10001) );
  NAND U11023 ( .A(n9999), .B(n9998), .Z(n10000) );
  NAND U11024 ( .A(n10001), .B(n10000), .Z(n10276) );
  XOR U11025 ( .A(n10277), .B(n10276), .Z(n10278) );
  XOR U11026 ( .A(n10279), .B(n10278), .Z(n10135) );
  XOR U11027 ( .A(n10134), .B(n10135), .Z(n10137) );
  XOR U11028 ( .A(n10131), .B(n10130), .Z(n10123) );
  XOR U11029 ( .A(n10122), .B(n10123), .Z(n10125) );
  AND U11030 ( .A(\stack[1][27] ), .B(o[28]), .Z(n10283) );
  NAND U11031 ( .A(n10003), .B(n10002), .Z(n10006) );
  NAND U11032 ( .A(n16290), .B(n10004), .Z(n10005) );
  NAND U11033 ( .A(n10006), .B(n10005), .Z(n10282) );
  XOR U11034 ( .A(n10283), .B(n10282), .Z(n10284) );
  XOR U11035 ( .A(n10285), .B(n10284), .Z(n10289) );
  XOR U11036 ( .A(n10288), .B(n10289), .Z(n10291) );
  AND U11037 ( .A(\stack[1][26] ), .B(o[29]), .Z(n10290) );
  XOR U11038 ( .A(n10291), .B(n10290), .Z(n10297) );
  AND U11039 ( .A(\stack[1][25] ), .B(o[30]), .Z(n10295) );
  NAND U11040 ( .A(n10008), .B(n10007), .Z(n10012) );
  NAND U11041 ( .A(n10010), .B(n10009), .Z(n10011) );
  NAND U11042 ( .A(n10012), .B(n10011), .Z(n10294) );
  XOR U11043 ( .A(n10295), .B(n10294), .Z(n10296) );
  XOR U11044 ( .A(n10297), .B(n10296), .Z(n10117) );
  XOR U11045 ( .A(n10116), .B(n10117), .Z(n10119) );
  AND U11046 ( .A(\stack[1][24] ), .B(o[31]), .Z(n10118) );
  XOR U11047 ( .A(n10119), .B(n10118), .Z(n10113) );
  AND U11048 ( .A(\stack[1][23] ), .B(o[32]), .Z(n10111) );
  NAND U11049 ( .A(n10014), .B(n10013), .Z(n10018) );
  NAND U11050 ( .A(n10016), .B(n10015), .Z(n10017) );
  NAND U11051 ( .A(n10018), .B(n10017), .Z(n10110) );
  XOR U11052 ( .A(n10111), .B(n10110), .Z(n10112) );
  XOR U11053 ( .A(n10113), .B(n10112), .Z(n10105) );
  XOR U11054 ( .A(n10104), .B(n10105), .Z(n10107) );
  AND U11055 ( .A(\stack[1][22] ), .B(o[33]), .Z(n10106) );
  XOR U11056 ( .A(n10107), .B(n10106), .Z(n10101) );
  AND U11057 ( .A(\stack[1][21] ), .B(o[34]), .Z(n10099) );
  NAND U11058 ( .A(n10020), .B(n10019), .Z(n10024) );
  NAND U11059 ( .A(n10022), .B(n10021), .Z(n10023) );
  NAND U11060 ( .A(n10024), .B(n10023), .Z(n10098) );
  XOR U11061 ( .A(n10099), .B(n10098), .Z(n10100) );
  XOR U11062 ( .A(n10101), .B(n10100), .Z(n10093) );
  XOR U11063 ( .A(n10092), .B(n10093), .Z(n10095) );
  AND U11064 ( .A(\stack[1][19] ), .B(o[36]), .Z(n10301) );
  NAND U11065 ( .A(n10026), .B(n10025), .Z(n10030) );
  NAND U11066 ( .A(n10028), .B(n10027), .Z(n10029) );
  NAND U11067 ( .A(n10030), .B(n10029), .Z(n10300) );
  XOR U11068 ( .A(n10301), .B(n10300), .Z(n10302) );
  XOR U11069 ( .A(n10303), .B(n10302), .Z(n10307) );
  XOR U11070 ( .A(n10306), .B(n10307), .Z(n10309) );
  AND U11071 ( .A(\stack[1][18] ), .B(o[37]), .Z(n10308) );
  XOR U11072 ( .A(n10309), .B(n10308), .Z(n10315) );
  AND U11073 ( .A(\stack[1][17] ), .B(o[38]), .Z(n10313) );
  NAND U11074 ( .A(n10032), .B(n10031), .Z(n10036) );
  NAND U11075 ( .A(n10034), .B(n10033), .Z(n10035) );
  NAND U11076 ( .A(n10036), .B(n10035), .Z(n10312) );
  XOR U11077 ( .A(n10313), .B(n10312), .Z(n10314) );
  XOR U11078 ( .A(n10315), .B(n10314), .Z(n10319) );
  XOR U11079 ( .A(n10318), .B(n10319), .Z(n10321) );
  AND U11080 ( .A(\stack[1][15] ), .B(o[40]), .Z(n10325) );
  NAND U11081 ( .A(n10038), .B(n10037), .Z(n10042) );
  NAND U11082 ( .A(n10040), .B(n10039), .Z(n10041) );
  NAND U11083 ( .A(n10042), .B(n10041), .Z(n10324) );
  XOR U11084 ( .A(n10325), .B(n10324), .Z(n10326) );
  XOR U11085 ( .A(n10327), .B(n10326), .Z(n10087) );
  XOR U11086 ( .A(n10086), .B(n10087), .Z(n10089) );
  AND U11087 ( .A(\stack[1][13] ), .B(o[42]), .Z(n10331) );
  NAND U11088 ( .A(n10044), .B(n10043), .Z(n10048) );
  NAND U11089 ( .A(n10046), .B(n10045), .Z(n10047) );
  NAND U11090 ( .A(n10048), .B(n10047), .Z(n10330) );
  XOR U11091 ( .A(n10331), .B(n10330), .Z(n10332) );
  XOR U11092 ( .A(n10333), .B(n10332), .Z(n10080) );
  AND U11093 ( .A(\stack[1][12] ), .B(o[43]), .Z(n10083) );
  AND U11094 ( .A(\stack[1][11] ), .B(o[44]), .Z(n10336) );
  NAND U11095 ( .A(n10050), .B(n10049), .Z(n10054) );
  NAND U11096 ( .A(n10052), .B(n10051), .Z(n10053) );
  NAND U11097 ( .A(n10054), .B(n10053), .Z(n10337) );
  XOR U11098 ( .A(n10339), .B(n10338), .Z(n10074) );
  XOR U11099 ( .A(n10077), .B(n10076), .Z(n10345) );
  AND U11100 ( .A(\stack[1][9] ), .B(o[46]), .Z(n10342) );
  NAND U11101 ( .A(n10056), .B(n10055), .Z(n10060) );
  NAND U11102 ( .A(n10058), .B(n10057), .Z(n10059) );
  NAND U11103 ( .A(n10060), .B(n10059), .Z(n10343) );
  XOR U11104 ( .A(n10345), .B(n10344), .Z(n10348) );
  AND U11105 ( .A(\stack[1][8] ), .B(o[47]), .Z(n10351) );
  AND U11106 ( .A(\stack[1][7] ), .B(o[48]), .Z(n10354) );
  NAND U11107 ( .A(n10062), .B(n10061), .Z(n10066) );
  NAND U11108 ( .A(n10064), .B(n10063), .Z(n10065) );
  NAND U11109 ( .A(n10066), .B(n10065), .Z(n10355) );
  XOR U11110 ( .A(n10357), .B(n10356), .Z(n10068) );
  NAND U11111 ( .A(n10067), .B(n10068), .Z(n10070) );
  AND U11112 ( .A(\stack[1][6] ), .B(o[49]), .Z(n12513) );
  NAND U11113 ( .A(n12513), .B(n12512), .Z(n10069) );
  AND U11114 ( .A(n10070), .B(n10069), .Z(n10073) );
  NAND U11115 ( .A(n10071), .B(n10073), .Z(n10361) );
  IV U11116 ( .A(n10071), .Z(n10072) );
  XNOR U11117 ( .A(n10073), .B(n10072), .Z(n12519) );
  NAND U11118 ( .A(n10075), .B(n10074), .Z(n10079) );
  NAND U11119 ( .A(n10077), .B(n10076), .Z(n10078) );
  NAND U11120 ( .A(n10079), .B(n10078), .Z(n10369) );
  AND U11121 ( .A(\stack[1][10] ), .B(o[46]), .Z(n10368) );
  NAND U11122 ( .A(n10081), .B(n10080), .Z(n10085) );
  NAND U11123 ( .A(n10083), .B(n10082), .Z(n10084) );
  NAND U11124 ( .A(n10085), .B(n10084), .Z(n10375) );
  AND U11125 ( .A(\stack[1][12] ), .B(o[44]), .Z(n10374) );
  NAND U11126 ( .A(n10087), .B(n10086), .Z(n10091) );
  NAND U11127 ( .A(n10089), .B(n10088), .Z(n10090) );
  NAND U11128 ( .A(n10091), .B(n10090), .Z(n10380) );
  AND U11129 ( .A(\stack[1][14] ), .B(o[42]), .Z(n10381) );
  XOR U11130 ( .A(n10380), .B(n10381), .Z(n10383) );
  NAND U11131 ( .A(n10093), .B(n10092), .Z(n10097) );
  NAND U11132 ( .A(n10095), .B(n10094), .Z(n10096) );
  AND U11133 ( .A(n10097), .B(n10096), .Z(n10399) );
  NAND U11134 ( .A(\stack[1][20] ), .B(o[36]), .Z(n10398) );
  XOR U11135 ( .A(n10399), .B(n10398), .Z(n10400) );
  NAND U11136 ( .A(n10099), .B(n10098), .Z(n10103) );
  NAND U11137 ( .A(n10101), .B(n10100), .Z(n10102) );
  NAND U11138 ( .A(n10103), .B(n10102), .Z(n10606) );
  NAND U11139 ( .A(n10105), .B(n10104), .Z(n10109) );
  NAND U11140 ( .A(n10107), .B(n10106), .Z(n10108) );
  AND U11141 ( .A(n10109), .B(n10108), .Z(n10405) );
  NAND U11142 ( .A(\stack[1][22] ), .B(o[34]), .Z(n10404) );
  XOR U11143 ( .A(n10405), .B(n10404), .Z(n10407) );
  NAND U11144 ( .A(n10111), .B(n10110), .Z(n10115) );
  NAND U11145 ( .A(n10113), .B(n10112), .Z(n10114) );
  NAND U11146 ( .A(n10115), .B(n10114), .Z(n10600) );
  NAND U11147 ( .A(n10117), .B(n10116), .Z(n10121) );
  NAND U11148 ( .A(n10119), .B(n10118), .Z(n10120) );
  AND U11149 ( .A(n10121), .B(n10120), .Z(n10411) );
  NAND U11150 ( .A(\stack[1][24] ), .B(o[32]), .Z(n10410) );
  XOR U11151 ( .A(n10411), .B(n10410), .Z(n10413) );
  AND U11152 ( .A(\stack[1][28] ), .B(o[28]), .Z(n16251) );
  NAND U11153 ( .A(n10123), .B(n10122), .Z(n10127) );
  NAND U11154 ( .A(n10125), .B(n10124), .Z(n10126) );
  NAND U11155 ( .A(n10127), .B(n10126), .Z(n10422) );
  XOR U11156 ( .A(n16251), .B(n10422), .Z(n10424) );
  NAND U11157 ( .A(n10129), .B(n10128), .Z(n10133) );
  NAND U11158 ( .A(n10131), .B(n10130), .Z(n10132) );
  NAND U11159 ( .A(n10133), .B(n10132), .Z(n10582) );
  NAND U11160 ( .A(n10135), .B(n10134), .Z(n10139) );
  NAND U11161 ( .A(n10137), .B(n10136), .Z(n10138) );
  AND U11162 ( .A(n10139), .B(n10138), .Z(n10576) );
  NAND U11163 ( .A(o[26]), .B(\stack[1][30] ), .Z(n10575) );
  XOR U11164 ( .A(n10576), .B(n10575), .Z(n10578) );
  NAND U11165 ( .A(n10141), .B(n10140), .Z(n10145) );
  NAND U11166 ( .A(n10143), .B(n10142), .Z(n10144) );
  NAND U11167 ( .A(n10145), .B(n10144), .Z(n10433) );
  AND U11168 ( .A(o[24]), .B(\stack[1][32] ), .Z(n10434) );
  XOR U11169 ( .A(n10433), .B(n10434), .Z(n10436) );
  NAND U11170 ( .A(n10147), .B(n10146), .Z(n10151) );
  NAND U11171 ( .A(n10149), .B(n10148), .Z(n10150) );
  NAND U11172 ( .A(n10151), .B(n10150), .Z(n10439) );
  AND U11173 ( .A(o[22]), .B(\stack[1][34] ), .Z(n10440) );
  XOR U11174 ( .A(n10439), .B(n10440), .Z(n10442) );
  NAND U11175 ( .A(n10153), .B(n10152), .Z(n10157) );
  NANDN U11176 ( .A(n10155), .B(n10154), .Z(n10156) );
  NAND U11177 ( .A(n10157), .B(n10156), .Z(n10451) );
  AND U11178 ( .A(o[20]), .B(\stack[1][36] ), .Z(n10452) );
  XOR U11179 ( .A(n10451), .B(n10452), .Z(n10454) );
  NAND U11180 ( .A(n10159), .B(n10158), .Z(n10163) );
  NAND U11181 ( .A(n10161), .B(n10160), .Z(n10162) );
  NAND U11182 ( .A(n10163), .B(n10162), .Z(n10563) );
  AND U11183 ( .A(o[19]), .B(\stack[1][37] ), .Z(n10564) );
  XOR U11184 ( .A(n10563), .B(n10564), .Z(n10566) );
  AND U11185 ( .A(o[18]), .B(\stack[1][38] ), .Z(n10560) );
  NAND U11186 ( .A(n10165), .B(n10164), .Z(n10169) );
  NAND U11187 ( .A(n10167), .B(n10166), .Z(n10168) );
  AND U11188 ( .A(n10169), .B(n10168), .Z(n10558) );
  NAND U11189 ( .A(o[17]), .B(\stack[1][39] ), .Z(n10459) );
  NAND U11190 ( .A(n10171), .B(n10170), .Z(n10175) );
  NAND U11191 ( .A(n10173), .B(n10172), .Z(n10174) );
  NAND U11192 ( .A(n10175), .B(n10174), .Z(n10547) );
  NAND U11193 ( .A(n10177), .B(n10176), .Z(n10181) );
  NAND U11194 ( .A(n10179), .B(n10178), .Z(n10180) );
  AND U11195 ( .A(n10181), .B(n10180), .Z(n10465) );
  AND U11196 ( .A(o[13]), .B(\stack[1][43] ), .Z(n10471) );
  NAND U11197 ( .A(n10183), .B(n10182), .Z(n10187) );
  NAND U11198 ( .A(n10185), .B(n10184), .Z(n10186) );
  NAND U11199 ( .A(n10187), .B(n10186), .Z(n10469) );
  NAND U11200 ( .A(n10189), .B(n10188), .Z(n10193) );
  NAND U11201 ( .A(n10191), .B(n10190), .Z(n10192) );
  AND U11202 ( .A(n10193), .B(n10192), .Z(n10475) );
  NAND U11203 ( .A(o[11]), .B(\stack[1][45] ), .Z(n10483) );
  NAND U11204 ( .A(n10195), .B(n10194), .Z(n10199) );
  NAND U11205 ( .A(n10197), .B(n10196), .Z(n10198) );
  AND U11206 ( .A(n10199), .B(n10198), .Z(n10481) );
  AND U11207 ( .A(o[10]), .B(\stack[1][46] ), .Z(n10490) );
  NAND U11208 ( .A(n10201), .B(n10200), .Z(n10205) );
  NAND U11209 ( .A(n10203), .B(n10202), .Z(n10204) );
  AND U11210 ( .A(n10205), .B(n10204), .Z(n10488) );
  NAND U11211 ( .A(o[9]), .B(\stack[1][47] ), .Z(n10495) );
  NAND U11212 ( .A(n10207), .B(n10206), .Z(n10211) );
  NAND U11213 ( .A(n10209), .B(n10208), .Z(n10210) );
  NAND U11214 ( .A(n10211), .B(n10210), .Z(n10535) );
  AND U11215 ( .A(o[6]), .B(\stack[1][50] ), .Z(n10502) );
  NAND U11216 ( .A(n10213), .B(n10212), .Z(n10217) );
  NAND U11217 ( .A(n10215), .B(n10214), .Z(n10216) );
  NAND U11218 ( .A(n10217), .B(n10216), .Z(n10527) );
  AND U11219 ( .A(o[4]), .B(\stack[1][52] ), .Z(n10508) );
  NANDN U11220 ( .A(n10218), .B(n10511), .Z(n10222) );
  NANDN U11221 ( .A(n10220), .B(n10219), .Z(n10221) );
  NAND U11222 ( .A(n10222), .B(n10221), .Z(n10521) );
  AND U11223 ( .A(o[2]), .B(\stack[1][54] ), .Z(n10512) );
  AND U11224 ( .A(n10223), .B(n10225), .Z(n10224) );
  AND U11225 ( .A(o[1]), .B(\stack[1][56] ), .Z(n10518) );
  NAND U11226 ( .A(n10516), .B(n10518), .Z(n10781) );
  XOR U11227 ( .A(n10224), .B(n10781), .Z(n10227) );
  AND U11228 ( .A(o[0]), .B(\stack[1][56] ), .Z(n10786) );
  OR U11229 ( .A(n10225), .B(n10786), .Z(n10226) );
  NAND U11230 ( .A(n10227), .B(n10226), .Z(n10513) );
  XNOR U11231 ( .A(n10512), .B(n10513), .Z(n10522) );
  XOR U11232 ( .A(n10521), .B(n10522), .Z(n10524) );
  AND U11233 ( .A(o[3]), .B(\stack[1][53] ), .Z(n10523) );
  XOR U11234 ( .A(n10524), .B(n10523), .Z(n10506) );
  NAND U11235 ( .A(n10229), .B(n10228), .Z(n10233) );
  NAND U11236 ( .A(n10231), .B(n10230), .Z(n10232) );
  NAND U11237 ( .A(n10233), .B(n10232), .Z(n10505) );
  XOR U11238 ( .A(n10506), .B(n10505), .Z(n10507) );
  XOR U11239 ( .A(n10508), .B(n10507), .Z(n10528) );
  XOR U11240 ( .A(n10527), .B(n10528), .Z(n10530) );
  AND U11241 ( .A(o[5]), .B(\stack[1][51] ), .Z(n10529) );
  XOR U11242 ( .A(n10530), .B(n10529), .Z(n10500) );
  NAND U11243 ( .A(n10235), .B(n10234), .Z(n10239) );
  NAND U11244 ( .A(n10237), .B(n10236), .Z(n10238) );
  NAND U11245 ( .A(n10239), .B(n10238), .Z(n10499) );
  XOR U11246 ( .A(n10500), .B(n10499), .Z(n10501) );
  XOR U11247 ( .A(n10502), .B(n10501), .Z(n10534) );
  AND U11248 ( .A(o[7]), .B(\stack[1][49] ), .Z(n10533) );
  XOR U11249 ( .A(n10534), .B(n10533), .Z(n10536) );
  XOR U11250 ( .A(n10535), .B(n10536), .Z(n10540) );
  AND U11251 ( .A(o[8]), .B(\stack[1][48] ), .Z(n10539) );
  XOR U11252 ( .A(n10540), .B(n10539), .Z(n10542) );
  NAND U11253 ( .A(n10241), .B(n10240), .Z(n10245) );
  NAND U11254 ( .A(n10243), .B(n10242), .Z(n10244) );
  NAND U11255 ( .A(n10245), .B(n10244), .Z(n10541) );
  XNOR U11256 ( .A(n10542), .B(n10541), .Z(n10494) );
  NAND U11257 ( .A(n10247), .B(n10246), .Z(n10251) );
  NAND U11258 ( .A(n10249), .B(n10248), .Z(n10250) );
  AND U11259 ( .A(n10251), .B(n10250), .Z(n10493) );
  XOR U11260 ( .A(n10495), .B(n10496), .Z(n10487) );
  XOR U11261 ( .A(n10488), .B(n10487), .Z(n10489) );
  XNOR U11262 ( .A(n10490), .B(n10489), .Z(n10482) );
  XNOR U11263 ( .A(n10483), .B(n10484), .Z(n10476) );
  AND U11264 ( .A(o[12]), .B(\stack[1][44] ), .Z(n10477) );
  XOR U11265 ( .A(n10478), .B(n10477), .Z(n10470) );
  XOR U11266 ( .A(n10469), .B(n10470), .Z(n10472) );
  NAND U11267 ( .A(o[14]), .B(\stack[1][42] ), .Z(n10463) );
  XOR U11268 ( .A(n10465), .B(n10466), .Z(n10546) );
  AND U11269 ( .A(o[15]), .B(\stack[1][41] ), .Z(n10545) );
  XOR U11270 ( .A(n10547), .B(n10548), .Z(n10552) );
  AND U11271 ( .A(o[16]), .B(\stack[1][40] ), .Z(n10551) );
  XOR U11272 ( .A(n10552), .B(n10551), .Z(n10554) );
  NAND U11273 ( .A(n10253), .B(n10252), .Z(n10257) );
  NAND U11274 ( .A(n10255), .B(n10254), .Z(n10256) );
  NAND U11275 ( .A(n10257), .B(n10256), .Z(n10553) );
  XNOR U11276 ( .A(n10554), .B(n10553), .Z(n10458) );
  NAND U11277 ( .A(n10259), .B(n10258), .Z(n10263) );
  NAND U11278 ( .A(n10261), .B(n10260), .Z(n10262) );
  AND U11279 ( .A(n10263), .B(n10262), .Z(n10457) );
  XOR U11280 ( .A(n10459), .B(n10460), .Z(n10557) );
  XOR U11281 ( .A(n10558), .B(n10557), .Z(n10559) );
  XOR U11282 ( .A(n10560), .B(n10559), .Z(n10565) );
  XOR U11283 ( .A(n10566), .B(n10565), .Z(n10453) );
  XOR U11284 ( .A(n10454), .B(n10453), .Z(n10448) );
  AND U11285 ( .A(o[21]), .B(\stack[1][35] ), .Z(n10446) );
  NAND U11286 ( .A(n10265), .B(n10264), .Z(n10269) );
  NAND U11287 ( .A(n10267), .B(n10266), .Z(n10268) );
  NAND U11288 ( .A(n10269), .B(n10268), .Z(n10445) );
  XOR U11289 ( .A(n10446), .B(n10445), .Z(n10447) );
  XOR U11290 ( .A(n10448), .B(n10447), .Z(n10441) );
  XOR U11291 ( .A(n10442), .B(n10441), .Z(n10570) );
  NAND U11292 ( .A(n10271), .B(n10270), .Z(n10275) );
  NAND U11293 ( .A(n10273), .B(n10272), .Z(n10274) );
  NAND U11294 ( .A(n10275), .B(n10274), .Z(n10569) );
  XOR U11295 ( .A(n10570), .B(n10569), .Z(n10572) );
  AND U11296 ( .A(o[23]), .B(\stack[1][33] ), .Z(n10571) );
  XOR U11297 ( .A(n10572), .B(n10571), .Z(n10435) );
  XOR U11298 ( .A(n10436), .B(n10435), .Z(n10428) );
  NAND U11299 ( .A(n10277), .B(n10276), .Z(n10281) );
  NAND U11300 ( .A(n10279), .B(n10278), .Z(n10280) );
  NAND U11301 ( .A(n10281), .B(n10280), .Z(n10427) );
  XOR U11302 ( .A(n10428), .B(n10427), .Z(n10430) );
  AND U11303 ( .A(o[25]), .B(\stack[1][31] ), .Z(n10429) );
  XNOR U11304 ( .A(n10430), .B(n10429), .Z(n10577) );
  XNOR U11305 ( .A(n10578), .B(n10577), .Z(n10581) );
  XOR U11306 ( .A(n10582), .B(n10581), .Z(n10584) );
  AND U11307 ( .A(\stack[1][29] ), .B(o[27]), .Z(n10583) );
  XOR U11308 ( .A(n10584), .B(n10583), .Z(n10423) );
  XOR U11309 ( .A(n10424), .B(n10423), .Z(n10588) );
  NAND U11310 ( .A(n10283), .B(n10282), .Z(n10287) );
  NAND U11311 ( .A(n10285), .B(n10284), .Z(n10286) );
  NAND U11312 ( .A(n10287), .B(n10286), .Z(n10587) );
  XOR U11313 ( .A(n10588), .B(n10587), .Z(n10590) );
  AND U11314 ( .A(\stack[1][27] ), .B(o[29]), .Z(n10589) );
  XOR U11315 ( .A(n10590), .B(n10589), .Z(n10418) );
  NAND U11316 ( .A(n10289), .B(n10288), .Z(n10293) );
  NAND U11317 ( .A(n10291), .B(n10290), .Z(n10292) );
  NAND U11318 ( .A(n10293), .B(n10292), .Z(n10416) );
  AND U11319 ( .A(\stack[1][26] ), .B(o[30]), .Z(n10417) );
  XOR U11320 ( .A(n10416), .B(n10417), .Z(n10419) );
  NAND U11321 ( .A(n10295), .B(n10294), .Z(n10299) );
  NAND U11322 ( .A(n10297), .B(n10296), .Z(n10298) );
  NAND U11323 ( .A(n10299), .B(n10298), .Z(n10593) );
  XOR U11324 ( .A(n10594), .B(n10593), .Z(n10596) );
  AND U11325 ( .A(\stack[1][25] ), .B(o[31]), .Z(n10595) );
  XNOR U11326 ( .A(n10596), .B(n10595), .Z(n10412) );
  XNOR U11327 ( .A(n10413), .B(n10412), .Z(n10599) );
  XOR U11328 ( .A(n10600), .B(n10599), .Z(n10602) );
  AND U11329 ( .A(\stack[1][23] ), .B(o[33]), .Z(n10601) );
  XNOR U11330 ( .A(n10602), .B(n10601), .Z(n10406) );
  XNOR U11331 ( .A(n10407), .B(n10406), .Z(n10605) );
  XOR U11332 ( .A(n10606), .B(n10605), .Z(n10608) );
  AND U11333 ( .A(\stack[1][21] ), .B(o[35]), .Z(n10607) );
  XNOR U11334 ( .A(n10608), .B(n10607), .Z(n10401) );
  NAND U11335 ( .A(n10301), .B(n10300), .Z(n10305) );
  NAND U11336 ( .A(n10303), .B(n10302), .Z(n10304) );
  NAND U11337 ( .A(n10305), .B(n10304), .Z(n10611) );
  AND U11338 ( .A(\stack[1][19] ), .B(o[37]), .Z(n10613) );
  XNOR U11339 ( .A(n10614), .B(n10613), .Z(n10395) );
  NAND U11340 ( .A(n10307), .B(n10306), .Z(n10311) );
  NAND U11341 ( .A(n10309), .B(n10308), .Z(n10310) );
  AND U11342 ( .A(n10311), .B(n10310), .Z(n10393) );
  NAND U11343 ( .A(\stack[1][18] ), .B(o[38]), .Z(n10392) );
  XOR U11344 ( .A(n10393), .B(n10392), .Z(n10394) );
  NAND U11345 ( .A(n10313), .B(n10312), .Z(n10317) );
  NAND U11346 ( .A(n10315), .B(n10314), .Z(n10316) );
  NAND U11347 ( .A(n10317), .B(n10316), .Z(n10617) );
  AND U11348 ( .A(\stack[1][17] ), .B(o[39]), .Z(n10619) );
  XNOR U11349 ( .A(n10620), .B(n10619), .Z(n10389) );
  NAND U11350 ( .A(n10319), .B(n10318), .Z(n10323) );
  NAND U11351 ( .A(n10321), .B(n10320), .Z(n10322) );
  AND U11352 ( .A(n10323), .B(n10322), .Z(n10387) );
  NAND U11353 ( .A(\stack[1][16] ), .B(o[40]), .Z(n10386) );
  XOR U11354 ( .A(n10387), .B(n10386), .Z(n10388) );
  NAND U11355 ( .A(n10325), .B(n10324), .Z(n10329) );
  NAND U11356 ( .A(n10327), .B(n10326), .Z(n10328) );
  NAND U11357 ( .A(n10329), .B(n10328), .Z(n10623) );
  AND U11358 ( .A(\stack[1][15] ), .B(o[41]), .Z(n10625) );
  XOR U11359 ( .A(n10626), .B(n10625), .Z(n10382) );
  XOR U11360 ( .A(n10383), .B(n10382), .Z(n10630) );
  NAND U11361 ( .A(n10331), .B(n10330), .Z(n10335) );
  NAND U11362 ( .A(n10333), .B(n10332), .Z(n10334) );
  NAND U11363 ( .A(n10335), .B(n10334), .Z(n10629) );
  XOR U11364 ( .A(n10630), .B(n10629), .Z(n10632) );
  AND U11365 ( .A(\stack[1][13] ), .B(o[43]), .Z(n10631) );
  XOR U11366 ( .A(n10632), .B(n10631), .Z(n10376) );
  XOR U11367 ( .A(n10377), .B(n10376), .Z(n10635) );
  NAND U11368 ( .A(n10337), .B(n10336), .Z(n10341) );
  NAND U11369 ( .A(n10339), .B(n10338), .Z(n10340) );
  NAND U11370 ( .A(n10341), .B(n10340), .Z(n10636) );
  AND U11371 ( .A(\stack[1][11] ), .B(o[45]), .Z(n10638) );
  XOR U11372 ( .A(n10371), .B(n10370), .Z(n10641) );
  NAND U11373 ( .A(n10343), .B(n10342), .Z(n10347) );
  NAND U11374 ( .A(n10345), .B(n10344), .Z(n10346) );
  NAND U11375 ( .A(n10347), .B(n10346), .Z(n10642) );
  AND U11376 ( .A(\stack[1][9] ), .B(o[47]), .Z(n10644) );
  NAND U11377 ( .A(n10349), .B(n10348), .Z(n10353) );
  NAND U11378 ( .A(n10351), .B(n10350), .Z(n10352) );
  NAND U11379 ( .A(n10353), .B(n10352), .Z(n10363) );
  AND U11380 ( .A(\stack[1][8] ), .B(o[48]), .Z(n10362) );
  XOR U11381 ( .A(n10365), .B(n10364), .Z(n10648) );
  NAND U11382 ( .A(n10355), .B(n10354), .Z(n10359) );
  NAND U11383 ( .A(n10357), .B(n10356), .Z(n10358) );
  NAND U11384 ( .A(n10359), .B(n10358), .Z(n10649) );
  AND U11385 ( .A(\stack[1][7] ), .B(o[49]), .Z(n10650) );
  XNOR U11386 ( .A(n10651), .B(n10650), .Z(n12518) );
  NAND U11387 ( .A(n12519), .B(n12518), .Z(n10360) );
  AND U11388 ( .A(n10361), .B(n10360), .Z(n10656) );
  NAND U11389 ( .A(n10363), .B(n10362), .Z(n10367) );
  NAND U11390 ( .A(n10365), .B(n10364), .Z(n10366) );
  NAND U11391 ( .A(n10367), .B(n10366), .Z(n10662) );
  NAND U11392 ( .A(n10369), .B(n10368), .Z(n10373) );
  NAND U11393 ( .A(n10371), .B(n10370), .Z(n10372) );
  NAND U11394 ( .A(n10373), .B(n10372), .Z(n10942) );
  NAND U11395 ( .A(n10375), .B(n10374), .Z(n10379) );
  NAND U11396 ( .A(n10377), .B(n10376), .Z(n10378) );
  NAND U11397 ( .A(n10379), .B(n10378), .Z(n10673) );
  NAND U11398 ( .A(n10381), .B(n10380), .Z(n10385) );
  NAND U11399 ( .A(n10383), .B(n10382), .Z(n10384) );
  NAND U11400 ( .A(n10385), .B(n10384), .Z(n10679) );
  AND U11401 ( .A(\stack[1][16] ), .B(o[41]), .Z(n10688) );
  NAND U11402 ( .A(n10387), .B(n10386), .Z(n10391) );
  NAND U11403 ( .A(n10389), .B(n10388), .Z(n10390) );
  AND U11404 ( .A(n10391), .B(n10390), .Z(n10686) );
  NAND U11405 ( .A(n10393), .B(n10392), .Z(n10397) );
  NAND U11406 ( .A(n10395), .B(n10394), .Z(n10396) );
  AND U11407 ( .A(n10397), .B(n10396), .Z(n10692) );
  AND U11408 ( .A(\stack[1][20] ), .B(o[37]), .Z(n10706) );
  NAND U11409 ( .A(n10399), .B(n10398), .Z(n10403) );
  NAND U11410 ( .A(n10401), .B(n10400), .Z(n10402) );
  AND U11411 ( .A(n10403), .B(n10402), .Z(n10704) );
  NAND U11412 ( .A(n10405), .B(n10404), .Z(n10409) );
  NAND U11413 ( .A(n10407), .B(n10406), .Z(n10408) );
  AND U11414 ( .A(n10409), .B(n10408), .Z(n10912) );
  AND U11415 ( .A(\stack[1][24] ), .B(o[33]), .Z(n10902) );
  NAND U11416 ( .A(n10411), .B(n10410), .Z(n10415) );
  NAND U11417 ( .A(n10413), .B(n10412), .Z(n10414) );
  AND U11418 ( .A(n10415), .B(n10414), .Z(n10900) );
  NAND U11419 ( .A(n10417), .B(n10416), .Z(n10421) );
  NAND U11420 ( .A(n10419), .B(n10418), .Z(n10420) );
  NAND U11421 ( .A(n10421), .B(n10420), .Z(n10709) );
  NAND U11422 ( .A(n16251), .B(n10422), .Z(n10426) );
  NAND U11423 ( .A(n10424), .B(n10423), .Z(n10425) );
  NAND U11424 ( .A(n10426), .B(n10425), .Z(n10715) );
  AND U11425 ( .A(o[27]), .B(\stack[1][30] ), .Z(n10724) );
  AND U11426 ( .A(o[26]), .B(\stack[1][31] ), .Z(n10876) );
  NAND U11427 ( .A(n10428), .B(n10427), .Z(n10432) );
  NAND U11428 ( .A(n10430), .B(n10429), .Z(n10431) );
  NAND U11429 ( .A(n10432), .B(n10431), .Z(n10875) );
  XOR U11430 ( .A(n10876), .B(n10875), .Z(n10878) );
  NAND U11431 ( .A(n10434), .B(n10433), .Z(n10438) );
  NAND U11432 ( .A(n10436), .B(n10435), .Z(n10437) );
  NAND U11433 ( .A(n10438), .B(n10437), .Z(n10727) );
  AND U11434 ( .A(o[23]), .B(\stack[1][34] ), .Z(n10735) );
  NAND U11435 ( .A(n10440), .B(n10439), .Z(n10444) );
  NAND U11436 ( .A(n10442), .B(n10441), .Z(n10443) );
  NAND U11437 ( .A(n10444), .B(n10443), .Z(n10733) );
  NAND U11438 ( .A(n10446), .B(n10445), .Z(n10450) );
  NAND U11439 ( .A(n10448), .B(n10447), .Z(n10449) );
  NAND U11440 ( .A(n10450), .B(n10449), .Z(n10865) );
  NAND U11441 ( .A(n10452), .B(n10451), .Z(n10456) );
  NAND U11442 ( .A(n10454), .B(n10453), .Z(n10455) );
  NAND U11443 ( .A(n10456), .B(n10455), .Z(n10857) );
  NAND U11444 ( .A(o[19]), .B(\stack[1][38] ), .Z(n10741) );
  NAND U11445 ( .A(n10458), .B(n10457), .Z(n10462) );
  NANDN U11446 ( .A(n10460), .B(n10459), .Z(n10461) );
  AND U11447 ( .A(n10462), .B(n10461), .Z(n10845) );
  NAND U11448 ( .A(o[17]), .B(\stack[1][40] ), .Z(n10747) );
  NAND U11449 ( .A(n10464), .B(n10463), .Z(n10468) );
  NANDN U11450 ( .A(n10466), .B(n10465), .Z(n10467) );
  AND U11451 ( .A(n10468), .B(n10467), .Z(n10836) );
  NAND U11452 ( .A(n10470), .B(n10469), .Z(n10474) );
  NAND U11453 ( .A(n10472), .B(n10471), .Z(n10473) );
  NAND U11454 ( .A(n10474), .B(n10473), .Z(n10753) );
  AND U11455 ( .A(o[13]), .B(\stack[1][44] ), .Z(n10829) );
  NAND U11456 ( .A(n10476), .B(n10475), .Z(n10480) );
  NAND U11457 ( .A(n10478), .B(n10477), .Z(n10479) );
  NAND U11458 ( .A(n10480), .B(n10479), .Z(n10827) );
  AND U11459 ( .A(o[12]), .B(\stack[1][45] ), .Z(n10824) );
  NAND U11460 ( .A(n10482), .B(n10481), .Z(n10486) );
  NAND U11461 ( .A(n10484), .B(n10483), .Z(n10485) );
  AND U11462 ( .A(n10486), .B(n10485), .Z(n10821) );
  NAND U11463 ( .A(o[11]), .B(\stack[1][46] ), .Z(n10759) );
  NAND U11464 ( .A(n10488), .B(n10487), .Z(n10492) );
  NAND U11465 ( .A(n10490), .B(n10489), .Z(n10491) );
  AND U11466 ( .A(n10492), .B(n10491), .Z(n10757) );
  NAND U11467 ( .A(n10494), .B(n10493), .Z(n10498) );
  NANDN U11468 ( .A(n10496), .B(n10495), .Z(n10497) );
  AND U11469 ( .A(n10498), .B(n10497), .Z(n10763) );
  NAND U11470 ( .A(o[9]), .B(\stack[1][48] ), .Z(n10771) );
  NAND U11471 ( .A(n10500), .B(n10499), .Z(n10504) );
  NAND U11472 ( .A(n10502), .B(n10501), .Z(n10503) );
  NAND U11473 ( .A(n10504), .B(n10503), .Z(n10811) );
  AND U11474 ( .A(o[6]), .B(\stack[1][51] ), .Z(n10778) );
  NAND U11475 ( .A(n10506), .B(n10505), .Z(n10510) );
  NAND U11476 ( .A(n10508), .B(n10507), .Z(n10509) );
  NAND U11477 ( .A(n10510), .B(n10509), .Z(n10803) );
  AND U11478 ( .A(o[4]), .B(\stack[1][53] ), .Z(n10800) );
  NANDN U11479 ( .A(n10511), .B(n10781), .Z(n10515) );
  NANDN U11480 ( .A(n10513), .B(n10512), .Z(n10514) );
  NAND U11481 ( .A(n10515), .B(n10514), .Z(n10791) );
  AND U11482 ( .A(o[2]), .B(\stack[1][55] ), .Z(n10782) );
  AND U11483 ( .A(n10516), .B(n10518), .Z(n10517) );
  AND U11484 ( .A(o[1]), .B(\stack[1][57] ), .Z(n10788) );
  NAND U11485 ( .A(n10786), .B(n10788), .Z(n11117) );
  XOR U11486 ( .A(n10517), .B(n11117), .Z(n10520) );
  AND U11487 ( .A(o[0]), .B(\stack[1][57] ), .Z(n11122) );
  OR U11488 ( .A(n10518), .B(n11122), .Z(n10519) );
  NAND U11489 ( .A(n10520), .B(n10519), .Z(n10783) );
  XNOR U11490 ( .A(n10782), .B(n10783), .Z(n10792) );
  XOR U11491 ( .A(n10791), .B(n10792), .Z(n10794) );
  AND U11492 ( .A(o[3]), .B(\stack[1][54] ), .Z(n10793) );
  XOR U11493 ( .A(n10794), .B(n10793), .Z(n10798) );
  NAND U11494 ( .A(n10522), .B(n10521), .Z(n10526) );
  NAND U11495 ( .A(n10524), .B(n10523), .Z(n10525) );
  NAND U11496 ( .A(n10526), .B(n10525), .Z(n10797) );
  XOR U11497 ( .A(n10798), .B(n10797), .Z(n10799) );
  XOR U11498 ( .A(n10800), .B(n10799), .Z(n10804) );
  XOR U11499 ( .A(n10803), .B(n10804), .Z(n10806) );
  AND U11500 ( .A(o[5]), .B(\stack[1][52] ), .Z(n10805) );
  XOR U11501 ( .A(n10806), .B(n10805), .Z(n10776) );
  NAND U11502 ( .A(n10528), .B(n10527), .Z(n10532) );
  NAND U11503 ( .A(n10530), .B(n10529), .Z(n10531) );
  NAND U11504 ( .A(n10532), .B(n10531), .Z(n10775) );
  XOR U11505 ( .A(n10776), .B(n10775), .Z(n10777) );
  XOR U11506 ( .A(n10778), .B(n10777), .Z(n10810) );
  AND U11507 ( .A(o[7]), .B(\stack[1][50] ), .Z(n10809) );
  XOR U11508 ( .A(n10810), .B(n10809), .Z(n10812) );
  XOR U11509 ( .A(n10811), .B(n10812), .Z(n10816) );
  AND U11510 ( .A(o[8]), .B(\stack[1][49] ), .Z(n10815) );
  XOR U11511 ( .A(n10816), .B(n10815), .Z(n10818) );
  NAND U11512 ( .A(n10534), .B(n10533), .Z(n10538) );
  NAND U11513 ( .A(n10536), .B(n10535), .Z(n10537) );
  NAND U11514 ( .A(n10538), .B(n10537), .Z(n10817) );
  XNOR U11515 ( .A(n10818), .B(n10817), .Z(n10770) );
  NAND U11516 ( .A(n10540), .B(n10539), .Z(n10544) );
  NAND U11517 ( .A(n10542), .B(n10541), .Z(n10543) );
  AND U11518 ( .A(n10544), .B(n10543), .Z(n10769) );
  XNOR U11519 ( .A(n10771), .B(n10772), .Z(n10764) );
  AND U11520 ( .A(o[10]), .B(\stack[1][47] ), .Z(n10765) );
  XNOR U11521 ( .A(n10766), .B(n10765), .Z(n10758) );
  XNOR U11522 ( .A(n10759), .B(n10760), .Z(n10822) );
  XOR U11523 ( .A(n10824), .B(n10823), .Z(n10828) );
  XOR U11524 ( .A(n10827), .B(n10828), .Z(n10830) );
  AND U11525 ( .A(o[14]), .B(\stack[1][43] ), .Z(n10751) );
  XOR U11526 ( .A(n10752), .B(n10751), .Z(n10754) );
  XOR U11527 ( .A(n10753), .B(n10754), .Z(n10834) );
  AND U11528 ( .A(o[15]), .B(\stack[1][42] ), .Z(n10833) );
  XOR U11529 ( .A(n10834), .B(n10833), .Z(n10835) );
  XOR U11530 ( .A(n10836), .B(n10835), .Z(n10840) );
  AND U11531 ( .A(o[16]), .B(\stack[1][41] ), .Z(n10839) );
  XOR U11532 ( .A(n10840), .B(n10839), .Z(n10842) );
  NAND U11533 ( .A(n10546), .B(n10545), .Z(n10550) );
  NAND U11534 ( .A(n10548), .B(n10547), .Z(n10549) );
  NAND U11535 ( .A(n10550), .B(n10549), .Z(n10841) );
  XNOR U11536 ( .A(n10842), .B(n10841), .Z(n10746) );
  NAND U11537 ( .A(n10552), .B(n10551), .Z(n10556) );
  NAND U11538 ( .A(n10554), .B(n10553), .Z(n10555) );
  AND U11539 ( .A(n10556), .B(n10555), .Z(n10745) );
  XNOR U11540 ( .A(n10747), .B(n10748), .Z(n10846) );
  AND U11541 ( .A(o[18]), .B(\stack[1][39] ), .Z(n10847) );
  XNOR U11542 ( .A(n10848), .B(n10847), .Z(n10740) );
  NAND U11543 ( .A(n10558), .B(n10557), .Z(n10562) );
  NAND U11544 ( .A(n10560), .B(n10559), .Z(n10561) );
  AND U11545 ( .A(n10562), .B(n10561), .Z(n10739) );
  XNOR U11546 ( .A(n10741), .B(n10742), .Z(n10854) );
  AND U11547 ( .A(o[20]), .B(\stack[1][37] ), .Z(n10852) );
  NAND U11548 ( .A(n10564), .B(n10563), .Z(n10568) );
  NAND U11549 ( .A(n10566), .B(n10565), .Z(n10567) );
  NAND U11550 ( .A(n10568), .B(n10567), .Z(n10851) );
  XOR U11551 ( .A(n10852), .B(n10851), .Z(n10853) );
  XOR U11552 ( .A(n10857), .B(n10858), .Z(n10860) );
  AND U11553 ( .A(o[21]), .B(\stack[1][36] ), .Z(n10859) );
  XOR U11554 ( .A(n10860), .B(n10859), .Z(n10864) );
  AND U11555 ( .A(o[22]), .B(\stack[1][35] ), .Z(n10863) );
  XOR U11556 ( .A(n10864), .B(n10863), .Z(n10866) );
  XOR U11557 ( .A(n10865), .B(n10866), .Z(n10734) );
  XNOR U11558 ( .A(n10735), .B(n10736), .Z(n10872) );
  AND U11559 ( .A(o[24]), .B(\stack[1][33] ), .Z(n10870) );
  NAND U11560 ( .A(n10570), .B(n10569), .Z(n10574) );
  NAND U11561 ( .A(n10572), .B(n10571), .Z(n10573) );
  NAND U11562 ( .A(n10574), .B(n10573), .Z(n10869) );
  XOR U11563 ( .A(n10870), .B(n10869), .Z(n10871) );
  XOR U11564 ( .A(n10872), .B(n10871), .Z(n10728) );
  XOR U11565 ( .A(n10727), .B(n10728), .Z(n10730) );
  AND U11566 ( .A(o[25]), .B(\stack[1][32] ), .Z(n10729) );
  XOR U11567 ( .A(n10730), .B(n10729), .Z(n10877) );
  XOR U11568 ( .A(n10878), .B(n10877), .Z(n10722) );
  NAND U11569 ( .A(n10576), .B(n10575), .Z(n10580) );
  NAND U11570 ( .A(n10578), .B(n10577), .Z(n10579) );
  AND U11571 ( .A(n10580), .B(n10579), .Z(n10721) );
  XOR U11572 ( .A(n10722), .B(n10721), .Z(n10723) );
  XOR U11573 ( .A(n10724), .B(n10723), .Z(n10884) );
  AND U11574 ( .A(\stack[1][29] ), .B(o[28]), .Z(n10882) );
  NAND U11575 ( .A(n10582), .B(n10581), .Z(n10586) );
  NAND U11576 ( .A(n10584), .B(n10583), .Z(n10585) );
  NAND U11577 ( .A(n10586), .B(n10585), .Z(n10881) );
  XOR U11578 ( .A(n10882), .B(n10881), .Z(n10883) );
  XOR U11579 ( .A(n10884), .B(n10883), .Z(n10716) );
  XOR U11580 ( .A(n10715), .B(n10716), .Z(n10718) );
  AND U11581 ( .A(\stack[1][28] ), .B(o[29]), .Z(n10717) );
  XOR U11582 ( .A(n10718), .B(n10717), .Z(n10890) );
  AND U11583 ( .A(\stack[1][27] ), .B(o[30]), .Z(n10888) );
  NAND U11584 ( .A(n10588), .B(n10587), .Z(n10592) );
  NAND U11585 ( .A(n10590), .B(n10589), .Z(n10591) );
  NAND U11586 ( .A(n10592), .B(n10591), .Z(n10887) );
  XOR U11587 ( .A(n10888), .B(n10887), .Z(n10889) );
  XOR U11588 ( .A(n10890), .B(n10889), .Z(n10710) );
  XOR U11589 ( .A(n10709), .B(n10710), .Z(n10712) );
  AND U11590 ( .A(\stack[1][26] ), .B(o[31]), .Z(n10711) );
  XOR U11591 ( .A(n10712), .B(n10711), .Z(n10896) );
  AND U11592 ( .A(\stack[1][25] ), .B(o[32]), .Z(n10894) );
  NAND U11593 ( .A(n10594), .B(n10593), .Z(n10598) );
  NAND U11594 ( .A(n10596), .B(n10595), .Z(n10597) );
  NAND U11595 ( .A(n10598), .B(n10597), .Z(n10893) );
  XOR U11596 ( .A(n10894), .B(n10893), .Z(n10895) );
  XOR U11597 ( .A(n10896), .B(n10895), .Z(n10899) );
  XOR U11598 ( .A(n10900), .B(n10899), .Z(n10901) );
  XOR U11599 ( .A(n10902), .B(n10901), .Z(n10908) );
  AND U11600 ( .A(\stack[1][23] ), .B(o[34]), .Z(n10906) );
  NAND U11601 ( .A(n10600), .B(n10599), .Z(n10604) );
  NAND U11602 ( .A(n10602), .B(n10601), .Z(n10603) );
  NAND U11603 ( .A(n10604), .B(n10603), .Z(n10905) );
  XOR U11604 ( .A(n10906), .B(n10905), .Z(n10907) );
  XOR U11605 ( .A(n10908), .B(n10907), .Z(n10911) );
  XOR U11606 ( .A(n10912), .B(n10911), .Z(n10914) );
  AND U11607 ( .A(\stack[1][22] ), .B(o[35]), .Z(n10913) );
  XOR U11608 ( .A(n10914), .B(n10913), .Z(n10920) );
  AND U11609 ( .A(\stack[1][21] ), .B(o[36]), .Z(n10918) );
  NAND U11610 ( .A(n10606), .B(n10605), .Z(n10610) );
  NAND U11611 ( .A(n10608), .B(n10607), .Z(n10609) );
  NAND U11612 ( .A(n10610), .B(n10609), .Z(n10917) );
  XOR U11613 ( .A(n10918), .B(n10917), .Z(n10919) );
  XOR U11614 ( .A(n10920), .B(n10919), .Z(n10703) );
  XOR U11615 ( .A(n10704), .B(n10703), .Z(n10705) );
  XOR U11616 ( .A(n10706), .B(n10705), .Z(n10700) );
  AND U11617 ( .A(\stack[1][19] ), .B(o[38]), .Z(n10698) );
  NAND U11618 ( .A(n10612), .B(n10611), .Z(n10616) );
  NAND U11619 ( .A(n10614), .B(n10613), .Z(n10615) );
  NAND U11620 ( .A(n10616), .B(n10615), .Z(n10697) );
  XOR U11621 ( .A(n10698), .B(n10697), .Z(n10699) );
  XOR U11622 ( .A(n10700), .B(n10699), .Z(n10691) );
  XOR U11623 ( .A(n10692), .B(n10691), .Z(n10694) );
  AND U11624 ( .A(\stack[1][18] ), .B(o[39]), .Z(n10693) );
  XOR U11625 ( .A(n10694), .B(n10693), .Z(n10926) );
  AND U11626 ( .A(\stack[1][17] ), .B(o[40]), .Z(n10924) );
  NAND U11627 ( .A(n10618), .B(n10617), .Z(n10622) );
  NAND U11628 ( .A(n10620), .B(n10619), .Z(n10621) );
  NAND U11629 ( .A(n10622), .B(n10621), .Z(n10923) );
  XOR U11630 ( .A(n10924), .B(n10923), .Z(n10925) );
  XOR U11631 ( .A(n10926), .B(n10925), .Z(n10685) );
  XOR U11632 ( .A(n10686), .B(n10685), .Z(n10687) );
  XOR U11633 ( .A(n10688), .B(n10687), .Z(n10932) );
  AND U11634 ( .A(\stack[1][15] ), .B(o[42]), .Z(n10930) );
  NAND U11635 ( .A(n10624), .B(n10623), .Z(n10628) );
  NAND U11636 ( .A(n10626), .B(n10625), .Z(n10627) );
  NAND U11637 ( .A(n10628), .B(n10627), .Z(n10929) );
  XOR U11638 ( .A(n10930), .B(n10929), .Z(n10931) );
  XOR U11639 ( .A(n10932), .B(n10931), .Z(n10680) );
  XOR U11640 ( .A(n10679), .B(n10680), .Z(n10682) );
  AND U11641 ( .A(\stack[1][14] ), .B(o[43]), .Z(n10681) );
  XOR U11642 ( .A(n10682), .B(n10681), .Z(n10938) );
  AND U11643 ( .A(\stack[1][13] ), .B(o[44]), .Z(n10936) );
  NAND U11644 ( .A(n10630), .B(n10629), .Z(n10634) );
  NAND U11645 ( .A(n10632), .B(n10631), .Z(n10633) );
  NAND U11646 ( .A(n10634), .B(n10633), .Z(n10935) );
  XOR U11647 ( .A(n10936), .B(n10935), .Z(n10937) );
  XOR U11648 ( .A(n10938), .B(n10937), .Z(n10674) );
  XOR U11649 ( .A(n10673), .B(n10674), .Z(n10676) );
  AND U11650 ( .A(\stack[1][12] ), .B(o[45]), .Z(n10675) );
  XOR U11651 ( .A(n10676), .B(n10675), .Z(n10670) );
  AND U11652 ( .A(\stack[1][11] ), .B(o[46]), .Z(n10668) );
  NAND U11653 ( .A(n10636), .B(n10635), .Z(n10640) );
  NAND U11654 ( .A(n10638), .B(n10637), .Z(n10639) );
  NAND U11655 ( .A(n10640), .B(n10639), .Z(n10667) );
  XOR U11656 ( .A(n10668), .B(n10667), .Z(n10669) );
  XOR U11657 ( .A(n10670), .B(n10669), .Z(n10941) );
  AND U11658 ( .A(\stack[1][10] ), .B(o[47]), .Z(n10944) );
  AND U11659 ( .A(\stack[1][9] ), .B(o[48]), .Z(n10947) );
  NAND U11660 ( .A(n10642), .B(n10641), .Z(n10646) );
  NAND U11661 ( .A(n10644), .B(n10643), .Z(n10645) );
  NAND U11662 ( .A(n10646), .B(n10645), .Z(n10948) );
  XOR U11663 ( .A(n10950), .B(n10949), .Z(n10661) );
  AND U11664 ( .A(\stack[1][8] ), .B(o[49]), .Z(n10664) );
  IV U11665 ( .A(n10664), .Z(n10647) );
  XNOR U11666 ( .A(n10663), .B(n10647), .Z(n10956) );
  AND U11667 ( .A(\stack[1][7] ), .B(o[50]), .Z(n10953) );
  NAND U11668 ( .A(n10649), .B(n10648), .Z(n10653) );
  NAND U11669 ( .A(n10651), .B(n10650), .Z(n10652) );
  NAND U11670 ( .A(n10653), .B(n10652), .Z(n10954) );
  IV U11671 ( .A(n10954), .Z(n10654) );
  XNOR U11672 ( .A(n10953), .B(n10654), .Z(n10955) );
  XOR U11673 ( .A(n10956), .B(n10955), .Z(n10655) );
  NAND U11674 ( .A(n10656), .B(n10655), .Z(n10658) );
  AND U11675 ( .A(\stack[1][6] ), .B(o[51]), .Z(n12525) );
  XOR U11676 ( .A(n10656), .B(n10655), .Z(n12524) );
  NAND U11677 ( .A(n12525), .B(n12524), .Z(n10657) );
  NAND U11678 ( .A(n10658), .B(n10657), .Z(n10659) );
  AND U11679 ( .A(\stack[1][6] ), .B(o[52]), .Z(n10660) );
  NAND U11680 ( .A(n10659), .B(n10660), .Z(n10960) );
  NAND U11681 ( .A(n10662), .B(n10661), .Z(n10666) );
  NAND U11682 ( .A(n10664), .B(n10663), .Z(n10665) );
  NAND U11683 ( .A(n10666), .B(n10665), .Z(n10962) );
  AND U11684 ( .A(\stack[1][8] ), .B(o[50]), .Z(n10961) );
  NAND U11685 ( .A(n10668), .B(n10667), .Z(n10672) );
  NAND U11686 ( .A(n10670), .B(n10669), .Z(n10671) );
  NAND U11687 ( .A(n10672), .B(n10671), .Z(n11248) );
  NAND U11688 ( .A(n10674), .B(n10673), .Z(n10678) );
  NAND U11689 ( .A(n10676), .B(n10675), .Z(n10677) );
  AND U11690 ( .A(n10678), .B(n10677), .Z(n10974) );
  NAND U11691 ( .A(\stack[1][12] ), .B(o[46]), .Z(n10973) );
  XOR U11692 ( .A(n10974), .B(n10973), .Z(n10976) );
  NAND U11693 ( .A(n10680), .B(n10679), .Z(n10684) );
  NAND U11694 ( .A(n10682), .B(n10681), .Z(n10683) );
  NAND U11695 ( .A(n10684), .B(n10683), .Z(n10979) );
  AND U11696 ( .A(\stack[1][14] ), .B(o[44]), .Z(n10980) );
  XOR U11697 ( .A(n10979), .B(n10980), .Z(n10982) );
  NAND U11698 ( .A(n10686), .B(n10685), .Z(n10690) );
  NAND U11699 ( .A(n10688), .B(n10687), .Z(n10689) );
  NAND U11700 ( .A(n10690), .B(n10689), .Z(n10985) );
  AND U11701 ( .A(\stack[1][16] ), .B(o[42]), .Z(n10986) );
  XOR U11702 ( .A(n10985), .B(n10986), .Z(n10988) );
  NAND U11703 ( .A(n10692), .B(n10691), .Z(n10696) );
  NAND U11704 ( .A(n10694), .B(n10693), .Z(n10695) );
  NAND U11705 ( .A(n10696), .B(n10695), .Z(n10991) );
  AND U11706 ( .A(\stack[1][18] ), .B(o[40]), .Z(n10992) );
  XOR U11707 ( .A(n10991), .B(n10992), .Z(n10994) );
  NAND U11708 ( .A(n10698), .B(n10697), .Z(n10702) );
  NAND U11709 ( .A(n10700), .B(n10699), .Z(n10701) );
  NAND U11710 ( .A(n10702), .B(n10701), .Z(n11224) );
  NAND U11711 ( .A(n10704), .B(n10703), .Z(n10708) );
  NAND U11712 ( .A(n10706), .B(n10705), .Z(n10707) );
  AND U11713 ( .A(n10708), .B(n10707), .Z(n10998) );
  NAND U11714 ( .A(\stack[1][20] ), .B(o[38]), .Z(n10997) );
  XOR U11715 ( .A(n10998), .B(n10997), .Z(n11000) );
  NAND U11716 ( .A(n10710), .B(n10709), .Z(n10714) );
  NAND U11717 ( .A(n10712), .B(n10711), .Z(n10713) );
  NAND U11718 ( .A(n10714), .B(n10713), .Z(n11015) );
  AND U11719 ( .A(\stack[1][26] ), .B(o[32]), .Z(n11016) );
  XOR U11720 ( .A(n11015), .B(n11016), .Z(n11018) );
  NAND U11721 ( .A(n10716), .B(n10715), .Z(n10720) );
  NAND U11722 ( .A(n10718), .B(n10717), .Z(n10719) );
  NAND U11723 ( .A(n10720), .B(n10719), .Z(n11021) );
  AND U11724 ( .A(\stack[1][28] ), .B(o[30]), .Z(n11022) );
  XOR U11725 ( .A(n11021), .B(n11022), .Z(n11024) );
  AND U11726 ( .A(\stack[1][29] ), .B(o[29]), .Z(n11030) );
  NAND U11727 ( .A(n10722), .B(n10721), .Z(n10726) );
  NAND U11728 ( .A(n10724), .B(n10723), .Z(n10725) );
  NAND U11729 ( .A(n10726), .B(n10725), .Z(n11033) );
  AND U11730 ( .A(o[28]), .B(\stack[1][30] ), .Z(n11034) );
  XOR U11731 ( .A(n11033), .B(n11034), .Z(n11036) );
  NAND U11732 ( .A(n10728), .B(n10727), .Z(n10732) );
  NAND U11733 ( .A(n10730), .B(n10729), .Z(n10731) );
  NAND U11734 ( .A(n10732), .B(n10731), .Z(n11039) );
  AND U11735 ( .A(o[26]), .B(\stack[1][32] ), .Z(n11040) );
  XOR U11736 ( .A(n11039), .B(n11040), .Z(n11042) );
  NAND U11737 ( .A(n10734), .B(n10733), .Z(n10738) );
  NANDN U11738 ( .A(n10736), .B(n10735), .Z(n10737) );
  NAND U11739 ( .A(n10738), .B(n10737), .Z(n11045) );
  AND U11740 ( .A(o[24]), .B(\stack[1][34] ), .Z(n11046) );
  XOR U11741 ( .A(n11045), .B(n11046), .Z(n11048) );
  AND U11742 ( .A(o[22]), .B(\stack[1][36] ), .Z(n11060) );
  NAND U11743 ( .A(o[20]), .B(\stack[1][38] ), .Z(n11065) );
  NAND U11744 ( .A(n10740), .B(n10739), .Z(n10744) );
  NAND U11745 ( .A(n10742), .B(n10741), .Z(n10743) );
  NAND U11746 ( .A(n10744), .B(n10743), .Z(n11063) );
  AND U11747 ( .A(o[18]), .B(\stack[1][40] ), .Z(n11178) );
  NAND U11748 ( .A(n10746), .B(n10745), .Z(n10750) );
  NAND U11749 ( .A(n10748), .B(n10747), .Z(n10749) );
  AND U11750 ( .A(n10750), .B(n10749), .Z(n11176) );
  NAND U11751 ( .A(o[17]), .B(\stack[1][41] ), .Z(n11077) );
  NAND U11752 ( .A(n10752), .B(n10751), .Z(n10756) );
  NAND U11753 ( .A(n10754), .B(n10753), .Z(n10755) );
  NAND U11754 ( .A(n10756), .B(n10755), .Z(n11165) );
  AND U11755 ( .A(o[13]), .B(\stack[1][45] ), .Z(n11159) );
  NAND U11756 ( .A(n10758), .B(n10757), .Z(n10762) );
  NAND U11757 ( .A(n10760), .B(n10759), .Z(n10761) );
  NAND U11758 ( .A(n10762), .B(n10761), .Z(n11151) );
  NAND U11759 ( .A(o[11]), .B(\stack[1][47] ), .Z(n11089) );
  NAND U11760 ( .A(n10764), .B(n10763), .Z(n10768) );
  NAND U11761 ( .A(n10766), .B(n10765), .Z(n10767) );
  AND U11762 ( .A(n10768), .B(n10767), .Z(n11087) );
  AND U11763 ( .A(o[10]), .B(\stack[1][48] ), .Z(n11096) );
  NAND U11764 ( .A(n10770), .B(n10769), .Z(n10774) );
  NAND U11765 ( .A(n10772), .B(n10771), .Z(n10773) );
  AND U11766 ( .A(n10774), .B(n10773), .Z(n11094) );
  NAND U11767 ( .A(o[9]), .B(\stack[1][49] ), .Z(n11101) );
  NAND U11768 ( .A(n10776), .B(n10775), .Z(n10780) );
  NAND U11769 ( .A(n10778), .B(n10777), .Z(n10779) );
  NAND U11770 ( .A(n10780), .B(n10779), .Z(n11141) );
  AND U11771 ( .A(o[6]), .B(\stack[1][52] ), .Z(n11108) );
  NAND U11772 ( .A(o[4]), .B(\stack[1][54] ), .Z(n11113) );
  NANDN U11773 ( .A(n10781), .B(n11117), .Z(n10785) );
  NANDN U11774 ( .A(n10783), .B(n10782), .Z(n10784) );
  NAND U11775 ( .A(n10785), .B(n10784), .Z(n11127) );
  AND U11776 ( .A(o[2]), .B(\stack[1][56] ), .Z(n11118) );
  AND U11777 ( .A(n10786), .B(n10788), .Z(n10787) );
  AND U11778 ( .A(o[1]), .B(\stack[1][58] ), .Z(n11124) );
  NAND U11779 ( .A(n11122), .B(n11124), .Z(n11403) );
  XOR U11780 ( .A(n10787), .B(n11403), .Z(n10790) );
  AND U11781 ( .A(o[0]), .B(\stack[1][58] ), .Z(n11408) );
  OR U11782 ( .A(n10788), .B(n11408), .Z(n10789) );
  NAND U11783 ( .A(n10790), .B(n10789), .Z(n11119) );
  XNOR U11784 ( .A(n11118), .B(n11119), .Z(n11128) );
  XOR U11785 ( .A(n11127), .B(n11128), .Z(n11130) );
  AND U11786 ( .A(o[3]), .B(\stack[1][55] ), .Z(n11129) );
  XNOR U11787 ( .A(n11130), .B(n11129), .Z(n11112) );
  NAND U11788 ( .A(n10792), .B(n10791), .Z(n10796) );
  NAND U11789 ( .A(n10794), .B(n10793), .Z(n10795) );
  AND U11790 ( .A(n10796), .B(n10795), .Z(n11111) );
  XNOR U11791 ( .A(n11113), .B(n11114), .Z(n11134) );
  NAND U11792 ( .A(n10798), .B(n10797), .Z(n10802) );
  NAND U11793 ( .A(n10800), .B(n10799), .Z(n10801) );
  NAND U11794 ( .A(n10802), .B(n10801), .Z(n11133) );
  AND U11795 ( .A(o[5]), .B(\stack[1][53] ), .Z(n11135) );
  XOR U11796 ( .A(n11136), .B(n11135), .Z(n11106) );
  NAND U11797 ( .A(n10804), .B(n10803), .Z(n10808) );
  NAND U11798 ( .A(n10806), .B(n10805), .Z(n10807) );
  NAND U11799 ( .A(n10808), .B(n10807), .Z(n11105) );
  XOR U11800 ( .A(n11106), .B(n11105), .Z(n11107) );
  XOR U11801 ( .A(n11108), .B(n11107), .Z(n11140) );
  AND U11802 ( .A(o[7]), .B(\stack[1][51] ), .Z(n11139) );
  XOR U11803 ( .A(n11140), .B(n11139), .Z(n11142) );
  XOR U11804 ( .A(n11141), .B(n11142), .Z(n11146) );
  AND U11805 ( .A(o[8]), .B(\stack[1][50] ), .Z(n11145) );
  XOR U11806 ( .A(n11146), .B(n11145), .Z(n11148) );
  NAND U11807 ( .A(n10810), .B(n10809), .Z(n10814) );
  NAND U11808 ( .A(n10812), .B(n10811), .Z(n10813) );
  NAND U11809 ( .A(n10814), .B(n10813), .Z(n11147) );
  XNOR U11810 ( .A(n11148), .B(n11147), .Z(n11100) );
  NAND U11811 ( .A(n10816), .B(n10815), .Z(n10820) );
  NAND U11812 ( .A(n10818), .B(n10817), .Z(n10819) );
  AND U11813 ( .A(n10820), .B(n10819), .Z(n11099) );
  XOR U11814 ( .A(n11101), .B(n11102), .Z(n11093) );
  XOR U11815 ( .A(n11094), .B(n11093), .Z(n11095) );
  XNOR U11816 ( .A(n11096), .B(n11095), .Z(n11088) );
  XOR U11817 ( .A(n11089), .B(n11090), .Z(n11152) );
  XOR U11818 ( .A(n11151), .B(n11152), .Z(n11154) );
  NAND U11819 ( .A(o[12]), .B(\stack[1][46] ), .Z(n11153) );
  XNOR U11820 ( .A(n11154), .B(n11153), .Z(n11158) );
  NAND U11821 ( .A(n10822), .B(n10821), .Z(n10826) );
  NAND U11822 ( .A(n10824), .B(n10823), .Z(n10825) );
  NAND U11823 ( .A(n10826), .B(n10825), .Z(n11157) );
  XNOR U11824 ( .A(n11159), .B(n11160), .Z(n11082) );
  AND U11825 ( .A(o[14]), .B(\stack[1][44] ), .Z(n11081) );
  XOR U11826 ( .A(n11082), .B(n11081), .Z(n11084) );
  NAND U11827 ( .A(n10828), .B(n10827), .Z(n10832) );
  NAND U11828 ( .A(n10830), .B(n10829), .Z(n10831) );
  NAND U11829 ( .A(n10832), .B(n10831), .Z(n11083) );
  XOR U11830 ( .A(n11084), .B(n11083), .Z(n11164) );
  AND U11831 ( .A(o[15]), .B(\stack[1][43] ), .Z(n11163) );
  XOR U11832 ( .A(n11164), .B(n11163), .Z(n11166) );
  XOR U11833 ( .A(n11165), .B(n11166), .Z(n11170) );
  AND U11834 ( .A(o[16]), .B(\stack[1][42] ), .Z(n11169) );
  XOR U11835 ( .A(n11170), .B(n11169), .Z(n11172) );
  NAND U11836 ( .A(n10834), .B(n10833), .Z(n10838) );
  NAND U11837 ( .A(n10836), .B(n10835), .Z(n10837) );
  NAND U11838 ( .A(n10838), .B(n10837), .Z(n11171) );
  XNOR U11839 ( .A(n11172), .B(n11171), .Z(n11076) );
  NAND U11840 ( .A(n10840), .B(n10839), .Z(n10844) );
  NAND U11841 ( .A(n10842), .B(n10841), .Z(n10843) );
  AND U11842 ( .A(n10844), .B(n10843), .Z(n11075) );
  XOR U11843 ( .A(n11077), .B(n11078), .Z(n11175) );
  XOR U11844 ( .A(n11176), .B(n11175), .Z(n11177) );
  XNOR U11845 ( .A(n11178), .B(n11177), .Z(n11070) );
  NAND U11846 ( .A(n10846), .B(n10845), .Z(n10850) );
  NAND U11847 ( .A(n10848), .B(n10847), .Z(n10849) );
  AND U11848 ( .A(n10850), .B(n10849), .Z(n11069) );
  NAND U11849 ( .A(o[19]), .B(\stack[1][39] ), .Z(n11071) );
  XOR U11850 ( .A(n11072), .B(n11071), .Z(n11064) );
  XOR U11851 ( .A(n11063), .B(n11064), .Z(n11066) );
  XNOR U11852 ( .A(n11065), .B(n11066), .Z(n11184) );
  AND U11853 ( .A(o[21]), .B(\stack[1][37] ), .Z(n11182) );
  NAND U11854 ( .A(n10852), .B(n10851), .Z(n10856) );
  NAND U11855 ( .A(n10854), .B(n10853), .Z(n10855) );
  NAND U11856 ( .A(n10856), .B(n10855), .Z(n11181) );
  XOR U11857 ( .A(n11182), .B(n11181), .Z(n11183) );
  NAND U11858 ( .A(n10858), .B(n10857), .Z(n10862) );
  NAND U11859 ( .A(n10860), .B(n10859), .Z(n10861) );
  NAND U11860 ( .A(n10862), .B(n10861), .Z(n11057) );
  XOR U11861 ( .A(n11058), .B(n11057), .Z(n11059) );
  XOR U11862 ( .A(n11060), .B(n11059), .Z(n11054) );
  AND U11863 ( .A(o[23]), .B(\stack[1][35] ), .Z(n11052) );
  NAND U11864 ( .A(n10864), .B(n10863), .Z(n10868) );
  NAND U11865 ( .A(n10866), .B(n10865), .Z(n10867) );
  NAND U11866 ( .A(n10868), .B(n10867), .Z(n11051) );
  XOR U11867 ( .A(n11052), .B(n11051), .Z(n11053) );
  XOR U11868 ( .A(n11054), .B(n11053), .Z(n11047) );
  XOR U11869 ( .A(n11048), .B(n11047), .Z(n11188) );
  NAND U11870 ( .A(n10870), .B(n10869), .Z(n10874) );
  NAND U11871 ( .A(n10872), .B(n10871), .Z(n10873) );
  NAND U11872 ( .A(n10874), .B(n10873), .Z(n11187) );
  XOR U11873 ( .A(n11188), .B(n11187), .Z(n11190) );
  AND U11874 ( .A(o[25]), .B(\stack[1][33] ), .Z(n11189) );
  XOR U11875 ( .A(n11190), .B(n11189), .Z(n11041) );
  XOR U11876 ( .A(n11042), .B(n11041), .Z(n11194) );
  NAND U11877 ( .A(n10876), .B(n10875), .Z(n10880) );
  NAND U11878 ( .A(n10878), .B(n10877), .Z(n10879) );
  NAND U11879 ( .A(n10880), .B(n10879), .Z(n11193) );
  XOR U11880 ( .A(n11194), .B(n11193), .Z(n11196) );
  AND U11881 ( .A(o[27]), .B(\stack[1][31] ), .Z(n11195) );
  XOR U11882 ( .A(n11196), .B(n11195), .Z(n11035) );
  XOR U11883 ( .A(n11036), .B(n11035), .Z(n11028) );
  NAND U11884 ( .A(n10882), .B(n10881), .Z(n10886) );
  NAND U11885 ( .A(n10884), .B(n10883), .Z(n10885) );
  NAND U11886 ( .A(n10886), .B(n10885), .Z(n11027) );
  XOR U11887 ( .A(n11028), .B(n11027), .Z(n11029) );
  XOR U11888 ( .A(n11030), .B(n11029), .Z(n11023) );
  XOR U11889 ( .A(n11024), .B(n11023), .Z(n11200) );
  NAND U11890 ( .A(n10888), .B(n10887), .Z(n10892) );
  NAND U11891 ( .A(n10890), .B(n10889), .Z(n10891) );
  NAND U11892 ( .A(n10892), .B(n10891), .Z(n11199) );
  XOR U11893 ( .A(n11200), .B(n11199), .Z(n11202) );
  AND U11894 ( .A(\stack[1][27] ), .B(o[31]), .Z(n11201) );
  XOR U11895 ( .A(n11202), .B(n11201), .Z(n11017) );
  XOR U11896 ( .A(n11018), .B(n11017), .Z(n11206) );
  NAND U11897 ( .A(n10894), .B(n10893), .Z(n10898) );
  NAND U11898 ( .A(n10896), .B(n10895), .Z(n10897) );
  NAND U11899 ( .A(n10898), .B(n10897), .Z(n11205) );
  XOR U11900 ( .A(n11206), .B(n11205), .Z(n11208) );
  AND U11901 ( .A(\stack[1][25] ), .B(o[33]), .Z(n11207) );
  XOR U11902 ( .A(n11208), .B(n11207), .Z(n11011) );
  NAND U11903 ( .A(n10900), .B(n10899), .Z(n10904) );
  NAND U11904 ( .A(n10902), .B(n10901), .Z(n10903) );
  NAND U11905 ( .A(n10904), .B(n10903), .Z(n11009) );
  AND U11906 ( .A(\stack[1][24] ), .B(o[34]), .Z(n11010) );
  XOR U11907 ( .A(n11009), .B(n11010), .Z(n11012) );
  NAND U11908 ( .A(n10906), .B(n10905), .Z(n10910) );
  NAND U11909 ( .A(n10908), .B(n10907), .Z(n10909) );
  NAND U11910 ( .A(n10910), .B(n10909), .Z(n11211) );
  XOR U11911 ( .A(n11212), .B(n11211), .Z(n11214) );
  AND U11912 ( .A(\stack[1][23] ), .B(o[35]), .Z(n11213) );
  XOR U11913 ( .A(n11214), .B(n11213), .Z(n11005) );
  NAND U11914 ( .A(n10912), .B(n10911), .Z(n10916) );
  NAND U11915 ( .A(n10914), .B(n10913), .Z(n10915) );
  NAND U11916 ( .A(n10916), .B(n10915), .Z(n11003) );
  AND U11917 ( .A(\stack[1][22] ), .B(o[36]), .Z(n11004) );
  XOR U11918 ( .A(n11003), .B(n11004), .Z(n11006) );
  NAND U11919 ( .A(n10918), .B(n10917), .Z(n10922) );
  NAND U11920 ( .A(n10920), .B(n10919), .Z(n10921) );
  NAND U11921 ( .A(n10922), .B(n10921), .Z(n11217) );
  XOR U11922 ( .A(n11218), .B(n11217), .Z(n11220) );
  AND U11923 ( .A(\stack[1][21] ), .B(o[37]), .Z(n11219) );
  XNOR U11924 ( .A(n11220), .B(n11219), .Z(n10999) );
  XNOR U11925 ( .A(n11000), .B(n10999), .Z(n11223) );
  XOR U11926 ( .A(n11224), .B(n11223), .Z(n11226) );
  AND U11927 ( .A(\stack[1][19] ), .B(o[39]), .Z(n11225) );
  XOR U11928 ( .A(n11226), .B(n11225), .Z(n10993) );
  XOR U11929 ( .A(n10994), .B(n10993), .Z(n11230) );
  NAND U11930 ( .A(n10924), .B(n10923), .Z(n10928) );
  NAND U11931 ( .A(n10926), .B(n10925), .Z(n10927) );
  NAND U11932 ( .A(n10928), .B(n10927), .Z(n11229) );
  XOR U11933 ( .A(n11230), .B(n11229), .Z(n11232) );
  AND U11934 ( .A(\stack[1][17] ), .B(o[41]), .Z(n11231) );
  XOR U11935 ( .A(n11232), .B(n11231), .Z(n10987) );
  XOR U11936 ( .A(n10988), .B(n10987), .Z(n11236) );
  NAND U11937 ( .A(n10930), .B(n10929), .Z(n10934) );
  NAND U11938 ( .A(n10932), .B(n10931), .Z(n10933) );
  NAND U11939 ( .A(n10934), .B(n10933), .Z(n11235) );
  XOR U11940 ( .A(n11236), .B(n11235), .Z(n11238) );
  AND U11941 ( .A(\stack[1][15] ), .B(o[43]), .Z(n11237) );
  XOR U11942 ( .A(n11238), .B(n11237), .Z(n10981) );
  XOR U11943 ( .A(n10982), .B(n10981), .Z(n11242) );
  NAND U11944 ( .A(n10936), .B(n10935), .Z(n10940) );
  NAND U11945 ( .A(n10938), .B(n10937), .Z(n10939) );
  NAND U11946 ( .A(n10940), .B(n10939), .Z(n11241) );
  XOR U11947 ( .A(n11242), .B(n11241), .Z(n11244) );
  AND U11948 ( .A(\stack[1][13] ), .B(o[45]), .Z(n11243) );
  XNOR U11949 ( .A(n11244), .B(n11243), .Z(n10975) );
  XNOR U11950 ( .A(n10976), .B(n10975), .Z(n11247) );
  XOR U11951 ( .A(n11248), .B(n11247), .Z(n11250) );
  AND U11952 ( .A(\stack[1][11] ), .B(o[47]), .Z(n11249) );
  XNOR U11953 ( .A(n11250), .B(n11249), .Z(n10970) );
  NAND U11954 ( .A(n10942), .B(n10941), .Z(n10946) );
  NAND U11955 ( .A(n10944), .B(n10943), .Z(n10945) );
  AND U11956 ( .A(n10946), .B(n10945), .Z(n10967) );
  NAND U11957 ( .A(\stack[1][10] ), .B(o[48]), .Z(n10968) );
  NAND U11958 ( .A(n10948), .B(n10947), .Z(n10952) );
  NAND U11959 ( .A(n10950), .B(n10949), .Z(n10951) );
  NAND U11960 ( .A(n10952), .B(n10951), .Z(n11253) );
  XOR U11961 ( .A(n11254), .B(n11253), .Z(n11255) );
  AND U11962 ( .A(\stack[1][9] ), .B(o[49]), .Z(n11256) );
  XOR U11963 ( .A(n10964), .B(n10963), .Z(n11259) );
  NAND U11964 ( .A(n10954), .B(n10953), .Z(n10958) );
  NAND U11965 ( .A(n10956), .B(n10955), .Z(n10957) );
  NAND U11966 ( .A(n10958), .B(n10957), .Z(n11260) );
  AND U11967 ( .A(\stack[1][7] ), .B(o[51]), .Z(n11262) );
  NAND U11968 ( .A(n12532), .B(n12531), .Z(n10959) );
  NAND U11969 ( .A(n10960), .B(n10959), .Z(n11265) );
  AND U11970 ( .A(\stack[1][8] ), .B(o[51]), .Z(n11572) );
  NAND U11971 ( .A(n10962), .B(n10961), .Z(n10966) );
  NAND U11972 ( .A(n10964), .B(n10963), .Z(n10965) );
  NAND U11973 ( .A(n10966), .B(n10965), .Z(n11570) );
  NAND U11974 ( .A(n10968), .B(n10967), .Z(n10972) );
  NAND U11975 ( .A(n10970), .B(n10969), .Z(n10971) );
  AND U11976 ( .A(n10972), .B(n10971), .Z(n11558) );
  NAND U11977 ( .A(n10974), .B(n10973), .Z(n10978) );
  NAND U11978 ( .A(n10976), .B(n10975), .Z(n10977) );
  AND U11979 ( .A(n10978), .B(n10977), .Z(n11272) );
  NAND U11980 ( .A(n10980), .B(n10979), .Z(n10984) );
  NAND U11981 ( .A(n10982), .B(n10981), .Z(n10983) );
  NAND U11982 ( .A(n10984), .B(n10983), .Z(n11539) );
  AND U11983 ( .A(\stack[1][16] ), .B(o[43]), .Z(n11285) );
  NAND U11984 ( .A(n10986), .B(n10985), .Z(n10990) );
  NAND U11985 ( .A(n10988), .B(n10987), .Z(n10989) );
  NAND U11986 ( .A(n10990), .B(n10989), .Z(n11283) );
  NAND U11987 ( .A(n10992), .B(n10991), .Z(n10996) );
  NAND U11988 ( .A(n10994), .B(n10993), .Z(n10995) );
  NAND U11989 ( .A(n10996), .B(n10995), .Z(n11295) );
  AND U11990 ( .A(\stack[1][20] ), .B(o[39]), .Z(n11304) );
  NAND U11991 ( .A(n10998), .B(n10997), .Z(n11002) );
  NAND U11992 ( .A(n11000), .B(n10999), .Z(n11001) );
  AND U11993 ( .A(n11002), .B(n11001), .Z(n11302) );
  AND U11994 ( .A(\stack[1][22] ), .B(o[37]), .Z(n11315) );
  NAND U11995 ( .A(n11004), .B(n11003), .Z(n11008) );
  NAND U11996 ( .A(n11006), .B(n11005), .Z(n11007) );
  NAND U11997 ( .A(n11008), .B(n11007), .Z(n11313) );
  AND U11998 ( .A(\stack[1][24] ), .B(o[35]), .Z(n11321) );
  NAND U11999 ( .A(n11010), .B(n11009), .Z(n11014) );
  NAND U12000 ( .A(n11012), .B(n11011), .Z(n11013) );
  NAND U12001 ( .A(n11014), .B(n11013), .Z(n11319) );
  NAND U12002 ( .A(n11016), .B(n11015), .Z(n11020) );
  NAND U12003 ( .A(n11018), .B(n11017), .Z(n11019) );
  NAND U12004 ( .A(n11020), .B(n11019), .Z(n11325) );
  AND U12005 ( .A(\stack[1][28] ), .B(o[31]), .Z(n11333) );
  NAND U12006 ( .A(n11022), .B(n11021), .Z(n11026) );
  NAND U12007 ( .A(n11024), .B(n11023), .Z(n11025) );
  NAND U12008 ( .A(n11026), .B(n11025), .Z(n11331) );
  AND U12009 ( .A(\stack[1][29] ), .B(o[30]), .Z(n11510) );
  NAND U12010 ( .A(n11028), .B(n11027), .Z(n11032) );
  NAND U12011 ( .A(n11030), .B(n11029), .Z(n11031) );
  NAND U12012 ( .A(n11032), .B(n11031), .Z(n11509) );
  XOR U12013 ( .A(n11510), .B(n11509), .Z(n11512) );
  AND U12014 ( .A(\stack[1][30] ), .B(o[29]), .Z(n11505) );
  NAND U12015 ( .A(n11034), .B(n11033), .Z(n11038) );
  NAND U12016 ( .A(n11036), .B(n11035), .Z(n11037) );
  NAND U12017 ( .A(n11038), .B(n11037), .Z(n11503) );
  NAND U12018 ( .A(n11040), .B(n11039), .Z(n11044) );
  NAND U12019 ( .A(n11042), .B(n11041), .Z(n11043) );
  NAND U12020 ( .A(n11044), .B(n11043), .Z(n11491) );
  NAND U12021 ( .A(n11046), .B(n11045), .Z(n11050) );
  NAND U12022 ( .A(n11048), .B(n11047), .Z(n11049) );
  NAND U12023 ( .A(n11050), .B(n11049), .Z(n11337) );
  NAND U12024 ( .A(n11052), .B(n11051), .Z(n11056) );
  NAND U12025 ( .A(n11054), .B(n11053), .Z(n11055) );
  NAND U12026 ( .A(n11056), .B(n11055), .Z(n11481) );
  NAND U12027 ( .A(n11058), .B(n11057), .Z(n11062) );
  NAND U12028 ( .A(n11060), .B(n11059), .Z(n11061) );
  NAND U12029 ( .A(n11062), .B(n11061), .Z(n11473) );
  NAND U12030 ( .A(o[21]), .B(\stack[1][38] ), .Z(n11345) );
  NAND U12031 ( .A(n11064), .B(n11063), .Z(n11068) );
  NAND U12032 ( .A(n11066), .B(n11065), .Z(n11067) );
  NAND U12033 ( .A(n11068), .B(n11067), .Z(n11344) );
  NAND U12034 ( .A(n11070), .B(n11069), .Z(n11074) );
  NAND U12035 ( .A(n11072), .B(n11071), .Z(n11073) );
  AND U12036 ( .A(n11074), .B(n11073), .Z(n11464) );
  AND U12037 ( .A(o[18]), .B(\stack[1][41] ), .Z(n11452) );
  NAND U12038 ( .A(n11076), .B(n11075), .Z(n11080) );
  NANDN U12039 ( .A(n11078), .B(n11077), .Z(n11079) );
  AND U12040 ( .A(n11080), .B(n11079), .Z(n11450) );
  NAND U12041 ( .A(o[17]), .B(\stack[1][42] ), .Z(n11351) );
  NAND U12042 ( .A(n11082), .B(n11081), .Z(n11086) );
  NAND U12043 ( .A(n11084), .B(n11083), .Z(n11085) );
  NAND U12044 ( .A(n11086), .B(n11085), .Z(n11439) );
  AND U12045 ( .A(o[13]), .B(\stack[1][46] ), .Z(n11364) );
  AND U12046 ( .A(o[12]), .B(\stack[1][47] ), .Z(n11370) );
  NAND U12047 ( .A(n11088), .B(n11087), .Z(n11092) );
  NAND U12048 ( .A(n11090), .B(n11089), .Z(n11091) );
  AND U12049 ( .A(n11092), .B(n11091), .Z(n11368) );
  NAND U12050 ( .A(o[11]), .B(\stack[1][48] ), .Z(n11375) );
  NAND U12051 ( .A(n11094), .B(n11093), .Z(n11098) );
  NAND U12052 ( .A(n11096), .B(n11095), .Z(n11097) );
  AND U12053 ( .A(n11098), .B(n11097), .Z(n11374) );
  AND U12054 ( .A(o[10]), .B(\stack[1][49] ), .Z(n11382) );
  NAND U12055 ( .A(n11100), .B(n11099), .Z(n11104) );
  NANDN U12056 ( .A(n11102), .B(n11101), .Z(n11103) );
  AND U12057 ( .A(n11104), .B(n11103), .Z(n11379) );
  NAND U12058 ( .A(o[9]), .B(\stack[1][50] ), .Z(n11387) );
  NAND U12059 ( .A(n11106), .B(n11105), .Z(n11110) );
  NAND U12060 ( .A(n11108), .B(n11107), .Z(n11109) );
  NAND U12061 ( .A(n11110), .B(n11109), .Z(n11427) );
  AND U12062 ( .A(o[6]), .B(\stack[1][53] ), .Z(n11394) );
  NAND U12063 ( .A(n11112), .B(n11111), .Z(n11116) );
  NAND U12064 ( .A(n11114), .B(n11113), .Z(n11115) );
  AND U12065 ( .A(n11116), .B(n11115), .Z(n11420) );
  AND U12066 ( .A(o[4]), .B(\stack[1][55] ), .Z(n11400) );
  NANDN U12067 ( .A(n11117), .B(n11403), .Z(n11121) );
  NANDN U12068 ( .A(n11119), .B(n11118), .Z(n11120) );
  NAND U12069 ( .A(n11121), .B(n11120), .Z(n11413) );
  AND U12070 ( .A(o[2]), .B(\stack[1][57] ), .Z(n11404) );
  AND U12071 ( .A(n11122), .B(n11124), .Z(n11123) );
  AND U12072 ( .A(o[1]), .B(\stack[1][59] ), .Z(n11410) );
  NAND U12073 ( .A(n11408), .B(n11410), .Z(n11762) );
  XOR U12074 ( .A(n11123), .B(n11762), .Z(n11126) );
  AND U12075 ( .A(o[0]), .B(\stack[1][59] ), .Z(n11767) );
  OR U12076 ( .A(n11124), .B(n11767), .Z(n11125) );
  NAND U12077 ( .A(n11126), .B(n11125), .Z(n11405) );
  XNOR U12078 ( .A(n11404), .B(n11405), .Z(n11414) );
  XOR U12079 ( .A(n11413), .B(n11414), .Z(n11416) );
  AND U12080 ( .A(o[3]), .B(\stack[1][56] ), .Z(n11415) );
  XOR U12081 ( .A(n11416), .B(n11415), .Z(n11398) );
  NAND U12082 ( .A(n11128), .B(n11127), .Z(n11132) );
  NAND U12083 ( .A(n11130), .B(n11129), .Z(n11131) );
  NAND U12084 ( .A(n11132), .B(n11131), .Z(n11397) );
  XOR U12085 ( .A(n11398), .B(n11397), .Z(n11399) );
  XOR U12086 ( .A(n11400), .B(n11399), .Z(n11419) );
  XOR U12087 ( .A(n11420), .B(n11419), .Z(n11422) );
  AND U12088 ( .A(o[5]), .B(\stack[1][54] ), .Z(n11421) );
  XOR U12089 ( .A(n11422), .B(n11421), .Z(n11392) );
  NAND U12090 ( .A(n11134), .B(n11133), .Z(n11138) );
  NAND U12091 ( .A(n11136), .B(n11135), .Z(n11137) );
  NAND U12092 ( .A(n11138), .B(n11137), .Z(n11391) );
  XOR U12093 ( .A(n11392), .B(n11391), .Z(n11393) );
  XOR U12094 ( .A(n11394), .B(n11393), .Z(n11426) );
  AND U12095 ( .A(o[7]), .B(\stack[1][52] ), .Z(n11425) );
  XOR U12096 ( .A(n11426), .B(n11425), .Z(n11428) );
  XOR U12097 ( .A(n11427), .B(n11428), .Z(n11432) );
  AND U12098 ( .A(o[8]), .B(\stack[1][51] ), .Z(n11431) );
  XOR U12099 ( .A(n11432), .B(n11431), .Z(n11434) );
  NAND U12100 ( .A(n11140), .B(n11139), .Z(n11144) );
  NAND U12101 ( .A(n11142), .B(n11141), .Z(n11143) );
  NAND U12102 ( .A(n11144), .B(n11143), .Z(n11433) );
  XNOR U12103 ( .A(n11434), .B(n11433), .Z(n11386) );
  NAND U12104 ( .A(n11146), .B(n11145), .Z(n11150) );
  NAND U12105 ( .A(n11148), .B(n11147), .Z(n11149) );
  AND U12106 ( .A(n11150), .B(n11149), .Z(n11385) );
  XNOR U12107 ( .A(n11387), .B(n11388), .Z(n11380) );
  XNOR U12108 ( .A(n11382), .B(n11381), .Z(n11373) );
  XOR U12109 ( .A(n11374), .B(n11373), .Z(n11376) );
  XNOR U12110 ( .A(n11375), .B(n11376), .Z(n11367) );
  XOR U12111 ( .A(n11368), .B(n11367), .Z(n11369) );
  XOR U12112 ( .A(n11370), .B(n11369), .Z(n11362) );
  NAND U12113 ( .A(n11152), .B(n11151), .Z(n11156) );
  NAND U12114 ( .A(n11154), .B(n11153), .Z(n11155) );
  AND U12115 ( .A(n11156), .B(n11155), .Z(n11361) );
  XOR U12116 ( .A(n11362), .B(n11361), .Z(n11363) );
  XOR U12117 ( .A(n11364), .B(n11363), .Z(n11356) );
  AND U12118 ( .A(o[14]), .B(\stack[1][45] ), .Z(n11355) );
  XOR U12119 ( .A(n11356), .B(n11355), .Z(n11358) );
  NAND U12120 ( .A(n11158), .B(n11157), .Z(n11162) );
  NANDN U12121 ( .A(n11160), .B(n11159), .Z(n11161) );
  NAND U12122 ( .A(n11162), .B(n11161), .Z(n11357) );
  XOR U12123 ( .A(n11358), .B(n11357), .Z(n11438) );
  AND U12124 ( .A(o[15]), .B(\stack[1][44] ), .Z(n11437) );
  XOR U12125 ( .A(n11438), .B(n11437), .Z(n11440) );
  XOR U12126 ( .A(n11439), .B(n11440), .Z(n11444) );
  AND U12127 ( .A(o[16]), .B(\stack[1][43] ), .Z(n11443) );
  XOR U12128 ( .A(n11444), .B(n11443), .Z(n11446) );
  NAND U12129 ( .A(n11164), .B(n11163), .Z(n11168) );
  NAND U12130 ( .A(n11166), .B(n11165), .Z(n11167) );
  NAND U12131 ( .A(n11168), .B(n11167), .Z(n11445) );
  XNOR U12132 ( .A(n11446), .B(n11445), .Z(n11350) );
  NAND U12133 ( .A(n11170), .B(n11169), .Z(n11174) );
  NAND U12134 ( .A(n11172), .B(n11171), .Z(n11173) );
  AND U12135 ( .A(n11174), .B(n11173), .Z(n11349) );
  XOR U12136 ( .A(n11351), .B(n11352), .Z(n11449) );
  XOR U12137 ( .A(n11450), .B(n11449), .Z(n11451) );
  XOR U12138 ( .A(n11452), .B(n11451), .Z(n11456) );
  AND U12139 ( .A(o[19]), .B(\stack[1][40] ), .Z(n11455) );
  XOR U12140 ( .A(n11456), .B(n11455), .Z(n11458) );
  NAND U12141 ( .A(n11176), .B(n11175), .Z(n11180) );
  NAND U12142 ( .A(n11178), .B(n11177), .Z(n11179) );
  NAND U12143 ( .A(n11180), .B(n11179), .Z(n11457) );
  XOR U12144 ( .A(n11458), .B(n11457), .Z(n11462) );
  AND U12145 ( .A(o[20]), .B(\stack[1][39] ), .Z(n11461) );
  XOR U12146 ( .A(n11462), .B(n11461), .Z(n11463) );
  XNOR U12147 ( .A(n11464), .B(n11463), .Z(n11343) );
  XOR U12148 ( .A(n11344), .B(n11343), .Z(n11346) );
  XNOR U12149 ( .A(n11345), .B(n11346), .Z(n11470) );
  AND U12150 ( .A(o[22]), .B(\stack[1][37] ), .Z(n11468) );
  NAND U12151 ( .A(n11182), .B(n11181), .Z(n11186) );
  NAND U12152 ( .A(n11184), .B(n11183), .Z(n11185) );
  NAND U12153 ( .A(n11186), .B(n11185), .Z(n11467) );
  XOR U12154 ( .A(n11468), .B(n11467), .Z(n11469) );
  XOR U12155 ( .A(n11473), .B(n11474), .Z(n11476) );
  AND U12156 ( .A(o[23]), .B(\stack[1][36] ), .Z(n11475) );
  XOR U12157 ( .A(n11476), .B(n11475), .Z(n11480) );
  AND U12158 ( .A(o[24]), .B(\stack[1][35] ), .Z(n11479) );
  XOR U12159 ( .A(n11480), .B(n11479), .Z(n11482) );
  XOR U12160 ( .A(n11481), .B(n11482), .Z(n11338) );
  XOR U12161 ( .A(n11337), .B(n11338), .Z(n11340) );
  AND U12162 ( .A(o[25]), .B(\stack[1][34] ), .Z(n11339) );
  XOR U12163 ( .A(n11340), .B(n11339), .Z(n11488) );
  AND U12164 ( .A(o[26]), .B(\stack[1][33] ), .Z(n11486) );
  NAND U12165 ( .A(n11188), .B(n11187), .Z(n11192) );
  NAND U12166 ( .A(n11190), .B(n11189), .Z(n11191) );
  NAND U12167 ( .A(n11192), .B(n11191), .Z(n11485) );
  XOR U12168 ( .A(n11486), .B(n11485), .Z(n11487) );
  XOR U12169 ( .A(n11488), .B(n11487), .Z(n11492) );
  XOR U12170 ( .A(n11491), .B(n11492), .Z(n11494) );
  AND U12171 ( .A(o[27]), .B(\stack[1][32] ), .Z(n11493) );
  XOR U12172 ( .A(n11494), .B(n11493), .Z(n11500) );
  AND U12173 ( .A(o[28]), .B(\stack[1][31] ), .Z(n11498) );
  NAND U12174 ( .A(n11194), .B(n11193), .Z(n11198) );
  NAND U12175 ( .A(n11196), .B(n11195), .Z(n11197) );
  NAND U12176 ( .A(n11198), .B(n11197), .Z(n11497) );
  XOR U12177 ( .A(n11498), .B(n11497), .Z(n11499) );
  XOR U12178 ( .A(n11500), .B(n11499), .Z(n11504) );
  XOR U12179 ( .A(n11503), .B(n11504), .Z(n11506) );
  XOR U12180 ( .A(n11512), .B(n11511), .Z(n11332) );
  XOR U12181 ( .A(n11331), .B(n11332), .Z(n11334) );
  AND U12182 ( .A(\stack[1][27] ), .B(o[32]), .Z(n11516) );
  NAND U12183 ( .A(n11200), .B(n11199), .Z(n11204) );
  NAND U12184 ( .A(n11202), .B(n11201), .Z(n11203) );
  NAND U12185 ( .A(n11204), .B(n11203), .Z(n11515) );
  XOR U12186 ( .A(n11516), .B(n11515), .Z(n11517) );
  XOR U12187 ( .A(n11518), .B(n11517), .Z(n11326) );
  XOR U12188 ( .A(n11325), .B(n11326), .Z(n11328) );
  AND U12189 ( .A(\stack[1][26] ), .B(o[33]), .Z(n11327) );
  XOR U12190 ( .A(n11328), .B(n11327), .Z(n11524) );
  AND U12191 ( .A(\stack[1][25] ), .B(o[34]), .Z(n11522) );
  NAND U12192 ( .A(n11206), .B(n11205), .Z(n11210) );
  NAND U12193 ( .A(n11208), .B(n11207), .Z(n11209) );
  NAND U12194 ( .A(n11210), .B(n11209), .Z(n11521) );
  XOR U12195 ( .A(n11522), .B(n11521), .Z(n11523) );
  XOR U12196 ( .A(n11524), .B(n11523), .Z(n11320) );
  XOR U12197 ( .A(n11319), .B(n11320), .Z(n11322) );
  AND U12198 ( .A(\stack[1][23] ), .B(o[36]), .Z(n11528) );
  NAND U12199 ( .A(n11212), .B(n11211), .Z(n11216) );
  NAND U12200 ( .A(n11214), .B(n11213), .Z(n11215) );
  NAND U12201 ( .A(n11216), .B(n11215), .Z(n11527) );
  XOR U12202 ( .A(n11528), .B(n11527), .Z(n11529) );
  XOR U12203 ( .A(n11530), .B(n11529), .Z(n11314) );
  XOR U12204 ( .A(n11313), .B(n11314), .Z(n11316) );
  AND U12205 ( .A(\stack[1][21] ), .B(o[38]), .Z(n11308) );
  NAND U12206 ( .A(n11218), .B(n11217), .Z(n11222) );
  NAND U12207 ( .A(n11220), .B(n11219), .Z(n11221) );
  NAND U12208 ( .A(n11222), .B(n11221), .Z(n11307) );
  XOR U12209 ( .A(n11308), .B(n11307), .Z(n11309) );
  XOR U12210 ( .A(n11310), .B(n11309), .Z(n11301) );
  XOR U12211 ( .A(n11302), .B(n11301), .Z(n11303) );
  XOR U12212 ( .A(n11304), .B(n11303), .Z(n11536) );
  AND U12213 ( .A(\stack[1][19] ), .B(o[40]), .Z(n11534) );
  NAND U12214 ( .A(n11224), .B(n11223), .Z(n11228) );
  NAND U12215 ( .A(n11226), .B(n11225), .Z(n11227) );
  NAND U12216 ( .A(n11228), .B(n11227), .Z(n11533) );
  XOR U12217 ( .A(n11534), .B(n11533), .Z(n11535) );
  XOR U12218 ( .A(n11536), .B(n11535), .Z(n11296) );
  XOR U12219 ( .A(n11295), .B(n11296), .Z(n11298) );
  AND U12220 ( .A(\stack[1][18] ), .B(o[41]), .Z(n11297) );
  XOR U12221 ( .A(n11298), .B(n11297), .Z(n11292) );
  AND U12222 ( .A(\stack[1][17] ), .B(o[42]), .Z(n11290) );
  NAND U12223 ( .A(n11230), .B(n11229), .Z(n11234) );
  NAND U12224 ( .A(n11232), .B(n11231), .Z(n11233) );
  NAND U12225 ( .A(n11234), .B(n11233), .Z(n11289) );
  XOR U12226 ( .A(n11290), .B(n11289), .Z(n11291) );
  XOR U12227 ( .A(n11292), .B(n11291), .Z(n11284) );
  XOR U12228 ( .A(n11283), .B(n11284), .Z(n11286) );
  AND U12229 ( .A(\stack[1][15] ), .B(o[44]), .Z(n11278) );
  NAND U12230 ( .A(n11236), .B(n11235), .Z(n11240) );
  NAND U12231 ( .A(n11238), .B(n11237), .Z(n11239) );
  NAND U12232 ( .A(n11240), .B(n11239), .Z(n11277) );
  XOR U12233 ( .A(n11278), .B(n11277), .Z(n11279) );
  XOR U12234 ( .A(n11280), .B(n11279), .Z(n11540) );
  XOR U12235 ( .A(n11539), .B(n11540), .Z(n11542) );
  AND U12236 ( .A(\stack[1][14] ), .B(o[45]), .Z(n11541) );
  XOR U12237 ( .A(n11542), .B(n11541), .Z(n11548) );
  AND U12238 ( .A(\stack[1][13] ), .B(o[46]), .Z(n11546) );
  NAND U12239 ( .A(n11242), .B(n11241), .Z(n11246) );
  NAND U12240 ( .A(n11244), .B(n11243), .Z(n11245) );
  NAND U12241 ( .A(n11246), .B(n11245), .Z(n11545) );
  XOR U12242 ( .A(n11546), .B(n11545), .Z(n11547) );
  XOR U12243 ( .A(n11548), .B(n11547), .Z(n11271) );
  XOR U12244 ( .A(n11272), .B(n11271), .Z(n11274) );
  AND U12245 ( .A(\stack[1][12] ), .B(o[47]), .Z(n11273) );
  XOR U12246 ( .A(n11274), .B(n11273), .Z(n11554) );
  AND U12247 ( .A(\stack[1][11] ), .B(o[48]), .Z(n11552) );
  NAND U12248 ( .A(n11248), .B(n11247), .Z(n11252) );
  NAND U12249 ( .A(n11250), .B(n11249), .Z(n11251) );
  NAND U12250 ( .A(n11252), .B(n11251), .Z(n11551) );
  XOR U12251 ( .A(n11552), .B(n11551), .Z(n11553) );
  XOR U12252 ( .A(n11554), .B(n11553), .Z(n11557) );
  XOR U12253 ( .A(n11558), .B(n11557), .Z(n11560) );
  AND U12254 ( .A(\stack[1][10] ), .B(o[49]), .Z(n11559) );
  XOR U12255 ( .A(n11560), .B(n11559), .Z(n11566) );
  AND U12256 ( .A(\stack[1][9] ), .B(o[50]), .Z(n11564) );
  NAND U12257 ( .A(n11254), .B(n11253), .Z(n11258) );
  NAND U12258 ( .A(n11256), .B(n11255), .Z(n11257) );
  NAND U12259 ( .A(n11258), .B(n11257), .Z(n11563) );
  XOR U12260 ( .A(n11564), .B(n11563), .Z(n11565) );
  XOR U12261 ( .A(n11566), .B(n11565), .Z(n11569) );
  XOR U12262 ( .A(n11572), .B(n11571), .Z(n11578) );
  AND U12263 ( .A(\stack[1][7] ), .B(o[52]), .Z(n11575) );
  NAND U12264 ( .A(n11260), .B(n11259), .Z(n11264) );
  NAND U12265 ( .A(n11262), .B(n11261), .Z(n11263) );
  NAND U12266 ( .A(n11264), .B(n11263), .Z(n11576) );
  XOR U12267 ( .A(n11578), .B(n11577), .Z(n11266) );
  NAND U12268 ( .A(n11265), .B(n11266), .Z(n11268) );
  AND U12269 ( .A(\stack[1][6] ), .B(o[53]), .Z(n12537) );
  NAND U12270 ( .A(n12537), .B(n12538), .Z(n11267) );
  NAND U12271 ( .A(n11268), .B(n11267), .Z(n11269) );
  AND U12272 ( .A(\stack[1][6] ), .B(o[54]), .Z(n11270) );
  NAND U12273 ( .A(n11269), .B(n11270), .Z(n11582) );
  NAND U12274 ( .A(n11272), .B(n11271), .Z(n11276) );
  NAND U12275 ( .A(n11274), .B(n11273), .Z(n11275) );
  NAND U12276 ( .A(n11276), .B(n11275), .Z(n11595) );
  AND U12277 ( .A(\stack[1][12] ), .B(o[48]), .Z(n11596) );
  XOR U12278 ( .A(n11595), .B(n11596), .Z(n11598) );
  NAND U12279 ( .A(n11278), .B(n11277), .Z(n11282) );
  NAND U12280 ( .A(n11280), .B(n11279), .Z(n11281) );
  NAND U12281 ( .A(n11282), .B(n11281), .Z(n11869) );
  NAND U12282 ( .A(n11284), .B(n11283), .Z(n11288) );
  NAND U12283 ( .A(n11286), .B(n11285), .Z(n11287) );
  AND U12284 ( .A(n11288), .B(n11287), .Z(n11608) );
  NAND U12285 ( .A(\stack[1][16] ), .B(o[44]), .Z(n11607) );
  XOR U12286 ( .A(n11608), .B(n11607), .Z(n11610) );
  NAND U12287 ( .A(n11290), .B(n11289), .Z(n11294) );
  NAND U12288 ( .A(n11292), .B(n11291), .Z(n11293) );
  NAND U12289 ( .A(n11294), .B(n11293), .Z(n11863) );
  NAND U12290 ( .A(n11296), .B(n11295), .Z(n11300) );
  NAND U12291 ( .A(n11298), .B(n11297), .Z(n11299) );
  AND U12292 ( .A(n11300), .B(n11299), .Z(n11614) );
  NAND U12293 ( .A(\stack[1][18] ), .B(o[42]), .Z(n11613) );
  XOR U12294 ( .A(n11614), .B(n11613), .Z(n11616) );
  NAND U12295 ( .A(n11302), .B(n11301), .Z(n11306) );
  NAND U12296 ( .A(n11304), .B(n11303), .Z(n11305) );
  NAND U12297 ( .A(n11306), .B(n11305), .Z(n11619) );
  AND U12298 ( .A(\stack[1][20] ), .B(o[40]), .Z(n11620) );
  XOR U12299 ( .A(n11619), .B(n11620), .Z(n11622) );
  NAND U12300 ( .A(n11308), .B(n11307), .Z(n11312) );
  NAND U12301 ( .A(n11310), .B(n11309), .Z(n11311) );
  NAND U12302 ( .A(n11312), .B(n11311), .Z(n11851) );
  NAND U12303 ( .A(n11314), .B(n11313), .Z(n11318) );
  NAND U12304 ( .A(n11316), .B(n11315), .Z(n11317) );
  AND U12305 ( .A(n11318), .B(n11317), .Z(n11626) );
  NAND U12306 ( .A(\stack[1][22] ), .B(o[38]), .Z(n11625) );
  XOR U12307 ( .A(n11626), .B(n11625), .Z(n11628) );
  NAND U12308 ( .A(n11320), .B(n11319), .Z(n11324) );
  NAND U12309 ( .A(n11322), .B(n11321), .Z(n11323) );
  NAND U12310 ( .A(n11324), .B(n11323), .Z(n11631) );
  AND U12311 ( .A(\stack[1][24] ), .B(o[36]), .Z(n11632) );
  XOR U12312 ( .A(n11631), .B(n11632), .Z(n11634) );
  NAND U12313 ( .A(n11326), .B(n11325), .Z(n11330) );
  NAND U12314 ( .A(n11328), .B(n11327), .Z(n11329) );
  NAND U12315 ( .A(n11330), .B(n11329), .Z(n11637) );
  AND U12316 ( .A(\stack[1][26] ), .B(o[34]), .Z(n11638) );
  XOR U12317 ( .A(n11637), .B(n11638), .Z(n11640) );
  NAND U12318 ( .A(n11332), .B(n11331), .Z(n11336) );
  NAND U12319 ( .A(n11334), .B(n11333), .Z(n11335) );
  NAND U12320 ( .A(n11336), .B(n11335), .Z(n11643) );
  AND U12321 ( .A(\stack[1][28] ), .B(o[32]), .Z(n11644) );
  XOR U12322 ( .A(n11643), .B(n11644), .Z(n11646) );
  NAND U12323 ( .A(n11338), .B(n11337), .Z(n11342) );
  NAND U12324 ( .A(n11340), .B(n11339), .Z(n11341) );
  NAND U12325 ( .A(n11342), .B(n11341), .Z(n11666) );
  AND U12326 ( .A(o[26]), .B(\stack[1][34] ), .Z(n11667) );
  XOR U12327 ( .A(n11666), .B(n11667), .Z(n11669) );
  AND U12328 ( .A(o[24]), .B(\stack[1][36] ), .Z(n11681) );
  NAND U12329 ( .A(o[22]), .B(\stack[1][38] ), .Z(n11686) );
  NAND U12330 ( .A(n11344), .B(n11343), .Z(n11348) );
  NAND U12331 ( .A(n11346), .B(n11345), .Z(n11347) );
  NAND U12332 ( .A(n11348), .B(n11347), .Z(n11684) );
  NAND U12333 ( .A(o[21]), .B(\stack[1][39] ), .Z(n11692) );
  AND U12334 ( .A(o[18]), .B(\stack[1][42] ), .Z(n11799) );
  NAND U12335 ( .A(n11350), .B(n11349), .Z(n11354) );
  NANDN U12336 ( .A(n11352), .B(n11351), .Z(n11353) );
  AND U12337 ( .A(n11354), .B(n11353), .Z(n11797) );
  NAND U12338 ( .A(o[17]), .B(\stack[1][43] ), .Z(n11698) );
  NAND U12339 ( .A(n11356), .B(n11355), .Z(n11360) );
  NAND U12340 ( .A(n11358), .B(n11357), .Z(n11359) );
  NAND U12341 ( .A(n11360), .B(n11359), .Z(n11704) );
  NAND U12342 ( .A(n11362), .B(n11361), .Z(n11366) );
  NAND U12343 ( .A(n11364), .B(n11363), .Z(n11365) );
  NAND U12344 ( .A(n11366), .B(n11365), .Z(n11710) );
  NAND U12345 ( .A(n11368), .B(n11367), .Z(n11372) );
  NAND U12346 ( .A(n11370), .B(n11369), .Z(n11371) );
  NAND U12347 ( .A(n11372), .B(n11371), .Z(n11714) );
  AND U12348 ( .A(o[12]), .B(\stack[1][48] ), .Z(n11723) );
  NAND U12349 ( .A(n11374), .B(n11373), .Z(n11378) );
  NAND U12350 ( .A(n11376), .B(n11375), .Z(n11377) );
  AND U12351 ( .A(n11378), .B(n11377), .Z(n11721) );
  NAND U12352 ( .A(o[11]), .B(\stack[1][49] ), .Z(n11728) );
  NAND U12353 ( .A(n11380), .B(n11379), .Z(n11384) );
  NAND U12354 ( .A(n11382), .B(n11381), .Z(n11383) );
  AND U12355 ( .A(n11384), .B(n11383), .Z(n11727) );
  NAND U12356 ( .A(n11386), .B(n11385), .Z(n11390) );
  NAND U12357 ( .A(n11388), .B(n11387), .Z(n11389) );
  AND U12358 ( .A(n11390), .B(n11389), .Z(n11732) );
  NAND U12359 ( .A(o[9]), .B(\stack[1][51] ), .Z(n11740) );
  NAND U12360 ( .A(n11392), .B(n11391), .Z(n11396) );
  NAND U12361 ( .A(n11394), .B(n11393), .Z(n11395) );
  NAND U12362 ( .A(n11396), .B(n11395), .Z(n11746) );
  AND U12363 ( .A(o[6]), .B(\stack[1][54] ), .Z(n11753) );
  NAND U12364 ( .A(n11398), .B(n11397), .Z(n11402) );
  NAND U12365 ( .A(n11400), .B(n11399), .Z(n11401) );
  NAND U12366 ( .A(n11402), .B(n11401), .Z(n11778) );
  NANDN U12367 ( .A(n11403), .B(n11762), .Z(n11407) );
  NANDN U12368 ( .A(n11405), .B(n11404), .Z(n11406) );
  NAND U12369 ( .A(n11407), .B(n11406), .Z(n11772) );
  AND U12370 ( .A(o[2]), .B(\stack[1][58] ), .Z(n11763) );
  AND U12371 ( .A(n11408), .B(n11410), .Z(n11409) );
  AND U12372 ( .A(o[1]), .B(\stack[1][60] ), .Z(n11769) );
  NAND U12373 ( .A(n11767), .B(n11769), .Z(n12046) );
  XOR U12374 ( .A(n11409), .B(n12046), .Z(n11412) );
  NAND U12375 ( .A(o[0]), .B(\stack[1][60] ), .Z(n12052) );
  NANDN U12376 ( .A(n11410), .B(n12052), .Z(n11411) );
  NAND U12377 ( .A(n11412), .B(n11411), .Z(n11764) );
  XNOR U12378 ( .A(n11763), .B(n11764), .Z(n11773) );
  XOR U12379 ( .A(n11772), .B(n11773), .Z(n11775) );
  AND U12380 ( .A(o[3]), .B(\stack[1][57] ), .Z(n11774) );
  XOR U12381 ( .A(n11775), .B(n11774), .Z(n11757) );
  NAND U12382 ( .A(n11414), .B(n11413), .Z(n11418) );
  NAND U12383 ( .A(n11416), .B(n11415), .Z(n11417) );
  NAND U12384 ( .A(n11418), .B(n11417), .Z(n11756) );
  XOR U12385 ( .A(n11757), .B(n11756), .Z(n11759) );
  AND U12386 ( .A(o[4]), .B(\stack[1][56] ), .Z(n11758) );
  XOR U12387 ( .A(n11759), .B(n11758), .Z(n11779) );
  XOR U12388 ( .A(n11778), .B(n11779), .Z(n11781) );
  AND U12389 ( .A(o[5]), .B(\stack[1][55] ), .Z(n11780) );
  XOR U12390 ( .A(n11781), .B(n11780), .Z(n11751) );
  NAND U12391 ( .A(n11420), .B(n11419), .Z(n11424) );
  NAND U12392 ( .A(n11422), .B(n11421), .Z(n11423) );
  NAND U12393 ( .A(n11424), .B(n11423), .Z(n11750) );
  XOR U12394 ( .A(n11751), .B(n11750), .Z(n11752) );
  XOR U12395 ( .A(n11753), .B(n11752), .Z(n11745) );
  AND U12396 ( .A(o[7]), .B(\stack[1][53] ), .Z(n11744) );
  XOR U12397 ( .A(n11745), .B(n11744), .Z(n11747) );
  XOR U12398 ( .A(n11746), .B(n11747), .Z(n11785) );
  AND U12399 ( .A(o[8]), .B(\stack[1][52] ), .Z(n11784) );
  XOR U12400 ( .A(n11785), .B(n11784), .Z(n11787) );
  NAND U12401 ( .A(n11426), .B(n11425), .Z(n11430) );
  NAND U12402 ( .A(n11428), .B(n11427), .Z(n11429) );
  NAND U12403 ( .A(n11430), .B(n11429), .Z(n11786) );
  XNOR U12404 ( .A(n11787), .B(n11786), .Z(n11739) );
  NAND U12405 ( .A(n11432), .B(n11431), .Z(n11436) );
  NAND U12406 ( .A(n11434), .B(n11433), .Z(n11435) );
  AND U12407 ( .A(n11436), .B(n11435), .Z(n11738) );
  XNOR U12408 ( .A(n11740), .B(n11741), .Z(n11733) );
  AND U12409 ( .A(o[10]), .B(\stack[1][50] ), .Z(n11734) );
  XNOR U12410 ( .A(n11735), .B(n11734), .Z(n11726) );
  XOR U12411 ( .A(n11727), .B(n11726), .Z(n11729) );
  XNOR U12412 ( .A(n11728), .B(n11729), .Z(n11720) );
  XOR U12413 ( .A(n11721), .B(n11720), .Z(n11722) );
  XOR U12414 ( .A(n11723), .B(n11722), .Z(n11715) );
  XOR U12415 ( .A(n11714), .B(n11715), .Z(n11717) );
  AND U12416 ( .A(o[13]), .B(\stack[1][47] ), .Z(n11716) );
  XOR U12417 ( .A(n11717), .B(n11716), .Z(n11709) );
  AND U12418 ( .A(o[14]), .B(\stack[1][46] ), .Z(n11708) );
  XOR U12419 ( .A(n11709), .B(n11708), .Z(n11711) );
  XOR U12420 ( .A(n11710), .B(n11711), .Z(n11703) );
  AND U12421 ( .A(o[15]), .B(\stack[1][45] ), .Z(n11702) );
  XOR U12422 ( .A(n11703), .B(n11702), .Z(n11705) );
  XOR U12423 ( .A(n11704), .B(n11705), .Z(n11791) );
  AND U12424 ( .A(o[16]), .B(\stack[1][44] ), .Z(n11790) );
  XOR U12425 ( .A(n11791), .B(n11790), .Z(n11793) );
  NAND U12426 ( .A(n11438), .B(n11437), .Z(n11442) );
  NAND U12427 ( .A(n11440), .B(n11439), .Z(n11441) );
  NAND U12428 ( .A(n11442), .B(n11441), .Z(n11792) );
  XNOR U12429 ( .A(n11793), .B(n11792), .Z(n11697) );
  NAND U12430 ( .A(n11444), .B(n11443), .Z(n11448) );
  NAND U12431 ( .A(n11446), .B(n11445), .Z(n11447) );
  AND U12432 ( .A(n11448), .B(n11447), .Z(n11696) );
  XOR U12433 ( .A(n11698), .B(n11699), .Z(n11796) );
  XOR U12434 ( .A(n11797), .B(n11796), .Z(n11798) );
  XOR U12435 ( .A(n11799), .B(n11798), .Z(n11803) );
  AND U12436 ( .A(o[19]), .B(\stack[1][41] ), .Z(n11802) );
  XOR U12437 ( .A(n11803), .B(n11802), .Z(n11805) );
  NAND U12438 ( .A(n11450), .B(n11449), .Z(n11454) );
  NAND U12439 ( .A(n11452), .B(n11451), .Z(n11453) );
  NAND U12440 ( .A(n11454), .B(n11453), .Z(n11804) );
  XOR U12441 ( .A(n11805), .B(n11804), .Z(n11809) );
  AND U12442 ( .A(o[20]), .B(\stack[1][40] ), .Z(n11808) );
  XOR U12443 ( .A(n11809), .B(n11808), .Z(n11811) );
  NAND U12444 ( .A(n11456), .B(n11455), .Z(n11460) );
  NAND U12445 ( .A(n11458), .B(n11457), .Z(n11459) );
  NAND U12446 ( .A(n11460), .B(n11459), .Z(n11810) );
  XNOR U12447 ( .A(n11811), .B(n11810), .Z(n11691) );
  NAND U12448 ( .A(n11462), .B(n11461), .Z(n11466) );
  NAND U12449 ( .A(n11464), .B(n11463), .Z(n11465) );
  AND U12450 ( .A(n11466), .B(n11465), .Z(n11690) );
  XOR U12451 ( .A(n11692), .B(n11693), .Z(n11685) );
  XOR U12452 ( .A(n11684), .B(n11685), .Z(n11687) );
  XNOR U12453 ( .A(n11686), .B(n11687), .Z(n11817) );
  AND U12454 ( .A(o[23]), .B(\stack[1][37] ), .Z(n11815) );
  NAND U12455 ( .A(n11468), .B(n11467), .Z(n11472) );
  NAND U12456 ( .A(n11470), .B(n11469), .Z(n11471) );
  NAND U12457 ( .A(n11472), .B(n11471), .Z(n11814) );
  XOR U12458 ( .A(n11815), .B(n11814), .Z(n11816) );
  NAND U12459 ( .A(n11474), .B(n11473), .Z(n11478) );
  NAND U12460 ( .A(n11476), .B(n11475), .Z(n11477) );
  NAND U12461 ( .A(n11478), .B(n11477), .Z(n11678) );
  XOR U12462 ( .A(n11679), .B(n11678), .Z(n11680) );
  XOR U12463 ( .A(n11681), .B(n11680), .Z(n11675) );
  AND U12464 ( .A(o[25]), .B(\stack[1][35] ), .Z(n11673) );
  NAND U12465 ( .A(n11480), .B(n11479), .Z(n11484) );
  NAND U12466 ( .A(n11482), .B(n11481), .Z(n11483) );
  NAND U12467 ( .A(n11484), .B(n11483), .Z(n11672) );
  XOR U12468 ( .A(n11673), .B(n11672), .Z(n11674) );
  XOR U12469 ( .A(n11675), .B(n11674), .Z(n11668) );
  XOR U12470 ( .A(n11669), .B(n11668), .Z(n11821) );
  NAND U12471 ( .A(n11486), .B(n11485), .Z(n11490) );
  NAND U12472 ( .A(n11488), .B(n11487), .Z(n11489) );
  NAND U12473 ( .A(n11490), .B(n11489), .Z(n11820) );
  XOR U12474 ( .A(n11821), .B(n11820), .Z(n11823) );
  AND U12475 ( .A(o[27]), .B(\stack[1][33] ), .Z(n11822) );
  XOR U12476 ( .A(n11823), .B(n11822), .Z(n11662) );
  NAND U12477 ( .A(n11492), .B(n11491), .Z(n11496) );
  NAND U12478 ( .A(n11494), .B(n11493), .Z(n11495) );
  NAND U12479 ( .A(n11496), .B(n11495), .Z(n11660) );
  AND U12480 ( .A(o[28]), .B(\stack[1][32] ), .Z(n11661) );
  XOR U12481 ( .A(n11660), .B(n11661), .Z(n11663) );
  NAND U12482 ( .A(n11498), .B(n11497), .Z(n11502) );
  NAND U12483 ( .A(n11500), .B(n11499), .Z(n11501) );
  NAND U12484 ( .A(n11502), .B(n11501), .Z(n11654) );
  XOR U12485 ( .A(n11655), .B(n11654), .Z(n11657) );
  AND U12486 ( .A(\stack[1][31] ), .B(o[29]), .Z(n11656) );
  XOR U12487 ( .A(n11657), .B(n11656), .Z(n11651) );
  AND U12488 ( .A(\stack[1][30] ), .B(o[30]), .Z(n16172) );
  NAND U12489 ( .A(n11504), .B(n11503), .Z(n11508) );
  NAND U12490 ( .A(n11506), .B(n11505), .Z(n11507) );
  NAND U12491 ( .A(n11508), .B(n11507), .Z(n11649) );
  XOR U12492 ( .A(n16172), .B(n11649), .Z(n11650) );
  XOR U12493 ( .A(n11651), .B(n11650), .Z(n11827) );
  NAND U12494 ( .A(n11510), .B(n11509), .Z(n11514) );
  NAND U12495 ( .A(n11512), .B(n11511), .Z(n11513) );
  NAND U12496 ( .A(n11514), .B(n11513), .Z(n11826) );
  XOR U12497 ( .A(n11827), .B(n11826), .Z(n11829) );
  AND U12498 ( .A(\stack[1][29] ), .B(o[31]), .Z(n11828) );
  XOR U12499 ( .A(n11829), .B(n11828), .Z(n11645) );
  XOR U12500 ( .A(n11646), .B(n11645), .Z(n11833) );
  NAND U12501 ( .A(n11516), .B(n11515), .Z(n11520) );
  NAND U12502 ( .A(n11518), .B(n11517), .Z(n11519) );
  NAND U12503 ( .A(n11520), .B(n11519), .Z(n11832) );
  XOR U12504 ( .A(n11833), .B(n11832), .Z(n11835) );
  AND U12505 ( .A(\stack[1][27] ), .B(o[33]), .Z(n11834) );
  XOR U12506 ( .A(n11835), .B(n11834), .Z(n11639) );
  XOR U12507 ( .A(n11640), .B(n11639), .Z(n11839) );
  NAND U12508 ( .A(n11522), .B(n11521), .Z(n11526) );
  NAND U12509 ( .A(n11524), .B(n11523), .Z(n11525) );
  NAND U12510 ( .A(n11526), .B(n11525), .Z(n11838) );
  XOR U12511 ( .A(n11839), .B(n11838), .Z(n11841) );
  AND U12512 ( .A(\stack[1][25] ), .B(o[35]), .Z(n11840) );
  XOR U12513 ( .A(n11841), .B(n11840), .Z(n11633) );
  XOR U12514 ( .A(n11634), .B(n11633), .Z(n11845) );
  NAND U12515 ( .A(n11528), .B(n11527), .Z(n11532) );
  NAND U12516 ( .A(n11530), .B(n11529), .Z(n11531) );
  NAND U12517 ( .A(n11532), .B(n11531), .Z(n11844) );
  XOR U12518 ( .A(n11845), .B(n11844), .Z(n11847) );
  AND U12519 ( .A(\stack[1][23] ), .B(o[37]), .Z(n11846) );
  XNOR U12520 ( .A(n11847), .B(n11846), .Z(n11627) );
  XNOR U12521 ( .A(n11628), .B(n11627), .Z(n11850) );
  XOR U12522 ( .A(n11851), .B(n11850), .Z(n11853) );
  AND U12523 ( .A(\stack[1][21] ), .B(o[39]), .Z(n11852) );
  XOR U12524 ( .A(n11853), .B(n11852), .Z(n11621) );
  XOR U12525 ( .A(n11622), .B(n11621), .Z(n11857) );
  NAND U12526 ( .A(n11534), .B(n11533), .Z(n11538) );
  NAND U12527 ( .A(n11536), .B(n11535), .Z(n11537) );
  NAND U12528 ( .A(n11538), .B(n11537), .Z(n11856) );
  XOR U12529 ( .A(n11857), .B(n11856), .Z(n11859) );
  AND U12530 ( .A(\stack[1][19] ), .B(o[41]), .Z(n11858) );
  XNOR U12531 ( .A(n11859), .B(n11858), .Z(n11615) );
  XNOR U12532 ( .A(n11616), .B(n11615), .Z(n11862) );
  XOR U12533 ( .A(n11863), .B(n11862), .Z(n11865) );
  AND U12534 ( .A(\stack[1][17] ), .B(o[43]), .Z(n11864) );
  XNOR U12535 ( .A(n11865), .B(n11864), .Z(n11609) );
  XNOR U12536 ( .A(n11610), .B(n11609), .Z(n11868) );
  XOR U12537 ( .A(n11869), .B(n11868), .Z(n11871) );
  AND U12538 ( .A(\stack[1][15] ), .B(o[45]), .Z(n11870) );
  XNOR U12539 ( .A(n11871), .B(n11870), .Z(n11604) );
  NAND U12540 ( .A(n11540), .B(n11539), .Z(n11544) );
  NAND U12541 ( .A(n11542), .B(n11541), .Z(n11543) );
  AND U12542 ( .A(n11544), .B(n11543), .Z(n11602) );
  NAND U12543 ( .A(\stack[1][14] ), .B(o[46]), .Z(n11601) );
  XOR U12544 ( .A(n11602), .B(n11601), .Z(n11603) );
  NAND U12545 ( .A(n11546), .B(n11545), .Z(n11550) );
  NAND U12546 ( .A(n11548), .B(n11547), .Z(n11549) );
  NAND U12547 ( .A(n11550), .B(n11549), .Z(n11874) );
  AND U12548 ( .A(\stack[1][13] ), .B(o[47]), .Z(n11876) );
  XOR U12549 ( .A(n11877), .B(n11876), .Z(n11597) );
  XOR U12550 ( .A(n11598), .B(n11597), .Z(n11881) );
  NAND U12551 ( .A(n11552), .B(n11551), .Z(n11556) );
  NAND U12552 ( .A(n11554), .B(n11553), .Z(n11555) );
  NAND U12553 ( .A(n11556), .B(n11555), .Z(n11880) );
  XOR U12554 ( .A(n11881), .B(n11880), .Z(n11883) );
  AND U12555 ( .A(\stack[1][11] ), .B(o[49]), .Z(n11882) );
  XOR U12556 ( .A(n11883), .B(n11882), .Z(n11591) );
  NAND U12557 ( .A(n11558), .B(n11557), .Z(n11562) );
  NAND U12558 ( .A(n11560), .B(n11559), .Z(n11561) );
  NAND U12559 ( .A(n11562), .B(n11561), .Z(n11589) );
  AND U12560 ( .A(\stack[1][10] ), .B(o[50]), .Z(n11590) );
  XOR U12561 ( .A(n11589), .B(n11590), .Z(n11592) );
  NAND U12562 ( .A(n11564), .B(n11563), .Z(n11568) );
  NAND U12563 ( .A(n11566), .B(n11565), .Z(n11567) );
  NAND U12564 ( .A(n11568), .B(n11567), .Z(n11886) );
  XOR U12565 ( .A(n11887), .B(n11886), .Z(n11889) );
  AND U12566 ( .A(\stack[1][9] ), .B(o[51]), .Z(n11888) );
  XNOR U12567 ( .A(n11889), .B(n11888), .Z(n11586) );
  NAND U12568 ( .A(n11570), .B(n11569), .Z(n11574) );
  NAND U12569 ( .A(n11572), .B(n11571), .Z(n11573) );
  AND U12570 ( .A(n11574), .B(n11573), .Z(n11583) );
  NAND U12571 ( .A(\stack[1][8] ), .B(o[52]), .Z(n11584) );
  NAND U12572 ( .A(n11576), .B(n11575), .Z(n11580) );
  NAND U12573 ( .A(n11578), .B(n11577), .Z(n11579) );
  NAND U12574 ( .A(n11580), .B(n11579), .Z(n11892) );
  XOR U12575 ( .A(n11893), .B(n11892), .Z(n11894) );
  AND U12576 ( .A(\stack[1][7] ), .B(o[53]), .Z(n11895) );
  NAND U12577 ( .A(n12544), .B(n12543), .Z(n11581) );
  NAND U12578 ( .A(n11582), .B(n11581), .Z(n11898) );
  AND U12579 ( .A(\stack[1][8] ), .B(o[53]), .Z(n11905) );
  NAND U12580 ( .A(n11584), .B(n11583), .Z(n11588) );
  NAND U12581 ( .A(n11586), .B(n11585), .Z(n11587) );
  AND U12582 ( .A(n11588), .B(n11587), .Z(n11903) );
  AND U12583 ( .A(\stack[1][10] ), .B(o[51]), .Z(n11910) );
  NAND U12584 ( .A(n11590), .B(n11589), .Z(n11594) );
  NAND U12585 ( .A(n11592), .B(n11591), .Z(n11593) );
  NAND U12586 ( .A(n11594), .B(n11593), .Z(n11908) );
  AND U12587 ( .A(\stack[1][12] ), .B(o[49]), .Z(n11916) );
  NAND U12588 ( .A(n11596), .B(n11595), .Z(n11600) );
  NAND U12589 ( .A(n11598), .B(n11597), .Z(n11599) );
  NAND U12590 ( .A(n11600), .B(n11599), .Z(n11914) );
  NAND U12591 ( .A(n11602), .B(n11601), .Z(n11606) );
  NAND U12592 ( .A(n11604), .B(n11603), .Z(n11605) );
  AND U12593 ( .A(n11606), .B(n11605), .Z(n12194) );
  NAND U12594 ( .A(n11608), .B(n11607), .Z(n11612) );
  NAND U12595 ( .A(n11610), .B(n11609), .Z(n11611) );
  AND U12596 ( .A(n11612), .B(n11611), .Z(n12182) );
  NAND U12597 ( .A(n11614), .B(n11613), .Z(n11618) );
  NAND U12598 ( .A(n11616), .B(n11615), .Z(n11617) );
  AND U12599 ( .A(n11618), .B(n11617), .Z(n11921) );
  NAND U12600 ( .A(n11620), .B(n11619), .Z(n11624) );
  NAND U12601 ( .A(n11622), .B(n11621), .Z(n11623) );
  NAND U12602 ( .A(n11624), .B(n11623), .Z(n12163) );
  AND U12603 ( .A(\stack[1][22] ), .B(o[39]), .Z(n11929) );
  NAND U12604 ( .A(n11626), .B(n11625), .Z(n11630) );
  NAND U12605 ( .A(n11628), .B(n11627), .Z(n11629) );
  AND U12606 ( .A(n11630), .B(n11629), .Z(n11927) );
  AND U12607 ( .A(\stack[1][24] ), .B(o[37]), .Z(n11934) );
  NAND U12608 ( .A(n11632), .B(n11631), .Z(n11636) );
  NAND U12609 ( .A(n11634), .B(n11633), .Z(n11635) );
  NAND U12610 ( .A(n11636), .B(n11635), .Z(n11932) );
  AND U12611 ( .A(\stack[1][26] ), .B(o[35]), .Z(n11940) );
  NAND U12612 ( .A(n11638), .B(n11637), .Z(n11642) );
  NAND U12613 ( .A(n11640), .B(n11639), .Z(n11641) );
  NAND U12614 ( .A(n11642), .B(n11641), .Z(n11938) );
  NAND U12615 ( .A(n11644), .B(n11643), .Z(n11648) );
  NAND U12616 ( .A(n11646), .B(n11645), .Z(n11647) );
  NAND U12617 ( .A(n11648), .B(n11647), .Z(n11944) );
  AND U12618 ( .A(\stack[1][30] ), .B(o[31]), .Z(n12129) );
  NAND U12619 ( .A(n16172), .B(n11649), .Z(n11653) );
  NAND U12620 ( .A(n11651), .B(n11650), .Z(n11652) );
  NAND U12621 ( .A(n11653), .B(n11652), .Z(n12127) );
  AND U12622 ( .A(\stack[1][31] ), .B(o[30]), .Z(n11951) );
  NAND U12623 ( .A(n11655), .B(n11654), .Z(n11659) );
  NAND U12624 ( .A(n11657), .B(n11656), .Z(n11658) );
  NAND U12625 ( .A(n11659), .B(n11658), .Z(n11950) );
  XOR U12626 ( .A(n11951), .B(n11950), .Z(n11953) );
  AND U12627 ( .A(o[29]), .B(\stack[1][32] ), .Z(n11958) );
  NAND U12628 ( .A(n11661), .B(n11660), .Z(n11665) );
  NAND U12629 ( .A(n11663), .B(n11662), .Z(n11664) );
  NAND U12630 ( .A(n11665), .B(n11664), .Z(n11956) );
  AND U12631 ( .A(o[27]), .B(\stack[1][34] ), .Z(n11964) );
  NAND U12632 ( .A(n11667), .B(n11666), .Z(n11671) );
  NAND U12633 ( .A(n11669), .B(n11668), .Z(n11670) );
  NAND U12634 ( .A(n11671), .B(n11670), .Z(n11962) );
  NAND U12635 ( .A(n11673), .B(n11672), .Z(n11677) );
  NAND U12636 ( .A(n11675), .B(n11674), .Z(n11676) );
  NAND U12637 ( .A(n11677), .B(n11676), .Z(n12117) );
  NAND U12638 ( .A(n11679), .B(n11678), .Z(n11683) );
  NAND U12639 ( .A(n11681), .B(n11680), .Z(n11682) );
  NAND U12640 ( .A(n11683), .B(n11682), .Z(n12109) );
  NAND U12641 ( .A(o[23]), .B(\stack[1][38] ), .Z(n12099) );
  NAND U12642 ( .A(n11685), .B(n11684), .Z(n11689) );
  NAND U12643 ( .A(n11687), .B(n11686), .Z(n11688) );
  NAND U12644 ( .A(n11689), .B(n11688), .Z(n12098) );
  AND U12645 ( .A(o[22]), .B(\stack[1][39] ), .Z(n11971) );
  NAND U12646 ( .A(n11691), .B(n11690), .Z(n11695) );
  NAND U12647 ( .A(n11693), .B(n11692), .Z(n11694) );
  AND U12648 ( .A(n11695), .B(n11694), .Z(n11968) );
  NAND U12649 ( .A(o[21]), .B(\stack[1][40] ), .Z(n11976) );
  AND U12650 ( .A(o[18]), .B(\stack[1][43] ), .Z(n12088) );
  NAND U12651 ( .A(n11697), .B(n11696), .Z(n11701) );
  NANDN U12652 ( .A(n11699), .B(n11698), .Z(n11700) );
  AND U12653 ( .A(n11701), .B(n11700), .Z(n12086) );
  NAND U12654 ( .A(o[17]), .B(\stack[1][44] ), .Z(n11988) );
  NAND U12655 ( .A(n11703), .B(n11702), .Z(n11707) );
  NAND U12656 ( .A(n11705), .B(n11704), .Z(n11706) );
  NAND U12657 ( .A(n11707), .B(n11706), .Z(n12081) );
  NAND U12658 ( .A(n11709), .B(n11708), .Z(n11713) );
  NAND U12659 ( .A(n11711), .B(n11710), .Z(n11712) );
  NAND U12660 ( .A(n11713), .B(n11712), .Z(n12075) );
  NAND U12661 ( .A(n11715), .B(n11714), .Z(n11719) );
  NAND U12662 ( .A(n11717), .B(n11716), .Z(n11718) );
  NAND U12663 ( .A(n11719), .B(n11718), .Z(n11994) );
  AND U12664 ( .A(o[13]), .B(\stack[1][48] ), .Z(n12000) );
  NAND U12665 ( .A(n11721), .B(n11720), .Z(n11725) );
  NAND U12666 ( .A(n11723), .B(n11722), .Z(n11724) );
  NAND U12667 ( .A(n11725), .B(n11724), .Z(n11998) );
  AND U12668 ( .A(o[12]), .B(\stack[1][49] ), .Z(n12007) );
  NAND U12669 ( .A(n11727), .B(n11726), .Z(n11731) );
  NAND U12670 ( .A(n11729), .B(n11728), .Z(n11730) );
  AND U12671 ( .A(n11731), .B(n11730), .Z(n12004) );
  NAND U12672 ( .A(n11733), .B(n11732), .Z(n11737) );
  NAND U12673 ( .A(n11735), .B(n11734), .Z(n11736) );
  AND U12674 ( .A(n11737), .B(n11736), .Z(n12010) );
  AND U12675 ( .A(o[10]), .B(\stack[1][51] ), .Z(n12019) );
  NAND U12676 ( .A(n11739), .B(n11738), .Z(n11743) );
  NAND U12677 ( .A(n11741), .B(n11740), .Z(n11742) );
  AND U12678 ( .A(n11743), .B(n11742), .Z(n12017) );
  NAND U12679 ( .A(o[9]), .B(\stack[1][52] ), .Z(n12024) );
  NAND U12680 ( .A(n11745), .B(n11744), .Z(n11749) );
  NAND U12681 ( .A(n11747), .B(n11746), .Z(n11748) );
  NAND U12682 ( .A(n11749), .B(n11748), .Z(n12069) );
  NAND U12683 ( .A(n11751), .B(n11750), .Z(n11755) );
  NAND U12684 ( .A(n11753), .B(n11752), .Z(n11754) );
  NAND U12685 ( .A(n11755), .B(n11754), .Z(n12030) );
  AND U12686 ( .A(o[6]), .B(\stack[1][55] ), .Z(n12037) );
  NAND U12687 ( .A(n11757), .B(n11756), .Z(n11761) );
  NAND U12688 ( .A(n11759), .B(n11758), .Z(n11760) );
  NAND U12689 ( .A(n11761), .B(n11760), .Z(n12040) );
  AND U12690 ( .A(o[4]), .B(\stack[1][57] ), .Z(n12064) );
  NANDN U12691 ( .A(n11762), .B(n12046), .Z(n11766) );
  NANDN U12692 ( .A(n11764), .B(n11763), .Z(n11765) );
  NAND U12693 ( .A(n11766), .B(n11765), .Z(n12055) );
  AND U12694 ( .A(o[2]), .B(\stack[1][59] ), .Z(n12047) );
  AND U12695 ( .A(n11767), .B(n11769), .Z(n11768) );
  AND U12696 ( .A(o[1]), .B(\stack[1][61] ), .Z(n12051) );
  XNOR U12697 ( .A(n11768), .B(n12683), .Z(n11771) );
  NAND U12698 ( .A(o[0]), .B(\stack[1][61] ), .Z(n12705) );
  NANDN U12699 ( .A(n11769), .B(n12705), .Z(n11770) );
  NAND U12700 ( .A(n11771), .B(n11770), .Z(n12048) );
  XNOR U12701 ( .A(n12047), .B(n12048), .Z(n12056) );
  XOR U12702 ( .A(n12055), .B(n12056), .Z(n12058) );
  AND U12703 ( .A(o[3]), .B(\stack[1][58] ), .Z(n12057) );
  XOR U12704 ( .A(n12058), .B(n12057), .Z(n12062) );
  NAND U12705 ( .A(n11773), .B(n11772), .Z(n11777) );
  NAND U12706 ( .A(n11775), .B(n11774), .Z(n11776) );
  NAND U12707 ( .A(n11777), .B(n11776), .Z(n12061) );
  XOR U12708 ( .A(n12062), .B(n12061), .Z(n12063) );
  XOR U12709 ( .A(n12064), .B(n12063), .Z(n12041) );
  XOR U12710 ( .A(n12040), .B(n12041), .Z(n12043) );
  AND U12711 ( .A(o[5]), .B(\stack[1][56] ), .Z(n12042) );
  XOR U12712 ( .A(n12043), .B(n12042), .Z(n12035) );
  NAND U12713 ( .A(n11779), .B(n11778), .Z(n11783) );
  NAND U12714 ( .A(n11781), .B(n11780), .Z(n11782) );
  NAND U12715 ( .A(n11783), .B(n11782), .Z(n12034) );
  XOR U12716 ( .A(n12035), .B(n12034), .Z(n12036) );
  XOR U12717 ( .A(n12037), .B(n12036), .Z(n12029) );
  AND U12718 ( .A(o[7]), .B(\stack[1][54] ), .Z(n12028) );
  XOR U12719 ( .A(n12029), .B(n12028), .Z(n12031) );
  XOR U12720 ( .A(n12030), .B(n12031), .Z(n12068) );
  AND U12721 ( .A(o[8]), .B(\stack[1][53] ), .Z(n12067) );
  XOR U12722 ( .A(n12068), .B(n12067), .Z(n12070) );
  XNOR U12723 ( .A(n12069), .B(n12070), .Z(n12023) );
  NAND U12724 ( .A(n11785), .B(n11784), .Z(n11789) );
  NAND U12725 ( .A(n11787), .B(n11786), .Z(n11788) );
  AND U12726 ( .A(n11789), .B(n11788), .Z(n12022) );
  XOR U12727 ( .A(n12024), .B(n12025), .Z(n12016) );
  XOR U12728 ( .A(n12017), .B(n12016), .Z(n12018) );
  XNOR U12729 ( .A(n12019), .B(n12018), .Z(n12011) );
  NAND U12730 ( .A(o[11]), .B(\stack[1][50] ), .Z(n12012) );
  XNOR U12731 ( .A(n12013), .B(n12012), .Z(n12005) );
  XOR U12732 ( .A(n12007), .B(n12006), .Z(n11999) );
  XOR U12733 ( .A(n11998), .B(n11999), .Z(n12001) );
  AND U12734 ( .A(o[14]), .B(\stack[1][47] ), .Z(n11992) );
  XOR U12735 ( .A(n11993), .B(n11992), .Z(n11995) );
  XOR U12736 ( .A(n11994), .B(n11995), .Z(n12074) );
  AND U12737 ( .A(o[15]), .B(\stack[1][46] ), .Z(n12073) );
  XOR U12738 ( .A(n12074), .B(n12073), .Z(n12076) );
  XOR U12739 ( .A(n12075), .B(n12076), .Z(n12080) );
  AND U12740 ( .A(o[16]), .B(\stack[1][45] ), .Z(n12079) );
  XOR U12741 ( .A(n12080), .B(n12079), .Z(n12082) );
  XNOR U12742 ( .A(n12081), .B(n12082), .Z(n11987) );
  NAND U12743 ( .A(n11791), .B(n11790), .Z(n11795) );
  NAND U12744 ( .A(n11793), .B(n11792), .Z(n11794) );
  AND U12745 ( .A(n11795), .B(n11794), .Z(n11986) );
  XOR U12746 ( .A(n11988), .B(n11989), .Z(n12085) );
  XOR U12747 ( .A(n12086), .B(n12085), .Z(n12087) );
  XOR U12748 ( .A(n12088), .B(n12087), .Z(n11981) );
  AND U12749 ( .A(o[19]), .B(\stack[1][42] ), .Z(n11980) );
  XOR U12750 ( .A(n11981), .B(n11980), .Z(n11983) );
  NAND U12751 ( .A(n11797), .B(n11796), .Z(n11801) );
  NAND U12752 ( .A(n11799), .B(n11798), .Z(n11800) );
  NAND U12753 ( .A(n11801), .B(n11800), .Z(n11982) );
  XOR U12754 ( .A(n11983), .B(n11982), .Z(n12092) );
  AND U12755 ( .A(o[20]), .B(\stack[1][41] ), .Z(n12091) );
  XOR U12756 ( .A(n12092), .B(n12091), .Z(n12094) );
  NAND U12757 ( .A(n11803), .B(n11802), .Z(n11807) );
  NAND U12758 ( .A(n11805), .B(n11804), .Z(n11806) );
  NAND U12759 ( .A(n11807), .B(n11806), .Z(n12093) );
  XNOR U12760 ( .A(n12094), .B(n12093), .Z(n11975) );
  NAND U12761 ( .A(n11809), .B(n11808), .Z(n11813) );
  NAND U12762 ( .A(n11811), .B(n11810), .Z(n11812) );
  AND U12763 ( .A(n11813), .B(n11812), .Z(n11974) );
  XNOR U12764 ( .A(n11976), .B(n11977), .Z(n11969) );
  XNOR U12765 ( .A(n11971), .B(n11970), .Z(n12097) );
  XOR U12766 ( .A(n12098), .B(n12097), .Z(n12100) );
  XNOR U12767 ( .A(n12099), .B(n12100), .Z(n12106) );
  AND U12768 ( .A(o[24]), .B(\stack[1][37] ), .Z(n12104) );
  NAND U12769 ( .A(n11815), .B(n11814), .Z(n11819) );
  NAND U12770 ( .A(n11817), .B(n11816), .Z(n11818) );
  NAND U12771 ( .A(n11819), .B(n11818), .Z(n12103) );
  XOR U12772 ( .A(n12104), .B(n12103), .Z(n12105) );
  XOR U12773 ( .A(n12109), .B(n12110), .Z(n12112) );
  AND U12774 ( .A(o[25]), .B(\stack[1][36] ), .Z(n12111) );
  XOR U12775 ( .A(n12112), .B(n12111), .Z(n12116) );
  AND U12776 ( .A(o[26]), .B(\stack[1][35] ), .Z(n12115) );
  XOR U12777 ( .A(n12116), .B(n12115), .Z(n12118) );
  XOR U12778 ( .A(n12117), .B(n12118), .Z(n11963) );
  XNOR U12779 ( .A(n11964), .B(n11965), .Z(n12124) );
  AND U12780 ( .A(o[28]), .B(\stack[1][33] ), .Z(n12122) );
  NAND U12781 ( .A(n11821), .B(n11820), .Z(n11825) );
  NAND U12782 ( .A(n11823), .B(n11822), .Z(n11824) );
  NAND U12783 ( .A(n11825), .B(n11824), .Z(n12121) );
  XOR U12784 ( .A(n12122), .B(n12121), .Z(n12123) );
  XOR U12785 ( .A(n12124), .B(n12123), .Z(n11957) );
  XOR U12786 ( .A(n11956), .B(n11957), .Z(n11959) );
  XOR U12787 ( .A(n11953), .B(n11952), .Z(n12128) );
  XOR U12788 ( .A(n12127), .B(n12128), .Z(n12130) );
  AND U12789 ( .A(\stack[1][29] ), .B(o[32]), .Z(n12134) );
  NAND U12790 ( .A(n11827), .B(n11826), .Z(n11831) );
  NAND U12791 ( .A(n11829), .B(n11828), .Z(n11830) );
  NAND U12792 ( .A(n11831), .B(n11830), .Z(n12133) );
  XOR U12793 ( .A(n12134), .B(n12133), .Z(n12135) );
  XOR U12794 ( .A(n12136), .B(n12135), .Z(n11945) );
  XOR U12795 ( .A(n11944), .B(n11945), .Z(n11947) );
  AND U12796 ( .A(\stack[1][28] ), .B(o[33]), .Z(n11946) );
  XOR U12797 ( .A(n11947), .B(n11946), .Z(n12142) );
  AND U12798 ( .A(\stack[1][27] ), .B(o[34]), .Z(n12140) );
  NAND U12799 ( .A(n11833), .B(n11832), .Z(n11837) );
  NAND U12800 ( .A(n11835), .B(n11834), .Z(n11836) );
  NAND U12801 ( .A(n11837), .B(n11836), .Z(n12139) );
  XOR U12802 ( .A(n12140), .B(n12139), .Z(n12141) );
  XOR U12803 ( .A(n12142), .B(n12141), .Z(n11939) );
  XOR U12804 ( .A(n11938), .B(n11939), .Z(n11941) );
  AND U12805 ( .A(\stack[1][25] ), .B(o[36]), .Z(n12146) );
  NAND U12806 ( .A(n11839), .B(n11838), .Z(n11843) );
  NAND U12807 ( .A(n11841), .B(n11840), .Z(n11842) );
  NAND U12808 ( .A(n11843), .B(n11842), .Z(n12145) );
  XOR U12809 ( .A(n12146), .B(n12145), .Z(n12147) );
  XOR U12810 ( .A(n12148), .B(n12147), .Z(n11933) );
  XOR U12811 ( .A(n11932), .B(n11933), .Z(n11935) );
  AND U12812 ( .A(\stack[1][23] ), .B(o[38]), .Z(n12152) );
  NAND U12813 ( .A(n11845), .B(n11844), .Z(n11849) );
  NAND U12814 ( .A(n11847), .B(n11846), .Z(n11848) );
  NAND U12815 ( .A(n11849), .B(n11848), .Z(n12151) );
  XOR U12816 ( .A(n12152), .B(n12151), .Z(n12153) );
  XOR U12817 ( .A(n12154), .B(n12153), .Z(n11926) );
  XOR U12818 ( .A(n11927), .B(n11926), .Z(n11928) );
  XOR U12819 ( .A(n11929), .B(n11928), .Z(n12160) );
  AND U12820 ( .A(\stack[1][21] ), .B(o[40]), .Z(n12158) );
  NAND U12821 ( .A(n11851), .B(n11850), .Z(n11855) );
  NAND U12822 ( .A(n11853), .B(n11852), .Z(n11854) );
  NAND U12823 ( .A(n11855), .B(n11854), .Z(n12157) );
  XOR U12824 ( .A(n12158), .B(n12157), .Z(n12159) );
  XOR U12825 ( .A(n12160), .B(n12159), .Z(n12164) );
  XOR U12826 ( .A(n12163), .B(n12164), .Z(n12166) );
  AND U12827 ( .A(\stack[1][20] ), .B(o[41]), .Z(n12165) );
  XOR U12828 ( .A(n12166), .B(n12165), .Z(n12172) );
  AND U12829 ( .A(\stack[1][19] ), .B(o[42]), .Z(n12170) );
  NAND U12830 ( .A(n11857), .B(n11856), .Z(n11861) );
  NAND U12831 ( .A(n11859), .B(n11858), .Z(n11860) );
  NAND U12832 ( .A(n11861), .B(n11860), .Z(n12169) );
  XOR U12833 ( .A(n12170), .B(n12169), .Z(n12171) );
  XOR U12834 ( .A(n12172), .B(n12171), .Z(n11920) );
  XOR U12835 ( .A(n11921), .B(n11920), .Z(n11923) );
  AND U12836 ( .A(\stack[1][18] ), .B(o[43]), .Z(n11922) );
  XOR U12837 ( .A(n11923), .B(n11922), .Z(n12178) );
  AND U12838 ( .A(\stack[1][17] ), .B(o[44]), .Z(n12176) );
  NAND U12839 ( .A(n11863), .B(n11862), .Z(n11867) );
  NAND U12840 ( .A(n11865), .B(n11864), .Z(n11866) );
  NAND U12841 ( .A(n11867), .B(n11866), .Z(n12175) );
  XOR U12842 ( .A(n12176), .B(n12175), .Z(n12177) );
  XOR U12843 ( .A(n12178), .B(n12177), .Z(n12181) );
  XOR U12844 ( .A(n12182), .B(n12181), .Z(n12184) );
  AND U12845 ( .A(\stack[1][16] ), .B(o[45]), .Z(n12183) );
  XOR U12846 ( .A(n12184), .B(n12183), .Z(n12190) );
  AND U12847 ( .A(\stack[1][15] ), .B(o[46]), .Z(n12188) );
  NAND U12848 ( .A(n11869), .B(n11868), .Z(n11873) );
  NAND U12849 ( .A(n11871), .B(n11870), .Z(n11872) );
  NAND U12850 ( .A(n11873), .B(n11872), .Z(n12187) );
  XOR U12851 ( .A(n12188), .B(n12187), .Z(n12189) );
  XOR U12852 ( .A(n12190), .B(n12189), .Z(n12193) );
  XOR U12853 ( .A(n12194), .B(n12193), .Z(n12196) );
  AND U12854 ( .A(\stack[1][14] ), .B(o[47]), .Z(n12195) );
  XOR U12855 ( .A(n12196), .B(n12195), .Z(n12202) );
  AND U12856 ( .A(\stack[1][13] ), .B(o[48]), .Z(n12200) );
  NAND U12857 ( .A(n11875), .B(n11874), .Z(n11879) );
  NAND U12858 ( .A(n11877), .B(n11876), .Z(n11878) );
  NAND U12859 ( .A(n11879), .B(n11878), .Z(n12199) );
  XOR U12860 ( .A(n12200), .B(n12199), .Z(n12201) );
  XOR U12861 ( .A(n12202), .B(n12201), .Z(n11915) );
  XOR U12862 ( .A(n11914), .B(n11915), .Z(n11917) );
  AND U12863 ( .A(\stack[1][11] ), .B(o[50]), .Z(n12206) );
  NAND U12864 ( .A(n11881), .B(n11880), .Z(n11885) );
  NAND U12865 ( .A(n11883), .B(n11882), .Z(n11884) );
  NAND U12866 ( .A(n11885), .B(n11884), .Z(n12205) );
  XOR U12867 ( .A(n12206), .B(n12205), .Z(n12207) );
  XOR U12868 ( .A(n12208), .B(n12207), .Z(n11909) );
  XOR U12869 ( .A(n11908), .B(n11909), .Z(n11911) );
  AND U12870 ( .A(\stack[1][9] ), .B(o[52]), .Z(n12212) );
  NAND U12871 ( .A(n11887), .B(n11886), .Z(n11891) );
  NAND U12872 ( .A(n11889), .B(n11888), .Z(n11890) );
  NAND U12873 ( .A(n11891), .B(n11890), .Z(n12211) );
  XOR U12874 ( .A(n12212), .B(n12211), .Z(n12213) );
  XOR U12875 ( .A(n12214), .B(n12213), .Z(n11902) );
  XOR U12876 ( .A(n11903), .B(n11902), .Z(n11904) );
  XOR U12877 ( .A(n11905), .B(n11904), .Z(n12220) );
  AND U12878 ( .A(\stack[1][7] ), .B(o[54]), .Z(n12218) );
  NAND U12879 ( .A(n11893), .B(n11892), .Z(n11897) );
  NAND U12880 ( .A(n11895), .B(n11894), .Z(n11896) );
  NAND U12881 ( .A(n11897), .B(n11896), .Z(n12217) );
  XOR U12882 ( .A(n12218), .B(n12217), .Z(n12219) );
  XOR U12883 ( .A(n12220), .B(n12219), .Z(n11899) );
  NAND U12884 ( .A(n11898), .B(n11899), .Z(n11901) );
  AND U12885 ( .A(\stack[1][6] ), .B(o[55]), .Z(n12549) );
  NAND U12886 ( .A(n12549), .B(n12550), .Z(n11900) );
  NAND U12887 ( .A(n11901), .B(n11900), .Z(n12561) );
  AND U12888 ( .A(\stack[1][6] ), .B(o[56]), .Z(n12562) );
  XOR U12889 ( .A(n12561), .B(n12562), .Z(n12560) );
  NAND U12890 ( .A(n11903), .B(n11902), .Z(n11907) );
  NAND U12891 ( .A(n11905), .B(n11904), .Z(n11906) );
  NAND U12892 ( .A(n11907), .B(n11906), .Z(n13114) );
  AND U12893 ( .A(\stack[1][8] ), .B(o[54]), .Z(n13115) );
  XOR U12894 ( .A(n13114), .B(n13115), .Z(n13113) );
  NAND U12895 ( .A(n11909), .B(n11908), .Z(n11913) );
  NAND U12896 ( .A(n11911), .B(n11910), .Z(n11912) );
  NAND U12897 ( .A(n11913), .B(n11912), .Z(n12567) );
  AND U12898 ( .A(\stack[1][10] ), .B(o[52]), .Z(n12568) );
  XOR U12899 ( .A(n12567), .B(n12568), .Z(n12566) );
  NAND U12900 ( .A(n11915), .B(n11914), .Z(n11919) );
  NAND U12901 ( .A(n11917), .B(n11916), .Z(n11918) );
  NAND U12902 ( .A(n11919), .B(n11918), .Z(n13078) );
  AND U12903 ( .A(\stack[1][12] ), .B(o[50]), .Z(n13079) );
  XOR U12904 ( .A(n13078), .B(n13079), .Z(n13077) );
  NAND U12905 ( .A(n11921), .B(n11920), .Z(n11925) );
  NAND U12906 ( .A(n11923), .B(n11922), .Z(n11924) );
  NAND U12907 ( .A(n11925), .B(n11924), .Z(n12585) );
  AND U12908 ( .A(\stack[1][18] ), .B(o[44]), .Z(n12586) );
  XOR U12909 ( .A(n12585), .B(n12586), .Z(n12584) );
  NAND U12910 ( .A(n11927), .B(n11926), .Z(n11931) );
  NAND U12911 ( .A(n11929), .B(n11928), .Z(n11930) );
  NAND U12912 ( .A(n11931), .B(n11930), .Z(n12591) );
  AND U12913 ( .A(\stack[1][22] ), .B(o[40]), .Z(n12592) );
  XOR U12914 ( .A(n12591), .B(n12592), .Z(n12590) );
  NAND U12915 ( .A(n11933), .B(n11932), .Z(n11937) );
  NAND U12916 ( .A(n11935), .B(n11934), .Z(n11936) );
  NAND U12917 ( .A(n11937), .B(n11936), .Z(n12597) );
  AND U12918 ( .A(\stack[1][24] ), .B(o[38]), .Z(n12598) );
  XOR U12919 ( .A(n12597), .B(n12598), .Z(n12596) );
  NAND U12920 ( .A(n11939), .B(n11938), .Z(n11943) );
  NAND U12921 ( .A(n11941), .B(n11940), .Z(n11942) );
  NAND U12922 ( .A(n11943), .B(n11942), .Z(n13004) );
  AND U12923 ( .A(\stack[1][26] ), .B(o[36]), .Z(n13005) );
  XOR U12924 ( .A(n13004), .B(n13005), .Z(n13007) );
  NAND U12925 ( .A(n11945), .B(n11944), .Z(n11949) );
  NAND U12926 ( .A(n11947), .B(n11946), .Z(n11948) );
  NAND U12927 ( .A(n11949), .B(n11948), .Z(n12603) );
  AND U12928 ( .A(\stack[1][28] ), .B(o[34]), .Z(n12604) );
  XOR U12929 ( .A(n12603), .B(n12604), .Z(n12602) );
  AND U12930 ( .A(\stack[1][31] ), .B(o[31]), .Z(n12968) );
  NAND U12931 ( .A(n11951), .B(n11950), .Z(n11955) );
  NAND U12932 ( .A(n11953), .B(n11952), .Z(n11954) );
  NAND U12933 ( .A(n11955), .B(n11954), .Z(n12970) );
  NAND U12934 ( .A(n11957), .B(n11956), .Z(n11961) );
  NAND U12935 ( .A(n11959), .B(n11958), .Z(n11960) );
  AND U12936 ( .A(n11961), .B(n11960), .Z(n12610) );
  NAND U12937 ( .A(o[30]), .B(\stack[1][32] ), .Z(n12609) );
  XOR U12938 ( .A(n12610), .B(n12609), .Z(n12607) );
  NAND U12939 ( .A(n11963), .B(n11962), .Z(n11967) );
  NANDN U12940 ( .A(n11965), .B(n11964), .Z(n11966) );
  NAND U12941 ( .A(n11967), .B(n11966), .Z(n12615) );
  AND U12942 ( .A(o[28]), .B(\stack[1][34] ), .Z(n12616) );
  XOR U12943 ( .A(n12615), .B(n12616), .Z(n12614) );
  AND U12944 ( .A(o[26]), .B(\stack[1][36] ), .Z(n12927) );
  NAND U12945 ( .A(o[24]), .B(\stack[1][38] ), .Z(n12619) );
  NAND U12946 ( .A(n11969), .B(n11968), .Z(n11973) );
  NAND U12947 ( .A(n11971), .B(n11970), .Z(n11972) );
  NAND U12948 ( .A(n11973), .B(n11972), .Z(n12908) );
  AND U12949 ( .A(o[22]), .B(\stack[1][40] ), .Z(n12915) );
  NAND U12950 ( .A(n11975), .B(n11974), .Z(n11979) );
  NAND U12951 ( .A(n11977), .B(n11976), .Z(n11978) );
  AND U12952 ( .A(n11979), .B(n11978), .Z(n12917) );
  NAND U12953 ( .A(o[21]), .B(\stack[1][41] ), .Z(n12625) );
  NAND U12954 ( .A(n11981), .B(n11980), .Z(n11985) );
  NAND U12955 ( .A(n11983), .B(n11982), .Z(n11984) );
  NAND U12956 ( .A(n11985), .B(n11984), .Z(n12890) );
  NAND U12957 ( .A(o[19]), .B(\stack[1][43] ), .Z(n12896) );
  NAND U12958 ( .A(n11987), .B(n11986), .Z(n11991) );
  NANDN U12959 ( .A(n11989), .B(n11988), .Z(n11990) );
  NAND U12960 ( .A(n11991), .B(n11990), .Z(n12633) );
  NAND U12961 ( .A(o[17]), .B(\stack[1][45] ), .Z(n12872) );
  NAND U12962 ( .A(n11993), .B(n11992), .Z(n11997) );
  NAND U12963 ( .A(n11995), .B(n11994), .Z(n11996) );
  NAND U12964 ( .A(n11997), .B(n11996), .Z(n12637) );
  NAND U12965 ( .A(n11999), .B(n11998), .Z(n12003) );
  NAND U12966 ( .A(n12001), .B(n12000), .Z(n12002) );
  NAND U12967 ( .A(n12003), .B(n12002), .Z(n12854) );
  AND U12968 ( .A(o[13]), .B(\stack[1][49] ), .Z(n12860) );
  NAND U12969 ( .A(n12005), .B(n12004), .Z(n12009) );
  NAND U12970 ( .A(n12007), .B(n12006), .Z(n12008) );
  NAND U12971 ( .A(n12009), .B(n12008), .Z(n12862) );
  AND U12972 ( .A(o[12]), .B(\stack[1][50] ), .Z(n12644) );
  NAND U12973 ( .A(n12011), .B(n12010), .Z(n12015) );
  NAND U12974 ( .A(n12013), .B(n12012), .Z(n12014) );
  AND U12975 ( .A(n12015), .B(n12014), .Z(n12645) );
  NAND U12976 ( .A(o[11]), .B(\stack[1][51] ), .Z(n12836) );
  NAND U12977 ( .A(n12017), .B(n12016), .Z(n12021) );
  NAND U12978 ( .A(n12019), .B(n12018), .Z(n12020) );
  AND U12979 ( .A(n12021), .B(n12020), .Z(n12839) );
  NAND U12980 ( .A(n12023), .B(n12022), .Z(n12027) );
  NANDN U12981 ( .A(n12025), .B(n12024), .Z(n12026) );
  AND U12982 ( .A(n12027), .B(n12026), .Z(n12843) );
  NAND U12983 ( .A(o[9]), .B(\stack[1][53] ), .Z(n12649) );
  NAND U12984 ( .A(n12029), .B(n12028), .Z(n12033) );
  NAND U12985 ( .A(n12031), .B(n12030), .Z(n12032) );
  NAND U12986 ( .A(n12033), .B(n12032), .Z(n12818) );
  NAND U12987 ( .A(n12035), .B(n12034), .Z(n12039) );
  NAND U12988 ( .A(n12037), .B(n12036), .Z(n12038) );
  NAND U12989 ( .A(n12039), .B(n12038), .Z(n12824) );
  AND U12990 ( .A(o[6]), .B(\stack[1][56] ), .Z(n12655) );
  NAND U12991 ( .A(n12041), .B(n12040), .Z(n12045) );
  NAND U12992 ( .A(n12043), .B(n12042), .Z(n12044) );
  NAND U12993 ( .A(n12045), .B(n12044), .Z(n12657) );
  NAND U12994 ( .A(o[5]), .B(\stack[1][57] ), .Z(n12770) );
  NAND U12995 ( .A(o[4]), .B(\stack[1][58] ), .Z(n12776) );
  OR U12996 ( .A(n12046), .B(n12683), .Z(n12050) );
  NANDN U12997 ( .A(n12048), .B(n12047), .Z(n12049) );
  NAND U12998 ( .A(n12050), .B(n12049), .Z(n12663) );
  AND U12999 ( .A(\stack[1][62] ), .B(o[0]), .Z(n12054) );
  NAND U13000 ( .A(n12052), .B(n12051), .Z(n12053) );
  XNOR U13001 ( .A(n12054), .B(n12053), .Z(n12682) );
  AND U13002 ( .A(o[2]), .B(\stack[1][60] ), .Z(n12681) );
  XOR U13003 ( .A(n12682), .B(n12681), .Z(n12664) );
  XOR U13004 ( .A(n12663), .B(n12664), .Z(n12662) );
  AND U13005 ( .A(o[3]), .B(\stack[1][59] ), .Z(n12661) );
  XNOR U13006 ( .A(n12662), .B(n12661), .Z(n12779) );
  NAND U13007 ( .A(n12056), .B(n12055), .Z(n12060) );
  NAND U13008 ( .A(n12058), .B(n12057), .Z(n12059) );
  AND U13009 ( .A(n12060), .B(n12059), .Z(n12778) );
  XOR U13010 ( .A(n12776), .B(n12777), .Z(n12773) );
  NAND U13011 ( .A(n12062), .B(n12061), .Z(n12066) );
  NAND U13012 ( .A(n12064), .B(n12063), .Z(n12065) );
  AND U13013 ( .A(n12066), .B(n12065), .Z(n12772) );
  XOR U13014 ( .A(n12773), .B(n12772), .Z(n12771) );
  XNOR U13015 ( .A(n12770), .B(n12771), .Z(n12658) );
  XNOR U13016 ( .A(n12655), .B(n12656), .Z(n12827) );
  AND U13017 ( .A(o[7]), .B(\stack[1][55] ), .Z(n12826) );
  XOR U13018 ( .A(n12827), .B(n12826), .Z(n12825) );
  XOR U13019 ( .A(n12824), .B(n12825), .Z(n12821) );
  AND U13020 ( .A(o[8]), .B(\stack[1][54] ), .Z(n12820) );
  XOR U13021 ( .A(n12821), .B(n12820), .Z(n12819) );
  XNOR U13022 ( .A(n12818), .B(n12819), .Z(n12652) );
  NAND U13023 ( .A(n12068), .B(n12067), .Z(n12072) );
  NAND U13024 ( .A(n12070), .B(n12069), .Z(n12071) );
  AND U13025 ( .A(n12072), .B(n12071), .Z(n12651) );
  XNOR U13026 ( .A(n12649), .B(n12650), .Z(n12842) );
  AND U13027 ( .A(o[10]), .B(\stack[1][52] ), .Z(n12844) );
  XNOR U13028 ( .A(n12845), .B(n12844), .Z(n12838) );
  XNOR U13029 ( .A(n12836), .B(n12837), .Z(n12646) );
  XOR U13030 ( .A(n12644), .B(n12643), .Z(n12863) );
  XOR U13031 ( .A(n12862), .B(n12863), .Z(n12861) );
  AND U13032 ( .A(o[14]), .B(\stack[1][48] ), .Z(n12856) );
  XOR U13033 ( .A(n12857), .B(n12856), .Z(n12855) );
  XOR U13034 ( .A(n12854), .B(n12855), .Z(n12640) );
  AND U13035 ( .A(o[15]), .B(\stack[1][47] ), .Z(n12639) );
  XOR U13036 ( .A(n12640), .B(n12639), .Z(n12638) );
  XOR U13037 ( .A(n12637), .B(n12638), .Z(n12881) );
  AND U13038 ( .A(o[16]), .B(\stack[1][46] ), .Z(n12880) );
  XOR U13039 ( .A(n12881), .B(n12880), .Z(n12879) );
  NAND U13040 ( .A(n12074), .B(n12073), .Z(n12078) );
  NAND U13041 ( .A(n12076), .B(n12075), .Z(n12077) );
  NAND U13042 ( .A(n12078), .B(n12077), .Z(n12878) );
  XNOR U13043 ( .A(n12879), .B(n12878), .Z(n12875) );
  NAND U13044 ( .A(n12080), .B(n12079), .Z(n12084) );
  NAND U13045 ( .A(n12082), .B(n12081), .Z(n12083) );
  AND U13046 ( .A(n12084), .B(n12083), .Z(n12874) );
  XOR U13047 ( .A(n12872), .B(n12873), .Z(n12634) );
  XOR U13048 ( .A(n12633), .B(n12634), .Z(n12632) );
  NAND U13049 ( .A(o[18]), .B(\stack[1][44] ), .Z(n12631) );
  XOR U13050 ( .A(n12632), .B(n12631), .Z(n12899) );
  NAND U13051 ( .A(n12086), .B(n12085), .Z(n12090) );
  NAND U13052 ( .A(n12088), .B(n12087), .Z(n12089) );
  AND U13053 ( .A(n12090), .B(n12089), .Z(n12898) );
  XOR U13054 ( .A(n12899), .B(n12898), .Z(n12897) );
  XNOR U13055 ( .A(n12896), .B(n12897), .Z(n12893) );
  AND U13056 ( .A(o[20]), .B(\stack[1][42] ), .Z(n12892) );
  XNOR U13057 ( .A(n12890), .B(n12891), .Z(n12628) );
  NAND U13058 ( .A(n12092), .B(n12091), .Z(n12096) );
  NAND U13059 ( .A(n12094), .B(n12093), .Z(n12095) );
  AND U13060 ( .A(n12096), .B(n12095), .Z(n12627) );
  XOR U13061 ( .A(n12625), .B(n12626), .Z(n12916) );
  XOR U13062 ( .A(n12917), .B(n12916), .Z(n12914) );
  XOR U13063 ( .A(n12915), .B(n12914), .Z(n12911) );
  AND U13064 ( .A(o[23]), .B(\stack[1][39] ), .Z(n12910) );
  XOR U13065 ( .A(n12911), .B(n12910), .Z(n12909) );
  XNOR U13066 ( .A(n12908), .B(n12909), .Z(n12622) );
  NAND U13067 ( .A(n12098), .B(n12097), .Z(n12102) );
  NAND U13068 ( .A(n12100), .B(n12099), .Z(n12101) );
  NAND U13069 ( .A(n12102), .B(n12101), .Z(n12621) );
  XNOR U13070 ( .A(n12619), .B(n12620), .Z(n12933) );
  AND U13071 ( .A(o[25]), .B(\stack[1][37] ), .Z(n12935) );
  NAND U13072 ( .A(n12104), .B(n12103), .Z(n12108) );
  NAND U13073 ( .A(n12106), .B(n12105), .Z(n12107) );
  NAND U13074 ( .A(n12108), .B(n12107), .Z(n12934) );
  XOR U13075 ( .A(n12935), .B(n12934), .Z(n12932) );
  NAND U13076 ( .A(n12110), .B(n12109), .Z(n12114) );
  NAND U13077 ( .A(n12112), .B(n12111), .Z(n12113) );
  NAND U13078 ( .A(n12114), .B(n12113), .Z(n12928) );
  XOR U13079 ( .A(n12929), .B(n12928), .Z(n12926) );
  XOR U13080 ( .A(n12927), .B(n12926), .Z(n12951) );
  AND U13081 ( .A(o[27]), .B(\stack[1][35] ), .Z(n12953) );
  NAND U13082 ( .A(n12116), .B(n12115), .Z(n12120) );
  NAND U13083 ( .A(n12118), .B(n12117), .Z(n12119) );
  NAND U13084 ( .A(n12120), .B(n12119), .Z(n12952) );
  XOR U13085 ( .A(n12953), .B(n12952), .Z(n12950) );
  XOR U13086 ( .A(n12951), .B(n12950), .Z(n12613) );
  XOR U13087 ( .A(n12614), .B(n12613), .Z(n12947) );
  NAND U13088 ( .A(n12122), .B(n12121), .Z(n12126) );
  NAND U13089 ( .A(n12124), .B(n12123), .Z(n12125) );
  NAND U13090 ( .A(n12126), .B(n12125), .Z(n12946) );
  XOR U13091 ( .A(n12947), .B(n12946), .Z(n12945) );
  AND U13092 ( .A(o[29]), .B(\stack[1][33] ), .Z(n12944) );
  XNOR U13093 ( .A(n12945), .B(n12944), .Z(n12608) );
  XNOR U13094 ( .A(n12968), .B(n12969), .Z(n12962) );
  NAND U13095 ( .A(n12128), .B(n12127), .Z(n12132) );
  NAND U13096 ( .A(n12130), .B(n12129), .Z(n12131) );
  NAND U13097 ( .A(n12132), .B(n12131), .Z(n12964) );
  AND U13098 ( .A(\stack[1][30] ), .B(o[32]), .Z(n12965) );
  XOR U13099 ( .A(n12964), .B(n12965), .Z(n12963) );
  NAND U13100 ( .A(n12134), .B(n12133), .Z(n12138) );
  NAND U13101 ( .A(n12136), .B(n12135), .Z(n12137) );
  NAND U13102 ( .A(n12138), .B(n12137), .Z(n12988) );
  XOR U13103 ( .A(n12989), .B(n12988), .Z(n12987) );
  AND U13104 ( .A(\stack[1][29] ), .B(o[33]), .Z(n12986) );
  XOR U13105 ( .A(n12987), .B(n12986), .Z(n12601) );
  XOR U13106 ( .A(n12602), .B(n12601), .Z(n12983) );
  NAND U13107 ( .A(n12140), .B(n12139), .Z(n12144) );
  NAND U13108 ( .A(n12142), .B(n12141), .Z(n12143) );
  NAND U13109 ( .A(n12144), .B(n12143), .Z(n12982) );
  XOR U13110 ( .A(n12983), .B(n12982), .Z(n12981) );
  AND U13111 ( .A(\stack[1][27] ), .B(o[35]), .Z(n12980) );
  XOR U13112 ( .A(n12981), .B(n12980), .Z(n13006) );
  XOR U13113 ( .A(n13007), .B(n13006), .Z(n13001) );
  NAND U13114 ( .A(n12146), .B(n12145), .Z(n12150) );
  NAND U13115 ( .A(n12148), .B(n12147), .Z(n12149) );
  NAND U13116 ( .A(n12150), .B(n12149), .Z(n13000) );
  XOR U13117 ( .A(n13001), .B(n13000), .Z(n12999) );
  AND U13118 ( .A(\stack[1][25] ), .B(o[37]), .Z(n12998) );
  XOR U13119 ( .A(n12999), .B(n12998), .Z(n12595) );
  XOR U13120 ( .A(n12596), .B(n12595), .Z(n13025) );
  NAND U13121 ( .A(n12152), .B(n12151), .Z(n12156) );
  NAND U13122 ( .A(n12154), .B(n12153), .Z(n12155) );
  NAND U13123 ( .A(n12156), .B(n12155), .Z(n13024) );
  XOR U13124 ( .A(n13025), .B(n13024), .Z(n13023) );
  AND U13125 ( .A(\stack[1][23] ), .B(o[39]), .Z(n13022) );
  XOR U13126 ( .A(n13023), .B(n13022), .Z(n12589) );
  XOR U13127 ( .A(n12590), .B(n12589), .Z(n13019) );
  NAND U13128 ( .A(n12158), .B(n12157), .Z(n12162) );
  NAND U13129 ( .A(n12160), .B(n12159), .Z(n12161) );
  NAND U13130 ( .A(n12162), .B(n12161), .Z(n13018) );
  XOR U13131 ( .A(n13019), .B(n13018), .Z(n13017) );
  AND U13132 ( .A(\stack[1][21] ), .B(o[41]), .Z(n13016) );
  XOR U13133 ( .A(n13017), .B(n13016), .Z(n13041) );
  AND U13134 ( .A(\stack[1][20] ), .B(o[42]), .Z(n13043) );
  NAND U13135 ( .A(n12164), .B(n12163), .Z(n12168) );
  NAND U13136 ( .A(n12166), .B(n12165), .Z(n12167) );
  NAND U13137 ( .A(n12168), .B(n12167), .Z(n13042) );
  XOR U13138 ( .A(n13043), .B(n13042), .Z(n13040) );
  XOR U13139 ( .A(n13041), .B(n13040), .Z(n13037) );
  NAND U13140 ( .A(n12170), .B(n12169), .Z(n12174) );
  NAND U13141 ( .A(n12172), .B(n12171), .Z(n12173) );
  NAND U13142 ( .A(n12174), .B(n12173), .Z(n13036) );
  XOR U13143 ( .A(n13037), .B(n13036), .Z(n13035) );
  AND U13144 ( .A(\stack[1][19] ), .B(o[43]), .Z(n13034) );
  XOR U13145 ( .A(n13035), .B(n13034), .Z(n12583) );
  XOR U13146 ( .A(n12584), .B(n12583), .Z(n12580) );
  NAND U13147 ( .A(n12176), .B(n12175), .Z(n12180) );
  NAND U13148 ( .A(n12178), .B(n12177), .Z(n12179) );
  NAND U13149 ( .A(n12180), .B(n12179), .Z(n12579) );
  XOR U13150 ( .A(n12580), .B(n12579), .Z(n12578) );
  AND U13151 ( .A(\stack[1][17] ), .B(o[45]), .Z(n12577) );
  XOR U13152 ( .A(n12578), .B(n12577), .Z(n13058) );
  NAND U13153 ( .A(n12182), .B(n12181), .Z(n12186) );
  NAND U13154 ( .A(n12184), .B(n12183), .Z(n12185) );
  NAND U13155 ( .A(n12186), .B(n12185), .Z(n13060) );
  AND U13156 ( .A(\stack[1][16] ), .B(o[46]), .Z(n13061) );
  XOR U13157 ( .A(n13060), .B(n13061), .Z(n13059) );
  NAND U13158 ( .A(n12188), .B(n12187), .Z(n12192) );
  NAND U13159 ( .A(n12190), .B(n12189), .Z(n12191) );
  NAND U13160 ( .A(n12192), .B(n12191), .Z(n13054) );
  XOR U13161 ( .A(n13055), .B(n13054), .Z(n13053) );
  AND U13162 ( .A(\stack[1][15] ), .B(o[47]), .Z(n13052) );
  XOR U13163 ( .A(n13053), .B(n13052), .Z(n12571) );
  NAND U13164 ( .A(n12194), .B(n12193), .Z(n12198) );
  NAND U13165 ( .A(n12196), .B(n12195), .Z(n12197) );
  NAND U13166 ( .A(n12198), .B(n12197), .Z(n12573) );
  AND U13167 ( .A(\stack[1][14] ), .B(o[48]), .Z(n12574) );
  XOR U13168 ( .A(n12573), .B(n12574), .Z(n12572) );
  NAND U13169 ( .A(n12200), .B(n12199), .Z(n12204) );
  NAND U13170 ( .A(n12202), .B(n12201), .Z(n12203) );
  NAND U13171 ( .A(n12204), .B(n12203), .Z(n13072) );
  XOR U13172 ( .A(n13073), .B(n13072), .Z(n13071) );
  AND U13173 ( .A(\stack[1][13] ), .B(o[49]), .Z(n13070) );
  XOR U13174 ( .A(n13071), .B(n13070), .Z(n13076) );
  XOR U13175 ( .A(n13077), .B(n13076), .Z(n13097) );
  NAND U13176 ( .A(n12206), .B(n12205), .Z(n12210) );
  NAND U13177 ( .A(n12208), .B(n12207), .Z(n12209) );
  NAND U13178 ( .A(n12210), .B(n12209), .Z(n13096) );
  XOR U13179 ( .A(n13097), .B(n13096), .Z(n13095) );
  AND U13180 ( .A(\stack[1][11] ), .B(o[51]), .Z(n13094) );
  XOR U13181 ( .A(n13095), .B(n13094), .Z(n12565) );
  XOR U13182 ( .A(n12566), .B(n12565), .Z(n13091) );
  NAND U13183 ( .A(n12212), .B(n12211), .Z(n12216) );
  NAND U13184 ( .A(n12214), .B(n12213), .Z(n12215) );
  NAND U13185 ( .A(n12216), .B(n12215), .Z(n13090) );
  XOR U13186 ( .A(n13091), .B(n13090), .Z(n13089) );
  AND U13187 ( .A(\stack[1][9] ), .B(o[53]), .Z(n13088) );
  XOR U13188 ( .A(n13089), .B(n13088), .Z(n13112) );
  XOR U13189 ( .A(n13113), .B(n13112), .Z(n13109) );
  NAND U13190 ( .A(n12218), .B(n12217), .Z(n12222) );
  NAND U13191 ( .A(n12220), .B(n12219), .Z(n12221) );
  NAND U13192 ( .A(n12222), .B(n12221), .Z(n13108) );
  XOR U13193 ( .A(n13109), .B(n13108), .Z(n13107) );
  AND U13194 ( .A(\stack[1][7] ), .B(o[55]), .Z(n13106) );
  XOR U13195 ( .A(n13107), .B(n13106), .Z(n12559) );
  XOR U13196 ( .A(n12560), .B(n12559), .Z(n12555) );
  XNOR U13197 ( .A(n12226), .B(n12225), .Z(n12414) );
  XNOR U13198 ( .A(n12228), .B(n12227), .Z(n12356) );
  XNOR U13199 ( .A(n12232), .B(n12231), .Z(n12288) );
  AND U13200 ( .A(o[0]), .B(\stack[1][5] ), .Z(n12233) );
  AND U13201 ( .A(o[1]), .B(\stack[1][6] ), .Z(n12238) );
  AND U13202 ( .A(n12233), .B(n12238), .Z(n12234) );
  NAND U13203 ( .A(n12234), .B(o[2]), .Z(n12240) );
  NAND U13204 ( .A(n12238), .B(o[0]), .Z(n12235) );
  XNOR U13205 ( .A(o[2]), .B(n12235), .Z(n12236) );
  AND U13206 ( .A(\stack[1][5] ), .B(n12236), .Z(n13140) );
  NAND U13207 ( .A(\stack[1][7] ), .B(o[0]), .Z(n12237) );
  XNOR U13208 ( .A(n12238), .B(n12237), .Z(n13141) );
  NAND U13209 ( .A(n13140), .B(n13141), .Z(n12239) );
  NAND U13210 ( .A(n12240), .B(n12239), .Z(n12243) );
  NAND U13211 ( .A(n12243), .B(n12244), .Z(n12246) );
  AND U13212 ( .A(\stack[1][5] ), .B(o[3]), .Z(n13146) );
  NAND U13213 ( .A(n13146), .B(n13147), .Z(n12245) );
  NAND U13214 ( .A(n12246), .B(n12245), .Z(n12247) );
  AND U13215 ( .A(\stack[1][5] ), .B(o[4]), .Z(n12248) );
  NAND U13216 ( .A(n12247), .B(n12248), .Z(n12252) );
  NAND U13217 ( .A(n13131), .B(n13130), .Z(n12251) );
  NAND U13218 ( .A(n12252), .B(n12251), .Z(n12255) );
  XOR U13219 ( .A(n12254), .B(n12253), .Z(n12256) );
  NAND U13220 ( .A(n12255), .B(n12256), .Z(n12258) );
  AND U13221 ( .A(\stack[1][5] ), .B(o[5]), .Z(n17136) );
  NAND U13222 ( .A(n17136), .B(n13155), .Z(n12257) );
  NAND U13223 ( .A(n12258), .B(n12257), .Z(n12261) );
  NAND U13224 ( .A(n12261), .B(n12262), .Z(n12264) );
  AND U13225 ( .A(\stack[1][5] ), .B(o[6]), .Z(n13161) );
  NAND U13226 ( .A(n13161), .B(n13160), .Z(n12263) );
  NAND U13227 ( .A(n12264), .B(n12263), .Z(n12266) );
  XOR U13228 ( .A(n17097), .B(n12265), .Z(n12267) );
  NAND U13229 ( .A(n12266), .B(n12267), .Z(n12269) );
  AND U13230 ( .A(\stack[1][5] ), .B(o[7]), .Z(n13166) );
  NAND U13231 ( .A(n13166), .B(n13167), .Z(n12268) );
  NAND U13232 ( .A(n12269), .B(n12268), .Z(n12272) );
  AND U13233 ( .A(\stack[1][5] ), .B(o[8]), .Z(n12273) );
  NAND U13234 ( .A(n12272), .B(n12273), .Z(n12275) );
  NAND U13235 ( .A(n13129), .B(n13128), .Z(n12274) );
  NAND U13236 ( .A(n12275), .B(n12274), .Z(n12278) );
  XOR U13237 ( .A(n12277), .B(n12276), .Z(n12279) );
  NAND U13238 ( .A(n12278), .B(n12279), .Z(n12281) );
  AND U13239 ( .A(\stack[1][5] ), .B(o[9]), .Z(n13176) );
  NAND U13240 ( .A(n13176), .B(n13177), .Z(n12280) );
  NAND U13241 ( .A(n12281), .B(n12280), .Z(n12284) );
  AND U13242 ( .A(o[10]), .B(\stack[1][5] ), .Z(n12285) );
  NAND U13243 ( .A(n12284), .B(n12285), .Z(n12287) );
  XNOR U13244 ( .A(n12283), .B(n12282), .Z(n13182) );
  NAND U13245 ( .A(n13182), .B(n13183), .Z(n12286) );
  AND U13246 ( .A(n12287), .B(n12286), .Z(n12289) );
  NAND U13247 ( .A(n12288), .B(n12289), .Z(n12291) );
  NAND U13248 ( .A(\stack[1][5] ), .B(o[11]), .Z(n13188) );
  NAND U13249 ( .A(n13189), .B(n13188), .Z(n12290) );
  AND U13250 ( .A(n12291), .B(n12290), .Z(n12294) );
  AND U13251 ( .A(\stack[1][5] ), .B(o[12]), .Z(n12295) );
  NAND U13252 ( .A(n12294), .B(n12295), .Z(n12297) );
  NAND U13253 ( .A(n13127), .B(n13126), .Z(n12296) );
  NAND U13254 ( .A(n12297), .B(n12296), .Z(n12300) );
  XNOR U13255 ( .A(n12299), .B(n12298), .Z(n12301) );
  NAND U13256 ( .A(n12300), .B(n12301), .Z(n12303) );
  AND U13257 ( .A(\stack[1][5] ), .B(o[13]), .Z(n13200) );
  NAND U13258 ( .A(n13201), .B(n13200), .Z(n12302) );
  NAND U13259 ( .A(n12303), .B(n12302), .Z(n12306) );
  AND U13260 ( .A(\stack[1][5] ), .B(o[14]), .Z(n12307) );
  NAND U13261 ( .A(n12306), .B(n12307), .Z(n12309) );
  XOR U13262 ( .A(n12305), .B(n12304), .Z(n13205) );
  NAND U13263 ( .A(n13205), .B(n13204), .Z(n12308) );
  NAND U13264 ( .A(n12309), .B(n12308), .Z(n12312) );
  XOR U13265 ( .A(n12311), .B(n12310), .Z(n12313) );
  NAND U13266 ( .A(n12312), .B(n12313), .Z(n12315) );
  AND U13267 ( .A(\stack[1][5] ), .B(o[15]), .Z(n13212) );
  NAND U13268 ( .A(n13212), .B(n13213), .Z(n12314) );
  NAND U13269 ( .A(n12315), .B(n12314), .Z(n12318) );
  AND U13270 ( .A(\stack[1][5] ), .B(o[16]), .Z(n12319) );
  NAND U13271 ( .A(n12318), .B(n12319), .Z(n12321) );
  XOR U13272 ( .A(n12317), .B(n12316), .Z(n13217) );
  NAND U13273 ( .A(n13217), .B(n13216), .Z(n12320) );
  NAND U13274 ( .A(n12321), .B(n12320), .Z(n12322) );
  NAND U13275 ( .A(n12323), .B(n12322), .Z(n12325) );
  XOR U13276 ( .A(n12323), .B(n12322), .Z(n13223) );
  AND U13277 ( .A(\stack[1][5] ), .B(o[17]), .Z(n13222) );
  NAND U13278 ( .A(n13223), .B(n13222), .Z(n12324) );
  NAND U13279 ( .A(n12325), .B(n12324), .Z(n12328) );
  AND U13280 ( .A(\stack[1][5] ), .B(o[18]), .Z(n12329) );
  NAND U13281 ( .A(n12328), .B(n12329), .Z(n12331) );
  NAND U13282 ( .A(n13229), .B(n13228), .Z(n12330) );
  NAND U13283 ( .A(n12331), .B(n12330), .Z(n12334) );
  XOR U13284 ( .A(n12333), .B(n12332), .Z(n12335) );
  NAND U13285 ( .A(n12334), .B(n12335), .Z(n12337) );
  AND U13286 ( .A(\stack[1][5] ), .B(o[19]), .Z(n13236) );
  NAND U13287 ( .A(n13236), .B(n13237), .Z(n12336) );
  NAND U13288 ( .A(n12337), .B(n12336), .Z(n12340) );
  AND U13289 ( .A(\stack[1][5] ), .B(o[20]), .Z(n12341) );
  NAND U13290 ( .A(n12340), .B(n12341), .Z(n12343) );
  NAND U13291 ( .A(n13241), .B(n13240), .Z(n12342) );
  NAND U13292 ( .A(n12343), .B(n12342), .Z(n12346) );
  XOR U13293 ( .A(n12345), .B(n12344), .Z(n12347) );
  NAND U13294 ( .A(n12346), .B(n12347), .Z(n12349) );
  AND U13295 ( .A(\stack[1][5] ), .B(o[21]), .Z(n13246) );
  NAND U13296 ( .A(n13247), .B(n13246), .Z(n12348) );
  NAND U13297 ( .A(n12349), .B(n12348), .Z(n12352) );
  AND U13298 ( .A(\stack[1][5] ), .B(o[22]), .Z(n12353) );
  NAND U13299 ( .A(n12352), .B(n12353), .Z(n12355) );
  XOR U13300 ( .A(n12351), .B(n12350), .Z(n13253) );
  NAND U13301 ( .A(n13253), .B(n13252), .Z(n12354) );
  NAND U13302 ( .A(n12355), .B(n12354), .Z(n12357) );
  NAND U13303 ( .A(n12356), .B(n12357), .Z(n12359) );
  AND U13304 ( .A(\stack[1][5] ), .B(o[23]), .Z(n13260) );
  NAND U13305 ( .A(n13260), .B(n13261), .Z(n12358) );
  NAND U13306 ( .A(n12359), .B(n12358), .Z(n12362) );
  AND U13307 ( .A(\stack[1][5] ), .B(o[24]), .Z(n12363) );
  NAND U13308 ( .A(n12362), .B(n12363), .Z(n12365) );
  NAND U13309 ( .A(n13265), .B(n13264), .Z(n12364) );
  NAND U13310 ( .A(n12365), .B(n12364), .Z(n12368) );
  XOR U13311 ( .A(n12367), .B(n12366), .Z(n12369) );
  NAND U13312 ( .A(n12368), .B(n12369), .Z(n12371) );
  AND U13313 ( .A(\stack[1][5] ), .B(o[25]), .Z(n13272) );
  NAND U13314 ( .A(n13272), .B(n13273), .Z(n12370) );
  NAND U13315 ( .A(n12371), .B(n12370), .Z(n12374) );
  AND U13316 ( .A(\stack[1][5] ), .B(o[26]), .Z(n12375) );
  NAND U13317 ( .A(n12374), .B(n12375), .Z(n12377) );
  NAND U13318 ( .A(n13277), .B(n13276), .Z(n12376) );
  NAND U13319 ( .A(n12377), .B(n12376), .Z(n12380) );
  XOR U13320 ( .A(n12379), .B(n12378), .Z(n12381) );
  NAND U13321 ( .A(n12380), .B(n12381), .Z(n12383) );
  AND U13322 ( .A(\stack[1][5] ), .B(o[27]), .Z(n13284) );
  NAND U13323 ( .A(n13285), .B(n13284), .Z(n12382) );
  NAND U13324 ( .A(n12383), .B(n12382), .Z(n12386) );
  AND U13325 ( .A(\stack[1][5] ), .B(o[28]), .Z(n12387) );
  NAND U13326 ( .A(n12386), .B(n12387), .Z(n12389) );
  NAND U13327 ( .A(n13289), .B(n13288), .Z(n12388) );
  NAND U13328 ( .A(n12389), .B(n12388), .Z(n12392) );
  XOR U13329 ( .A(n12391), .B(n12390), .Z(n12393) );
  NAND U13330 ( .A(n12392), .B(n12393), .Z(n12395) );
  AND U13331 ( .A(\stack[1][5] ), .B(o[29]), .Z(n13294) );
  NAND U13332 ( .A(n13294), .B(n13295), .Z(n12394) );
  NAND U13333 ( .A(n12395), .B(n12394), .Z(n12398) );
  AND U13334 ( .A(\stack[1][5] ), .B(o[30]), .Z(n12399) );
  NAND U13335 ( .A(n12398), .B(n12399), .Z(n12401) );
  XOR U13336 ( .A(n12397), .B(n12396), .Z(n13301) );
  NAND U13337 ( .A(n13301), .B(n13300), .Z(n12400) );
  NAND U13338 ( .A(n12401), .B(n12400), .Z(n12404) );
  XOR U13339 ( .A(n12403), .B(n12402), .Z(n12405) );
  NAND U13340 ( .A(n12404), .B(n12405), .Z(n12407) );
  AND U13341 ( .A(\stack[1][5] ), .B(o[31]), .Z(n13308) );
  NAND U13342 ( .A(n13308), .B(n13309), .Z(n12406) );
  NAND U13343 ( .A(n12407), .B(n12406), .Z(n12410) );
  AND U13344 ( .A(\stack[1][5] ), .B(o[32]), .Z(n12411) );
  NAND U13345 ( .A(n12410), .B(n12411), .Z(n12413) );
  NAND U13346 ( .A(n13313), .B(n13312), .Z(n12412) );
  NAND U13347 ( .A(n12413), .B(n12412), .Z(n12415) );
  NAND U13348 ( .A(n12414), .B(n12415), .Z(n12417) );
  AND U13349 ( .A(\stack[1][5] ), .B(o[33]), .Z(n13320) );
  NAND U13350 ( .A(n13320), .B(n13321), .Z(n12416) );
  NAND U13351 ( .A(n12417), .B(n12416), .Z(n12420) );
  AND U13352 ( .A(\stack[1][5] ), .B(o[34]), .Z(n12421) );
  NAND U13353 ( .A(n12420), .B(n12421), .Z(n12423) );
  NAND U13354 ( .A(n13325), .B(n13324), .Z(n12422) );
  NAND U13355 ( .A(n12423), .B(n12422), .Z(n12426) );
  XOR U13356 ( .A(n12425), .B(n12424), .Z(n12427) );
  NAND U13357 ( .A(n12426), .B(n12427), .Z(n12429) );
  AND U13358 ( .A(\stack[1][5] ), .B(o[35]), .Z(n13332) );
  NAND U13359 ( .A(n13332), .B(n13333), .Z(n12428) );
  NAND U13360 ( .A(n12429), .B(n12428), .Z(n12432) );
  AND U13361 ( .A(\stack[1][5] ), .B(o[36]), .Z(n12433) );
  NAND U13362 ( .A(n12432), .B(n12433), .Z(n12435) );
  XOR U13363 ( .A(n12431), .B(n12430), .Z(n13337) );
  NAND U13364 ( .A(n13337), .B(n13336), .Z(n12434) );
  NAND U13365 ( .A(n12435), .B(n12434), .Z(n12438) );
  XOR U13366 ( .A(n12437), .B(n12436), .Z(n12439) );
  NAND U13367 ( .A(n12438), .B(n12439), .Z(n12441) );
  AND U13368 ( .A(\stack[1][5] ), .B(o[37]), .Z(n13344) );
  NAND U13369 ( .A(n13345), .B(n13344), .Z(n12440) );
  NAND U13370 ( .A(n12441), .B(n12440), .Z(n12444) );
  AND U13371 ( .A(\stack[1][5] ), .B(o[38]), .Z(n12445) );
  NAND U13372 ( .A(n12444), .B(n12445), .Z(n12447) );
  XOR U13373 ( .A(n12443), .B(n12442), .Z(n13349) );
  NAND U13374 ( .A(n13349), .B(n13348), .Z(n12446) );
  NAND U13375 ( .A(n12447), .B(n12446), .Z(n12450) );
  XNOR U13376 ( .A(n12449), .B(n12448), .Z(n12451) );
  NAND U13377 ( .A(n12450), .B(n12451), .Z(n12453) );
  AND U13378 ( .A(\stack[1][5] ), .B(o[39]), .Z(n13356) );
  NAND U13379 ( .A(n13356), .B(n13357), .Z(n12452) );
  NAND U13380 ( .A(n12453), .B(n12452), .Z(n12456) );
  AND U13381 ( .A(\stack[1][5] ), .B(o[40]), .Z(n12457) );
  NAND U13382 ( .A(n12456), .B(n12457), .Z(n12459) );
  NAND U13383 ( .A(n13361), .B(n13360), .Z(n12458) );
  NAND U13384 ( .A(n12459), .B(n12458), .Z(n12462) );
  XOR U13385 ( .A(n12461), .B(n12460), .Z(n12463) );
  NAND U13386 ( .A(n12462), .B(n12463), .Z(n12465) );
  AND U13387 ( .A(\stack[1][5] ), .B(o[41]), .Z(n13368) );
  NAND U13388 ( .A(n13368), .B(n13369), .Z(n12464) );
  NAND U13389 ( .A(n12465), .B(n12464), .Z(n12468) );
  AND U13390 ( .A(\stack[1][5] ), .B(o[42]), .Z(n12469) );
  NAND U13391 ( .A(n12468), .B(n12469), .Z(n12471) );
  NAND U13392 ( .A(n13373), .B(n13372), .Z(n12470) );
  NAND U13393 ( .A(n12471), .B(n12470), .Z(n12474) );
  XOR U13394 ( .A(n12473), .B(n12472), .Z(n12475) );
  NAND U13395 ( .A(n12474), .B(n12475), .Z(n12477) );
  AND U13396 ( .A(\stack[1][5] ), .B(o[43]), .Z(n13380) );
  NAND U13397 ( .A(n13381), .B(n13380), .Z(n12476) );
  NAND U13398 ( .A(n12477), .B(n12476), .Z(n12480) );
  AND U13399 ( .A(\stack[1][5] ), .B(o[44]), .Z(n12481) );
  NAND U13400 ( .A(n12480), .B(n12481), .Z(n12483) );
  XOR U13401 ( .A(n12479), .B(n12478), .Z(n13385) );
  NAND U13402 ( .A(n13385), .B(n13384), .Z(n12482) );
  NAND U13403 ( .A(n12483), .B(n12482), .Z(n12484) );
  NAND U13404 ( .A(n12485), .B(n12484), .Z(n12487) );
  AND U13405 ( .A(\stack[1][5] ), .B(o[45]), .Z(n13392) );
  XOR U13406 ( .A(n12485), .B(n12484), .Z(n13393) );
  NAND U13407 ( .A(n13392), .B(n13393), .Z(n12486) );
  NAND U13408 ( .A(n12487), .B(n12486), .Z(n12490) );
  AND U13409 ( .A(\stack[1][5] ), .B(o[46]), .Z(n12491) );
  NAND U13410 ( .A(n12490), .B(n12491), .Z(n12493) );
  NAND U13411 ( .A(n13397), .B(n13396), .Z(n12492) );
  NAND U13412 ( .A(n12493), .B(n12492), .Z(n12496) );
  XNOR U13413 ( .A(n12495), .B(n12494), .Z(n12497) );
  NAND U13414 ( .A(n12496), .B(n12497), .Z(n12499) );
  AND U13415 ( .A(\stack[1][5] ), .B(o[47]), .Z(n13402) );
  NAND U13416 ( .A(n13403), .B(n13402), .Z(n12498) );
  NAND U13417 ( .A(n12499), .B(n12498), .Z(n12502) );
  AND U13418 ( .A(\stack[1][5] ), .B(o[48]), .Z(n12503) );
  NAND U13419 ( .A(n12502), .B(n12503), .Z(n12505) );
  XOR U13420 ( .A(n12501), .B(n12500), .Z(n13409) );
  NAND U13421 ( .A(n13409), .B(n13408), .Z(n12504) );
  NAND U13422 ( .A(n12505), .B(n12504), .Z(n12508) );
  XOR U13423 ( .A(n12507), .B(n12506), .Z(n12509) );
  NAND U13424 ( .A(n12508), .B(n12509), .Z(n12511) );
  AND U13425 ( .A(\stack[1][5] ), .B(o[49]), .Z(n13416) );
  NAND U13426 ( .A(n13416), .B(n13418), .Z(n12510) );
  NAND U13427 ( .A(n12511), .B(n12510), .Z(n12514) );
  AND U13428 ( .A(\stack[1][5] ), .B(o[50]), .Z(n12515) );
  NAND U13429 ( .A(n12514), .B(n12515), .Z(n12517) );
  XOR U13430 ( .A(n12513), .B(n12512), .Z(n13422) );
  NAND U13431 ( .A(n13422), .B(n13421), .Z(n12516) );
  NAND U13432 ( .A(n12517), .B(n12516), .Z(n12520) );
  XNOR U13433 ( .A(n12519), .B(n12518), .Z(n12521) );
  NAND U13434 ( .A(n12520), .B(n12521), .Z(n12523) );
  AND U13435 ( .A(\stack[1][5] ), .B(o[51]), .Z(n13430) );
  NAND U13436 ( .A(n13431), .B(n13430), .Z(n12522) );
  NAND U13437 ( .A(n12523), .B(n12522), .Z(n12526) );
  AND U13438 ( .A(\stack[1][5] ), .B(o[52]), .Z(n12528) );
  NAND U13439 ( .A(n12526), .B(n12528), .Z(n12530) );
  XOR U13440 ( .A(n12525), .B(n12524), .Z(n13435) );
  IV U13441 ( .A(n12526), .Z(n12527) );
  XNOR U13442 ( .A(n12528), .B(n12527), .Z(n13434) );
  NAND U13443 ( .A(n13435), .B(n13434), .Z(n12529) );
  NAND U13444 ( .A(n12530), .B(n12529), .Z(n12533) );
  XOR U13445 ( .A(n12532), .B(n12531), .Z(n12534) );
  NAND U13446 ( .A(n12533), .B(n12534), .Z(n12536) );
  AND U13447 ( .A(\stack[1][5] ), .B(o[53]), .Z(n13443) );
  NAND U13448 ( .A(n13443), .B(n13445), .Z(n12535) );
  NAND U13449 ( .A(n12536), .B(n12535), .Z(n12539) );
  AND U13450 ( .A(\stack[1][5] ), .B(o[54]), .Z(n12540) );
  NAND U13451 ( .A(n12539), .B(n12540), .Z(n12542) );
  NAND U13452 ( .A(n13449), .B(n13448), .Z(n12541) );
  NAND U13453 ( .A(n12542), .B(n12541), .Z(n12545) );
  XOR U13454 ( .A(n12544), .B(n12543), .Z(n12546) );
  NAND U13455 ( .A(n12545), .B(n12546), .Z(n12548) );
  AND U13456 ( .A(\stack[1][5] ), .B(o[55]), .Z(n13456) );
  NAND U13457 ( .A(n13456), .B(n13458), .Z(n12547) );
  NAND U13458 ( .A(n12548), .B(n12547), .Z(n12551) );
  AND U13459 ( .A(\stack[1][5] ), .B(o[56]), .Z(n12552) );
  NAND U13460 ( .A(n12551), .B(n12552), .Z(n12554) );
  NAND U13461 ( .A(n13462), .B(n13461), .Z(n12553) );
  NAND U13462 ( .A(n12554), .B(n12553), .Z(n12556) );
  NAND U13463 ( .A(n13124), .B(n13125), .Z(n12558) );
  NAND U13464 ( .A(n12556), .B(n12555), .Z(n12557) );
  AND U13465 ( .A(n12558), .B(n12557), .Z(n14909) );
  NAND U13466 ( .A(n12560), .B(n12559), .Z(n12564) );
  NAND U13467 ( .A(n12562), .B(n12561), .Z(n12563) );
  AND U13468 ( .A(n12564), .B(n12563), .Z(n13825) );
  NAND U13469 ( .A(n12566), .B(n12565), .Z(n12570) );
  NAND U13470 ( .A(n12568), .B(n12567), .Z(n12569) );
  AND U13471 ( .A(n12570), .B(n12569), .Z(n13123) );
  NAND U13472 ( .A(n12572), .B(n12571), .Z(n12576) );
  NAND U13473 ( .A(n12574), .B(n12573), .Z(n12575) );
  AND U13474 ( .A(n12576), .B(n12575), .Z(n13105) );
  NAND U13475 ( .A(n12578), .B(n12577), .Z(n12582) );
  NAND U13476 ( .A(n12580), .B(n12579), .Z(n12581) );
  AND U13477 ( .A(n12582), .B(n12581), .Z(n13087) );
  NAND U13478 ( .A(n12584), .B(n12583), .Z(n12588) );
  NAND U13479 ( .A(n12586), .B(n12585), .Z(n12587) );
  AND U13480 ( .A(n12588), .B(n12587), .Z(n13069) );
  NAND U13481 ( .A(n12590), .B(n12589), .Z(n12594) );
  NAND U13482 ( .A(n12592), .B(n12591), .Z(n12593) );
  AND U13483 ( .A(n12594), .B(n12593), .Z(n13051) );
  NAND U13484 ( .A(n12596), .B(n12595), .Z(n12600) );
  NAND U13485 ( .A(n12598), .B(n12597), .Z(n12599) );
  AND U13486 ( .A(n12600), .B(n12599), .Z(n13033) );
  NAND U13487 ( .A(n12602), .B(n12601), .Z(n12606) );
  NAND U13488 ( .A(n12604), .B(n12603), .Z(n12605) );
  AND U13489 ( .A(n12606), .B(n12605), .Z(n13015) );
  NAND U13490 ( .A(n12608), .B(n12607), .Z(n12612) );
  NAND U13491 ( .A(n12610), .B(n12609), .Z(n12611) );
  AND U13492 ( .A(n12612), .B(n12611), .Z(n12997) );
  NAND U13493 ( .A(n12614), .B(n12613), .Z(n12618) );
  NAND U13494 ( .A(n12616), .B(n12615), .Z(n12617) );
  AND U13495 ( .A(n12618), .B(n12617), .Z(n12979) );
  NAND U13496 ( .A(n12620), .B(n12619), .Z(n12624) );
  NAND U13497 ( .A(n12622), .B(n12621), .Z(n12623) );
  AND U13498 ( .A(n12624), .B(n12623), .Z(n12961) );
  NANDN U13499 ( .A(n12626), .B(n12625), .Z(n12630) );
  NAND U13500 ( .A(n12628), .B(n12627), .Z(n12629) );
  AND U13501 ( .A(n12630), .B(n12629), .Z(n12943) );
  NAND U13502 ( .A(n12632), .B(n12631), .Z(n12636) );
  NAND U13503 ( .A(n12634), .B(n12633), .Z(n12635) );
  AND U13504 ( .A(n12636), .B(n12635), .Z(n12925) );
  NAND U13505 ( .A(n12638), .B(n12637), .Z(n12642) );
  NAND U13506 ( .A(n12640), .B(n12639), .Z(n12641) );
  AND U13507 ( .A(n12642), .B(n12641), .Z(n12907) );
  NAND U13508 ( .A(n12644), .B(n12643), .Z(n12648) );
  NAND U13509 ( .A(n12646), .B(n12645), .Z(n12647) );
  AND U13510 ( .A(n12648), .B(n12647), .Z(n12889) );
  NAND U13511 ( .A(n12650), .B(n12649), .Z(n12654) );
  NAND U13512 ( .A(n12652), .B(n12651), .Z(n12653) );
  AND U13513 ( .A(n12654), .B(n12653), .Z(n12871) );
  NANDN U13514 ( .A(n12656), .B(n12655), .Z(n12660) );
  NAND U13515 ( .A(n12658), .B(n12657), .Z(n12659) );
  AND U13516 ( .A(n12660), .B(n12659), .Z(n12853) );
  NAND U13517 ( .A(n12662), .B(n12661), .Z(n12666) );
  NAND U13518 ( .A(n12664), .B(n12663), .Z(n12665) );
  AND U13519 ( .A(n12666), .B(n12665), .Z(n12835) );
  AND U13520 ( .A(o[45]), .B(\stack[1][18] ), .Z(n12668) );
  NAND U13521 ( .A(o[46]), .B(\stack[1][17] ), .Z(n12667) );
  XNOR U13522 ( .A(n12668), .B(n12667), .Z(n12672) );
  AND U13523 ( .A(o[41]), .B(\stack[1][22] ), .Z(n12670) );
  NAND U13524 ( .A(o[42]), .B(\stack[1][21] ), .Z(n12669) );
  XNOR U13525 ( .A(n12670), .B(n12669), .Z(n12671) );
  XOR U13526 ( .A(n12672), .B(n12671), .Z(n12680) );
  AND U13527 ( .A(o[47]), .B(\stack[1][16] ), .Z(n12674) );
  NAND U13528 ( .A(o[53]), .B(\stack[1][10] ), .Z(n12673) );
  XNOR U13529 ( .A(n12674), .B(n12673), .Z(n12678) );
  AND U13530 ( .A(o[54]), .B(\stack[1][9] ), .Z(n12676) );
  NAND U13531 ( .A(o[58]), .B(\stack[1][5] ), .Z(n12675) );
  XNOR U13532 ( .A(n12676), .B(n12675), .Z(n12677) );
  XNOR U13533 ( .A(n12678), .B(n12677), .Z(n12679) );
  XNOR U13534 ( .A(n12680), .B(n12679), .Z(n12687) );
  NAND U13535 ( .A(n12682), .B(n12681), .Z(n12685) );
  NANDN U13536 ( .A(\stack[1][62] ), .B(n12683), .Z(n12684) );
  NAND U13537 ( .A(n12685), .B(n12684), .Z(n12686) );
  XNOR U13538 ( .A(n12687), .B(n12686), .Z(n12737) );
  AND U13539 ( .A(o[49]), .B(\stack[1][14] ), .Z(n12689) );
  NAND U13540 ( .A(o[51]), .B(\stack[1][12] ), .Z(n12688) );
  XNOR U13541 ( .A(n12689), .B(n12688), .Z(n12693) );
  AND U13542 ( .A(o[39]), .B(\stack[1][24] ), .Z(n12691) );
  NAND U13543 ( .A(o[40]), .B(\stack[1][23] ), .Z(n12690) );
  XNOR U13544 ( .A(n12691), .B(n12690), .Z(n12692) );
  XOR U13545 ( .A(n12693), .B(n12692), .Z(n12701) );
  AND U13546 ( .A(o[52]), .B(\stack[1][11] ), .Z(n12695) );
  NAND U13547 ( .A(o[55]), .B(\stack[1][8] ), .Z(n12694) );
  XNOR U13548 ( .A(n12695), .B(n12694), .Z(n12699) );
  AND U13549 ( .A(o[48]), .B(\stack[1][15] ), .Z(n12697) );
  NAND U13550 ( .A(o[50]), .B(\stack[1][13] ), .Z(n12696) );
  XNOR U13551 ( .A(n12697), .B(n12696), .Z(n12698) );
  XNOR U13552 ( .A(n12699), .B(n12698), .Z(n12700) );
  XNOR U13553 ( .A(n12701), .B(n12700), .Z(n12727) );
  AND U13554 ( .A(\stack[1][0] ), .B(o[63]), .Z(n12725) );
  AND U13555 ( .A(o[60]), .B(\stack[1][3] ), .Z(n12703) );
  NAND U13556 ( .A(o[59]), .B(\stack[1][4] ), .Z(n12702) );
  XNOR U13557 ( .A(n12703), .B(n12702), .Z(n12707) );
  AND U13558 ( .A(\stack[1][62] ), .B(o[1]), .Z(n12704) );
  NAND U13559 ( .A(n12705), .B(n12704), .Z(n12706) );
  XNOR U13560 ( .A(n12707), .B(n12706), .Z(n12723) );
  AND U13561 ( .A(o[31]), .B(\stack[1][32] ), .Z(n12709) );
  NAND U13562 ( .A(o[33]), .B(\stack[1][30] ), .Z(n12708) );
  XNOR U13563 ( .A(n12709), .B(n12708), .Z(n12713) );
  AND U13564 ( .A(\stack[1][40] ), .B(o[23]), .Z(n12711) );
  NAND U13565 ( .A(\stack[1][46] ), .B(o[17]), .Z(n12710) );
  XNOR U13566 ( .A(n12711), .B(n12710), .Z(n12712) );
  XOR U13567 ( .A(n12713), .B(n12712), .Z(n12721) );
  AND U13568 ( .A(o[37]), .B(\stack[1][26] ), .Z(n12715) );
  NAND U13569 ( .A(o[38]), .B(\stack[1][25] ), .Z(n12714) );
  XNOR U13570 ( .A(n12715), .B(n12714), .Z(n12719) );
  AND U13571 ( .A(o[34]), .B(\stack[1][29] ), .Z(n12717) );
  NAND U13572 ( .A(o[35]), .B(\stack[1][28] ), .Z(n12716) );
  XNOR U13573 ( .A(n12717), .B(n12716), .Z(n12718) );
  XNOR U13574 ( .A(n12719), .B(n12718), .Z(n12720) );
  XNOR U13575 ( .A(n12721), .B(n12720), .Z(n12722) );
  XNOR U13576 ( .A(n12723), .B(n12722), .Z(n12724) );
  XNOR U13577 ( .A(n12725), .B(n12724), .Z(n12726) );
  XOR U13578 ( .A(n12727), .B(n12726), .Z(n12735) );
  AND U13579 ( .A(o[62]), .B(\stack[1][1] ), .Z(n12729) );
  NAND U13580 ( .A(o[61]), .B(\stack[1][2] ), .Z(n12728) );
  XNOR U13581 ( .A(n12729), .B(n12728), .Z(n12733) );
  AND U13582 ( .A(o[56]), .B(\stack[1][7] ), .Z(n12731) );
  NAND U13583 ( .A(o[57]), .B(\stack[1][6] ), .Z(n12730) );
  XNOR U13584 ( .A(n12731), .B(n12730), .Z(n12732) );
  XNOR U13585 ( .A(n12733), .B(n12732), .Z(n12734) );
  XNOR U13586 ( .A(n12735), .B(n12734), .Z(n12736) );
  XOR U13587 ( .A(n12737), .B(n12736), .Z(n12769) );
  AND U13588 ( .A(o[36]), .B(\stack[1][27] ), .Z(n12739) );
  NAND U13589 ( .A(o[43]), .B(\stack[1][20] ), .Z(n12738) );
  XNOR U13590 ( .A(n12739), .B(n12738), .Z(n12743) );
  AND U13591 ( .A(\stack[1][34] ), .B(o[29]), .Z(n12741) );
  NAND U13592 ( .A(o[44]), .B(\stack[1][19] ), .Z(n12740) );
  XNOR U13593 ( .A(n12741), .B(n12740), .Z(n12742) );
  XOR U13594 ( .A(n12743), .B(n12742), .Z(n12751) );
  AND U13595 ( .A(\stack[1][33] ), .B(o[30]), .Z(n12745) );
  NAND U13596 ( .A(o[32]), .B(\stack[1][31] ), .Z(n12744) );
  XNOR U13597 ( .A(n12745), .B(n12744), .Z(n12749) );
  AND U13598 ( .A(\stack[1][35] ), .B(o[28]), .Z(n12747) );
  NAND U13599 ( .A(\stack[1][37] ), .B(o[26]), .Z(n12746) );
  XNOR U13600 ( .A(n12747), .B(n12746), .Z(n12748) );
  XNOR U13601 ( .A(n12749), .B(n12748), .Z(n12750) );
  XNOR U13602 ( .A(n12751), .B(n12750), .Z(n12767) );
  AND U13603 ( .A(\stack[1][36] ), .B(o[27]), .Z(n12753) );
  NAND U13604 ( .A(\stack[1][41] ), .B(o[22]), .Z(n12752) );
  XNOR U13605 ( .A(n12753), .B(n12752), .Z(n12757) );
  AND U13606 ( .A(\stack[1][38] ), .B(o[25]), .Z(n12755) );
  NAND U13607 ( .A(\stack[1][39] ), .B(o[24]), .Z(n12754) );
  XNOR U13608 ( .A(n12755), .B(n12754), .Z(n12756) );
  XOR U13609 ( .A(n12757), .B(n12756), .Z(n12765) );
  AND U13610 ( .A(\stack[1][43] ), .B(o[20]), .Z(n12759) );
  NAND U13611 ( .A(\stack[1][51] ), .B(o[12]), .Z(n12758) );
  XNOR U13612 ( .A(n12759), .B(n12758), .Z(n12763) );
  AND U13613 ( .A(\stack[1][42] ), .B(o[21]), .Z(n12761) );
  NAND U13614 ( .A(\stack[1][49] ), .B(o[14]), .Z(n12760) );
  XNOR U13615 ( .A(n12761), .B(n12760), .Z(n12762) );
  XNOR U13616 ( .A(n12763), .B(n12762), .Z(n12764) );
  XNOR U13617 ( .A(n12765), .B(n12764), .Z(n12766) );
  XNOR U13618 ( .A(n12767), .B(n12766), .Z(n12768) );
  XNOR U13619 ( .A(n12769), .B(n12768), .Z(n12785) );
  NAND U13620 ( .A(n12771), .B(n12770), .Z(n12775) );
  NAND U13621 ( .A(n12773), .B(n12772), .Z(n12774) );
  AND U13622 ( .A(n12775), .B(n12774), .Z(n12783) );
  NAND U13623 ( .A(n12777), .B(n12776), .Z(n12781) );
  NAND U13624 ( .A(n12779), .B(n12778), .Z(n12780) );
  NAND U13625 ( .A(n12781), .B(n12780), .Z(n12782) );
  XNOR U13626 ( .A(n12783), .B(n12782), .Z(n12784) );
  XOR U13627 ( .A(n12785), .B(n12784), .Z(n12817) );
  AND U13628 ( .A(\stack[1][54] ), .B(o[9]), .Z(n12787) );
  NAND U13629 ( .A(\stack[1][58] ), .B(o[5]), .Z(n12786) );
  XNOR U13630 ( .A(n12787), .B(n12786), .Z(n12791) );
  AND U13631 ( .A(\stack[1][56] ), .B(o[7]), .Z(n12789) );
  NAND U13632 ( .A(\stack[1][59] ), .B(o[4]), .Z(n12788) );
  XNOR U13633 ( .A(n12789), .B(n12788), .Z(n12790) );
  XOR U13634 ( .A(n12791), .B(n12790), .Z(n12799) );
  AND U13635 ( .A(\stack[1][57] ), .B(o[6]), .Z(n12793) );
  NAND U13636 ( .A(o[0]), .B(\stack[1][63] ), .Z(n12792) );
  XNOR U13637 ( .A(n12793), .B(n12792), .Z(n12797) );
  AND U13638 ( .A(\stack[1][50] ), .B(o[13]), .Z(n12795) );
  NAND U13639 ( .A(\stack[1][53] ), .B(o[10]), .Z(n12794) );
  XNOR U13640 ( .A(n12795), .B(n12794), .Z(n12796) );
  XNOR U13641 ( .A(n12797), .B(n12796), .Z(n12798) );
  XNOR U13642 ( .A(n12799), .B(n12798), .Z(n12815) );
  AND U13643 ( .A(\stack[1][52] ), .B(o[11]), .Z(n12801) );
  NAND U13644 ( .A(\stack[1][55] ), .B(o[8]), .Z(n12800) );
  XNOR U13645 ( .A(n12801), .B(n12800), .Z(n12805) );
  AND U13646 ( .A(\stack[1][60] ), .B(o[3]), .Z(n12803) );
  NAND U13647 ( .A(\stack[1][61] ), .B(o[2]), .Z(n12802) );
  XNOR U13648 ( .A(n12803), .B(n12802), .Z(n12804) );
  XOR U13649 ( .A(n12805), .B(n12804), .Z(n12813) );
  AND U13650 ( .A(\stack[1][45] ), .B(o[18]), .Z(n12807) );
  NAND U13651 ( .A(\stack[1][47] ), .B(o[16]), .Z(n12806) );
  XNOR U13652 ( .A(n12807), .B(n12806), .Z(n12811) );
  AND U13653 ( .A(\stack[1][44] ), .B(o[19]), .Z(n12809) );
  NAND U13654 ( .A(\stack[1][48] ), .B(o[15]), .Z(n12808) );
  XNOR U13655 ( .A(n12809), .B(n12808), .Z(n12810) );
  XNOR U13656 ( .A(n12811), .B(n12810), .Z(n12812) );
  XNOR U13657 ( .A(n12813), .B(n12812), .Z(n12814) );
  XNOR U13658 ( .A(n12815), .B(n12814), .Z(n12816) );
  XNOR U13659 ( .A(n12817), .B(n12816), .Z(n12833) );
  NAND U13660 ( .A(n12819), .B(n12818), .Z(n12823) );
  NAND U13661 ( .A(n12821), .B(n12820), .Z(n12822) );
  AND U13662 ( .A(n12823), .B(n12822), .Z(n12831) );
  NAND U13663 ( .A(n12825), .B(n12824), .Z(n12829) );
  NAND U13664 ( .A(n12827), .B(n12826), .Z(n12828) );
  NAND U13665 ( .A(n12829), .B(n12828), .Z(n12830) );
  XNOR U13666 ( .A(n12831), .B(n12830), .Z(n12832) );
  XNOR U13667 ( .A(n12833), .B(n12832), .Z(n12834) );
  XNOR U13668 ( .A(n12835), .B(n12834), .Z(n12851) );
  NAND U13669 ( .A(n12837), .B(n12836), .Z(n12841) );
  AND U13670 ( .A(n12839), .B(n12838), .Z(n12840) );
  ANDN U13671 ( .B(n12841), .A(n12840), .Z(n12849) );
  AND U13672 ( .A(n12843), .B(n12842), .Z(n12847) );
  AND U13673 ( .A(n12845), .B(n12844), .Z(n12846) );
  OR U13674 ( .A(n12847), .B(n12846), .Z(n12848) );
  XNOR U13675 ( .A(n12849), .B(n12848), .Z(n12850) );
  XNOR U13676 ( .A(n12851), .B(n12850), .Z(n12852) );
  XNOR U13677 ( .A(n12853), .B(n12852), .Z(n12869) );
  NAND U13678 ( .A(n12855), .B(n12854), .Z(n12859) );
  NAND U13679 ( .A(n12857), .B(n12856), .Z(n12858) );
  AND U13680 ( .A(n12859), .B(n12858), .Z(n12867) );
  NAND U13681 ( .A(n12861), .B(n12860), .Z(n12865) );
  NAND U13682 ( .A(n12863), .B(n12862), .Z(n12864) );
  NAND U13683 ( .A(n12865), .B(n12864), .Z(n12866) );
  XNOR U13684 ( .A(n12867), .B(n12866), .Z(n12868) );
  XNOR U13685 ( .A(n12869), .B(n12868), .Z(n12870) );
  XNOR U13686 ( .A(n12871), .B(n12870), .Z(n12887) );
  NAND U13687 ( .A(n12873), .B(n12872), .Z(n12877) );
  NAND U13688 ( .A(n12875), .B(n12874), .Z(n12876) );
  AND U13689 ( .A(n12877), .B(n12876), .Z(n12885) );
  NAND U13690 ( .A(n12879), .B(n12878), .Z(n12883) );
  NAND U13691 ( .A(n12881), .B(n12880), .Z(n12882) );
  NAND U13692 ( .A(n12883), .B(n12882), .Z(n12884) );
  XNOR U13693 ( .A(n12885), .B(n12884), .Z(n12886) );
  XNOR U13694 ( .A(n12887), .B(n12886), .Z(n12888) );
  XNOR U13695 ( .A(n12889), .B(n12888), .Z(n12905) );
  NAND U13696 ( .A(n12891), .B(n12890), .Z(n12895) );
  NAND U13697 ( .A(n12893), .B(n12892), .Z(n12894) );
  AND U13698 ( .A(n12895), .B(n12894), .Z(n12903) );
  NAND U13699 ( .A(n12897), .B(n12896), .Z(n12901) );
  NAND U13700 ( .A(n12899), .B(n12898), .Z(n12900) );
  NAND U13701 ( .A(n12901), .B(n12900), .Z(n12902) );
  XNOR U13702 ( .A(n12903), .B(n12902), .Z(n12904) );
  XNOR U13703 ( .A(n12905), .B(n12904), .Z(n12906) );
  XNOR U13704 ( .A(n12907), .B(n12906), .Z(n12923) );
  NAND U13705 ( .A(n12909), .B(n12908), .Z(n12913) );
  NAND U13706 ( .A(n12911), .B(n12910), .Z(n12912) );
  AND U13707 ( .A(n12913), .B(n12912), .Z(n12921) );
  NAND U13708 ( .A(n12915), .B(n12914), .Z(n12919) );
  NAND U13709 ( .A(n12917), .B(n12916), .Z(n12918) );
  NAND U13710 ( .A(n12919), .B(n12918), .Z(n12920) );
  XNOR U13711 ( .A(n12921), .B(n12920), .Z(n12922) );
  XNOR U13712 ( .A(n12923), .B(n12922), .Z(n12924) );
  XNOR U13713 ( .A(n12925), .B(n12924), .Z(n12941) );
  NAND U13714 ( .A(n12927), .B(n12926), .Z(n12931) );
  NAND U13715 ( .A(n12929), .B(n12928), .Z(n12930) );
  AND U13716 ( .A(n12931), .B(n12930), .Z(n12939) );
  NAND U13717 ( .A(n12933), .B(n12932), .Z(n12937) );
  NAND U13718 ( .A(n12935), .B(n12934), .Z(n12936) );
  NAND U13719 ( .A(n12937), .B(n12936), .Z(n12938) );
  XNOR U13720 ( .A(n12939), .B(n12938), .Z(n12940) );
  XNOR U13721 ( .A(n12941), .B(n12940), .Z(n12942) );
  XNOR U13722 ( .A(n12943), .B(n12942), .Z(n12959) );
  NAND U13723 ( .A(n12945), .B(n12944), .Z(n12949) );
  NAND U13724 ( .A(n12947), .B(n12946), .Z(n12948) );
  AND U13725 ( .A(n12949), .B(n12948), .Z(n12957) );
  NAND U13726 ( .A(n12951), .B(n12950), .Z(n12955) );
  NAND U13727 ( .A(n12953), .B(n12952), .Z(n12954) );
  NAND U13728 ( .A(n12955), .B(n12954), .Z(n12956) );
  XNOR U13729 ( .A(n12957), .B(n12956), .Z(n12958) );
  XNOR U13730 ( .A(n12959), .B(n12958), .Z(n12960) );
  XNOR U13731 ( .A(n12961), .B(n12960), .Z(n12977) );
  NAND U13732 ( .A(n12963), .B(n12962), .Z(n12967) );
  NAND U13733 ( .A(n12965), .B(n12964), .Z(n12966) );
  AND U13734 ( .A(n12967), .B(n12966), .Z(n12975) );
  NANDN U13735 ( .A(n12969), .B(n12968), .Z(n12973) );
  NAND U13736 ( .A(n12971), .B(n12970), .Z(n12972) );
  NAND U13737 ( .A(n12973), .B(n12972), .Z(n12974) );
  XNOR U13738 ( .A(n12975), .B(n12974), .Z(n12976) );
  XNOR U13739 ( .A(n12977), .B(n12976), .Z(n12978) );
  XNOR U13740 ( .A(n12979), .B(n12978), .Z(n12995) );
  NAND U13741 ( .A(n12981), .B(n12980), .Z(n12985) );
  NAND U13742 ( .A(n12983), .B(n12982), .Z(n12984) );
  AND U13743 ( .A(n12985), .B(n12984), .Z(n12993) );
  NAND U13744 ( .A(n12987), .B(n12986), .Z(n12991) );
  NAND U13745 ( .A(n12989), .B(n12988), .Z(n12990) );
  NAND U13746 ( .A(n12991), .B(n12990), .Z(n12992) );
  XNOR U13747 ( .A(n12993), .B(n12992), .Z(n12994) );
  XNOR U13748 ( .A(n12995), .B(n12994), .Z(n12996) );
  XNOR U13749 ( .A(n12997), .B(n12996), .Z(n13013) );
  NAND U13750 ( .A(n12999), .B(n12998), .Z(n13003) );
  AND U13751 ( .A(n13001), .B(n13000), .Z(n13002) );
  ANDN U13752 ( .B(n13003), .A(n13002), .Z(n13011) );
  AND U13753 ( .A(n13005), .B(n13004), .Z(n13009) );
  AND U13754 ( .A(n13007), .B(n13006), .Z(n13008) );
  OR U13755 ( .A(n13009), .B(n13008), .Z(n13010) );
  XNOR U13756 ( .A(n13011), .B(n13010), .Z(n13012) );
  XNOR U13757 ( .A(n13013), .B(n13012), .Z(n13014) );
  XNOR U13758 ( .A(n13015), .B(n13014), .Z(n13031) );
  NAND U13759 ( .A(n13017), .B(n13016), .Z(n13021) );
  NAND U13760 ( .A(n13019), .B(n13018), .Z(n13020) );
  AND U13761 ( .A(n13021), .B(n13020), .Z(n13029) );
  NAND U13762 ( .A(n13023), .B(n13022), .Z(n13027) );
  NAND U13763 ( .A(n13025), .B(n13024), .Z(n13026) );
  NAND U13764 ( .A(n13027), .B(n13026), .Z(n13028) );
  XNOR U13765 ( .A(n13029), .B(n13028), .Z(n13030) );
  XNOR U13766 ( .A(n13031), .B(n13030), .Z(n13032) );
  XNOR U13767 ( .A(n13033), .B(n13032), .Z(n13049) );
  NAND U13768 ( .A(n13035), .B(n13034), .Z(n13039) );
  NAND U13769 ( .A(n13037), .B(n13036), .Z(n13038) );
  AND U13770 ( .A(n13039), .B(n13038), .Z(n13047) );
  NAND U13771 ( .A(n13041), .B(n13040), .Z(n13045) );
  NAND U13772 ( .A(n13043), .B(n13042), .Z(n13044) );
  NAND U13773 ( .A(n13045), .B(n13044), .Z(n13046) );
  XNOR U13774 ( .A(n13047), .B(n13046), .Z(n13048) );
  XNOR U13775 ( .A(n13049), .B(n13048), .Z(n13050) );
  XNOR U13776 ( .A(n13051), .B(n13050), .Z(n13067) );
  NAND U13777 ( .A(n13053), .B(n13052), .Z(n13057) );
  NAND U13778 ( .A(n13055), .B(n13054), .Z(n13056) );
  AND U13779 ( .A(n13057), .B(n13056), .Z(n13065) );
  NAND U13780 ( .A(n13059), .B(n13058), .Z(n13063) );
  NAND U13781 ( .A(n13061), .B(n13060), .Z(n13062) );
  NAND U13782 ( .A(n13063), .B(n13062), .Z(n13064) );
  XNOR U13783 ( .A(n13065), .B(n13064), .Z(n13066) );
  XNOR U13784 ( .A(n13067), .B(n13066), .Z(n13068) );
  XNOR U13785 ( .A(n13069), .B(n13068), .Z(n13085) );
  NAND U13786 ( .A(n13071), .B(n13070), .Z(n13075) );
  NAND U13787 ( .A(n13073), .B(n13072), .Z(n13074) );
  AND U13788 ( .A(n13075), .B(n13074), .Z(n13083) );
  NAND U13789 ( .A(n13077), .B(n13076), .Z(n13081) );
  NAND U13790 ( .A(n13079), .B(n13078), .Z(n13080) );
  NAND U13791 ( .A(n13081), .B(n13080), .Z(n13082) );
  XNOR U13792 ( .A(n13083), .B(n13082), .Z(n13084) );
  XNOR U13793 ( .A(n13085), .B(n13084), .Z(n13086) );
  XNOR U13794 ( .A(n13087), .B(n13086), .Z(n13103) );
  NAND U13795 ( .A(n13089), .B(n13088), .Z(n13093) );
  NAND U13796 ( .A(n13091), .B(n13090), .Z(n13092) );
  AND U13797 ( .A(n13093), .B(n13092), .Z(n13101) );
  NAND U13798 ( .A(n13095), .B(n13094), .Z(n13099) );
  NAND U13799 ( .A(n13097), .B(n13096), .Z(n13098) );
  NAND U13800 ( .A(n13099), .B(n13098), .Z(n13100) );
  XNOR U13801 ( .A(n13101), .B(n13100), .Z(n13102) );
  XNOR U13802 ( .A(n13103), .B(n13102), .Z(n13104) );
  XNOR U13803 ( .A(n13105), .B(n13104), .Z(n13121) );
  NAND U13804 ( .A(n13107), .B(n13106), .Z(n13111) );
  NAND U13805 ( .A(n13109), .B(n13108), .Z(n13110) );
  AND U13806 ( .A(n13111), .B(n13110), .Z(n13119) );
  NAND U13807 ( .A(n13113), .B(n13112), .Z(n13117) );
  NAND U13808 ( .A(n13115), .B(n13114), .Z(n13116) );
  NAND U13809 ( .A(n13117), .B(n13116), .Z(n13118) );
  XNOR U13810 ( .A(n13119), .B(n13118), .Z(n13120) );
  XNOR U13811 ( .A(n13121), .B(n13120), .Z(n13122) );
  XNOR U13812 ( .A(n13123), .B(n13122), .Z(n13823) );
  NAND U13813 ( .A(\stack[1][4] ), .B(o[52]), .Z(n13427) );
  NAND U13814 ( .A(\stack[1][4] ), .B(o[48]), .Z(n13404) );
  NAND U13815 ( .A(\stack[1][4] ), .B(o[44]), .Z(n13378) );
  NAND U13816 ( .A(\stack[1][4] ), .B(o[38]), .Z(n13342) );
  NAND U13817 ( .A(\stack[1][4] ), .B(o[28]), .Z(n13282) );
  NAND U13818 ( .A(\stack[1][4] ), .B(o[22]), .Z(n13248) );
  NAND U13819 ( .A(\stack[1][4] ), .B(o[18]), .Z(n13224) );
  XNOR U13820 ( .A(n13127), .B(n13126), .Z(n13194) );
  XNOR U13821 ( .A(n13129), .B(n13128), .Z(n13172) );
  AND U13822 ( .A(\stack[1][4] ), .B(o[5]), .Z(n13151) );
  XOR U13823 ( .A(n13131), .B(n13130), .Z(n13152) );
  NAND U13824 ( .A(n13151), .B(n13152), .Z(n13154) );
  AND U13825 ( .A(\stack[1][5] ), .B(o[1]), .Z(n13137) );
  AND U13826 ( .A(o[0]), .B(\stack[1][4] ), .Z(n13132) );
  AND U13827 ( .A(n13137), .B(n13132), .Z(n13133) );
  NAND U13828 ( .A(n13133), .B(o[2]), .Z(n13139) );
  NAND U13829 ( .A(n13137), .B(o[0]), .Z(n13134) );
  XNOR U13830 ( .A(o[2]), .B(n13134), .Z(n13135) );
  AND U13831 ( .A(\stack[1][4] ), .B(n13135), .Z(n13484) );
  NAND U13832 ( .A(\stack[1][6] ), .B(o[0]), .Z(n13136) );
  XNOR U13833 ( .A(n13137), .B(n13136), .Z(n13485) );
  NAND U13834 ( .A(n13484), .B(n13485), .Z(n13138) );
  NAND U13835 ( .A(n13139), .B(n13138), .Z(n13142) );
  NAND U13836 ( .A(n13142), .B(n13143), .Z(n13145) );
  AND U13837 ( .A(\stack[1][4] ), .B(o[3]), .Z(n13492) );
  NAND U13838 ( .A(n13492), .B(n13493), .Z(n13144) );
  NAND U13839 ( .A(n13145), .B(n13144), .Z(n13148) );
  AND U13840 ( .A(\stack[1][4] ), .B(o[4]), .Z(n17175) );
  NAND U13841 ( .A(n13148), .B(n17175), .Z(n13150) );
  NAND U13842 ( .A(n13497), .B(n13496), .Z(n13149) );
  NAND U13843 ( .A(n13150), .B(n13149), .Z(n13502) );
  NAND U13844 ( .A(n13502), .B(n13503), .Z(n13153) );
  NAND U13845 ( .A(n13154), .B(n13153), .Z(n13156) );
  XOR U13846 ( .A(n17136), .B(n13155), .Z(n13157) );
  NAND U13847 ( .A(n13156), .B(n13157), .Z(n13159) );
  AND U13848 ( .A(\stack[1][4] ), .B(o[6]), .Z(n13509) );
  NAND U13849 ( .A(n13509), .B(n13508), .Z(n13158) );
  NAND U13850 ( .A(n13159), .B(n13158), .Z(n13162) );
  XOR U13851 ( .A(n13161), .B(n13160), .Z(n13163) );
  NAND U13852 ( .A(n13162), .B(n13163), .Z(n13165) );
  AND U13853 ( .A(\stack[1][4] ), .B(o[7]), .Z(n13514) );
  NAND U13854 ( .A(n13514), .B(n13515), .Z(n13164) );
  NAND U13855 ( .A(n13165), .B(n13164), .Z(n13168) );
  AND U13856 ( .A(\stack[1][4] ), .B(o[8]), .Z(n13169) );
  NAND U13857 ( .A(n13168), .B(n13169), .Z(n13171) );
  NAND U13858 ( .A(n13521), .B(n13520), .Z(n13170) );
  AND U13859 ( .A(n13171), .B(n13170), .Z(n13173) );
  NAND U13860 ( .A(n13172), .B(n13173), .Z(n13175) );
  NAND U13861 ( .A(\stack[1][4] ), .B(o[9]), .Z(n13526) );
  NAND U13862 ( .A(n13527), .B(n13526), .Z(n13174) );
  AND U13863 ( .A(n13175), .B(n13174), .Z(n13178) );
  AND U13864 ( .A(o[10]), .B(\stack[1][4] ), .Z(n13179) );
  NAND U13865 ( .A(n13178), .B(n13179), .Z(n13181) );
  NAND U13866 ( .A(n13476), .B(n13475), .Z(n13180) );
  NAND U13867 ( .A(n13181), .B(n13180), .Z(n13184) );
  NAND U13868 ( .A(n13184), .B(n13185), .Z(n13187) );
  AND U13869 ( .A(\stack[1][4] ), .B(o[11]), .Z(n13537) );
  NAND U13870 ( .A(n13537), .B(n13536), .Z(n13186) );
  NAND U13871 ( .A(n13187), .B(n13186), .Z(n13190) );
  AND U13872 ( .A(\stack[1][4] ), .B(o[12]), .Z(n13191) );
  NAND U13873 ( .A(n13190), .B(n13191), .Z(n13193) );
  XNOR U13874 ( .A(n13189), .B(n13188), .Z(n13542) );
  NAND U13875 ( .A(n13542), .B(n13543), .Z(n13192) );
  AND U13876 ( .A(n13193), .B(n13192), .Z(n13195) );
  NAND U13877 ( .A(n13194), .B(n13195), .Z(n13197) );
  NAND U13878 ( .A(\stack[1][4] ), .B(o[13]), .Z(n13548) );
  NAND U13879 ( .A(n13549), .B(n13548), .Z(n13196) );
  NAND U13880 ( .A(n13197), .B(n13196), .Z(n13198) );
  NAND U13881 ( .A(\stack[1][4] ), .B(o[14]), .Z(n13199) );
  NAND U13882 ( .A(n13198), .B(n13199), .Z(n13203) );
  XNOR U13883 ( .A(n13201), .B(n13200), .Z(n13554) );
  NAND U13884 ( .A(n13555), .B(n13554), .Z(n13202) );
  AND U13885 ( .A(n13203), .B(n13202), .Z(n13207) );
  XOR U13886 ( .A(n13205), .B(n13204), .Z(n13206) );
  NAND U13887 ( .A(n13207), .B(n13206), .Z(n13209) );
  AND U13888 ( .A(\stack[1][4] ), .B(o[15]), .Z(n13561) );
  XOR U13889 ( .A(n13207), .B(n13206), .Z(n13560) );
  NAND U13890 ( .A(n13561), .B(n13560), .Z(n13208) );
  NAND U13891 ( .A(n13209), .B(n13208), .Z(n13210) );
  AND U13892 ( .A(\stack[1][4] ), .B(o[16]), .Z(n13211) );
  NAND U13893 ( .A(n13210), .B(n13211), .Z(n13215) );
  NAND U13894 ( .A(n13567), .B(n13566), .Z(n13214) );
  NAND U13895 ( .A(n13215), .B(n13214), .Z(n13218) );
  XOR U13896 ( .A(n13217), .B(n13216), .Z(n13219) );
  NAND U13897 ( .A(n13218), .B(n13219), .Z(n13221) );
  AND U13898 ( .A(\stack[1][4] ), .B(o[17]), .Z(n13572) );
  NAND U13899 ( .A(n13572), .B(n13573), .Z(n13220) );
  AND U13900 ( .A(n13221), .B(n13220), .Z(n13225) );
  NAND U13901 ( .A(n13224), .B(n13225), .Z(n13227) );
  XNOR U13902 ( .A(n13223), .B(n13222), .Z(n13473) );
  NAND U13903 ( .A(n13473), .B(n13474), .Z(n13226) );
  AND U13904 ( .A(n13227), .B(n13226), .Z(n13231) );
  XOR U13905 ( .A(n13229), .B(n13228), .Z(n13230) );
  NAND U13906 ( .A(n13231), .B(n13230), .Z(n13233) );
  AND U13907 ( .A(\stack[1][4] ), .B(o[19]), .Z(n13583) );
  XOR U13908 ( .A(n13231), .B(n13230), .Z(n13582) );
  NAND U13909 ( .A(n13583), .B(n13582), .Z(n13232) );
  NAND U13910 ( .A(n13233), .B(n13232), .Z(n13234) );
  AND U13911 ( .A(\stack[1][4] ), .B(o[20]), .Z(n13235) );
  NAND U13912 ( .A(n13234), .B(n13235), .Z(n13239) );
  NAND U13913 ( .A(n13589), .B(n13588), .Z(n13238) );
  NAND U13914 ( .A(n13239), .B(n13238), .Z(n13242) );
  XOR U13915 ( .A(n13241), .B(n13240), .Z(n13243) );
  NAND U13916 ( .A(n13242), .B(n13243), .Z(n13245) );
  AND U13917 ( .A(\stack[1][4] ), .B(o[21]), .Z(n13594) );
  NAND U13918 ( .A(n13594), .B(n13595), .Z(n13244) );
  AND U13919 ( .A(n13245), .B(n13244), .Z(n13249) );
  NAND U13920 ( .A(n13248), .B(n13249), .Z(n13251) );
  XNOR U13921 ( .A(n13247), .B(n13246), .Z(n13471) );
  NAND U13922 ( .A(n13471), .B(n13472), .Z(n13250) );
  AND U13923 ( .A(n13251), .B(n13250), .Z(n13255) );
  XOR U13924 ( .A(n13253), .B(n13252), .Z(n13254) );
  NAND U13925 ( .A(n13255), .B(n13254), .Z(n13257) );
  AND U13926 ( .A(\stack[1][4] ), .B(o[23]), .Z(n13605) );
  XOR U13927 ( .A(n13255), .B(n13254), .Z(n13604) );
  NAND U13928 ( .A(n13605), .B(n13604), .Z(n13256) );
  NAND U13929 ( .A(n13257), .B(n13256), .Z(n13258) );
  AND U13930 ( .A(\stack[1][4] ), .B(o[24]), .Z(n13259) );
  NAND U13931 ( .A(n13258), .B(n13259), .Z(n13263) );
  NAND U13932 ( .A(n13611), .B(n13610), .Z(n13262) );
  NAND U13933 ( .A(n13263), .B(n13262), .Z(n13266) );
  XOR U13934 ( .A(n13265), .B(n13264), .Z(n13267) );
  NAND U13935 ( .A(n13266), .B(n13267), .Z(n13269) );
  AND U13936 ( .A(\stack[1][4] ), .B(o[25]), .Z(n13616) );
  NAND U13937 ( .A(n13616), .B(n13617), .Z(n13268) );
  NAND U13938 ( .A(n13269), .B(n13268), .Z(n13270) );
  AND U13939 ( .A(\stack[1][4] ), .B(o[26]), .Z(n13271) );
  NAND U13940 ( .A(n13270), .B(n13271), .Z(n13275) );
  NAND U13941 ( .A(n13623), .B(n13622), .Z(n13274) );
  NAND U13942 ( .A(n13275), .B(n13274), .Z(n13278) );
  XOR U13943 ( .A(n13277), .B(n13276), .Z(n13279) );
  NAND U13944 ( .A(n13278), .B(n13279), .Z(n13281) );
  AND U13945 ( .A(\stack[1][4] ), .B(o[27]), .Z(n13628) );
  NAND U13946 ( .A(n13628), .B(n13629), .Z(n13280) );
  AND U13947 ( .A(n13281), .B(n13280), .Z(n13283) );
  NAND U13948 ( .A(n13282), .B(n13283), .Z(n13287) );
  XNOR U13949 ( .A(n13285), .B(n13284), .Z(n13634) );
  NAND U13950 ( .A(n13635), .B(n13634), .Z(n13286) );
  AND U13951 ( .A(n13287), .B(n13286), .Z(n13291) );
  XOR U13952 ( .A(n13289), .B(n13288), .Z(n13290) );
  NAND U13953 ( .A(n13291), .B(n13290), .Z(n13293) );
  AND U13954 ( .A(\stack[1][4] ), .B(o[29]), .Z(n13640) );
  XOR U13955 ( .A(n13291), .B(n13290), .Z(n13641) );
  NAND U13956 ( .A(n13640), .B(n13641), .Z(n13292) );
  NAND U13957 ( .A(n13293), .B(n13292), .Z(n13296) );
  AND U13958 ( .A(\stack[1][4] ), .B(o[30]), .Z(n13297) );
  NAND U13959 ( .A(n13296), .B(n13297), .Z(n13299) );
  NAND U13960 ( .A(n13647), .B(n13646), .Z(n13298) );
  NAND U13961 ( .A(n13299), .B(n13298), .Z(n13302) );
  XOR U13962 ( .A(n13301), .B(n13300), .Z(n13303) );
  NAND U13963 ( .A(n13302), .B(n13303), .Z(n13305) );
  AND U13964 ( .A(\stack[1][4] ), .B(o[31]), .Z(n13652) );
  NAND U13965 ( .A(n13652), .B(n13653), .Z(n13304) );
  NAND U13966 ( .A(n13305), .B(n13304), .Z(n13306) );
  AND U13967 ( .A(\stack[1][4] ), .B(o[32]), .Z(n13307) );
  NAND U13968 ( .A(n13306), .B(n13307), .Z(n13311) );
  NAND U13969 ( .A(n13659), .B(n13658), .Z(n13310) );
  NAND U13970 ( .A(n13311), .B(n13310), .Z(n13314) );
  XOR U13971 ( .A(n13313), .B(n13312), .Z(n13315) );
  NAND U13972 ( .A(n13314), .B(n13315), .Z(n13317) );
  AND U13973 ( .A(\stack[1][4] ), .B(o[33]), .Z(n13664) );
  NAND U13974 ( .A(n13664), .B(n13665), .Z(n13316) );
  NAND U13975 ( .A(n13317), .B(n13316), .Z(n13318) );
  AND U13976 ( .A(\stack[1][4] ), .B(o[34]), .Z(n13319) );
  NAND U13977 ( .A(n13318), .B(n13319), .Z(n13323) );
  NAND U13978 ( .A(n13671), .B(n13670), .Z(n13322) );
  NAND U13979 ( .A(n13323), .B(n13322), .Z(n13326) );
  XOR U13980 ( .A(n13325), .B(n13324), .Z(n13327) );
  NAND U13981 ( .A(n13326), .B(n13327), .Z(n13329) );
  AND U13982 ( .A(\stack[1][4] ), .B(o[35]), .Z(n13676) );
  NAND U13983 ( .A(n13676), .B(n13677), .Z(n13328) );
  NAND U13984 ( .A(n13329), .B(n13328), .Z(n13330) );
  AND U13985 ( .A(\stack[1][4] ), .B(o[36]), .Z(n13331) );
  NAND U13986 ( .A(n13330), .B(n13331), .Z(n13335) );
  NAND U13987 ( .A(n13683), .B(n13682), .Z(n13334) );
  NAND U13988 ( .A(n13335), .B(n13334), .Z(n13338) );
  XOR U13989 ( .A(n13337), .B(n13336), .Z(n13339) );
  NAND U13990 ( .A(n13338), .B(n13339), .Z(n13341) );
  AND U13991 ( .A(\stack[1][4] ), .B(o[37]), .Z(n13688) );
  NAND U13992 ( .A(n13688), .B(n13689), .Z(n13340) );
  AND U13993 ( .A(n13341), .B(n13340), .Z(n13343) );
  NAND U13994 ( .A(n13342), .B(n13343), .Z(n13347) );
  XNOR U13995 ( .A(n13345), .B(n13344), .Z(n13694) );
  NAND U13996 ( .A(n13695), .B(n13694), .Z(n13346) );
  AND U13997 ( .A(n13347), .B(n13346), .Z(n13351) );
  XOR U13998 ( .A(n13349), .B(n13348), .Z(n13350) );
  NAND U13999 ( .A(n13351), .B(n13350), .Z(n13353) );
  AND U14000 ( .A(\stack[1][4] ), .B(o[39]), .Z(n13700) );
  XOR U14001 ( .A(n13351), .B(n13350), .Z(n13701) );
  NAND U14002 ( .A(n13700), .B(n13701), .Z(n13352) );
  NAND U14003 ( .A(n13353), .B(n13352), .Z(n13354) );
  AND U14004 ( .A(\stack[1][4] ), .B(o[40]), .Z(n13355) );
  NAND U14005 ( .A(n13354), .B(n13355), .Z(n13359) );
  NAND U14006 ( .A(n13707), .B(n13706), .Z(n13358) );
  NAND U14007 ( .A(n13359), .B(n13358), .Z(n13362) );
  XOR U14008 ( .A(n13361), .B(n13360), .Z(n13363) );
  NAND U14009 ( .A(n13362), .B(n13363), .Z(n13365) );
  AND U14010 ( .A(\stack[1][4] ), .B(o[41]), .Z(n13713) );
  NAND U14011 ( .A(n13713), .B(n13712), .Z(n13364) );
  NAND U14012 ( .A(n13365), .B(n13364), .Z(n13366) );
  AND U14013 ( .A(\stack[1][4] ), .B(o[42]), .Z(n13367) );
  NAND U14014 ( .A(n13366), .B(n13367), .Z(n13371) );
  NAND U14015 ( .A(n13719), .B(n13718), .Z(n13370) );
  NAND U14016 ( .A(n13371), .B(n13370), .Z(n13374) );
  XOR U14017 ( .A(n13373), .B(n13372), .Z(n13375) );
  NAND U14018 ( .A(n13374), .B(n13375), .Z(n13377) );
  AND U14019 ( .A(\stack[1][4] ), .B(o[43]), .Z(n13725) );
  NAND U14020 ( .A(n13725), .B(n13724), .Z(n13376) );
  AND U14021 ( .A(n13377), .B(n13376), .Z(n13379) );
  NAND U14022 ( .A(n13378), .B(n13379), .Z(n13383) );
  XNOR U14023 ( .A(n13381), .B(n13380), .Z(n13730) );
  NAND U14024 ( .A(n13731), .B(n13730), .Z(n13382) );
  AND U14025 ( .A(n13383), .B(n13382), .Z(n13387) );
  XOR U14026 ( .A(n13385), .B(n13384), .Z(n13386) );
  NAND U14027 ( .A(n13387), .B(n13386), .Z(n13389) );
  AND U14028 ( .A(\stack[1][4] ), .B(o[45]), .Z(n13737) );
  XOR U14029 ( .A(n13387), .B(n13386), .Z(n13736) );
  NAND U14030 ( .A(n13737), .B(n13736), .Z(n13388) );
  NAND U14031 ( .A(n13389), .B(n13388), .Z(n13390) );
  AND U14032 ( .A(\stack[1][4] ), .B(o[46]), .Z(n13391) );
  NAND U14033 ( .A(n13390), .B(n13391), .Z(n13395) );
  NAND U14034 ( .A(n13743), .B(n13742), .Z(n13394) );
  NAND U14035 ( .A(n13395), .B(n13394), .Z(n13398) );
  XOR U14036 ( .A(n13397), .B(n13396), .Z(n13399) );
  NAND U14037 ( .A(n13398), .B(n13399), .Z(n13401) );
  AND U14038 ( .A(\stack[1][4] ), .B(o[47]), .Z(n13748) );
  NAND U14039 ( .A(n13748), .B(n13749), .Z(n13400) );
  AND U14040 ( .A(n13401), .B(n13400), .Z(n13405) );
  NAND U14041 ( .A(n13404), .B(n13405), .Z(n13407) );
  XNOR U14042 ( .A(n13403), .B(n13402), .Z(n13469) );
  NAND U14043 ( .A(n13469), .B(n13470), .Z(n13406) );
  AND U14044 ( .A(n13407), .B(n13406), .Z(n13411) );
  XOR U14045 ( .A(n13409), .B(n13408), .Z(n13410) );
  NAND U14046 ( .A(n13411), .B(n13410), .Z(n13413) );
  AND U14047 ( .A(\stack[1][4] ), .B(o[49]), .Z(n13759) );
  XOR U14048 ( .A(n13411), .B(n13410), .Z(n13758) );
  NAND U14049 ( .A(n13759), .B(n13758), .Z(n13412) );
  NAND U14050 ( .A(n13413), .B(n13412), .Z(n13414) );
  AND U14051 ( .A(\stack[1][4] ), .B(o[50]), .Z(n13415) );
  NAND U14052 ( .A(n13414), .B(n13415), .Z(n13420) );
  IV U14053 ( .A(n13416), .Z(n13417) );
  XNOR U14054 ( .A(n13418), .B(n13417), .Z(n13764) );
  NAND U14055 ( .A(n13765), .B(n13764), .Z(n13419) );
  NAND U14056 ( .A(n13420), .B(n13419), .Z(n13423) );
  XOR U14057 ( .A(n13422), .B(n13421), .Z(n13424) );
  NAND U14058 ( .A(n13423), .B(n13424), .Z(n13426) );
  AND U14059 ( .A(\stack[1][4] ), .B(o[51]), .Z(n13770) );
  NAND U14060 ( .A(n13770), .B(n13771), .Z(n13425) );
  AND U14061 ( .A(n13426), .B(n13425), .Z(n13429) );
  NAND U14062 ( .A(n13427), .B(n13429), .Z(n13433) );
  IV U14063 ( .A(n13427), .Z(n13428) );
  XNOR U14064 ( .A(n13429), .B(n13428), .Z(n13468) );
  XNOR U14065 ( .A(n13431), .B(n13430), .Z(n13467) );
  NAND U14066 ( .A(n13468), .B(n13467), .Z(n13432) );
  AND U14067 ( .A(n13433), .B(n13432), .Z(n13437) );
  XOR U14068 ( .A(n13435), .B(n13434), .Z(n13436) );
  NAND U14069 ( .A(n13437), .B(n13436), .Z(n13439) );
  AND U14070 ( .A(\stack[1][4] ), .B(o[53]), .Z(n13780) );
  XOR U14071 ( .A(n13437), .B(n13436), .Z(n13781) );
  NAND U14072 ( .A(n13780), .B(n13781), .Z(n13438) );
  NAND U14073 ( .A(n13439), .B(n13438), .Z(n13440) );
  AND U14074 ( .A(\stack[1][4] ), .B(o[54]), .Z(n13441) );
  NAND U14075 ( .A(n13440), .B(n13441), .Z(n13447) );
  IV U14076 ( .A(n13440), .Z(n13442) );
  XNOR U14077 ( .A(n13442), .B(n13441), .Z(n13787) );
  IV U14078 ( .A(n13443), .Z(n13444) );
  XNOR U14079 ( .A(n13445), .B(n13444), .Z(n13786) );
  NAND U14080 ( .A(n13787), .B(n13786), .Z(n13446) );
  NAND U14081 ( .A(n13447), .B(n13446), .Z(n13450) );
  XOR U14082 ( .A(n13449), .B(n13448), .Z(n13451) );
  NAND U14083 ( .A(n13450), .B(n13451), .Z(n13453) );
  AND U14084 ( .A(\stack[1][4] ), .B(o[55]), .Z(n13792) );
  NAND U14085 ( .A(n13792), .B(n13793), .Z(n13452) );
  NAND U14086 ( .A(n13453), .B(n13452), .Z(n13454) );
  AND U14087 ( .A(\stack[1][4] ), .B(o[56]), .Z(n13455) );
  NAND U14088 ( .A(n13454), .B(n13455), .Z(n13460) );
  IV U14089 ( .A(n13456), .Z(n13457) );
  XNOR U14090 ( .A(n13458), .B(n13457), .Z(n13798) );
  NAND U14091 ( .A(n13799), .B(n13798), .Z(n13459) );
  NAND U14092 ( .A(n13460), .B(n13459), .Z(n13463) );
  XOR U14093 ( .A(n13462), .B(n13461), .Z(n13464) );
  NAND U14094 ( .A(n13463), .B(n13464), .Z(n13466) );
  AND U14095 ( .A(\stack[1][4] ), .B(o[57]), .Z(n13805) );
  NAND U14096 ( .A(n13805), .B(n13804), .Z(n13465) );
  AND U14097 ( .A(n13466), .B(n13465), .Z(n13817) );
  NAND U14098 ( .A(\stack[1][4] ), .B(o[58]), .Z(n13816) );
  XOR U14099 ( .A(n13817), .B(n13816), .Z(n13814) );
  XNOR U14100 ( .A(n13468), .B(n13467), .Z(n13776) );
  XNOR U14101 ( .A(n13476), .B(n13475), .Z(n13532) );
  AND U14102 ( .A(o[0]), .B(\stack[1][3] ), .Z(n14190) );
  AND U14103 ( .A(o[1]), .B(\stack[1][4] ), .Z(n13481) );
  AND U14104 ( .A(n14190), .B(n13481), .Z(n13477) );
  NAND U14105 ( .A(o[2]), .B(n13477), .Z(n13483) );
  NAND U14106 ( .A(n13481), .B(o[0]), .Z(n13478) );
  XNOR U14107 ( .A(o[2]), .B(n13478), .Z(n13479) );
  AND U14108 ( .A(\stack[1][3] ), .B(n13479), .Z(n13839) );
  NAND U14109 ( .A(\stack[1][5] ), .B(o[0]), .Z(n13480) );
  XNOR U14110 ( .A(n13481), .B(n13480), .Z(n13840) );
  NAND U14111 ( .A(n13839), .B(n13840), .Z(n13482) );
  NAND U14112 ( .A(n13483), .B(n13482), .Z(n13486) );
  NAND U14113 ( .A(n13486), .B(n13487), .Z(n13489) );
  AND U14114 ( .A(\stack[1][3] ), .B(o[3]), .Z(n17214) );
  NAND U14115 ( .A(n17214), .B(n13845), .Z(n13488) );
  NAND U14116 ( .A(n13489), .B(n13488), .Z(n13490) );
  AND U14117 ( .A(\stack[1][3] ), .B(o[4]), .Z(n13491) );
  NAND U14118 ( .A(n13490), .B(n13491), .Z(n13495) );
  NAND U14119 ( .A(n13831), .B(n13830), .Z(n13494) );
  NAND U14120 ( .A(n13495), .B(n13494), .Z(n13498) );
  XOR U14121 ( .A(n13497), .B(n13496), .Z(n13499) );
  NAND U14122 ( .A(n13498), .B(n13499), .Z(n13501) );
  AND U14123 ( .A(\stack[1][3] ), .B(o[5]), .Z(n13854) );
  NAND U14124 ( .A(n13854), .B(n13855), .Z(n13500) );
  NAND U14125 ( .A(n13501), .B(n13500), .Z(n13504) );
  NAND U14126 ( .A(n13504), .B(n13505), .Z(n13507) );
  AND U14127 ( .A(\stack[1][3] ), .B(o[6]), .Z(n13861) );
  NAND U14128 ( .A(n13861), .B(n13860), .Z(n13506) );
  NAND U14129 ( .A(n13507), .B(n13506), .Z(n13510) );
  XOR U14130 ( .A(n13509), .B(n13508), .Z(n13511) );
  NAND U14131 ( .A(n13510), .B(n13511), .Z(n13513) );
  AND U14132 ( .A(\stack[1][3] ), .B(o[7]), .Z(n13866) );
  NAND U14133 ( .A(n13866), .B(n13867), .Z(n13512) );
  NAND U14134 ( .A(n13513), .B(n13512), .Z(n13516) );
  AND U14135 ( .A(\stack[1][3] ), .B(o[8]), .Z(n13517) );
  NAND U14136 ( .A(n13516), .B(n13517), .Z(n13519) );
  NAND U14137 ( .A(n13829), .B(n13828), .Z(n13518) );
  NAND U14138 ( .A(n13519), .B(n13518), .Z(n13522) );
  XOR U14139 ( .A(n13521), .B(n13520), .Z(n13523) );
  NAND U14140 ( .A(n13522), .B(n13523), .Z(n13525) );
  AND U14141 ( .A(\stack[1][3] ), .B(o[9]), .Z(n13876) );
  NAND U14142 ( .A(n13876), .B(n13877), .Z(n13524) );
  NAND U14143 ( .A(n13525), .B(n13524), .Z(n13528) );
  AND U14144 ( .A(o[10]), .B(\stack[1][3] ), .Z(n13529) );
  NAND U14145 ( .A(n13528), .B(n13529), .Z(n13531) );
  XNOR U14146 ( .A(n13527), .B(n13526), .Z(n13882) );
  NAND U14147 ( .A(n13882), .B(n13883), .Z(n13530) );
  AND U14148 ( .A(n13531), .B(n13530), .Z(n13533) );
  NAND U14149 ( .A(n13532), .B(n13533), .Z(n13535) );
  NAND U14150 ( .A(\stack[1][3] ), .B(o[11]), .Z(n13888) );
  NAND U14151 ( .A(n13889), .B(n13888), .Z(n13534) );
  AND U14152 ( .A(n13535), .B(n13534), .Z(n13538) );
  AND U14153 ( .A(\stack[1][3] ), .B(o[12]), .Z(n13539) );
  NAND U14154 ( .A(n13538), .B(n13539), .Z(n13541) );
  XOR U14155 ( .A(n13537), .B(n13536), .Z(n13827) );
  NAND U14156 ( .A(n13827), .B(n13826), .Z(n13540) );
  NAND U14157 ( .A(n13541), .B(n13540), .Z(n13544) );
  NAND U14158 ( .A(n13544), .B(n13545), .Z(n13547) );
  AND U14159 ( .A(\stack[1][3] ), .B(o[13]), .Z(n13898) );
  NAND U14160 ( .A(n13898), .B(n13899), .Z(n13546) );
  NAND U14161 ( .A(n13547), .B(n13546), .Z(n13550) );
  AND U14162 ( .A(\stack[1][3] ), .B(o[14]), .Z(n13551) );
  NAND U14163 ( .A(n13550), .B(n13551), .Z(n13553) );
  XNOR U14164 ( .A(n13549), .B(n13548), .Z(n13904) );
  NAND U14165 ( .A(n13904), .B(n13905), .Z(n13552) );
  NAND U14166 ( .A(n13553), .B(n13552), .Z(n13556) );
  XNOR U14167 ( .A(n13555), .B(n13554), .Z(n13557) );
  NAND U14168 ( .A(n13556), .B(n13557), .Z(n13559) );
  AND U14169 ( .A(\stack[1][3] ), .B(o[15]), .Z(n13910) );
  NAND U14170 ( .A(n13911), .B(n13910), .Z(n13558) );
  NAND U14171 ( .A(n13559), .B(n13558), .Z(n13562) );
  AND U14172 ( .A(\stack[1][3] ), .B(o[16]), .Z(n13563) );
  NAND U14173 ( .A(n13562), .B(n13563), .Z(n13565) );
  XOR U14174 ( .A(n13561), .B(n13560), .Z(n13917) );
  NAND U14175 ( .A(n13917), .B(n13916), .Z(n13564) );
  NAND U14176 ( .A(n13565), .B(n13564), .Z(n13568) );
  XOR U14177 ( .A(n13567), .B(n13566), .Z(n13569) );
  NAND U14178 ( .A(n13568), .B(n13569), .Z(n13571) );
  AND U14179 ( .A(\stack[1][3] ), .B(o[17]), .Z(n13922) );
  NAND U14180 ( .A(n13922), .B(n13923), .Z(n13570) );
  NAND U14181 ( .A(n13571), .B(n13570), .Z(n13574) );
  AND U14182 ( .A(\stack[1][3] ), .B(o[18]), .Z(n13575) );
  NAND U14183 ( .A(n13574), .B(n13575), .Z(n13577) );
  NAND U14184 ( .A(n13929), .B(n13928), .Z(n13576) );
  NAND U14185 ( .A(n13577), .B(n13576), .Z(n13578) );
  NAND U14186 ( .A(n13579), .B(n13578), .Z(n13581) );
  AND U14187 ( .A(\stack[1][3] ), .B(o[19]), .Z(n13936) );
  XOR U14188 ( .A(n13579), .B(n13578), .Z(n13937) );
  NAND U14189 ( .A(n13936), .B(n13937), .Z(n13580) );
  NAND U14190 ( .A(n13581), .B(n13580), .Z(n13584) );
  AND U14191 ( .A(\stack[1][3] ), .B(o[20]), .Z(n13585) );
  NAND U14192 ( .A(n13584), .B(n13585), .Z(n13587) );
  XOR U14193 ( .A(n13583), .B(n13582), .Z(n13941) );
  NAND U14194 ( .A(n13941), .B(n13940), .Z(n13586) );
  NAND U14195 ( .A(n13587), .B(n13586), .Z(n13590) );
  XOR U14196 ( .A(n13589), .B(n13588), .Z(n13591) );
  NAND U14197 ( .A(n13590), .B(n13591), .Z(n13593) );
  AND U14198 ( .A(\stack[1][3] ), .B(o[21]), .Z(n13948) );
  NAND U14199 ( .A(n13948), .B(n13949), .Z(n13592) );
  NAND U14200 ( .A(n13593), .B(n13592), .Z(n13596) );
  AND U14201 ( .A(\stack[1][3] ), .B(o[22]), .Z(n13597) );
  NAND U14202 ( .A(n13596), .B(n13597), .Z(n13599) );
  NAND U14203 ( .A(n13953), .B(n13952), .Z(n13598) );
  NAND U14204 ( .A(n13599), .B(n13598), .Z(n13600) );
  NAND U14205 ( .A(n13601), .B(n13600), .Z(n13603) );
  XOR U14206 ( .A(n13601), .B(n13600), .Z(n13959) );
  AND U14207 ( .A(\stack[1][3] ), .B(o[23]), .Z(n13958) );
  NAND U14208 ( .A(n13959), .B(n13958), .Z(n13602) );
  NAND U14209 ( .A(n13603), .B(n13602), .Z(n13606) );
  AND U14210 ( .A(\stack[1][3] ), .B(o[24]), .Z(n13607) );
  NAND U14211 ( .A(n13606), .B(n13607), .Z(n13609) );
  XOR U14212 ( .A(n13605), .B(n13604), .Z(n13965) );
  NAND U14213 ( .A(n13965), .B(n13964), .Z(n13608) );
  NAND U14214 ( .A(n13609), .B(n13608), .Z(n13612) );
  XOR U14215 ( .A(n13611), .B(n13610), .Z(n13613) );
  NAND U14216 ( .A(n13612), .B(n13613), .Z(n13615) );
  AND U14217 ( .A(\stack[1][3] ), .B(o[25]), .Z(n13972) );
  NAND U14218 ( .A(n13972), .B(n13973), .Z(n13614) );
  NAND U14219 ( .A(n13615), .B(n13614), .Z(n13618) );
  AND U14220 ( .A(\stack[1][3] ), .B(o[26]), .Z(n13619) );
  NAND U14221 ( .A(n13618), .B(n13619), .Z(n13621) );
  NAND U14222 ( .A(n13977), .B(n13976), .Z(n13620) );
  NAND U14223 ( .A(n13621), .B(n13620), .Z(n13624) );
  XOR U14224 ( .A(n13623), .B(n13622), .Z(n13625) );
  NAND U14225 ( .A(n13624), .B(n13625), .Z(n13627) );
  AND U14226 ( .A(\stack[1][3] ), .B(o[27]), .Z(n13984) );
  NAND U14227 ( .A(n13984), .B(n13985), .Z(n13626) );
  NAND U14228 ( .A(n13627), .B(n13626), .Z(n13630) );
  AND U14229 ( .A(\stack[1][3] ), .B(o[28]), .Z(n13631) );
  NAND U14230 ( .A(n13630), .B(n13631), .Z(n13633) );
  NAND U14231 ( .A(n13989), .B(n13988), .Z(n13632) );
  NAND U14232 ( .A(n13633), .B(n13632), .Z(n13636) );
  XNOR U14233 ( .A(n13635), .B(n13634), .Z(n13637) );
  NAND U14234 ( .A(n13636), .B(n13637), .Z(n13639) );
  AND U14235 ( .A(\stack[1][3] ), .B(o[29]), .Z(n13994) );
  NAND U14236 ( .A(n13995), .B(n13994), .Z(n13638) );
  NAND U14237 ( .A(n13639), .B(n13638), .Z(n13642) );
  AND U14238 ( .A(\stack[1][3] ), .B(o[30]), .Z(n13643) );
  NAND U14239 ( .A(n13642), .B(n13643), .Z(n13645) );
  NAND U14240 ( .A(n14001), .B(n14000), .Z(n13644) );
  NAND U14241 ( .A(n13645), .B(n13644), .Z(n13648) );
  XOR U14242 ( .A(n13647), .B(n13646), .Z(n13649) );
  NAND U14243 ( .A(n13648), .B(n13649), .Z(n13651) );
  AND U14244 ( .A(\stack[1][3] ), .B(o[31]), .Z(n14006) );
  NAND U14245 ( .A(n14006), .B(n14007), .Z(n13650) );
  NAND U14246 ( .A(n13651), .B(n13650), .Z(n13654) );
  AND U14247 ( .A(\stack[1][3] ), .B(o[32]), .Z(n13655) );
  NAND U14248 ( .A(n13654), .B(n13655), .Z(n13657) );
  NAND U14249 ( .A(n14013), .B(n14012), .Z(n13656) );
  NAND U14250 ( .A(n13657), .B(n13656), .Z(n13660) );
  XOR U14251 ( .A(n13659), .B(n13658), .Z(n13661) );
  NAND U14252 ( .A(n13660), .B(n13661), .Z(n13663) );
  AND U14253 ( .A(\stack[1][3] ), .B(o[33]), .Z(n14020) );
  NAND U14254 ( .A(n14020), .B(n14021), .Z(n13662) );
  NAND U14255 ( .A(n13663), .B(n13662), .Z(n13666) );
  AND U14256 ( .A(\stack[1][3] ), .B(o[34]), .Z(n13667) );
  NAND U14257 ( .A(n13666), .B(n13667), .Z(n13669) );
  NAND U14258 ( .A(n14025), .B(n14024), .Z(n13668) );
  NAND U14259 ( .A(n13669), .B(n13668), .Z(n13672) );
  XOR U14260 ( .A(n13671), .B(n13670), .Z(n13673) );
  NAND U14261 ( .A(n13672), .B(n13673), .Z(n13675) );
  AND U14262 ( .A(\stack[1][3] ), .B(o[35]), .Z(n14032) );
  NAND U14263 ( .A(n14032), .B(n14033), .Z(n13674) );
  NAND U14264 ( .A(n13675), .B(n13674), .Z(n13678) );
  AND U14265 ( .A(\stack[1][3] ), .B(o[36]), .Z(n13679) );
  NAND U14266 ( .A(n13678), .B(n13679), .Z(n13681) );
  NAND U14267 ( .A(n14037), .B(n14036), .Z(n13680) );
  NAND U14268 ( .A(n13681), .B(n13680), .Z(n13684) );
  XOR U14269 ( .A(n13683), .B(n13682), .Z(n13685) );
  NAND U14270 ( .A(n13684), .B(n13685), .Z(n13687) );
  AND U14271 ( .A(\stack[1][3] ), .B(o[37]), .Z(n14042) );
  NAND U14272 ( .A(n14042), .B(n14043), .Z(n13686) );
  NAND U14273 ( .A(n13687), .B(n13686), .Z(n13690) );
  AND U14274 ( .A(\stack[1][3] ), .B(o[38]), .Z(n13691) );
  NAND U14275 ( .A(n13690), .B(n13691), .Z(n13693) );
  NAND U14276 ( .A(n14049), .B(n14048), .Z(n13692) );
  NAND U14277 ( .A(n13693), .B(n13692), .Z(n13696) );
  XNOR U14278 ( .A(n13695), .B(n13694), .Z(n13697) );
  NAND U14279 ( .A(n13696), .B(n13697), .Z(n13699) );
  AND U14280 ( .A(\stack[1][3] ), .B(o[39]), .Z(n14056) );
  NAND U14281 ( .A(n14057), .B(n14056), .Z(n13698) );
  NAND U14282 ( .A(n13699), .B(n13698), .Z(n13702) );
  AND U14283 ( .A(\stack[1][3] ), .B(o[40]), .Z(n13703) );
  NAND U14284 ( .A(n13702), .B(n13703), .Z(n13705) );
  NAND U14285 ( .A(n14061), .B(n14060), .Z(n13704) );
  NAND U14286 ( .A(n13705), .B(n13704), .Z(n13708) );
  XOR U14287 ( .A(n13707), .B(n13706), .Z(n13709) );
  NAND U14288 ( .A(n13708), .B(n13709), .Z(n13711) );
  AND U14289 ( .A(\stack[1][3] ), .B(o[41]), .Z(n14068) );
  NAND U14290 ( .A(n14068), .B(n14069), .Z(n13710) );
  NAND U14291 ( .A(n13711), .B(n13710), .Z(n13714) );
  AND U14292 ( .A(\stack[1][3] ), .B(o[42]), .Z(n13715) );
  NAND U14293 ( .A(n13714), .B(n13715), .Z(n13717) );
  XOR U14294 ( .A(n13713), .B(n13712), .Z(n14073) );
  NAND U14295 ( .A(n14073), .B(n14072), .Z(n13716) );
  NAND U14296 ( .A(n13717), .B(n13716), .Z(n13720) );
  XOR U14297 ( .A(n13719), .B(n13718), .Z(n13721) );
  NAND U14298 ( .A(n13720), .B(n13721), .Z(n13723) );
  AND U14299 ( .A(\stack[1][3] ), .B(o[43]), .Z(n14080) );
  NAND U14300 ( .A(n14080), .B(n14081), .Z(n13722) );
  NAND U14301 ( .A(n13723), .B(n13722), .Z(n13726) );
  AND U14302 ( .A(\stack[1][3] ), .B(o[44]), .Z(n13727) );
  NAND U14303 ( .A(n13726), .B(n13727), .Z(n13729) );
  XOR U14304 ( .A(n13725), .B(n13724), .Z(n14085) );
  NAND U14305 ( .A(n14085), .B(n14084), .Z(n13728) );
  NAND U14306 ( .A(n13729), .B(n13728), .Z(n13732) );
  XNOR U14307 ( .A(n13731), .B(n13730), .Z(n13733) );
  NAND U14308 ( .A(n13732), .B(n13733), .Z(n13735) );
  AND U14309 ( .A(\stack[1][3] ), .B(o[45]), .Z(n14090) );
  NAND U14310 ( .A(n14091), .B(n14090), .Z(n13734) );
  NAND U14311 ( .A(n13735), .B(n13734), .Z(n13738) );
  AND U14312 ( .A(\stack[1][3] ), .B(o[46]), .Z(n13739) );
  NAND U14313 ( .A(n13738), .B(n13739), .Z(n13741) );
  XOR U14314 ( .A(n13737), .B(n13736), .Z(n14097) );
  NAND U14315 ( .A(n14097), .B(n14096), .Z(n13740) );
  NAND U14316 ( .A(n13741), .B(n13740), .Z(n13744) );
  XOR U14317 ( .A(n13743), .B(n13742), .Z(n13745) );
  NAND U14318 ( .A(n13744), .B(n13745), .Z(n13747) );
  AND U14319 ( .A(\stack[1][3] ), .B(o[47]), .Z(n14104) );
  NAND U14320 ( .A(n14104), .B(n14105), .Z(n13746) );
  NAND U14321 ( .A(n13747), .B(n13746), .Z(n13750) );
  AND U14322 ( .A(\stack[1][3] ), .B(o[48]), .Z(n13751) );
  NAND U14323 ( .A(n13750), .B(n13751), .Z(n13753) );
  NAND U14324 ( .A(n14109), .B(n14108), .Z(n13752) );
  NAND U14325 ( .A(n13753), .B(n13752), .Z(n13754) );
  NAND U14326 ( .A(n13755), .B(n13754), .Z(n13757) );
  AND U14327 ( .A(\stack[1][3] ), .B(o[49]), .Z(n14116) );
  XOR U14328 ( .A(n13755), .B(n13754), .Z(n14117) );
  NAND U14329 ( .A(n14116), .B(n14117), .Z(n13756) );
  NAND U14330 ( .A(n13757), .B(n13756), .Z(n13760) );
  AND U14331 ( .A(\stack[1][3] ), .B(o[50]), .Z(n13761) );
  NAND U14332 ( .A(n13760), .B(n13761), .Z(n13763) );
  XOR U14333 ( .A(n13759), .B(n13758), .Z(n14121) );
  NAND U14334 ( .A(n14121), .B(n14120), .Z(n13762) );
  NAND U14335 ( .A(n13763), .B(n13762), .Z(n13766) );
  XOR U14336 ( .A(n13765), .B(n13764), .Z(n13767) );
  NAND U14337 ( .A(n13766), .B(n13767), .Z(n13769) );
  AND U14338 ( .A(\stack[1][3] ), .B(o[51]), .Z(n14128) );
  NAND U14339 ( .A(n14128), .B(n14129), .Z(n13768) );
  NAND U14340 ( .A(n13769), .B(n13768), .Z(n13772) );
  AND U14341 ( .A(\stack[1][3] ), .B(o[52]), .Z(n13773) );
  NAND U14342 ( .A(n13772), .B(n13773), .Z(n13775) );
  NAND U14343 ( .A(n14133), .B(n14132), .Z(n13774) );
  NAND U14344 ( .A(n13775), .B(n13774), .Z(n13777) );
  NAND U14345 ( .A(n13776), .B(n13777), .Z(n13779) );
  AND U14346 ( .A(\stack[1][3] ), .B(o[53]), .Z(n14140) );
  NAND U14347 ( .A(n14140), .B(n14141), .Z(n13778) );
  NAND U14348 ( .A(n13779), .B(n13778), .Z(n13782) );
  AND U14349 ( .A(\stack[1][3] ), .B(o[54]), .Z(n13783) );
  NAND U14350 ( .A(n13782), .B(n13783), .Z(n13785) );
  NAND U14351 ( .A(n14145), .B(n14144), .Z(n13784) );
  NAND U14352 ( .A(n13785), .B(n13784), .Z(n13788) );
  XOR U14353 ( .A(n13787), .B(n13786), .Z(n13789) );
  NAND U14354 ( .A(n13788), .B(n13789), .Z(n13791) );
  AND U14355 ( .A(\stack[1][3] ), .B(o[55]), .Z(n14152) );
  NAND U14356 ( .A(n14152), .B(n14153), .Z(n13790) );
  NAND U14357 ( .A(n13791), .B(n13790), .Z(n13794) );
  AND U14358 ( .A(\stack[1][3] ), .B(o[56]), .Z(n13795) );
  NAND U14359 ( .A(n13794), .B(n13795), .Z(n13797) );
  NAND U14360 ( .A(n14157), .B(n14156), .Z(n13796) );
  NAND U14361 ( .A(n13797), .B(n13796), .Z(n13800) );
  XOR U14362 ( .A(n13799), .B(n13798), .Z(n13801) );
  NAND U14363 ( .A(n13800), .B(n13801), .Z(n13803) );
  AND U14364 ( .A(\stack[1][3] ), .B(o[57]), .Z(n14162) );
  NAND U14365 ( .A(n14163), .B(n14162), .Z(n13802) );
  NAND U14366 ( .A(n13803), .B(n13802), .Z(n13806) );
  AND U14367 ( .A(\stack[1][3] ), .B(o[58]), .Z(n13807) );
  NAND U14368 ( .A(n13806), .B(n13807), .Z(n13809) );
  XOR U14369 ( .A(n13805), .B(n13804), .Z(n14169) );
  NAND U14370 ( .A(n14169), .B(n14168), .Z(n13808) );
  NAND U14371 ( .A(n13809), .B(n13808), .Z(n13810) );
  XOR U14372 ( .A(n13811), .B(n13810), .Z(n14175) );
  AND U14373 ( .A(\stack[1][3] ), .B(o[59]), .Z(n14174) );
  NAND U14374 ( .A(n14175), .B(n14174), .Z(n13813) );
  NAND U14375 ( .A(n13811), .B(n13810), .Z(n13812) );
  AND U14376 ( .A(n13813), .B(n13812), .Z(n13821) );
  NAND U14377 ( .A(n13815), .B(n13814), .Z(n13819) );
  NAND U14378 ( .A(n13817), .B(n13816), .Z(n13818) );
  NAND U14379 ( .A(n13819), .B(n13818), .Z(n13820) );
  XNOR U14380 ( .A(n13821), .B(n13820), .Z(n13822) );
  XNOR U14381 ( .A(n13823), .B(n13822), .Z(n13824) );
  XNOR U14382 ( .A(n13825), .B(n13824), .Z(n14907) );
  NAND U14383 ( .A(\stack[1][2] ), .B(o[58]), .Z(n14164) );
  NAND U14384 ( .A(\stack[1][2] ), .B(o[46]), .Z(n14092) );
  NAND U14385 ( .A(\stack[1][2] ), .B(o[40]), .Z(n14054) );
  NAND U14386 ( .A(\stack[1][2] ), .B(o[30]), .Z(n13996) );
  NAND U14387 ( .A(\stack[1][2] ), .B(o[24]), .Z(n13960) );
  NAND U14388 ( .A(\stack[1][2] ), .B(o[16]), .Z(n13912) );
  AND U14389 ( .A(\stack[1][2] ), .B(o[14]), .Z(n13900) );
  XNOR U14390 ( .A(n13827), .B(n13826), .Z(n13894) );
  XNOR U14391 ( .A(n13829), .B(n13828), .Z(n13872) );
  AND U14392 ( .A(\stack[1][2] ), .B(o[5]), .Z(n13850) );
  XOR U14393 ( .A(n13831), .B(n13830), .Z(n13851) );
  NAND U14394 ( .A(n13850), .B(n13851), .Z(n13853) );
  AND U14395 ( .A(\stack[1][2] ), .B(o[0]), .Z(n14590) );
  AND U14396 ( .A(\stack[1][3] ), .B(o[1]), .Z(n13834) );
  AND U14397 ( .A(n14590), .B(n13834), .Z(n13832) );
  NAND U14398 ( .A(o[2]), .B(n13832), .Z(n13838) );
  NAND U14399 ( .A(\stack[1][4] ), .B(o[0]), .Z(n13833) );
  XNOR U14400 ( .A(n13834), .B(n13833), .Z(n14196) );
  NAND U14401 ( .A(o[0]), .B(n13834), .Z(n13835) );
  XNOR U14402 ( .A(o[2]), .B(n13835), .Z(n13836) );
  AND U14403 ( .A(\stack[1][2] ), .B(n13836), .Z(n14197) );
  NAND U14404 ( .A(n14196), .B(n14197), .Z(n13837) );
  NAND U14405 ( .A(n13838), .B(n13837), .Z(n13841) );
  NAND U14406 ( .A(n13841), .B(n13842), .Z(n13844) );
  AND U14407 ( .A(\stack[1][2] ), .B(o[3]), .Z(n14203) );
  NAND U14408 ( .A(n14203), .B(n14202), .Z(n13843) );
  NAND U14409 ( .A(n13844), .B(n13843), .Z(n13846) );
  AND U14410 ( .A(\stack[1][2] ), .B(o[4]), .Z(n13847) );
  NAND U14411 ( .A(n13846), .B(n13847), .Z(n13849) );
  XOR U14412 ( .A(n17214), .B(n13845), .Z(n14209) );
  NAND U14413 ( .A(n14209), .B(n14208), .Z(n13848) );
  NAND U14414 ( .A(n13849), .B(n13848), .Z(n14214) );
  NAND U14415 ( .A(n14214), .B(n14215), .Z(n13852) );
  NAND U14416 ( .A(n13853), .B(n13852), .Z(n13856) );
  NAND U14417 ( .A(n13856), .B(n13857), .Z(n13859) );
  AND U14418 ( .A(\stack[1][2] ), .B(o[6]), .Z(n14221) );
  NAND U14419 ( .A(n14221), .B(n14220), .Z(n13858) );
  NAND U14420 ( .A(n13859), .B(n13858), .Z(n13862) );
  XOR U14421 ( .A(n13861), .B(n13860), .Z(n13863) );
  NAND U14422 ( .A(n13862), .B(n13863), .Z(n13865) );
  AND U14423 ( .A(\stack[1][2] ), .B(o[7]), .Z(n14226) );
  NAND U14424 ( .A(n14226), .B(n14227), .Z(n13864) );
  NAND U14425 ( .A(n13865), .B(n13864), .Z(n13868) );
  AND U14426 ( .A(\stack[1][2] ), .B(o[8]), .Z(n13869) );
  NAND U14427 ( .A(n13868), .B(n13869), .Z(n13871) );
  NAND U14428 ( .A(n14233), .B(n14232), .Z(n13870) );
  AND U14429 ( .A(n13871), .B(n13870), .Z(n13873) );
  NAND U14430 ( .A(n13872), .B(n13873), .Z(n13875) );
  NAND U14431 ( .A(\stack[1][2] ), .B(o[9]), .Z(n14238) );
  NAND U14432 ( .A(n14239), .B(n14238), .Z(n13874) );
  AND U14433 ( .A(n13875), .B(n13874), .Z(n13878) );
  AND U14434 ( .A(\stack[1][2] ), .B(o[10]), .Z(n13879) );
  NAND U14435 ( .A(n13878), .B(n13879), .Z(n13881) );
  NAND U14436 ( .A(n14187), .B(n14186), .Z(n13880) );
  NAND U14437 ( .A(n13881), .B(n13880), .Z(n13884) );
  NAND U14438 ( .A(n13884), .B(n13885), .Z(n13887) );
  AND U14439 ( .A(\stack[1][2] ), .B(o[11]), .Z(n14249) );
  NAND U14440 ( .A(n14249), .B(n14248), .Z(n13886) );
  NAND U14441 ( .A(n13887), .B(n13886), .Z(n13890) );
  AND U14442 ( .A(\stack[1][2] ), .B(o[12]), .Z(n13891) );
  NAND U14443 ( .A(n13890), .B(n13891), .Z(n13893) );
  XNOR U14444 ( .A(n13889), .B(n13888), .Z(n14254) );
  NAND U14445 ( .A(n14254), .B(n14255), .Z(n13892) );
  AND U14446 ( .A(n13893), .B(n13892), .Z(n13895) );
  NAND U14447 ( .A(n13894), .B(n13895), .Z(n13897) );
  NAND U14448 ( .A(\stack[1][2] ), .B(o[13]), .Z(n14260) );
  NAND U14449 ( .A(n14261), .B(n14260), .Z(n13896) );
  AND U14450 ( .A(n13897), .B(n13896), .Z(n13901) );
  NAND U14451 ( .A(n13900), .B(n13901), .Z(n13903) );
  NAND U14452 ( .A(n14267), .B(n14266), .Z(n13902) );
  NAND U14453 ( .A(n13903), .B(n13902), .Z(n13906) );
  NAND U14454 ( .A(n13906), .B(n13907), .Z(n13909) );
  AND U14455 ( .A(\stack[1][2] ), .B(o[15]), .Z(n14272) );
  NAND U14456 ( .A(n14272), .B(n14273), .Z(n13908) );
  AND U14457 ( .A(n13909), .B(n13908), .Z(n13913) );
  NAND U14458 ( .A(n13912), .B(n13913), .Z(n13915) );
  XNOR U14459 ( .A(n13911), .B(n13910), .Z(n14184) );
  NAND U14460 ( .A(n14184), .B(n14185), .Z(n13914) );
  AND U14461 ( .A(n13915), .B(n13914), .Z(n13919) );
  XOR U14462 ( .A(n13917), .B(n13916), .Z(n13918) );
  NAND U14463 ( .A(n13919), .B(n13918), .Z(n13921) );
  AND U14464 ( .A(\stack[1][2] ), .B(o[17]), .Z(n14282) );
  XOR U14465 ( .A(n13919), .B(n13918), .Z(n14283) );
  NAND U14466 ( .A(n14282), .B(n14283), .Z(n13920) );
  NAND U14467 ( .A(n13921), .B(n13920), .Z(n13924) );
  AND U14468 ( .A(\stack[1][2] ), .B(o[18]), .Z(n13925) );
  NAND U14469 ( .A(n13924), .B(n13925), .Z(n13927) );
  NAND U14470 ( .A(n14289), .B(n14288), .Z(n13926) );
  NAND U14471 ( .A(n13927), .B(n13926), .Z(n13930) );
  XOR U14472 ( .A(n13929), .B(n13928), .Z(n13931) );
  NAND U14473 ( .A(n13930), .B(n13931), .Z(n13933) );
  AND U14474 ( .A(\stack[1][2] ), .B(o[19]), .Z(n14295) );
  NAND U14475 ( .A(n14295), .B(n14294), .Z(n13932) );
  NAND U14476 ( .A(n13933), .B(n13932), .Z(n13934) );
  AND U14477 ( .A(\stack[1][2] ), .B(o[20]), .Z(n13935) );
  NAND U14478 ( .A(n13934), .B(n13935), .Z(n13939) );
  NAND U14479 ( .A(n14301), .B(n14300), .Z(n13938) );
  NAND U14480 ( .A(n13939), .B(n13938), .Z(n13942) );
  XOR U14481 ( .A(n13941), .B(n13940), .Z(n13943) );
  NAND U14482 ( .A(n13942), .B(n13943), .Z(n13945) );
  AND U14483 ( .A(\stack[1][2] ), .B(o[21]), .Z(n14307) );
  NAND U14484 ( .A(n14307), .B(n14306), .Z(n13944) );
  NAND U14485 ( .A(n13945), .B(n13944), .Z(n13946) );
  AND U14486 ( .A(\stack[1][2] ), .B(o[22]), .Z(n13947) );
  NAND U14487 ( .A(n13946), .B(n13947), .Z(n13951) );
  NAND U14488 ( .A(n14313), .B(n14312), .Z(n13950) );
  NAND U14489 ( .A(n13951), .B(n13950), .Z(n13954) );
  XOR U14490 ( .A(n13953), .B(n13952), .Z(n13955) );
  NAND U14491 ( .A(n13954), .B(n13955), .Z(n13957) );
  AND U14492 ( .A(\stack[1][2] ), .B(o[23]), .Z(n14318) );
  NAND U14493 ( .A(n14318), .B(n14319), .Z(n13956) );
  AND U14494 ( .A(n13957), .B(n13956), .Z(n13961) );
  NAND U14495 ( .A(n13960), .B(n13961), .Z(n13963) );
  XNOR U14496 ( .A(n13959), .B(n13958), .Z(n14182) );
  NAND U14497 ( .A(n14182), .B(n14183), .Z(n13962) );
  AND U14498 ( .A(n13963), .B(n13962), .Z(n13967) );
  XOR U14499 ( .A(n13965), .B(n13964), .Z(n13966) );
  NAND U14500 ( .A(n13967), .B(n13966), .Z(n13969) );
  AND U14501 ( .A(\stack[1][2] ), .B(o[25]), .Z(n14328) );
  XOR U14502 ( .A(n13967), .B(n13966), .Z(n14329) );
  NAND U14503 ( .A(n14328), .B(n14329), .Z(n13968) );
  NAND U14504 ( .A(n13969), .B(n13968), .Z(n13970) );
  AND U14505 ( .A(\stack[1][2] ), .B(o[26]), .Z(n13971) );
  NAND U14506 ( .A(n13970), .B(n13971), .Z(n13975) );
  NAND U14507 ( .A(n14335), .B(n14334), .Z(n13974) );
  NAND U14508 ( .A(n13975), .B(n13974), .Z(n13978) );
  XOR U14509 ( .A(n13977), .B(n13976), .Z(n13979) );
  NAND U14510 ( .A(n13978), .B(n13979), .Z(n13981) );
  AND U14511 ( .A(\stack[1][2] ), .B(o[27]), .Z(n14341) );
  NAND U14512 ( .A(n14341), .B(n14340), .Z(n13980) );
  NAND U14513 ( .A(n13981), .B(n13980), .Z(n13982) );
  AND U14514 ( .A(\stack[1][2] ), .B(o[28]), .Z(n13983) );
  NAND U14515 ( .A(n13982), .B(n13983), .Z(n13987) );
  NAND U14516 ( .A(n14347), .B(n14346), .Z(n13986) );
  NAND U14517 ( .A(n13987), .B(n13986), .Z(n13990) );
  XOR U14518 ( .A(n13989), .B(n13988), .Z(n13991) );
  NAND U14519 ( .A(n13990), .B(n13991), .Z(n13993) );
  AND U14520 ( .A(\stack[1][2] ), .B(o[29]), .Z(n14352) );
  NAND U14521 ( .A(n14352), .B(n14353), .Z(n13992) );
  AND U14522 ( .A(n13993), .B(n13992), .Z(n13997) );
  NAND U14523 ( .A(n13996), .B(n13997), .Z(n13999) );
  XNOR U14524 ( .A(n13995), .B(n13994), .Z(n14180) );
  NAND U14525 ( .A(n14180), .B(n14181), .Z(n13998) );
  AND U14526 ( .A(n13999), .B(n13998), .Z(n14003) );
  XOR U14527 ( .A(n14001), .B(n14000), .Z(n14002) );
  NAND U14528 ( .A(n14003), .B(n14002), .Z(n14005) );
  AND U14529 ( .A(\stack[1][2] ), .B(o[31]), .Z(n14362) );
  XOR U14530 ( .A(n14003), .B(n14002), .Z(n14363) );
  NAND U14531 ( .A(n14362), .B(n14363), .Z(n14004) );
  NAND U14532 ( .A(n14005), .B(n14004), .Z(n14008) );
  AND U14533 ( .A(\stack[1][2] ), .B(o[32]), .Z(n14009) );
  NAND U14534 ( .A(n14008), .B(n14009), .Z(n14011) );
  NAND U14535 ( .A(n14369), .B(n14368), .Z(n14010) );
  NAND U14536 ( .A(n14011), .B(n14010), .Z(n14014) );
  XOR U14537 ( .A(n14013), .B(n14012), .Z(n14015) );
  NAND U14538 ( .A(n14014), .B(n14015), .Z(n14017) );
  AND U14539 ( .A(\stack[1][2] ), .B(o[33]), .Z(n14375) );
  NAND U14540 ( .A(n14375), .B(n14374), .Z(n14016) );
  NAND U14541 ( .A(n14017), .B(n14016), .Z(n14018) );
  AND U14542 ( .A(\stack[1][2] ), .B(o[34]), .Z(n14019) );
  NAND U14543 ( .A(n14018), .B(n14019), .Z(n14023) );
  NAND U14544 ( .A(n14381), .B(n14380), .Z(n14022) );
  NAND U14545 ( .A(n14023), .B(n14022), .Z(n14026) );
  XOR U14546 ( .A(n14025), .B(n14024), .Z(n14027) );
  NAND U14547 ( .A(n14026), .B(n14027), .Z(n14029) );
  AND U14548 ( .A(\stack[1][2] ), .B(o[35]), .Z(n14387) );
  NAND U14549 ( .A(n14387), .B(n14386), .Z(n14028) );
  NAND U14550 ( .A(n14029), .B(n14028), .Z(n14030) );
  AND U14551 ( .A(\stack[1][2] ), .B(o[36]), .Z(n14031) );
  NAND U14552 ( .A(n14030), .B(n14031), .Z(n14035) );
  NAND U14553 ( .A(n14393), .B(n14392), .Z(n14034) );
  NAND U14554 ( .A(n14035), .B(n14034), .Z(n14038) );
  XOR U14555 ( .A(n14037), .B(n14036), .Z(n14039) );
  NAND U14556 ( .A(n14038), .B(n14039), .Z(n14041) );
  AND U14557 ( .A(\stack[1][2] ), .B(o[37]), .Z(n14398) );
  NAND U14558 ( .A(n14398), .B(n14399), .Z(n14040) );
  NAND U14559 ( .A(n14041), .B(n14040), .Z(n14044) );
  AND U14560 ( .A(\stack[1][2] ), .B(o[38]), .Z(n14045) );
  NAND U14561 ( .A(n14044), .B(n14045), .Z(n14047) );
  NAND U14562 ( .A(n14405), .B(n14404), .Z(n14046) );
  NAND U14563 ( .A(n14047), .B(n14046), .Z(n14050) );
  XOR U14564 ( .A(n14049), .B(n14048), .Z(n14051) );
  NAND U14565 ( .A(n14050), .B(n14051), .Z(n14053) );
  AND U14566 ( .A(\stack[1][2] ), .B(o[39]), .Z(n14411) );
  NAND U14567 ( .A(n14411), .B(n14410), .Z(n14052) );
  AND U14568 ( .A(n14053), .B(n14052), .Z(n14055) );
  NAND U14569 ( .A(n14054), .B(n14055), .Z(n14059) );
  XNOR U14570 ( .A(n14057), .B(n14056), .Z(n14416) );
  NAND U14571 ( .A(n14417), .B(n14416), .Z(n14058) );
  AND U14572 ( .A(n14059), .B(n14058), .Z(n14063) );
  XOR U14573 ( .A(n14061), .B(n14060), .Z(n14062) );
  NAND U14574 ( .A(n14063), .B(n14062), .Z(n14065) );
  AND U14575 ( .A(\stack[1][2] ), .B(o[41]), .Z(n14422) );
  XOR U14576 ( .A(n14063), .B(n14062), .Z(n14423) );
  NAND U14577 ( .A(n14422), .B(n14423), .Z(n14064) );
  NAND U14578 ( .A(n14065), .B(n14064), .Z(n14066) );
  AND U14579 ( .A(\stack[1][2] ), .B(o[42]), .Z(n14067) );
  NAND U14580 ( .A(n14066), .B(n14067), .Z(n14071) );
  NAND U14581 ( .A(n14429), .B(n14428), .Z(n14070) );
  NAND U14582 ( .A(n14071), .B(n14070), .Z(n14074) );
  XOR U14583 ( .A(n14073), .B(n14072), .Z(n14075) );
  NAND U14584 ( .A(n14074), .B(n14075), .Z(n14077) );
  AND U14585 ( .A(\stack[1][2] ), .B(o[43]), .Z(n14434) );
  NAND U14586 ( .A(n14434), .B(n14435), .Z(n14076) );
  NAND U14587 ( .A(n14077), .B(n14076), .Z(n14078) );
  AND U14588 ( .A(\stack[1][2] ), .B(o[44]), .Z(n14079) );
  NAND U14589 ( .A(n14078), .B(n14079), .Z(n14083) );
  NAND U14590 ( .A(n14441), .B(n14440), .Z(n14082) );
  NAND U14591 ( .A(n14083), .B(n14082), .Z(n14086) );
  XOR U14592 ( .A(n14085), .B(n14084), .Z(n14087) );
  NAND U14593 ( .A(n14086), .B(n14087), .Z(n14089) );
  AND U14594 ( .A(\stack[1][2] ), .B(o[45]), .Z(n14447) );
  NAND U14595 ( .A(n14447), .B(n14446), .Z(n14088) );
  AND U14596 ( .A(n14089), .B(n14088), .Z(n14093) );
  NAND U14597 ( .A(n14092), .B(n14093), .Z(n14095) );
  XNOR U14598 ( .A(n14091), .B(n14090), .Z(n14178) );
  NAND U14599 ( .A(n14178), .B(n14179), .Z(n14094) );
  AND U14600 ( .A(n14095), .B(n14094), .Z(n14099) );
  XOR U14601 ( .A(n14097), .B(n14096), .Z(n14098) );
  NAND U14602 ( .A(n14099), .B(n14098), .Z(n14101) );
  AND U14603 ( .A(\stack[1][2] ), .B(o[47]), .Z(n14457) );
  XOR U14604 ( .A(n14099), .B(n14098), .Z(n14456) );
  NAND U14605 ( .A(n14457), .B(n14456), .Z(n14100) );
  NAND U14606 ( .A(n14101), .B(n14100), .Z(n14102) );
  AND U14607 ( .A(\stack[1][2] ), .B(o[48]), .Z(n14103) );
  NAND U14608 ( .A(n14102), .B(n14103), .Z(n14107) );
  NAND U14609 ( .A(n14463), .B(n14462), .Z(n14106) );
  NAND U14610 ( .A(n14107), .B(n14106), .Z(n14110) );
  XOR U14611 ( .A(n14109), .B(n14108), .Z(n14111) );
  NAND U14612 ( .A(n14110), .B(n14111), .Z(n14113) );
  AND U14613 ( .A(\stack[1][2] ), .B(o[49]), .Z(n14468) );
  NAND U14614 ( .A(n14468), .B(n14469), .Z(n14112) );
  NAND U14615 ( .A(n14113), .B(n14112), .Z(n14114) );
  AND U14616 ( .A(\stack[1][2] ), .B(o[50]), .Z(n14115) );
  NAND U14617 ( .A(n14114), .B(n14115), .Z(n14119) );
  NAND U14618 ( .A(n14475), .B(n14474), .Z(n14118) );
  NAND U14619 ( .A(n14119), .B(n14118), .Z(n14122) );
  XOR U14620 ( .A(n14121), .B(n14120), .Z(n14123) );
  NAND U14621 ( .A(n14122), .B(n14123), .Z(n14125) );
  AND U14622 ( .A(\stack[1][2] ), .B(o[51]), .Z(n14481) );
  NAND U14623 ( .A(n14481), .B(n14480), .Z(n14124) );
  NAND U14624 ( .A(n14125), .B(n14124), .Z(n14126) );
  AND U14625 ( .A(\stack[1][2] ), .B(o[52]), .Z(n14127) );
  NAND U14626 ( .A(n14126), .B(n14127), .Z(n14131) );
  NAND U14627 ( .A(n14487), .B(n14486), .Z(n14130) );
  NAND U14628 ( .A(n14131), .B(n14130), .Z(n14134) );
  XOR U14629 ( .A(n14133), .B(n14132), .Z(n14135) );
  NAND U14630 ( .A(n14134), .B(n14135), .Z(n14137) );
  AND U14631 ( .A(\stack[1][2] ), .B(o[53]), .Z(n14492) );
  NAND U14632 ( .A(n14492), .B(n14493), .Z(n14136) );
  NAND U14633 ( .A(n14137), .B(n14136), .Z(n14138) );
  AND U14634 ( .A(\stack[1][2] ), .B(o[54]), .Z(n14139) );
  NAND U14635 ( .A(n14138), .B(n14139), .Z(n14143) );
  NAND U14636 ( .A(n14499), .B(n14498), .Z(n14142) );
  NAND U14637 ( .A(n14143), .B(n14142), .Z(n14146) );
  XOR U14638 ( .A(n14145), .B(n14144), .Z(n14147) );
  NAND U14639 ( .A(n14146), .B(n14147), .Z(n14149) );
  AND U14640 ( .A(\stack[1][2] ), .B(o[55]), .Z(n14505) );
  NAND U14641 ( .A(n14505), .B(n14504), .Z(n14148) );
  NAND U14642 ( .A(n14149), .B(n14148), .Z(n14150) );
  AND U14643 ( .A(\stack[1][2] ), .B(o[56]), .Z(n14151) );
  NAND U14644 ( .A(n14150), .B(n14151), .Z(n14155) );
  NAND U14645 ( .A(n14511), .B(n14510), .Z(n14154) );
  NAND U14646 ( .A(n14155), .B(n14154), .Z(n14158) );
  XOR U14647 ( .A(n14157), .B(n14156), .Z(n14159) );
  NAND U14648 ( .A(n14158), .B(n14159), .Z(n14161) );
  AND U14649 ( .A(\stack[1][2] ), .B(o[57]), .Z(n14516) );
  NAND U14650 ( .A(n14516), .B(n14517), .Z(n14160) );
  AND U14651 ( .A(n14161), .B(n14160), .Z(n14165) );
  NAND U14652 ( .A(n14164), .B(n14165), .Z(n14167) );
  XNOR U14653 ( .A(n14163), .B(n14162), .Z(n14176) );
  NAND U14654 ( .A(n14176), .B(n14177), .Z(n14166) );
  AND U14655 ( .A(n14167), .B(n14166), .Z(n14171) );
  XOR U14656 ( .A(n14169), .B(n14168), .Z(n14170) );
  NAND U14657 ( .A(n14171), .B(n14170), .Z(n14173) );
  AND U14658 ( .A(\stack[1][2] ), .B(o[59]), .Z(n14527) );
  XOR U14659 ( .A(n14171), .B(n14170), .Z(n14526) );
  NAND U14660 ( .A(n14527), .B(n14526), .Z(n14172) );
  AND U14661 ( .A(n14173), .B(n14172), .Z(n14913) );
  NAND U14662 ( .A(\stack[1][2] ), .B(o[60]), .Z(n14912) );
  XOR U14663 ( .A(n14913), .B(n14912), .Z(n14911) );
  XNOR U14664 ( .A(n14175), .B(n14174), .Z(n14910) );
  XNOR U14665 ( .A(n14911), .B(n14910), .Z(n14901) );
  XNOR U14666 ( .A(n14187), .B(n14186), .Z(n14244) );
  AND U14667 ( .A(o[0]), .B(\stack[1][1] ), .Z(n17292) );
  AND U14668 ( .A(\stack[1][2] ), .B(o[1]), .Z(n14191) );
  AND U14669 ( .A(n17292), .B(n14191), .Z(n14188) );
  NAND U14670 ( .A(o[2]), .B(n14188), .Z(n14195) );
  NAND U14671 ( .A(o[1]), .B(\stack[1][2] ), .Z(n14189) );
  XNOR U14672 ( .A(n14190), .B(n14189), .Z(n14597) );
  NAND U14673 ( .A(n14191), .B(o[0]), .Z(n14192) );
  XNOR U14674 ( .A(o[2]), .B(n14192), .Z(n14193) );
  AND U14675 ( .A(\stack[1][1] ), .B(n14193), .Z(n14596) );
  NAND U14676 ( .A(n14597), .B(n14596), .Z(n14194) );
  NAND U14677 ( .A(n14195), .B(n14194), .Z(n14198) );
  NAND U14678 ( .A(n14198), .B(n14199), .Z(n14201) );
  AND U14679 ( .A(o[3]), .B(\stack[1][1] ), .Z(n14584) );
  NAND U14680 ( .A(n14585), .B(n14584), .Z(n14200) );
  NAND U14681 ( .A(n14201), .B(n14200), .Z(n14204) );
  AND U14682 ( .A(o[4]), .B(\stack[1][1] ), .Z(n14205) );
  NAND U14683 ( .A(n14204), .B(n14205), .Z(n14207) );
  XOR U14684 ( .A(n14203), .B(n14202), .Z(n14607) );
  NAND U14685 ( .A(n14607), .B(n14606), .Z(n14206) );
  NAND U14686 ( .A(n14207), .B(n14206), .Z(n14210) );
  XOR U14687 ( .A(n14209), .B(n14208), .Z(n14211) );
  NAND U14688 ( .A(n14210), .B(n14211), .Z(n14213) );
  AND U14689 ( .A(o[5]), .B(\stack[1][1] ), .Z(n14582) );
  NAND U14690 ( .A(n14583), .B(n14582), .Z(n14212) );
  NAND U14691 ( .A(n14213), .B(n14212), .Z(n14216) );
  NAND U14692 ( .A(n14216), .B(n14217), .Z(n14219) );
  AND U14693 ( .A(o[6]), .B(\stack[1][1] ), .Z(n14617) );
  NAND U14694 ( .A(n14617), .B(n14616), .Z(n14218) );
  NAND U14695 ( .A(n14219), .B(n14218), .Z(n14222) );
  XOR U14696 ( .A(n14221), .B(n14220), .Z(n14223) );
  NAND U14697 ( .A(n14222), .B(n14223), .Z(n14225) );
  AND U14698 ( .A(o[7]), .B(\stack[1][1] ), .Z(n14620) );
  NAND U14699 ( .A(n14621), .B(n14620), .Z(n14224) );
  NAND U14700 ( .A(n14225), .B(n14224), .Z(n14228) );
  AND U14701 ( .A(o[8]), .B(\stack[1][1] ), .Z(n14229) );
  NAND U14702 ( .A(n14228), .B(n14229), .Z(n14231) );
  NAND U14703 ( .A(n14629), .B(n14628), .Z(n14230) );
  NAND U14704 ( .A(n14231), .B(n14230), .Z(n14234) );
  XOR U14705 ( .A(n14233), .B(n14232), .Z(n14235) );
  NAND U14706 ( .A(n14234), .B(n14235), .Z(n14237) );
  AND U14707 ( .A(o[9]), .B(\stack[1][1] ), .Z(n14580) );
  NAND U14708 ( .A(n14581), .B(n14580), .Z(n14236) );
  NAND U14709 ( .A(n14237), .B(n14236), .Z(n14240) );
  AND U14710 ( .A(o[10]), .B(\stack[1][1] ), .Z(n14241) );
  NAND U14711 ( .A(n14240), .B(n14241), .Z(n14243) );
  XOR U14712 ( .A(n14239), .B(n14238), .Z(n14639) );
  NANDN U14713 ( .A(n14639), .B(n14638), .Z(n14242) );
  AND U14714 ( .A(n14243), .B(n14242), .Z(n14245) );
  NAND U14715 ( .A(n14244), .B(n14245), .Z(n14247) );
  NAND U14716 ( .A(o[11]), .B(\stack[1][1] ), .Z(n14642) );
  NAND U14717 ( .A(n14642), .B(n14643), .Z(n14246) );
  AND U14718 ( .A(n14247), .B(n14246), .Z(n14250) );
  AND U14719 ( .A(o[12]), .B(\stack[1][1] ), .Z(n14251) );
  NAND U14720 ( .A(n14250), .B(n14251), .Z(n14253) );
  XOR U14721 ( .A(n14249), .B(n14248), .Z(n14651) );
  NAND U14722 ( .A(n14651), .B(n14650), .Z(n14252) );
  NAND U14723 ( .A(n14253), .B(n14252), .Z(n14256) );
  NAND U14724 ( .A(n14256), .B(n14257), .Z(n14259) );
  AND U14725 ( .A(o[13]), .B(\stack[1][1] ), .Z(n14578) );
  NAND U14726 ( .A(n14579), .B(n14578), .Z(n14258) );
  NAND U14727 ( .A(n14259), .B(n14258), .Z(n14262) );
  AND U14728 ( .A(o[14]), .B(\stack[1][1] ), .Z(n14263) );
  NAND U14729 ( .A(n14262), .B(n14263), .Z(n14265) );
  XOR U14730 ( .A(n14261), .B(n14260), .Z(n14661) );
  NANDN U14731 ( .A(n14661), .B(n14660), .Z(n14264) );
  NAND U14732 ( .A(n14265), .B(n14264), .Z(n14268) );
  XOR U14733 ( .A(n14267), .B(n14266), .Z(n14269) );
  NAND U14734 ( .A(n14268), .B(n14269), .Z(n14271) );
  AND U14735 ( .A(o[15]), .B(\stack[1][1] ), .Z(n14576) );
  NAND U14736 ( .A(n14577), .B(n14576), .Z(n14270) );
  NAND U14737 ( .A(n14271), .B(n14270), .Z(n14274) );
  AND U14738 ( .A(o[16]), .B(\stack[1][1] ), .Z(n14275) );
  NAND U14739 ( .A(n14274), .B(n14275), .Z(n14277) );
  NAND U14740 ( .A(n14671), .B(n14670), .Z(n14276) );
  NAND U14741 ( .A(n14277), .B(n14276), .Z(n14278) );
  NAND U14742 ( .A(n14279), .B(n14278), .Z(n14281) );
  XOR U14743 ( .A(n14279), .B(n14278), .Z(n14575) );
  AND U14744 ( .A(o[17]), .B(\stack[1][1] ), .Z(n14574) );
  NAND U14745 ( .A(n14575), .B(n14574), .Z(n14280) );
  NAND U14746 ( .A(n14281), .B(n14280), .Z(n14284) );
  AND U14747 ( .A(o[18]), .B(\stack[1][1] ), .Z(n14285) );
  NAND U14748 ( .A(n14284), .B(n14285), .Z(n14287) );
  NAND U14749 ( .A(n14681), .B(n14680), .Z(n14286) );
  NAND U14750 ( .A(n14287), .B(n14286), .Z(n14290) );
  XOR U14751 ( .A(n14289), .B(n14288), .Z(n14291) );
  NAND U14752 ( .A(n14290), .B(n14291), .Z(n14293) );
  AND U14753 ( .A(o[19]), .B(\stack[1][1] ), .Z(n14572) );
  NAND U14754 ( .A(n14573), .B(n14572), .Z(n14292) );
  NAND U14755 ( .A(n14293), .B(n14292), .Z(n14296) );
  AND U14756 ( .A(o[20]), .B(\stack[1][1] ), .Z(n14297) );
  NAND U14757 ( .A(n14296), .B(n14297), .Z(n14299) );
  XOR U14758 ( .A(n14295), .B(n14294), .Z(n14691) );
  NAND U14759 ( .A(n14691), .B(n14690), .Z(n14298) );
  NAND U14760 ( .A(n14299), .B(n14298), .Z(n14302) );
  XOR U14761 ( .A(n14301), .B(n14300), .Z(n14303) );
  NAND U14762 ( .A(n14302), .B(n14303), .Z(n14305) );
  AND U14763 ( .A(o[21]), .B(\stack[1][1] ), .Z(n14570) );
  NAND U14764 ( .A(n14571), .B(n14570), .Z(n14304) );
  NAND U14765 ( .A(n14305), .B(n14304), .Z(n14308) );
  AND U14766 ( .A(o[22]), .B(\stack[1][1] ), .Z(n14309) );
  NAND U14767 ( .A(n14308), .B(n14309), .Z(n14311) );
  XOR U14768 ( .A(n14307), .B(n14306), .Z(n14701) );
  NAND U14769 ( .A(n14701), .B(n14700), .Z(n14310) );
  NAND U14770 ( .A(n14311), .B(n14310), .Z(n14314) );
  XOR U14771 ( .A(n14313), .B(n14312), .Z(n14315) );
  NAND U14772 ( .A(n14314), .B(n14315), .Z(n14317) );
  AND U14773 ( .A(o[23]), .B(\stack[1][1] ), .Z(n14568) );
  NAND U14774 ( .A(n14569), .B(n14568), .Z(n14316) );
  NAND U14775 ( .A(n14317), .B(n14316), .Z(n14320) );
  AND U14776 ( .A(o[24]), .B(\stack[1][1] ), .Z(n14321) );
  NAND U14777 ( .A(n14320), .B(n14321), .Z(n14323) );
  NAND U14778 ( .A(n14711), .B(n14710), .Z(n14322) );
  NAND U14779 ( .A(n14323), .B(n14322), .Z(n14324) );
  NAND U14780 ( .A(n14325), .B(n14324), .Z(n14327) );
  XOR U14781 ( .A(n14325), .B(n14324), .Z(n14567) );
  AND U14782 ( .A(o[25]), .B(\stack[1][1] ), .Z(n14566) );
  NAND U14783 ( .A(n14567), .B(n14566), .Z(n14326) );
  NAND U14784 ( .A(n14327), .B(n14326), .Z(n14330) );
  AND U14785 ( .A(o[26]), .B(\stack[1][1] ), .Z(n14331) );
  NAND U14786 ( .A(n14330), .B(n14331), .Z(n14333) );
  NAND U14787 ( .A(n14721), .B(n14720), .Z(n14332) );
  NAND U14788 ( .A(n14333), .B(n14332), .Z(n14336) );
  XOR U14789 ( .A(n14335), .B(n14334), .Z(n14337) );
  NAND U14790 ( .A(n14336), .B(n14337), .Z(n14339) );
  AND U14791 ( .A(o[27]), .B(\stack[1][1] ), .Z(n14564) );
  NAND U14792 ( .A(n14565), .B(n14564), .Z(n14338) );
  NAND U14793 ( .A(n14339), .B(n14338), .Z(n14342) );
  AND U14794 ( .A(o[28]), .B(\stack[1][1] ), .Z(n14343) );
  NAND U14795 ( .A(n14342), .B(n14343), .Z(n14345) );
  XOR U14796 ( .A(n14341), .B(n14340), .Z(n14731) );
  NAND U14797 ( .A(n14731), .B(n14730), .Z(n14344) );
  NAND U14798 ( .A(n14345), .B(n14344), .Z(n14348) );
  XOR U14799 ( .A(n14347), .B(n14346), .Z(n14349) );
  NAND U14800 ( .A(n14348), .B(n14349), .Z(n14351) );
  AND U14801 ( .A(o[29]), .B(\stack[1][1] ), .Z(n14562) );
  NAND U14802 ( .A(n14563), .B(n14562), .Z(n14350) );
  NAND U14803 ( .A(n14351), .B(n14350), .Z(n14354) );
  AND U14804 ( .A(o[30]), .B(\stack[1][1] ), .Z(n14355) );
  NAND U14805 ( .A(n14354), .B(n14355), .Z(n14357) );
  NAND U14806 ( .A(n14741), .B(n14740), .Z(n14356) );
  NAND U14807 ( .A(n14357), .B(n14356), .Z(n14358) );
  NAND U14808 ( .A(n14359), .B(n14358), .Z(n14361) );
  XOR U14809 ( .A(n14359), .B(n14358), .Z(n14561) );
  AND U14810 ( .A(o[31]), .B(\stack[1][1] ), .Z(n14560) );
  NAND U14811 ( .A(n14561), .B(n14560), .Z(n14360) );
  NAND U14812 ( .A(n14361), .B(n14360), .Z(n14364) );
  AND U14813 ( .A(o[32]), .B(\stack[1][1] ), .Z(n14365) );
  NAND U14814 ( .A(n14364), .B(n14365), .Z(n14367) );
  NAND U14815 ( .A(n14751), .B(n14750), .Z(n14366) );
  NAND U14816 ( .A(n14367), .B(n14366), .Z(n14370) );
  XOR U14817 ( .A(n14369), .B(n14368), .Z(n14371) );
  NAND U14818 ( .A(n14370), .B(n14371), .Z(n14373) );
  AND U14819 ( .A(o[33]), .B(\stack[1][1] ), .Z(n14558) );
  NAND U14820 ( .A(n14559), .B(n14558), .Z(n14372) );
  NAND U14821 ( .A(n14373), .B(n14372), .Z(n14376) );
  AND U14822 ( .A(o[34]), .B(\stack[1][1] ), .Z(n14377) );
  NAND U14823 ( .A(n14376), .B(n14377), .Z(n14379) );
  XOR U14824 ( .A(n14375), .B(n14374), .Z(n14761) );
  NAND U14825 ( .A(n14761), .B(n14760), .Z(n14378) );
  NAND U14826 ( .A(n14379), .B(n14378), .Z(n14382) );
  XOR U14827 ( .A(n14381), .B(n14380), .Z(n14383) );
  NAND U14828 ( .A(n14382), .B(n14383), .Z(n14385) );
  AND U14829 ( .A(o[35]), .B(\stack[1][1] ), .Z(n14556) );
  NAND U14830 ( .A(n14557), .B(n14556), .Z(n14384) );
  NAND U14831 ( .A(n14385), .B(n14384), .Z(n14388) );
  AND U14832 ( .A(o[36]), .B(\stack[1][1] ), .Z(n14389) );
  NAND U14833 ( .A(n14388), .B(n14389), .Z(n14391) );
  XOR U14834 ( .A(n14387), .B(n14386), .Z(n14771) );
  NAND U14835 ( .A(n14771), .B(n14770), .Z(n14390) );
  NAND U14836 ( .A(n14391), .B(n14390), .Z(n14394) );
  XOR U14837 ( .A(n14393), .B(n14392), .Z(n14395) );
  NAND U14838 ( .A(n14394), .B(n14395), .Z(n14397) );
  AND U14839 ( .A(o[37]), .B(\stack[1][1] ), .Z(n14554) );
  NAND U14840 ( .A(n14555), .B(n14554), .Z(n14396) );
  NAND U14841 ( .A(n14397), .B(n14396), .Z(n14400) );
  AND U14842 ( .A(o[38]), .B(\stack[1][1] ), .Z(n14401) );
  NAND U14843 ( .A(n14400), .B(n14401), .Z(n14403) );
  NAND U14844 ( .A(n14781), .B(n14780), .Z(n14402) );
  NAND U14845 ( .A(n14403), .B(n14402), .Z(n14406) );
  XOR U14846 ( .A(n14405), .B(n14404), .Z(n14407) );
  NAND U14847 ( .A(n14406), .B(n14407), .Z(n14409) );
  AND U14848 ( .A(o[39]), .B(\stack[1][1] ), .Z(n14552) );
  NAND U14849 ( .A(n14553), .B(n14552), .Z(n14408) );
  NAND U14850 ( .A(n14409), .B(n14408), .Z(n14412) );
  AND U14851 ( .A(o[40]), .B(\stack[1][1] ), .Z(n14413) );
  NAND U14852 ( .A(n14412), .B(n14413), .Z(n14415) );
  XOR U14853 ( .A(n14411), .B(n14410), .Z(n14791) );
  NAND U14854 ( .A(n14791), .B(n14790), .Z(n14414) );
  NAND U14855 ( .A(n14415), .B(n14414), .Z(n14418) );
  XNOR U14856 ( .A(n14417), .B(n14416), .Z(n14419) );
  NAND U14857 ( .A(n14418), .B(n14419), .Z(n14421) );
  AND U14858 ( .A(o[41]), .B(\stack[1][1] ), .Z(n14550) );
  NAND U14859 ( .A(n14551), .B(n14550), .Z(n14420) );
  NAND U14860 ( .A(n14421), .B(n14420), .Z(n14424) );
  AND U14861 ( .A(o[42]), .B(\stack[1][1] ), .Z(n14425) );
  NAND U14862 ( .A(n14424), .B(n14425), .Z(n14427) );
  NAND U14863 ( .A(n14801), .B(n14800), .Z(n14426) );
  NAND U14864 ( .A(n14427), .B(n14426), .Z(n14430) );
  XOR U14865 ( .A(n14429), .B(n14428), .Z(n14431) );
  NAND U14866 ( .A(n14430), .B(n14431), .Z(n14433) );
  AND U14867 ( .A(o[43]), .B(\stack[1][1] ), .Z(n14548) );
  NAND U14868 ( .A(n14549), .B(n14548), .Z(n14432) );
  NAND U14869 ( .A(n14433), .B(n14432), .Z(n14436) );
  AND U14870 ( .A(o[44]), .B(\stack[1][1] ), .Z(n14437) );
  NAND U14871 ( .A(n14436), .B(n14437), .Z(n14439) );
  NAND U14872 ( .A(n14811), .B(n14810), .Z(n14438) );
  NAND U14873 ( .A(n14439), .B(n14438), .Z(n14442) );
  XOR U14874 ( .A(n14441), .B(n14440), .Z(n14443) );
  NAND U14875 ( .A(n14442), .B(n14443), .Z(n14445) );
  AND U14876 ( .A(o[45]), .B(\stack[1][1] ), .Z(n14546) );
  NAND U14877 ( .A(n14547), .B(n14546), .Z(n14444) );
  NAND U14878 ( .A(n14445), .B(n14444), .Z(n14448) );
  AND U14879 ( .A(o[46]), .B(\stack[1][1] ), .Z(n14449) );
  NAND U14880 ( .A(n14448), .B(n14449), .Z(n14451) );
  XOR U14881 ( .A(n14447), .B(n14446), .Z(n14821) );
  NAND U14882 ( .A(n14821), .B(n14820), .Z(n14450) );
  NAND U14883 ( .A(n14451), .B(n14450), .Z(n14452) );
  NAND U14884 ( .A(n14453), .B(n14452), .Z(n14455) );
  XOR U14885 ( .A(n14453), .B(n14452), .Z(n14545) );
  AND U14886 ( .A(o[47]), .B(\stack[1][1] ), .Z(n14544) );
  NAND U14887 ( .A(n14545), .B(n14544), .Z(n14454) );
  NAND U14888 ( .A(n14455), .B(n14454), .Z(n14458) );
  AND U14889 ( .A(o[48]), .B(\stack[1][1] ), .Z(n14459) );
  NAND U14890 ( .A(n14458), .B(n14459), .Z(n14461) );
  XOR U14891 ( .A(n14457), .B(n14456), .Z(n14831) );
  NAND U14892 ( .A(n14831), .B(n14830), .Z(n14460) );
  NAND U14893 ( .A(n14461), .B(n14460), .Z(n14464) );
  XOR U14894 ( .A(n14463), .B(n14462), .Z(n14465) );
  NAND U14895 ( .A(n14464), .B(n14465), .Z(n14467) );
  AND U14896 ( .A(o[49]), .B(\stack[1][1] ), .Z(n14542) );
  NAND U14897 ( .A(n14543), .B(n14542), .Z(n14466) );
  NAND U14898 ( .A(n14467), .B(n14466), .Z(n14470) );
  AND U14899 ( .A(o[50]), .B(\stack[1][1] ), .Z(n14471) );
  NAND U14900 ( .A(n14470), .B(n14471), .Z(n14473) );
  NAND U14901 ( .A(n14841), .B(n14840), .Z(n14472) );
  NAND U14902 ( .A(n14473), .B(n14472), .Z(n14476) );
  XOR U14903 ( .A(n14475), .B(n14474), .Z(n14477) );
  NAND U14904 ( .A(n14476), .B(n14477), .Z(n14479) );
  AND U14905 ( .A(o[51]), .B(\stack[1][1] ), .Z(n14540) );
  NAND U14906 ( .A(n14541), .B(n14540), .Z(n14478) );
  NAND U14907 ( .A(n14479), .B(n14478), .Z(n14482) );
  AND U14908 ( .A(o[52]), .B(\stack[1][1] ), .Z(n14483) );
  NAND U14909 ( .A(n14482), .B(n14483), .Z(n14485) );
  XOR U14910 ( .A(n14481), .B(n14480), .Z(n14851) );
  NAND U14911 ( .A(n14851), .B(n14850), .Z(n14484) );
  NAND U14912 ( .A(n14485), .B(n14484), .Z(n14488) );
  XOR U14913 ( .A(n14487), .B(n14486), .Z(n14489) );
  NAND U14914 ( .A(n14488), .B(n14489), .Z(n14491) );
  AND U14915 ( .A(o[53]), .B(\stack[1][1] ), .Z(n14538) );
  NAND U14916 ( .A(n14539), .B(n14538), .Z(n14490) );
  NAND U14917 ( .A(n14491), .B(n14490), .Z(n14494) );
  AND U14918 ( .A(o[54]), .B(\stack[1][1] ), .Z(n14495) );
  NAND U14919 ( .A(n14494), .B(n14495), .Z(n14497) );
  NAND U14920 ( .A(n14861), .B(n14860), .Z(n14496) );
  NAND U14921 ( .A(n14497), .B(n14496), .Z(n14500) );
  XOR U14922 ( .A(n14499), .B(n14498), .Z(n14501) );
  NAND U14923 ( .A(n14500), .B(n14501), .Z(n14503) );
  AND U14924 ( .A(o[55]), .B(\stack[1][1] ), .Z(n14536) );
  NAND U14925 ( .A(n14537), .B(n14536), .Z(n14502) );
  NAND U14926 ( .A(n14503), .B(n14502), .Z(n14506) );
  AND U14927 ( .A(o[56]), .B(\stack[1][1] ), .Z(n14507) );
  NAND U14928 ( .A(n14506), .B(n14507), .Z(n14509) );
  XOR U14929 ( .A(n14505), .B(n14504), .Z(n14871) );
  NAND U14930 ( .A(n14871), .B(n14870), .Z(n14508) );
  NAND U14931 ( .A(n14509), .B(n14508), .Z(n14512) );
  XOR U14932 ( .A(n14511), .B(n14510), .Z(n14513) );
  NAND U14933 ( .A(n14512), .B(n14513), .Z(n14515) );
  AND U14934 ( .A(o[57]), .B(\stack[1][1] ), .Z(n14534) );
  NAND U14935 ( .A(n14535), .B(n14534), .Z(n14514) );
  NAND U14936 ( .A(n14515), .B(n14514), .Z(n14518) );
  AND U14937 ( .A(o[58]), .B(\stack[1][1] ), .Z(n14519) );
  NAND U14938 ( .A(n14518), .B(n14519), .Z(n14521) );
  NAND U14939 ( .A(n14881), .B(n14880), .Z(n14520) );
  NAND U14940 ( .A(n14521), .B(n14520), .Z(n14522) );
  NAND U14941 ( .A(n14523), .B(n14522), .Z(n14525) );
  XOR U14942 ( .A(n14523), .B(n14522), .Z(n14533) );
  AND U14943 ( .A(o[59]), .B(\stack[1][1] ), .Z(n14532) );
  NAND U14944 ( .A(n14533), .B(n14532), .Z(n14524) );
  NAND U14945 ( .A(n14525), .B(n14524), .Z(n14528) );
  AND U14946 ( .A(o[60]), .B(\stack[1][1] ), .Z(n14529) );
  NAND U14947 ( .A(n14528), .B(n14529), .Z(n14531) );
  XOR U14948 ( .A(n14527), .B(n14526), .Z(n14891) );
  NAND U14949 ( .A(n14891), .B(n14890), .Z(n14530) );
  NAND U14950 ( .A(n14531), .B(n14530), .Z(n14900) );
  AND U14951 ( .A(\stack[1][1] ), .B(o[61]), .Z(n14898) );
  XNOR U14952 ( .A(n14899), .B(n14898), .Z(n14895) );
  NAND U14953 ( .A(o[61]), .B(\stack[1][0] ), .Z(n14888) );
  XNOR U14954 ( .A(n14533), .B(n14532), .Z(n14884) );
  NAND U14955 ( .A(o[59]), .B(\stack[1][0] ), .Z(n14878) );
  XNOR U14956 ( .A(n14535), .B(n14534), .Z(n14874) );
  NAND U14957 ( .A(o[57]), .B(\stack[1][0] ), .Z(n14868) );
  XNOR U14958 ( .A(n14537), .B(n14536), .Z(n14864) );
  NAND U14959 ( .A(o[55]), .B(\stack[1][0] ), .Z(n14858) );
  XNOR U14960 ( .A(n14539), .B(n14538), .Z(n14854) );
  NAND U14961 ( .A(o[53]), .B(\stack[1][0] ), .Z(n14848) );
  XNOR U14962 ( .A(n14541), .B(n14540), .Z(n14844) );
  NAND U14963 ( .A(o[51]), .B(\stack[1][0] ), .Z(n14838) );
  XNOR U14964 ( .A(n14543), .B(n14542), .Z(n14834) );
  NAND U14965 ( .A(o[49]), .B(\stack[1][0] ), .Z(n14828) );
  XNOR U14966 ( .A(n14545), .B(n14544), .Z(n14824) );
  NAND U14967 ( .A(o[47]), .B(\stack[1][0] ), .Z(n14818) );
  XNOR U14968 ( .A(n14547), .B(n14546), .Z(n14814) );
  NAND U14969 ( .A(o[45]), .B(\stack[1][0] ), .Z(n14808) );
  XNOR U14970 ( .A(n14549), .B(n14548), .Z(n14804) );
  NAND U14971 ( .A(o[43]), .B(\stack[1][0] ), .Z(n14798) );
  XNOR U14972 ( .A(n14551), .B(n14550), .Z(n14794) );
  NAND U14973 ( .A(o[41]), .B(\stack[1][0] ), .Z(n14788) );
  XNOR U14974 ( .A(n14553), .B(n14552), .Z(n14784) );
  NAND U14975 ( .A(o[39]), .B(\stack[1][0] ), .Z(n14778) );
  XNOR U14976 ( .A(n14555), .B(n14554), .Z(n14774) );
  NAND U14977 ( .A(o[37]), .B(\stack[1][0] ), .Z(n14768) );
  XNOR U14978 ( .A(n14557), .B(n14556), .Z(n14764) );
  NAND U14979 ( .A(o[35]), .B(\stack[1][0] ), .Z(n14758) );
  XNOR U14980 ( .A(n14559), .B(n14558), .Z(n14754) );
  NAND U14981 ( .A(o[33]), .B(\stack[1][0] ), .Z(n14748) );
  XNOR U14982 ( .A(n14561), .B(n14560), .Z(n14744) );
  NAND U14983 ( .A(o[31]), .B(\stack[1][0] ), .Z(n14738) );
  XNOR U14984 ( .A(n14563), .B(n14562), .Z(n14734) );
  NAND U14985 ( .A(o[29]), .B(\stack[1][0] ), .Z(n14728) );
  XNOR U14986 ( .A(n14565), .B(n14564), .Z(n14724) );
  NAND U14987 ( .A(o[27]), .B(\stack[1][0] ), .Z(n14718) );
  XNOR U14988 ( .A(n14567), .B(n14566), .Z(n14714) );
  NAND U14989 ( .A(o[25]), .B(\stack[1][0] ), .Z(n14708) );
  XNOR U14990 ( .A(n14569), .B(n14568), .Z(n14704) );
  NAND U14991 ( .A(o[23]), .B(\stack[1][0] ), .Z(n14698) );
  XNOR U14992 ( .A(n14571), .B(n14570), .Z(n14694) );
  NAND U14993 ( .A(o[21]), .B(\stack[1][0] ), .Z(n14688) );
  XNOR U14994 ( .A(n14573), .B(n14572), .Z(n14684) );
  NAND U14995 ( .A(o[19]), .B(\stack[1][0] ), .Z(n14678) );
  XNOR U14996 ( .A(n14575), .B(n14574), .Z(n14674) );
  NAND U14997 ( .A(o[17]), .B(\stack[1][0] ), .Z(n14668) );
  XNOR U14998 ( .A(n14577), .B(n14576), .Z(n14664) );
  NAND U14999 ( .A(o[15]), .B(\stack[1][0] ), .Z(n14658) );
  XNOR U15000 ( .A(n14579), .B(n14578), .Z(n14654) );
  NAND U15001 ( .A(o[13]), .B(\stack[1][0] ), .Z(n14648) );
  NAND U15002 ( .A(o[11]), .B(\stack[1][0] ), .Z(n14636) );
  XNOR U15003 ( .A(n14581), .B(n14580), .Z(n14632) );
  NAND U15004 ( .A(o[9]), .B(\stack[1][0] ), .Z(n14626) );
  NAND U15005 ( .A(o[7]), .B(\stack[1][0] ), .Z(n14614) );
  XNOR U15006 ( .A(n14583), .B(n14582), .Z(n14610) );
  NAND U15007 ( .A(o[5]), .B(\stack[1][0] ), .Z(n14604) );
  XNOR U15008 ( .A(n14585), .B(n14584), .Z(n14600) );
  NAND U15009 ( .A(o[3]), .B(\stack[1][0] ), .Z(n14594) );
  AND U15010 ( .A(o[1]), .B(\stack[1][0] ), .Z(n17291) );
  NAND U15011 ( .A(n17292), .B(n17291), .Z(n14587) );
  NAND U15012 ( .A(o[2]), .B(\stack[1][0] ), .Z(n14586) );
  AND U15013 ( .A(n14587), .B(n14586), .Z(n14593) );
  NAND U15014 ( .A(n17292), .B(o[1]), .Z(n14588) );
  XNOR U15015 ( .A(o[2]), .B(n14588), .Z(n14589) );
  AND U15016 ( .A(\stack[1][0] ), .B(n14589), .Z(n17260) );
  AND U15017 ( .A(\stack[1][1] ), .B(o[1]), .Z(n14591) );
  XNOR U15018 ( .A(n14591), .B(n14590), .Z(n17261) );
  NAND U15019 ( .A(n17260), .B(n17261), .Z(n14592) );
  NANDN U15020 ( .A(n14593), .B(n14592), .Z(n14595) );
  NAND U15021 ( .A(n14594), .B(n14595), .Z(n14599) );
  XNOR U15022 ( .A(n14597), .B(n14596), .Z(n17219) );
  NAND U15023 ( .A(n17218), .B(n17219), .Z(n14598) );
  NAND U15024 ( .A(n14599), .B(n14598), .Z(n14601) );
  NAND U15025 ( .A(n14600), .B(n14601), .Z(n14603) );
  NAND U15026 ( .A(o[4]), .B(\stack[1][0] ), .Z(n17180) );
  NAND U15027 ( .A(n17179), .B(n17180), .Z(n14602) );
  NAND U15028 ( .A(n14603), .B(n14602), .Z(n14605) );
  NAND U15029 ( .A(n14604), .B(n14605), .Z(n14609) );
  XNOR U15030 ( .A(n14607), .B(n14606), .Z(n17141) );
  NAND U15031 ( .A(n17140), .B(n17141), .Z(n14608) );
  NAND U15032 ( .A(n14609), .B(n14608), .Z(n14611) );
  NAND U15033 ( .A(n14610), .B(n14611), .Z(n14613) );
  NAND U15034 ( .A(o[6]), .B(\stack[1][0] ), .Z(n17102) );
  NAND U15035 ( .A(n17101), .B(n17102), .Z(n14612) );
  NAND U15036 ( .A(n14613), .B(n14612), .Z(n14615) );
  NAND U15037 ( .A(n14614), .B(n14615), .Z(n14619) );
  XNOR U15038 ( .A(n14617), .B(n14616), .Z(n17063) );
  NAND U15039 ( .A(n17062), .B(n17063), .Z(n14618) );
  NAND U15040 ( .A(n14619), .B(n14618), .Z(n14622) );
  XNOR U15041 ( .A(n14621), .B(n14620), .Z(n14623) );
  NAND U15042 ( .A(n14622), .B(n14623), .Z(n14625) );
  NAND U15043 ( .A(o[8]), .B(\stack[1][0] ), .Z(n17025) );
  NAND U15044 ( .A(n17024), .B(n17025), .Z(n14624) );
  NAND U15045 ( .A(n14625), .B(n14624), .Z(n14627) );
  NAND U15046 ( .A(n14626), .B(n14627), .Z(n14631) );
  XNOR U15047 ( .A(n14629), .B(n14628), .Z(n16986) );
  NAND U15048 ( .A(n16985), .B(n16986), .Z(n14630) );
  NAND U15049 ( .A(n14631), .B(n14630), .Z(n14633) );
  NAND U15050 ( .A(n14632), .B(n14633), .Z(n14635) );
  NAND U15051 ( .A(o[10]), .B(\stack[1][0] ), .Z(n16948) );
  NAND U15052 ( .A(n16947), .B(n16948), .Z(n14634) );
  NAND U15053 ( .A(n14635), .B(n14634), .Z(n14637) );
  NAND U15054 ( .A(n14636), .B(n14637), .Z(n14641) );
  XOR U15055 ( .A(n14639), .B(n14638), .Z(n16911) );
  NAND U15056 ( .A(n16910), .B(n16911), .Z(n14640) );
  NAND U15057 ( .A(n14641), .B(n14640), .Z(n14644) );
  NAND U15058 ( .A(n14644), .B(n14645), .Z(n14647) );
  NAND U15059 ( .A(o[12]), .B(\stack[1][0] ), .Z(n16871) );
  NAND U15060 ( .A(n16870), .B(n16871), .Z(n14646) );
  NAND U15061 ( .A(n14647), .B(n14646), .Z(n14649) );
  NAND U15062 ( .A(n14648), .B(n14649), .Z(n14653) );
  XNOR U15063 ( .A(n14651), .B(n14650), .Z(n16832) );
  NAND U15064 ( .A(n16831), .B(n16832), .Z(n14652) );
  NAND U15065 ( .A(n14653), .B(n14652), .Z(n14655) );
  NAND U15066 ( .A(n14654), .B(n14655), .Z(n14657) );
  NAND U15067 ( .A(o[14]), .B(\stack[1][0] ), .Z(n16793) );
  NAND U15068 ( .A(n16792), .B(n16793), .Z(n14656) );
  NAND U15069 ( .A(n14657), .B(n14656), .Z(n14659) );
  NAND U15070 ( .A(n14658), .B(n14659), .Z(n14663) );
  XOR U15071 ( .A(n14661), .B(n14660), .Z(n16755) );
  NAND U15072 ( .A(n16754), .B(n16755), .Z(n14662) );
  NAND U15073 ( .A(n14663), .B(n14662), .Z(n14665) );
  NAND U15074 ( .A(n14664), .B(n14665), .Z(n14667) );
  NAND U15075 ( .A(o[16]), .B(\stack[1][0] ), .Z(n16717) );
  NAND U15076 ( .A(n16716), .B(n16717), .Z(n14666) );
  NAND U15077 ( .A(n14667), .B(n14666), .Z(n14669) );
  NAND U15078 ( .A(n14668), .B(n14669), .Z(n14673) );
  XNOR U15079 ( .A(n14671), .B(n14670), .Z(n16678) );
  NAND U15080 ( .A(n16677), .B(n16678), .Z(n14672) );
  NAND U15081 ( .A(n14673), .B(n14672), .Z(n14675) );
  NAND U15082 ( .A(n14674), .B(n14675), .Z(n14677) );
  NAND U15083 ( .A(o[18]), .B(\stack[1][0] ), .Z(n16640) );
  NAND U15084 ( .A(n16639), .B(n16640), .Z(n14676) );
  NAND U15085 ( .A(n14677), .B(n14676), .Z(n14679) );
  NAND U15086 ( .A(n14678), .B(n14679), .Z(n14683) );
  XNOR U15087 ( .A(n14681), .B(n14680), .Z(n16601) );
  NAND U15088 ( .A(n16600), .B(n16601), .Z(n14682) );
  NAND U15089 ( .A(n14683), .B(n14682), .Z(n14685) );
  NAND U15090 ( .A(n14684), .B(n14685), .Z(n14687) );
  NAND U15091 ( .A(o[20]), .B(\stack[1][0] ), .Z(n16563) );
  NAND U15092 ( .A(n16562), .B(n16563), .Z(n14686) );
  NAND U15093 ( .A(n14687), .B(n14686), .Z(n14689) );
  NAND U15094 ( .A(n14688), .B(n14689), .Z(n14693) );
  XNOR U15095 ( .A(n14691), .B(n14690), .Z(n16524) );
  NAND U15096 ( .A(n16523), .B(n16524), .Z(n14692) );
  NAND U15097 ( .A(n14693), .B(n14692), .Z(n14695) );
  NAND U15098 ( .A(n14694), .B(n14695), .Z(n14697) );
  NAND U15099 ( .A(o[22]), .B(\stack[1][0] ), .Z(n16485) );
  NAND U15100 ( .A(n16484), .B(n16485), .Z(n14696) );
  NAND U15101 ( .A(n14697), .B(n14696), .Z(n14699) );
  NAND U15102 ( .A(n14698), .B(n14699), .Z(n14703) );
  XNOR U15103 ( .A(n14701), .B(n14700), .Z(n16447) );
  NAND U15104 ( .A(n16446), .B(n16447), .Z(n14702) );
  NAND U15105 ( .A(n14703), .B(n14702), .Z(n14705) );
  NAND U15106 ( .A(n14704), .B(n14705), .Z(n14707) );
  NAND U15107 ( .A(o[24]), .B(\stack[1][0] ), .Z(n16409) );
  NAND U15108 ( .A(n16408), .B(n16409), .Z(n14706) );
  NAND U15109 ( .A(n14707), .B(n14706), .Z(n14709) );
  NAND U15110 ( .A(n14708), .B(n14709), .Z(n14713) );
  XNOR U15111 ( .A(n14711), .B(n14710), .Z(n16371) );
  NAND U15112 ( .A(n16370), .B(n16371), .Z(n14712) );
  NAND U15113 ( .A(n14713), .B(n14712), .Z(n14715) );
  NAND U15114 ( .A(n14714), .B(n14715), .Z(n14717) );
  NAND U15115 ( .A(o[26]), .B(\stack[1][0] ), .Z(n16332) );
  NAND U15116 ( .A(n16331), .B(n16332), .Z(n14716) );
  NAND U15117 ( .A(n14717), .B(n14716), .Z(n14719) );
  NAND U15118 ( .A(n14718), .B(n14719), .Z(n14723) );
  XNOR U15119 ( .A(n14721), .B(n14720), .Z(n16293) );
  NAND U15120 ( .A(n16292), .B(n16293), .Z(n14722) );
  NAND U15121 ( .A(n14723), .B(n14722), .Z(n14725) );
  NAND U15122 ( .A(n14724), .B(n14725), .Z(n14727) );
  NAND U15123 ( .A(o[28]), .B(\stack[1][0] ), .Z(n16254) );
  NAND U15124 ( .A(n16253), .B(n16254), .Z(n14726) );
  NAND U15125 ( .A(n14727), .B(n14726), .Z(n14729) );
  NAND U15126 ( .A(n14728), .B(n14729), .Z(n14733) );
  XNOR U15127 ( .A(n14731), .B(n14730), .Z(n16215) );
  NAND U15128 ( .A(n16214), .B(n16215), .Z(n14732) );
  NAND U15129 ( .A(n14733), .B(n14732), .Z(n14735) );
  NAND U15130 ( .A(n14734), .B(n14735), .Z(n14737) );
  NAND U15131 ( .A(o[30]), .B(\stack[1][0] ), .Z(n16177) );
  NAND U15132 ( .A(n16176), .B(n16177), .Z(n14736) );
  NAND U15133 ( .A(n14737), .B(n14736), .Z(n14739) );
  NAND U15134 ( .A(n14738), .B(n14739), .Z(n14743) );
  XNOR U15135 ( .A(n14741), .B(n14740), .Z(n16138) );
  NAND U15136 ( .A(n16137), .B(n16138), .Z(n14742) );
  NAND U15137 ( .A(n14743), .B(n14742), .Z(n14745) );
  NAND U15138 ( .A(n14744), .B(n14745), .Z(n14747) );
  NAND U15139 ( .A(o[32]), .B(\stack[1][0] ), .Z(n16100) );
  NAND U15140 ( .A(n16099), .B(n16100), .Z(n14746) );
  NAND U15141 ( .A(n14747), .B(n14746), .Z(n14749) );
  NAND U15142 ( .A(n14748), .B(n14749), .Z(n14753) );
  XNOR U15143 ( .A(n14751), .B(n14750), .Z(n16063) );
  NAND U15144 ( .A(n16062), .B(n16063), .Z(n14752) );
  NAND U15145 ( .A(n14753), .B(n14752), .Z(n14755) );
  NAND U15146 ( .A(n14754), .B(n14755), .Z(n14757) );
  NAND U15147 ( .A(o[34]), .B(\stack[1][0] ), .Z(n16024) );
  NAND U15148 ( .A(n16023), .B(n16024), .Z(n14756) );
  NAND U15149 ( .A(n14757), .B(n14756), .Z(n14759) );
  NAND U15150 ( .A(n14758), .B(n14759), .Z(n14763) );
  XNOR U15151 ( .A(n14761), .B(n14760), .Z(n15987) );
  NAND U15152 ( .A(n15986), .B(n15987), .Z(n14762) );
  NAND U15153 ( .A(n14763), .B(n14762), .Z(n14765) );
  NAND U15154 ( .A(n14764), .B(n14765), .Z(n14767) );
  NAND U15155 ( .A(o[36]), .B(\stack[1][0] ), .Z(n15948) );
  NAND U15156 ( .A(n15947), .B(n15948), .Z(n14766) );
  NAND U15157 ( .A(n14767), .B(n14766), .Z(n14769) );
  NAND U15158 ( .A(n14768), .B(n14769), .Z(n14773) );
  XNOR U15159 ( .A(n14771), .B(n14770), .Z(n15911) );
  NAND U15160 ( .A(n15910), .B(n15911), .Z(n14772) );
  NAND U15161 ( .A(n14773), .B(n14772), .Z(n14775) );
  NAND U15162 ( .A(n14774), .B(n14775), .Z(n14777) );
  NAND U15163 ( .A(o[38]), .B(\stack[1][0] ), .Z(n15873) );
  NAND U15164 ( .A(n15872), .B(n15873), .Z(n14776) );
  NAND U15165 ( .A(n14777), .B(n14776), .Z(n14779) );
  NAND U15166 ( .A(n14778), .B(n14779), .Z(n14783) );
  XNOR U15167 ( .A(n14781), .B(n14780), .Z(n15835) );
  NAND U15168 ( .A(n15834), .B(n15835), .Z(n14782) );
  NAND U15169 ( .A(n14783), .B(n14782), .Z(n14785) );
  NAND U15170 ( .A(n14784), .B(n14785), .Z(n14787) );
  NAND U15171 ( .A(o[40]), .B(\stack[1][0] ), .Z(n15797) );
  NAND U15172 ( .A(n15796), .B(n15797), .Z(n14786) );
  NAND U15173 ( .A(n14787), .B(n14786), .Z(n14789) );
  NAND U15174 ( .A(n14788), .B(n14789), .Z(n14793) );
  XNOR U15175 ( .A(n14791), .B(n14790), .Z(n15759) );
  NAND U15176 ( .A(n15758), .B(n15759), .Z(n14792) );
  NAND U15177 ( .A(n14793), .B(n14792), .Z(n14795) );
  NAND U15178 ( .A(n14794), .B(n14795), .Z(n14797) );
  NAND U15179 ( .A(o[42]), .B(\stack[1][0] ), .Z(n15721) );
  NAND U15180 ( .A(n15720), .B(n15721), .Z(n14796) );
  NAND U15181 ( .A(n14797), .B(n14796), .Z(n14799) );
  NAND U15182 ( .A(n14798), .B(n14799), .Z(n14803) );
  XNOR U15183 ( .A(n14801), .B(n14800), .Z(n15683) );
  NAND U15184 ( .A(n15682), .B(n15683), .Z(n14802) );
  NAND U15185 ( .A(n14803), .B(n14802), .Z(n14805) );
  NAND U15186 ( .A(n14804), .B(n14805), .Z(n14807) );
  NAND U15187 ( .A(o[44]), .B(\stack[1][0] ), .Z(n15645) );
  NAND U15188 ( .A(n15644), .B(n15645), .Z(n14806) );
  NAND U15189 ( .A(n14807), .B(n14806), .Z(n14809) );
  NAND U15190 ( .A(n14808), .B(n14809), .Z(n14813) );
  XNOR U15191 ( .A(n14811), .B(n14810), .Z(n15607) );
  NAND U15192 ( .A(n15606), .B(n15607), .Z(n14812) );
  NAND U15193 ( .A(n14813), .B(n14812), .Z(n14815) );
  NAND U15194 ( .A(n14814), .B(n14815), .Z(n14817) );
  NAND U15195 ( .A(o[46]), .B(\stack[1][0] ), .Z(n15569) );
  NAND U15196 ( .A(n15568), .B(n15569), .Z(n14816) );
  NAND U15197 ( .A(n14817), .B(n14816), .Z(n14819) );
  NAND U15198 ( .A(n14818), .B(n14819), .Z(n14823) );
  XNOR U15199 ( .A(n14821), .B(n14820), .Z(n15531) );
  NAND U15200 ( .A(n15530), .B(n15531), .Z(n14822) );
  NAND U15201 ( .A(n14823), .B(n14822), .Z(n14825) );
  NAND U15202 ( .A(n14824), .B(n14825), .Z(n14827) );
  NAND U15203 ( .A(o[48]), .B(\stack[1][0] ), .Z(n15493) );
  NAND U15204 ( .A(n15492), .B(n15493), .Z(n14826) );
  NAND U15205 ( .A(n14827), .B(n14826), .Z(n14829) );
  NAND U15206 ( .A(n14828), .B(n14829), .Z(n14833) );
  XNOR U15207 ( .A(n14831), .B(n14830), .Z(n15455) );
  NAND U15208 ( .A(n15454), .B(n15455), .Z(n14832) );
  NAND U15209 ( .A(n14833), .B(n14832), .Z(n14835) );
  NAND U15210 ( .A(n14834), .B(n14835), .Z(n14837) );
  NAND U15211 ( .A(o[50]), .B(\stack[1][0] ), .Z(n15417) );
  NAND U15212 ( .A(n15416), .B(n15417), .Z(n14836) );
  NAND U15213 ( .A(n14837), .B(n14836), .Z(n14839) );
  NAND U15214 ( .A(n14838), .B(n14839), .Z(n14843) );
  XNOR U15215 ( .A(n14841), .B(n14840), .Z(n15379) );
  NAND U15216 ( .A(n15378), .B(n15379), .Z(n14842) );
  NAND U15217 ( .A(n14843), .B(n14842), .Z(n14845) );
  NAND U15218 ( .A(n14844), .B(n14845), .Z(n14847) );
  NAND U15219 ( .A(o[52]), .B(\stack[1][0] ), .Z(n15341) );
  NAND U15220 ( .A(n15340), .B(n15341), .Z(n14846) );
  NAND U15221 ( .A(n14847), .B(n14846), .Z(n14849) );
  NAND U15222 ( .A(n14848), .B(n14849), .Z(n14853) );
  XNOR U15223 ( .A(n14851), .B(n14850), .Z(n15303) );
  NAND U15224 ( .A(n15302), .B(n15303), .Z(n14852) );
  NAND U15225 ( .A(n14853), .B(n14852), .Z(n14855) );
  NAND U15226 ( .A(n14854), .B(n14855), .Z(n14857) );
  NAND U15227 ( .A(o[54]), .B(\stack[1][0] ), .Z(n15265) );
  NAND U15228 ( .A(n15264), .B(n15265), .Z(n14856) );
  NAND U15229 ( .A(n14857), .B(n14856), .Z(n14859) );
  NAND U15230 ( .A(n14858), .B(n14859), .Z(n14863) );
  XNOR U15231 ( .A(n14861), .B(n14860), .Z(n15227) );
  NAND U15232 ( .A(n15226), .B(n15227), .Z(n14862) );
  NAND U15233 ( .A(n14863), .B(n14862), .Z(n14865) );
  NAND U15234 ( .A(n14864), .B(n14865), .Z(n14867) );
  NAND U15235 ( .A(o[56]), .B(\stack[1][0] ), .Z(n15189) );
  NAND U15236 ( .A(n15188), .B(n15189), .Z(n14866) );
  NAND U15237 ( .A(n14867), .B(n14866), .Z(n14869) );
  NAND U15238 ( .A(n14868), .B(n14869), .Z(n14873) );
  XNOR U15239 ( .A(n14871), .B(n14870), .Z(n15151) );
  NAND U15240 ( .A(n15150), .B(n15151), .Z(n14872) );
  NAND U15241 ( .A(n14873), .B(n14872), .Z(n14875) );
  NAND U15242 ( .A(n14874), .B(n14875), .Z(n14877) );
  NAND U15243 ( .A(o[58]), .B(\stack[1][0] ), .Z(n15113) );
  NAND U15244 ( .A(n15112), .B(n15113), .Z(n14876) );
  NAND U15245 ( .A(n14877), .B(n14876), .Z(n14879) );
  NAND U15246 ( .A(n14878), .B(n14879), .Z(n14883) );
  XNOR U15247 ( .A(n14881), .B(n14880), .Z(n15075) );
  NAND U15248 ( .A(n15074), .B(n15075), .Z(n14882) );
  NAND U15249 ( .A(n14883), .B(n14882), .Z(n14885) );
  NAND U15250 ( .A(n14884), .B(n14885), .Z(n14887) );
  NAND U15251 ( .A(o[60]), .B(\stack[1][0] ), .Z(n15037) );
  NAND U15252 ( .A(n15036), .B(n15037), .Z(n14886) );
  NAND U15253 ( .A(n14887), .B(n14886), .Z(n14889) );
  NAND U15254 ( .A(n14888), .B(n14889), .Z(n14893) );
  XNOR U15255 ( .A(n14891), .B(n14890), .Z(n14999) );
  NAND U15256 ( .A(n14998), .B(n14999), .Z(n14892) );
  NAND U15257 ( .A(n14893), .B(n14892), .Z(n14894) );
  NAND U15258 ( .A(\stack[1][0] ), .B(o[62]), .Z(n14961) );
  NAND U15259 ( .A(n14960), .B(n14961), .Z(n14897) );
  NAND U15260 ( .A(n14895), .B(n14894), .Z(n14896) );
  AND U15261 ( .A(n14897), .B(n14896), .Z(n14905) );
  NAND U15262 ( .A(n14899), .B(n14898), .Z(n14903) );
  NAND U15263 ( .A(n14901), .B(n14900), .Z(n14902) );
  NAND U15264 ( .A(n14903), .B(n14902), .Z(n14904) );
  XNOR U15265 ( .A(n14905), .B(n14904), .Z(n14906) );
  XNOR U15266 ( .A(n14907), .B(n14906), .Z(n14908) );
  XNOR U15267 ( .A(n14909), .B(n14908), .Z(n14917) );
  AND U15268 ( .A(n14911), .B(n14910), .Z(n14915) );
  AND U15269 ( .A(n14913), .B(n14912), .Z(n14914) );
  OR U15270 ( .A(n14915), .B(n14914), .Z(n14916) );
  XNOR U15271 ( .A(n14917), .B(n14916), .Z(n14918) );
  NANDN U15272 ( .A(n17294), .B(n14918), .Z(n14922) );
  NAND U15273 ( .A(x[63]), .B(n17311), .Z(n14920) );
  AND U15274 ( .A(opcode[2]), .B(n17314), .Z(n17318) );
  NAND U15275 ( .A(\stack[1][63] ), .B(n17318), .Z(n14919) );
  AND U15276 ( .A(n14920), .B(n14919), .Z(n14921) );
  AND U15277 ( .A(n14922), .B(n14921), .Z(n14923) );
  XNOR U15278 ( .A(opcode[0]), .B(opcode[2]), .Z(n14925) );
  XNOR U15279 ( .A(opcode[2]), .B(opcode[1]), .Z(n14924) );
  NAND U15280 ( .A(n14925), .B(n14924), .Z(n17317) );
  AND U15281 ( .A(opcode[2]), .B(n3163), .Z(n17313) );
  NAND U15282 ( .A(\stack[1][63] ), .B(n17313), .Z(n14926) );
  NAND U15283 ( .A(n17317), .B(n14926), .Z(n14927) );
  NAND U15284 ( .A(o[63]), .B(n14927), .Z(n14928) );
  NAND U15285 ( .A(n14929), .B(n14928), .Z(n2132) );
  NAND U15286 ( .A(\stack[6][62] ), .B(n17311), .Z(n14931) );
  NANDN U15287 ( .A(n17311), .B(\stack[7][62] ), .Z(n14930) );
  NAND U15288 ( .A(n14931), .B(n14930), .Z(n2133) );
  NAND U15289 ( .A(\stack[5][62] ), .B(n17311), .Z(n14933) );
  NAND U15290 ( .A(n17305), .B(\stack[7][62] ), .Z(n14932) );
  AND U15291 ( .A(n14933), .B(n14932), .Z(n14935) );
  NAND U15292 ( .A(n17308), .B(\stack[6][62] ), .Z(n14934) );
  NAND U15293 ( .A(n14935), .B(n14934), .Z(n2134) );
  NAND U15294 ( .A(\stack[4][62] ), .B(n17311), .Z(n14937) );
  NAND U15295 ( .A(n17305), .B(\stack[6][62] ), .Z(n14936) );
  AND U15296 ( .A(n14937), .B(n14936), .Z(n14939) );
  NAND U15297 ( .A(n17308), .B(\stack[5][62] ), .Z(n14938) );
  NAND U15298 ( .A(n14939), .B(n14938), .Z(n2135) );
  NAND U15299 ( .A(\stack[3][62] ), .B(n17311), .Z(n14941) );
  NAND U15300 ( .A(n17305), .B(\stack[5][62] ), .Z(n14940) );
  AND U15301 ( .A(n14941), .B(n14940), .Z(n14943) );
  NAND U15302 ( .A(n17308), .B(\stack[4][62] ), .Z(n14942) );
  NAND U15303 ( .A(n14943), .B(n14942), .Z(n2136) );
  NAND U15304 ( .A(\stack[2][62] ), .B(n17311), .Z(n14945) );
  NAND U15305 ( .A(n17305), .B(\stack[4][62] ), .Z(n14944) );
  AND U15306 ( .A(n14945), .B(n14944), .Z(n14947) );
  NAND U15307 ( .A(n17308), .B(\stack[3][62] ), .Z(n14946) );
  NAND U15308 ( .A(n14947), .B(n14946), .Z(n2137) );
  NAND U15309 ( .A(n17311), .B(\stack[1][62] ), .Z(n14949) );
  NAND U15310 ( .A(n17305), .B(\stack[3][62] ), .Z(n14948) );
  AND U15311 ( .A(n14949), .B(n14948), .Z(n14951) );
  NAND U15312 ( .A(n17308), .B(\stack[2][62] ), .Z(n14950) );
  NAND U15313 ( .A(n14951), .B(n14950), .Z(n2138) );
  NAND U15314 ( .A(n17311), .B(o[62]), .Z(n14953) );
  NAND U15315 ( .A(n17305), .B(\stack[2][62] ), .Z(n14952) );
  AND U15316 ( .A(n14953), .B(n14952), .Z(n14955) );
  NAND U15317 ( .A(\stack[1][62] ), .B(n17308), .Z(n14954) );
  NAND U15318 ( .A(n14955), .B(n14954), .Z(n2139) );
  NAND U15319 ( .A(\stack[1][62] ), .B(n17313), .Z(n14956) );
  NAND U15320 ( .A(n17317), .B(n14956), .Z(n14957) );
  AND U15321 ( .A(o[62]), .B(n14957), .Z(n14966) );
  NAND U15322 ( .A(x[62]), .B(n17311), .Z(n14959) );
  NAND U15323 ( .A(\stack[1][62] ), .B(n17318), .Z(n14958) );
  AND U15324 ( .A(n14959), .B(n14958), .Z(n14964) );
  XNOR U15325 ( .A(n14961), .B(n14960), .Z(n14962) );
  NANDN U15326 ( .A(n17294), .B(n14962), .Z(n14963) );
  NAND U15327 ( .A(n14964), .B(n14963), .Z(n14965) );
  NOR U15328 ( .A(n14966), .B(n14965), .Z(n14967) );
  NAND U15329 ( .A(\stack[6][61] ), .B(n17311), .Z(n14969) );
  NANDN U15330 ( .A(n17311), .B(\stack[7][61] ), .Z(n14968) );
  NAND U15331 ( .A(n14969), .B(n14968), .Z(n2141) );
  NAND U15332 ( .A(\stack[5][61] ), .B(n17311), .Z(n14971) );
  NAND U15333 ( .A(n17305), .B(\stack[7][61] ), .Z(n14970) );
  AND U15334 ( .A(n14971), .B(n14970), .Z(n14973) );
  NAND U15335 ( .A(n17308), .B(\stack[6][61] ), .Z(n14972) );
  NAND U15336 ( .A(n14973), .B(n14972), .Z(n2142) );
  NAND U15337 ( .A(\stack[4][61] ), .B(n17311), .Z(n14975) );
  NAND U15338 ( .A(n17305), .B(\stack[6][61] ), .Z(n14974) );
  AND U15339 ( .A(n14975), .B(n14974), .Z(n14977) );
  NAND U15340 ( .A(n17308), .B(\stack[5][61] ), .Z(n14976) );
  NAND U15341 ( .A(n14977), .B(n14976), .Z(n2143) );
  NAND U15342 ( .A(\stack[3][61] ), .B(n17311), .Z(n14979) );
  NAND U15343 ( .A(n17305), .B(\stack[5][61] ), .Z(n14978) );
  AND U15344 ( .A(n14979), .B(n14978), .Z(n14981) );
  NAND U15345 ( .A(n17308), .B(\stack[4][61] ), .Z(n14980) );
  NAND U15346 ( .A(n14981), .B(n14980), .Z(n2144) );
  NAND U15347 ( .A(\stack[2][61] ), .B(n17311), .Z(n14983) );
  NAND U15348 ( .A(n17305), .B(\stack[4][61] ), .Z(n14982) );
  AND U15349 ( .A(n14983), .B(n14982), .Z(n14985) );
  NAND U15350 ( .A(n17308), .B(\stack[3][61] ), .Z(n14984) );
  NAND U15351 ( .A(n14985), .B(n14984), .Z(n2145) );
  NAND U15352 ( .A(n17311), .B(\stack[1][61] ), .Z(n14987) );
  NAND U15353 ( .A(n17305), .B(\stack[3][61] ), .Z(n14986) );
  AND U15354 ( .A(n14987), .B(n14986), .Z(n14989) );
  NAND U15355 ( .A(n17308), .B(\stack[2][61] ), .Z(n14988) );
  NAND U15356 ( .A(n14989), .B(n14988), .Z(n2146) );
  NAND U15357 ( .A(n17311), .B(o[61]), .Z(n14991) );
  NAND U15358 ( .A(n17305), .B(\stack[2][61] ), .Z(n14990) );
  AND U15359 ( .A(n14991), .B(n14990), .Z(n14993) );
  NAND U15360 ( .A(\stack[1][61] ), .B(n17308), .Z(n14992) );
  NAND U15361 ( .A(n14993), .B(n14992), .Z(n2147) );
  NAND U15362 ( .A(\stack[1][61] ), .B(n17313), .Z(n14994) );
  NAND U15363 ( .A(n17317), .B(n14994), .Z(n14995) );
  AND U15364 ( .A(o[61]), .B(n14995), .Z(n15004) );
  NAND U15365 ( .A(x[61]), .B(n17311), .Z(n14997) );
  NAND U15366 ( .A(\stack[1][61] ), .B(n17318), .Z(n14996) );
  AND U15367 ( .A(n14997), .B(n14996), .Z(n15002) );
  XNOR U15368 ( .A(n14999), .B(n14998), .Z(n15000) );
  NANDN U15369 ( .A(n17294), .B(n15000), .Z(n15001) );
  NAND U15370 ( .A(n15002), .B(n15001), .Z(n15003) );
  NOR U15371 ( .A(n15004), .B(n15003), .Z(n15005) );
  NAND U15372 ( .A(\stack[6][60] ), .B(n17311), .Z(n15007) );
  NANDN U15373 ( .A(n17311), .B(\stack[7][60] ), .Z(n15006) );
  NAND U15374 ( .A(n15007), .B(n15006), .Z(n2149) );
  NAND U15375 ( .A(\stack[5][60] ), .B(n17311), .Z(n15009) );
  NAND U15376 ( .A(n17305), .B(\stack[7][60] ), .Z(n15008) );
  AND U15377 ( .A(n15009), .B(n15008), .Z(n15011) );
  NAND U15378 ( .A(n17308), .B(\stack[6][60] ), .Z(n15010) );
  NAND U15379 ( .A(n15011), .B(n15010), .Z(n2150) );
  NAND U15380 ( .A(\stack[4][60] ), .B(n17311), .Z(n15013) );
  NAND U15381 ( .A(n17305), .B(\stack[6][60] ), .Z(n15012) );
  AND U15382 ( .A(n15013), .B(n15012), .Z(n15015) );
  NAND U15383 ( .A(n17308), .B(\stack[5][60] ), .Z(n15014) );
  NAND U15384 ( .A(n15015), .B(n15014), .Z(n2151) );
  NAND U15385 ( .A(\stack[3][60] ), .B(n17311), .Z(n15017) );
  NAND U15386 ( .A(n17305), .B(\stack[5][60] ), .Z(n15016) );
  AND U15387 ( .A(n15017), .B(n15016), .Z(n15019) );
  NAND U15388 ( .A(n17308), .B(\stack[4][60] ), .Z(n15018) );
  NAND U15389 ( .A(n15019), .B(n15018), .Z(n2152) );
  NAND U15390 ( .A(\stack[2][60] ), .B(n17311), .Z(n15021) );
  NAND U15391 ( .A(n17305), .B(\stack[4][60] ), .Z(n15020) );
  AND U15392 ( .A(n15021), .B(n15020), .Z(n15023) );
  NAND U15393 ( .A(n17308), .B(\stack[3][60] ), .Z(n15022) );
  NAND U15394 ( .A(n15023), .B(n15022), .Z(n2153) );
  NAND U15395 ( .A(n17311), .B(\stack[1][60] ), .Z(n15025) );
  NAND U15396 ( .A(n17305), .B(\stack[3][60] ), .Z(n15024) );
  AND U15397 ( .A(n15025), .B(n15024), .Z(n15027) );
  NAND U15398 ( .A(n17308), .B(\stack[2][60] ), .Z(n15026) );
  NAND U15399 ( .A(n15027), .B(n15026), .Z(n2154) );
  NAND U15400 ( .A(n17311), .B(o[60]), .Z(n15029) );
  NAND U15401 ( .A(n17305), .B(\stack[2][60] ), .Z(n15028) );
  AND U15402 ( .A(n15029), .B(n15028), .Z(n15031) );
  NAND U15403 ( .A(\stack[1][60] ), .B(n17308), .Z(n15030) );
  NAND U15404 ( .A(n15031), .B(n15030), .Z(n2155) );
  NAND U15405 ( .A(\stack[1][60] ), .B(n17313), .Z(n15032) );
  NAND U15406 ( .A(n17317), .B(n15032), .Z(n15033) );
  AND U15407 ( .A(o[60]), .B(n15033), .Z(n15042) );
  NAND U15408 ( .A(x[60]), .B(n17311), .Z(n15035) );
  NAND U15409 ( .A(\stack[1][60] ), .B(n17318), .Z(n15034) );
  AND U15410 ( .A(n15035), .B(n15034), .Z(n15040) );
  XNOR U15411 ( .A(n15037), .B(n15036), .Z(n15038) );
  NANDN U15412 ( .A(n17294), .B(n15038), .Z(n15039) );
  NAND U15413 ( .A(n15040), .B(n15039), .Z(n15041) );
  NOR U15414 ( .A(n15042), .B(n15041), .Z(n15043) );
  NAND U15415 ( .A(\stack[6][59] ), .B(n17311), .Z(n15045) );
  NANDN U15416 ( .A(n17311), .B(\stack[7][59] ), .Z(n15044) );
  NAND U15417 ( .A(n15045), .B(n15044), .Z(n2157) );
  NAND U15418 ( .A(\stack[5][59] ), .B(n17311), .Z(n15047) );
  NAND U15419 ( .A(n17305), .B(\stack[7][59] ), .Z(n15046) );
  AND U15420 ( .A(n15047), .B(n15046), .Z(n15049) );
  NAND U15421 ( .A(n17308), .B(\stack[6][59] ), .Z(n15048) );
  NAND U15422 ( .A(n15049), .B(n15048), .Z(n2158) );
  NAND U15423 ( .A(\stack[4][59] ), .B(n17311), .Z(n15051) );
  NAND U15424 ( .A(n17305), .B(\stack[6][59] ), .Z(n15050) );
  AND U15425 ( .A(n15051), .B(n15050), .Z(n15053) );
  NAND U15426 ( .A(n17308), .B(\stack[5][59] ), .Z(n15052) );
  NAND U15427 ( .A(n15053), .B(n15052), .Z(n2159) );
  NAND U15428 ( .A(\stack[3][59] ), .B(n17311), .Z(n15055) );
  NAND U15429 ( .A(n17305), .B(\stack[5][59] ), .Z(n15054) );
  AND U15430 ( .A(n15055), .B(n15054), .Z(n15057) );
  NAND U15431 ( .A(n17308), .B(\stack[4][59] ), .Z(n15056) );
  NAND U15432 ( .A(n15057), .B(n15056), .Z(n2160) );
  NAND U15433 ( .A(\stack[2][59] ), .B(n17311), .Z(n15059) );
  NAND U15434 ( .A(n17305), .B(\stack[4][59] ), .Z(n15058) );
  AND U15435 ( .A(n15059), .B(n15058), .Z(n15061) );
  NAND U15436 ( .A(n17308), .B(\stack[3][59] ), .Z(n15060) );
  NAND U15437 ( .A(n15061), .B(n15060), .Z(n2161) );
  NAND U15438 ( .A(n17311), .B(\stack[1][59] ), .Z(n15063) );
  NAND U15439 ( .A(n17305), .B(\stack[3][59] ), .Z(n15062) );
  AND U15440 ( .A(n15063), .B(n15062), .Z(n15065) );
  NAND U15441 ( .A(n17308), .B(\stack[2][59] ), .Z(n15064) );
  NAND U15442 ( .A(n15065), .B(n15064), .Z(n2162) );
  NAND U15443 ( .A(n17311), .B(o[59]), .Z(n15067) );
  NAND U15444 ( .A(n17305), .B(\stack[2][59] ), .Z(n15066) );
  AND U15445 ( .A(n15067), .B(n15066), .Z(n15069) );
  NAND U15446 ( .A(\stack[1][59] ), .B(n17308), .Z(n15068) );
  NAND U15447 ( .A(n15069), .B(n15068), .Z(n2163) );
  NAND U15448 ( .A(\stack[1][59] ), .B(n17313), .Z(n15070) );
  NAND U15449 ( .A(n17317), .B(n15070), .Z(n15071) );
  AND U15450 ( .A(o[59]), .B(n15071), .Z(n15080) );
  NAND U15451 ( .A(x[59]), .B(n17311), .Z(n15073) );
  NAND U15452 ( .A(\stack[1][59] ), .B(n17318), .Z(n15072) );
  AND U15453 ( .A(n15073), .B(n15072), .Z(n15078) );
  XNOR U15454 ( .A(n15075), .B(n15074), .Z(n15076) );
  NANDN U15455 ( .A(n17294), .B(n15076), .Z(n15077) );
  NAND U15456 ( .A(n15078), .B(n15077), .Z(n15079) );
  NOR U15457 ( .A(n15080), .B(n15079), .Z(n15081) );
  NAND U15458 ( .A(\stack[6][58] ), .B(n17311), .Z(n15083) );
  NANDN U15459 ( .A(n17311), .B(\stack[7][58] ), .Z(n15082) );
  NAND U15460 ( .A(n15083), .B(n15082), .Z(n2165) );
  NAND U15461 ( .A(\stack[5][58] ), .B(n17311), .Z(n15085) );
  NAND U15462 ( .A(n17305), .B(\stack[7][58] ), .Z(n15084) );
  AND U15463 ( .A(n15085), .B(n15084), .Z(n15087) );
  NAND U15464 ( .A(n17308), .B(\stack[6][58] ), .Z(n15086) );
  NAND U15465 ( .A(n15087), .B(n15086), .Z(n2166) );
  NAND U15466 ( .A(\stack[4][58] ), .B(n17311), .Z(n15089) );
  NAND U15467 ( .A(n17305), .B(\stack[6][58] ), .Z(n15088) );
  AND U15468 ( .A(n15089), .B(n15088), .Z(n15091) );
  NAND U15469 ( .A(n17308), .B(\stack[5][58] ), .Z(n15090) );
  NAND U15470 ( .A(n15091), .B(n15090), .Z(n2167) );
  NAND U15471 ( .A(\stack[3][58] ), .B(n17311), .Z(n15093) );
  NAND U15472 ( .A(n17305), .B(\stack[5][58] ), .Z(n15092) );
  AND U15473 ( .A(n15093), .B(n15092), .Z(n15095) );
  NAND U15474 ( .A(n17308), .B(\stack[4][58] ), .Z(n15094) );
  NAND U15475 ( .A(n15095), .B(n15094), .Z(n2168) );
  NAND U15476 ( .A(\stack[2][58] ), .B(n17311), .Z(n15097) );
  NAND U15477 ( .A(n17305), .B(\stack[4][58] ), .Z(n15096) );
  AND U15478 ( .A(n15097), .B(n15096), .Z(n15099) );
  NAND U15479 ( .A(n17308), .B(\stack[3][58] ), .Z(n15098) );
  NAND U15480 ( .A(n15099), .B(n15098), .Z(n2169) );
  NAND U15481 ( .A(n17311), .B(\stack[1][58] ), .Z(n15101) );
  NAND U15482 ( .A(n17305), .B(\stack[3][58] ), .Z(n15100) );
  AND U15483 ( .A(n15101), .B(n15100), .Z(n15103) );
  NAND U15484 ( .A(n17308), .B(\stack[2][58] ), .Z(n15102) );
  NAND U15485 ( .A(n15103), .B(n15102), .Z(n2170) );
  NAND U15486 ( .A(n17311), .B(o[58]), .Z(n15105) );
  NAND U15487 ( .A(n17305), .B(\stack[2][58] ), .Z(n15104) );
  AND U15488 ( .A(n15105), .B(n15104), .Z(n15107) );
  NAND U15489 ( .A(\stack[1][58] ), .B(n17308), .Z(n15106) );
  NAND U15490 ( .A(n15107), .B(n15106), .Z(n2171) );
  NAND U15491 ( .A(\stack[1][58] ), .B(n17313), .Z(n15108) );
  NAND U15492 ( .A(n17317), .B(n15108), .Z(n15109) );
  AND U15493 ( .A(o[58]), .B(n15109), .Z(n15118) );
  NAND U15494 ( .A(x[58]), .B(n17311), .Z(n15111) );
  NAND U15495 ( .A(\stack[1][58] ), .B(n17318), .Z(n15110) );
  AND U15496 ( .A(n15111), .B(n15110), .Z(n15116) );
  XNOR U15497 ( .A(n15113), .B(n15112), .Z(n15114) );
  NANDN U15498 ( .A(n17294), .B(n15114), .Z(n15115) );
  NAND U15499 ( .A(n15116), .B(n15115), .Z(n15117) );
  NOR U15500 ( .A(n15118), .B(n15117), .Z(n15119) );
  NAND U15501 ( .A(\stack[6][57] ), .B(n17311), .Z(n15121) );
  NANDN U15502 ( .A(n17311), .B(\stack[7][57] ), .Z(n15120) );
  NAND U15503 ( .A(n15121), .B(n15120), .Z(n2173) );
  NAND U15504 ( .A(\stack[5][57] ), .B(n17311), .Z(n15123) );
  NAND U15505 ( .A(n17305), .B(\stack[7][57] ), .Z(n15122) );
  AND U15506 ( .A(n15123), .B(n15122), .Z(n15125) );
  NAND U15507 ( .A(n17308), .B(\stack[6][57] ), .Z(n15124) );
  NAND U15508 ( .A(n15125), .B(n15124), .Z(n2174) );
  NAND U15509 ( .A(\stack[4][57] ), .B(n17311), .Z(n15127) );
  NAND U15510 ( .A(n17305), .B(\stack[6][57] ), .Z(n15126) );
  AND U15511 ( .A(n15127), .B(n15126), .Z(n15129) );
  NAND U15512 ( .A(n17308), .B(\stack[5][57] ), .Z(n15128) );
  NAND U15513 ( .A(n15129), .B(n15128), .Z(n2175) );
  NAND U15514 ( .A(\stack[3][57] ), .B(n17311), .Z(n15131) );
  NAND U15515 ( .A(n17305), .B(\stack[5][57] ), .Z(n15130) );
  AND U15516 ( .A(n15131), .B(n15130), .Z(n15133) );
  NAND U15517 ( .A(n17308), .B(\stack[4][57] ), .Z(n15132) );
  NAND U15518 ( .A(n15133), .B(n15132), .Z(n2176) );
  NAND U15519 ( .A(\stack[2][57] ), .B(n17311), .Z(n15135) );
  NAND U15520 ( .A(n17305), .B(\stack[4][57] ), .Z(n15134) );
  AND U15521 ( .A(n15135), .B(n15134), .Z(n15137) );
  NAND U15522 ( .A(n17308), .B(\stack[3][57] ), .Z(n15136) );
  NAND U15523 ( .A(n15137), .B(n15136), .Z(n2177) );
  NAND U15524 ( .A(n17311), .B(\stack[1][57] ), .Z(n15139) );
  NAND U15525 ( .A(n17305), .B(\stack[3][57] ), .Z(n15138) );
  AND U15526 ( .A(n15139), .B(n15138), .Z(n15141) );
  NAND U15527 ( .A(n17308), .B(\stack[2][57] ), .Z(n15140) );
  NAND U15528 ( .A(n15141), .B(n15140), .Z(n2178) );
  NAND U15529 ( .A(n17311), .B(o[57]), .Z(n15143) );
  NAND U15530 ( .A(n17305), .B(\stack[2][57] ), .Z(n15142) );
  AND U15531 ( .A(n15143), .B(n15142), .Z(n15145) );
  NAND U15532 ( .A(\stack[1][57] ), .B(n17308), .Z(n15144) );
  NAND U15533 ( .A(n15145), .B(n15144), .Z(n2179) );
  NAND U15534 ( .A(\stack[1][57] ), .B(n17313), .Z(n15146) );
  NAND U15535 ( .A(n17317), .B(n15146), .Z(n15147) );
  AND U15536 ( .A(o[57]), .B(n15147), .Z(n15156) );
  NAND U15537 ( .A(x[57]), .B(n17311), .Z(n15149) );
  NAND U15538 ( .A(\stack[1][57] ), .B(n17318), .Z(n15148) );
  AND U15539 ( .A(n15149), .B(n15148), .Z(n15154) );
  XNOR U15540 ( .A(n15151), .B(n15150), .Z(n15152) );
  NANDN U15541 ( .A(n17294), .B(n15152), .Z(n15153) );
  NAND U15542 ( .A(n15154), .B(n15153), .Z(n15155) );
  NOR U15543 ( .A(n15156), .B(n15155), .Z(n15157) );
  NAND U15544 ( .A(\stack[6][56] ), .B(n17311), .Z(n15159) );
  NANDN U15545 ( .A(n17311), .B(\stack[7][56] ), .Z(n15158) );
  NAND U15546 ( .A(n15159), .B(n15158), .Z(n2181) );
  NAND U15547 ( .A(\stack[5][56] ), .B(n17311), .Z(n15161) );
  NAND U15548 ( .A(n17305), .B(\stack[7][56] ), .Z(n15160) );
  AND U15549 ( .A(n15161), .B(n15160), .Z(n15163) );
  NAND U15550 ( .A(n17308), .B(\stack[6][56] ), .Z(n15162) );
  NAND U15551 ( .A(n15163), .B(n15162), .Z(n2182) );
  NAND U15552 ( .A(\stack[4][56] ), .B(n17311), .Z(n15165) );
  NAND U15553 ( .A(n17305), .B(\stack[6][56] ), .Z(n15164) );
  AND U15554 ( .A(n15165), .B(n15164), .Z(n15167) );
  NAND U15555 ( .A(n17308), .B(\stack[5][56] ), .Z(n15166) );
  NAND U15556 ( .A(n15167), .B(n15166), .Z(n2183) );
  NAND U15557 ( .A(\stack[3][56] ), .B(n17311), .Z(n15169) );
  NAND U15558 ( .A(n17305), .B(\stack[5][56] ), .Z(n15168) );
  AND U15559 ( .A(n15169), .B(n15168), .Z(n15171) );
  NAND U15560 ( .A(n17308), .B(\stack[4][56] ), .Z(n15170) );
  NAND U15561 ( .A(n15171), .B(n15170), .Z(n2184) );
  NAND U15562 ( .A(\stack[2][56] ), .B(n17311), .Z(n15173) );
  NAND U15563 ( .A(n17305), .B(\stack[4][56] ), .Z(n15172) );
  AND U15564 ( .A(n15173), .B(n15172), .Z(n15175) );
  NAND U15565 ( .A(n17308), .B(\stack[3][56] ), .Z(n15174) );
  NAND U15566 ( .A(n15175), .B(n15174), .Z(n2185) );
  NAND U15567 ( .A(n17311), .B(\stack[1][56] ), .Z(n15177) );
  NAND U15568 ( .A(n17305), .B(\stack[3][56] ), .Z(n15176) );
  AND U15569 ( .A(n15177), .B(n15176), .Z(n15179) );
  NAND U15570 ( .A(n17308), .B(\stack[2][56] ), .Z(n15178) );
  NAND U15571 ( .A(n15179), .B(n15178), .Z(n2186) );
  NAND U15572 ( .A(n17311), .B(o[56]), .Z(n15181) );
  NAND U15573 ( .A(n17305), .B(\stack[2][56] ), .Z(n15180) );
  AND U15574 ( .A(n15181), .B(n15180), .Z(n15183) );
  NAND U15575 ( .A(\stack[1][56] ), .B(n17308), .Z(n15182) );
  NAND U15576 ( .A(n15183), .B(n15182), .Z(n2187) );
  NAND U15577 ( .A(\stack[1][56] ), .B(n17313), .Z(n15184) );
  NAND U15578 ( .A(n17317), .B(n15184), .Z(n15185) );
  AND U15579 ( .A(o[56]), .B(n15185), .Z(n15194) );
  NAND U15580 ( .A(x[56]), .B(n17311), .Z(n15187) );
  NAND U15581 ( .A(\stack[1][56] ), .B(n17318), .Z(n15186) );
  AND U15582 ( .A(n15187), .B(n15186), .Z(n15192) );
  XNOR U15583 ( .A(n15189), .B(n15188), .Z(n15190) );
  NANDN U15584 ( .A(n17294), .B(n15190), .Z(n15191) );
  NAND U15585 ( .A(n15192), .B(n15191), .Z(n15193) );
  NOR U15586 ( .A(n15194), .B(n15193), .Z(n15195) );
  NAND U15587 ( .A(\stack[6][55] ), .B(n17311), .Z(n15197) );
  NANDN U15588 ( .A(n17311), .B(\stack[7][55] ), .Z(n15196) );
  NAND U15589 ( .A(n15197), .B(n15196), .Z(n2189) );
  NAND U15590 ( .A(\stack[5][55] ), .B(n17311), .Z(n15199) );
  NAND U15591 ( .A(n17305), .B(\stack[7][55] ), .Z(n15198) );
  AND U15592 ( .A(n15199), .B(n15198), .Z(n15201) );
  NAND U15593 ( .A(n17308), .B(\stack[6][55] ), .Z(n15200) );
  NAND U15594 ( .A(n15201), .B(n15200), .Z(n2190) );
  NAND U15595 ( .A(\stack[4][55] ), .B(n17311), .Z(n15203) );
  NAND U15596 ( .A(n17305), .B(\stack[6][55] ), .Z(n15202) );
  AND U15597 ( .A(n15203), .B(n15202), .Z(n15205) );
  NAND U15598 ( .A(n17308), .B(\stack[5][55] ), .Z(n15204) );
  NAND U15599 ( .A(n15205), .B(n15204), .Z(n2191) );
  NAND U15600 ( .A(\stack[3][55] ), .B(n17311), .Z(n15207) );
  NAND U15601 ( .A(n17305), .B(\stack[5][55] ), .Z(n15206) );
  AND U15602 ( .A(n15207), .B(n15206), .Z(n15209) );
  NAND U15603 ( .A(n17308), .B(\stack[4][55] ), .Z(n15208) );
  NAND U15604 ( .A(n15209), .B(n15208), .Z(n2192) );
  NAND U15605 ( .A(\stack[2][55] ), .B(n17311), .Z(n15211) );
  NAND U15606 ( .A(n17305), .B(\stack[4][55] ), .Z(n15210) );
  AND U15607 ( .A(n15211), .B(n15210), .Z(n15213) );
  NAND U15608 ( .A(n17308), .B(\stack[3][55] ), .Z(n15212) );
  NAND U15609 ( .A(n15213), .B(n15212), .Z(n2193) );
  NAND U15610 ( .A(n17311), .B(\stack[1][55] ), .Z(n15215) );
  NAND U15611 ( .A(n17305), .B(\stack[3][55] ), .Z(n15214) );
  AND U15612 ( .A(n15215), .B(n15214), .Z(n15217) );
  NAND U15613 ( .A(n17308), .B(\stack[2][55] ), .Z(n15216) );
  NAND U15614 ( .A(n15217), .B(n15216), .Z(n2194) );
  NAND U15615 ( .A(n17311), .B(o[55]), .Z(n15219) );
  NAND U15616 ( .A(n17305), .B(\stack[2][55] ), .Z(n15218) );
  AND U15617 ( .A(n15219), .B(n15218), .Z(n15221) );
  NAND U15618 ( .A(\stack[1][55] ), .B(n17308), .Z(n15220) );
  NAND U15619 ( .A(n15221), .B(n15220), .Z(n2195) );
  NAND U15620 ( .A(\stack[1][55] ), .B(n17313), .Z(n15222) );
  NAND U15621 ( .A(n17317), .B(n15222), .Z(n15223) );
  AND U15622 ( .A(o[55]), .B(n15223), .Z(n15232) );
  NAND U15623 ( .A(x[55]), .B(n17311), .Z(n15225) );
  NAND U15624 ( .A(\stack[1][55] ), .B(n17318), .Z(n15224) );
  AND U15625 ( .A(n15225), .B(n15224), .Z(n15230) );
  XNOR U15626 ( .A(n15227), .B(n15226), .Z(n15228) );
  NANDN U15627 ( .A(n17294), .B(n15228), .Z(n15229) );
  NAND U15628 ( .A(n15230), .B(n15229), .Z(n15231) );
  NOR U15629 ( .A(n15232), .B(n15231), .Z(n15233) );
  NAND U15630 ( .A(\stack[6][54] ), .B(n17311), .Z(n15235) );
  NANDN U15631 ( .A(n17311), .B(\stack[7][54] ), .Z(n15234) );
  NAND U15632 ( .A(n15235), .B(n15234), .Z(n2197) );
  NAND U15633 ( .A(\stack[5][54] ), .B(n17311), .Z(n15237) );
  NAND U15634 ( .A(n17305), .B(\stack[7][54] ), .Z(n15236) );
  AND U15635 ( .A(n15237), .B(n15236), .Z(n15239) );
  NAND U15636 ( .A(n17308), .B(\stack[6][54] ), .Z(n15238) );
  NAND U15637 ( .A(n15239), .B(n15238), .Z(n2198) );
  NAND U15638 ( .A(\stack[4][54] ), .B(n17311), .Z(n15241) );
  NAND U15639 ( .A(n17305), .B(\stack[6][54] ), .Z(n15240) );
  AND U15640 ( .A(n15241), .B(n15240), .Z(n15243) );
  NAND U15641 ( .A(n17308), .B(\stack[5][54] ), .Z(n15242) );
  NAND U15642 ( .A(n15243), .B(n15242), .Z(n2199) );
  NAND U15643 ( .A(\stack[3][54] ), .B(n17311), .Z(n15245) );
  NAND U15644 ( .A(n17305), .B(\stack[5][54] ), .Z(n15244) );
  AND U15645 ( .A(n15245), .B(n15244), .Z(n15247) );
  NAND U15646 ( .A(n17308), .B(\stack[4][54] ), .Z(n15246) );
  NAND U15647 ( .A(n15247), .B(n15246), .Z(n2200) );
  NAND U15648 ( .A(\stack[2][54] ), .B(n17311), .Z(n15249) );
  NAND U15649 ( .A(n17305), .B(\stack[4][54] ), .Z(n15248) );
  AND U15650 ( .A(n15249), .B(n15248), .Z(n15251) );
  NAND U15651 ( .A(n17308), .B(\stack[3][54] ), .Z(n15250) );
  NAND U15652 ( .A(n15251), .B(n15250), .Z(n2201) );
  NAND U15653 ( .A(n17311), .B(\stack[1][54] ), .Z(n15253) );
  NAND U15654 ( .A(n17305), .B(\stack[3][54] ), .Z(n15252) );
  AND U15655 ( .A(n15253), .B(n15252), .Z(n15255) );
  NAND U15656 ( .A(n17308), .B(\stack[2][54] ), .Z(n15254) );
  NAND U15657 ( .A(n15255), .B(n15254), .Z(n2202) );
  NAND U15658 ( .A(n17311), .B(o[54]), .Z(n15257) );
  NAND U15659 ( .A(n17305), .B(\stack[2][54] ), .Z(n15256) );
  AND U15660 ( .A(n15257), .B(n15256), .Z(n15259) );
  NAND U15661 ( .A(\stack[1][54] ), .B(n17308), .Z(n15258) );
  NAND U15662 ( .A(n15259), .B(n15258), .Z(n2203) );
  NAND U15663 ( .A(\stack[1][54] ), .B(n17313), .Z(n15260) );
  NAND U15664 ( .A(n17317), .B(n15260), .Z(n15261) );
  AND U15665 ( .A(o[54]), .B(n15261), .Z(n15270) );
  NAND U15666 ( .A(x[54]), .B(n17311), .Z(n15263) );
  NAND U15667 ( .A(\stack[1][54] ), .B(n17318), .Z(n15262) );
  AND U15668 ( .A(n15263), .B(n15262), .Z(n15268) );
  XNOR U15669 ( .A(n15265), .B(n15264), .Z(n15266) );
  NANDN U15670 ( .A(n17294), .B(n15266), .Z(n15267) );
  NAND U15671 ( .A(n15268), .B(n15267), .Z(n15269) );
  NOR U15672 ( .A(n15270), .B(n15269), .Z(n15271) );
  NAND U15673 ( .A(\stack[6][53] ), .B(n17311), .Z(n15273) );
  NANDN U15674 ( .A(n17311), .B(\stack[7][53] ), .Z(n15272) );
  NAND U15675 ( .A(n15273), .B(n15272), .Z(n2205) );
  NAND U15676 ( .A(\stack[5][53] ), .B(n17311), .Z(n15275) );
  NAND U15677 ( .A(n17305), .B(\stack[7][53] ), .Z(n15274) );
  AND U15678 ( .A(n15275), .B(n15274), .Z(n15277) );
  NAND U15679 ( .A(n17308), .B(\stack[6][53] ), .Z(n15276) );
  NAND U15680 ( .A(n15277), .B(n15276), .Z(n2206) );
  NAND U15681 ( .A(\stack[4][53] ), .B(n17311), .Z(n15279) );
  NAND U15682 ( .A(n17305), .B(\stack[6][53] ), .Z(n15278) );
  AND U15683 ( .A(n15279), .B(n15278), .Z(n15281) );
  NAND U15684 ( .A(n17308), .B(\stack[5][53] ), .Z(n15280) );
  NAND U15685 ( .A(n15281), .B(n15280), .Z(n2207) );
  NAND U15686 ( .A(\stack[3][53] ), .B(n17311), .Z(n15283) );
  NAND U15687 ( .A(n17305), .B(\stack[5][53] ), .Z(n15282) );
  AND U15688 ( .A(n15283), .B(n15282), .Z(n15285) );
  NAND U15689 ( .A(n17308), .B(\stack[4][53] ), .Z(n15284) );
  NAND U15690 ( .A(n15285), .B(n15284), .Z(n2208) );
  NAND U15691 ( .A(\stack[2][53] ), .B(n17311), .Z(n15287) );
  NAND U15692 ( .A(n17305), .B(\stack[4][53] ), .Z(n15286) );
  AND U15693 ( .A(n15287), .B(n15286), .Z(n15289) );
  NAND U15694 ( .A(n17308), .B(\stack[3][53] ), .Z(n15288) );
  NAND U15695 ( .A(n15289), .B(n15288), .Z(n2209) );
  NAND U15696 ( .A(n17311), .B(\stack[1][53] ), .Z(n15291) );
  NAND U15697 ( .A(n17305), .B(\stack[3][53] ), .Z(n15290) );
  AND U15698 ( .A(n15291), .B(n15290), .Z(n15293) );
  NAND U15699 ( .A(n17308), .B(\stack[2][53] ), .Z(n15292) );
  NAND U15700 ( .A(n15293), .B(n15292), .Z(n2210) );
  NAND U15701 ( .A(n17311), .B(o[53]), .Z(n15295) );
  NAND U15702 ( .A(n17305), .B(\stack[2][53] ), .Z(n15294) );
  AND U15703 ( .A(n15295), .B(n15294), .Z(n15297) );
  NAND U15704 ( .A(\stack[1][53] ), .B(n17308), .Z(n15296) );
  NAND U15705 ( .A(n15297), .B(n15296), .Z(n2211) );
  NAND U15706 ( .A(\stack[1][53] ), .B(n17313), .Z(n15298) );
  NAND U15707 ( .A(n17317), .B(n15298), .Z(n15299) );
  AND U15708 ( .A(o[53]), .B(n15299), .Z(n15308) );
  NAND U15709 ( .A(x[53]), .B(n17311), .Z(n15301) );
  NAND U15710 ( .A(\stack[1][53] ), .B(n17318), .Z(n15300) );
  AND U15711 ( .A(n15301), .B(n15300), .Z(n15306) );
  XNOR U15712 ( .A(n15303), .B(n15302), .Z(n15304) );
  NANDN U15713 ( .A(n17294), .B(n15304), .Z(n15305) );
  NAND U15714 ( .A(n15306), .B(n15305), .Z(n15307) );
  NOR U15715 ( .A(n15308), .B(n15307), .Z(n15309) );
  NAND U15716 ( .A(\stack[6][52] ), .B(n17311), .Z(n15311) );
  NANDN U15717 ( .A(n17311), .B(\stack[7][52] ), .Z(n15310) );
  NAND U15718 ( .A(n15311), .B(n15310), .Z(n2213) );
  NAND U15719 ( .A(\stack[5][52] ), .B(n17311), .Z(n15313) );
  NAND U15720 ( .A(n17305), .B(\stack[7][52] ), .Z(n15312) );
  AND U15721 ( .A(n15313), .B(n15312), .Z(n15315) );
  NAND U15722 ( .A(n17308), .B(\stack[6][52] ), .Z(n15314) );
  NAND U15723 ( .A(n15315), .B(n15314), .Z(n2214) );
  NAND U15724 ( .A(\stack[4][52] ), .B(n17311), .Z(n15317) );
  NAND U15725 ( .A(n17305), .B(\stack[6][52] ), .Z(n15316) );
  AND U15726 ( .A(n15317), .B(n15316), .Z(n15319) );
  NAND U15727 ( .A(n17308), .B(\stack[5][52] ), .Z(n15318) );
  NAND U15728 ( .A(n15319), .B(n15318), .Z(n2215) );
  NAND U15729 ( .A(\stack[3][52] ), .B(n17311), .Z(n15321) );
  NAND U15730 ( .A(n17305), .B(\stack[5][52] ), .Z(n15320) );
  AND U15731 ( .A(n15321), .B(n15320), .Z(n15323) );
  NAND U15732 ( .A(n17308), .B(\stack[4][52] ), .Z(n15322) );
  NAND U15733 ( .A(n15323), .B(n15322), .Z(n2216) );
  NAND U15734 ( .A(\stack[2][52] ), .B(n17311), .Z(n15325) );
  NAND U15735 ( .A(n17305), .B(\stack[4][52] ), .Z(n15324) );
  AND U15736 ( .A(n15325), .B(n15324), .Z(n15327) );
  NAND U15737 ( .A(n17308), .B(\stack[3][52] ), .Z(n15326) );
  NAND U15738 ( .A(n15327), .B(n15326), .Z(n2217) );
  NAND U15739 ( .A(n17311), .B(\stack[1][52] ), .Z(n15329) );
  NAND U15740 ( .A(n17305), .B(\stack[3][52] ), .Z(n15328) );
  AND U15741 ( .A(n15329), .B(n15328), .Z(n15331) );
  NAND U15742 ( .A(n17308), .B(\stack[2][52] ), .Z(n15330) );
  NAND U15743 ( .A(n15331), .B(n15330), .Z(n2218) );
  NAND U15744 ( .A(n17311), .B(o[52]), .Z(n15333) );
  NAND U15745 ( .A(n17305), .B(\stack[2][52] ), .Z(n15332) );
  AND U15746 ( .A(n15333), .B(n15332), .Z(n15335) );
  NAND U15747 ( .A(\stack[1][52] ), .B(n17308), .Z(n15334) );
  NAND U15748 ( .A(n15335), .B(n15334), .Z(n2219) );
  NAND U15749 ( .A(\stack[1][52] ), .B(n17313), .Z(n15336) );
  NAND U15750 ( .A(n17317), .B(n15336), .Z(n15337) );
  AND U15751 ( .A(o[52]), .B(n15337), .Z(n15346) );
  NAND U15752 ( .A(x[52]), .B(n17311), .Z(n15339) );
  NAND U15753 ( .A(\stack[1][52] ), .B(n17318), .Z(n15338) );
  AND U15754 ( .A(n15339), .B(n15338), .Z(n15344) );
  XNOR U15755 ( .A(n15341), .B(n15340), .Z(n15342) );
  NANDN U15756 ( .A(n17294), .B(n15342), .Z(n15343) );
  NAND U15757 ( .A(n15344), .B(n15343), .Z(n15345) );
  NOR U15758 ( .A(n15346), .B(n15345), .Z(n15347) );
  NAND U15759 ( .A(\stack[6][51] ), .B(n17311), .Z(n15349) );
  NANDN U15760 ( .A(n17311), .B(\stack[7][51] ), .Z(n15348) );
  NAND U15761 ( .A(n15349), .B(n15348), .Z(n2221) );
  NAND U15762 ( .A(\stack[5][51] ), .B(n17311), .Z(n15351) );
  NAND U15763 ( .A(n17305), .B(\stack[7][51] ), .Z(n15350) );
  AND U15764 ( .A(n15351), .B(n15350), .Z(n15353) );
  NAND U15765 ( .A(n17308), .B(\stack[6][51] ), .Z(n15352) );
  NAND U15766 ( .A(n15353), .B(n15352), .Z(n2222) );
  NAND U15767 ( .A(\stack[4][51] ), .B(n17311), .Z(n15355) );
  NAND U15768 ( .A(n17305), .B(\stack[6][51] ), .Z(n15354) );
  AND U15769 ( .A(n15355), .B(n15354), .Z(n15357) );
  NAND U15770 ( .A(n17308), .B(\stack[5][51] ), .Z(n15356) );
  NAND U15771 ( .A(n15357), .B(n15356), .Z(n2223) );
  NAND U15772 ( .A(\stack[3][51] ), .B(n17311), .Z(n15359) );
  NAND U15773 ( .A(n17305), .B(\stack[5][51] ), .Z(n15358) );
  AND U15774 ( .A(n15359), .B(n15358), .Z(n15361) );
  NAND U15775 ( .A(n17308), .B(\stack[4][51] ), .Z(n15360) );
  NAND U15776 ( .A(n15361), .B(n15360), .Z(n2224) );
  NAND U15777 ( .A(\stack[2][51] ), .B(n17311), .Z(n15363) );
  NAND U15778 ( .A(n17305), .B(\stack[4][51] ), .Z(n15362) );
  AND U15779 ( .A(n15363), .B(n15362), .Z(n15365) );
  NAND U15780 ( .A(n17308), .B(\stack[3][51] ), .Z(n15364) );
  NAND U15781 ( .A(n15365), .B(n15364), .Z(n2225) );
  NAND U15782 ( .A(n17311), .B(\stack[1][51] ), .Z(n15367) );
  NAND U15783 ( .A(n17305), .B(\stack[3][51] ), .Z(n15366) );
  AND U15784 ( .A(n15367), .B(n15366), .Z(n15369) );
  NAND U15785 ( .A(n17308), .B(\stack[2][51] ), .Z(n15368) );
  NAND U15786 ( .A(n15369), .B(n15368), .Z(n2226) );
  NAND U15787 ( .A(n17311), .B(o[51]), .Z(n15371) );
  NAND U15788 ( .A(n17305), .B(\stack[2][51] ), .Z(n15370) );
  AND U15789 ( .A(n15371), .B(n15370), .Z(n15373) );
  NAND U15790 ( .A(\stack[1][51] ), .B(n17308), .Z(n15372) );
  NAND U15791 ( .A(n15373), .B(n15372), .Z(n2227) );
  NAND U15792 ( .A(\stack[1][51] ), .B(n17313), .Z(n15374) );
  NAND U15793 ( .A(n17317), .B(n15374), .Z(n15375) );
  AND U15794 ( .A(o[51]), .B(n15375), .Z(n15384) );
  NAND U15795 ( .A(x[51]), .B(n17311), .Z(n15377) );
  NAND U15796 ( .A(\stack[1][51] ), .B(n17318), .Z(n15376) );
  AND U15797 ( .A(n15377), .B(n15376), .Z(n15382) );
  XNOR U15798 ( .A(n15379), .B(n15378), .Z(n15380) );
  NANDN U15799 ( .A(n17294), .B(n15380), .Z(n15381) );
  NAND U15800 ( .A(n15382), .B(n15381), .Z(n15383) );
  NOR U15801 ( .A(n15384), .B(n15383), .Z(n15385) );
  NAND U15802 ( .A(\stack[6][50] ), .B(n17311), .Z(n15387) );
  NANDN U15803 ( .A(n17311), .B(\stack[7][50] ), .Z(n15386) );
  NAND U15804 ( .A(n15387), .B(n15386), .Z(n2229) );
  NAND U15805 ( .A(\stack[5][50] ), .B(n17311), .Z(n15389) );
  NAND U15806 ( .A(n17305), .B(\stack[7][50] ), .Z(n15388) );
  AND U15807 ( .A(n15389), .B(n15388), .Z(n15391) );
  NAND U15808 ( .A(n17308), .B(\stack[6][50] ), .Z(n15390) );
  NAND U15809 ( .A(n15391), .B(n15390), .Z(n2230) );
  NAND U15810 ( .A(\stack[4][50] ), .B(n17311), .Z(n15393) );
  NAND U15811 ( .A(n17305), .B(\stack[6][50] ), .Z(n15392) );
  AND U15812 ( .A(n15393), .B(n15392), .Z(n15395) );
  NAND U15813 ( .A(n17308), .B(\stack[5][50] ), .Z(n15394) );
  NAND U15814 ( .A(n15395), .B(n15394), .Z(n2231) );
  NAND U15815 ( .A(\stack[3][50] ), .B(n17311), .Z(n15397) );
  NAND U15816 ( .A(n17305), .B(\stack[5][50] ), .Z(n15396) );
  AND U15817 ( .A(n15397), .B(n15396), .Z(n15399) );
  NAND U15818 ( .A(n17308), .B(\stack[4][50] ), .Z(n15398) );
  NAND U15819 ( .A(n15399), .B(n15398), .Z(n2232) );
  NAND U15820 ( .A(\stack[2][50] ), .B(n17311), .Z(n15401) );
  NAND U15821 ( .A(n17305), .B(\stack[4][50] ), .Z(n15400) );
  AND U15822 ( .A(n15401), .B(n15400), .Z(n15403) );
  NAND U15823 ( .A(n17308), .B(\stack[3][50] ), .Z(n15402) );
  NAND U15824 ( .A(n15403), .B(n15402), .Z(n2233) );
  NAND U15825 ( .A(n17311), .B(\stack[1][50] ), .Z(n15405) );
  NAND U15826 ( .A(n17305), .B(\stack[3][50] ), .Z(n15404) );
  AND U15827 ( .A(n15405), .B(n15404), .Z(n15407) );
  NAND U15828 ( .A(n17308), .B(\stack[2][50] ), .Z(n15406) );
  NAND U15829 ( .A(n15407), .B(n15406), .Z(n2234) );
  NAND U15830 ( .A(n17311), .B(o[50]), .Z(n15409) );
  NAND U15831 ( .A(n17305), .B(\stack[2][50] ), .Z(n15408) );
  AND U15832 ( .A(n15409), .B(n15408), .Z(n15411) );
  NAND U15833 ( .A(\stack[1][50] ), .B(n17308), .Z(n15410) );
  NAND U15834 ( .A(n15411), .B(n15410), .Z(n2235) );
  NAND U15835 ( .A(\stack[1][50] ), .B(n17313), .Z(n15412) );
  NAND U15836 ( .A(n17317), .B(n15412), .Z(n15413) );
  AND U15837 ( .A(o[50]), .B(n15413), .Z(n15422) );
  NAND U15838 ( .A(x[50]), .B(n17311), .Z(n15415) );
  NAND U15839 ( .A(\stack[1][50] ), .B(n17318), .Z(n15414) );
  AND U15840 ( .A(n15415), .B(n15414), .Z(n15420) );
  XNOR U15841 ( .A(n15417), .B(n15416), .Z(n15418) );
  NANDN U15842 ( .A(n17294), .B(n15418), .Z(n15419) );
  NAND U15843 ( .A(n15420), .B(n15419), .Z(n15421) );
  NOR U15844 ( .A(n15422), .B(n15421), .Z(n15423) );
  NAND U15845 ( .A(\stack[6][49] ), .B(n17311), .Z(n15425) );
  NANDN U15846 ( .A(n17311), .B(\stack[7][49] ), .Z(n15424) );
  NAND U15847 ( .A(n15425), .B(n15424), .Z(n2237) );
  NAND U15848 ( .A(\stack[5][49] ), .B(n17311), .Z(n15427) );
  NAND U15849 ( .A(n17305), .B(\stack[7][49] ), .Z(n15426) );
  AND U15850 ( .A(n15427), .B(n15426), .Z(n15429) );
  NAND U15851 ( .A(n17308), .B(\stack[6][49] ), .Z(n15428) );
  NAND U15852 ( .A(n15429), .B(n15428), .Z(n2238) );
  NAND U15853 ( .A(\stack[4][49] ), .B(n17311), .Z(n15431) );
  NAND U15854 ( .A(n17305), .B(\stack[6][49] ), .Z(n15430) );
  AND U15855 ( .A(n15431), .B(n15430), .Z(n15433) );
  NAND U15856 ( .A(n17308), .B(\stack[5][49] ), .Z(n15432) );
  NAND U15857 ( .A(n15433), .B(n15432), .Z(n2239) );
  NAND U15858 ( .A(\stack[3][49] ), .B(n17311), .Z(n15435) );
  NAND U15859 ( .A(n17305), .B(\stack[5][49] ), .Z(n15434) );
  AND U15860 ( .A(n15435), .B(n15434), .Z(n15437) );
  NAND U15861 ( .A(n17308), .B(\stack[4][49] ), .Z(n15436) );
  NAND U15862 ( .A(n15437), .B(n15436), .Z(n2240) );
  NAND U15863 ( .A(\stack[2][49] ), .B(n17311), .Z(n15439) );
  NAND U15864 ( .A(n17305), .B(\stack[4][49] ), .Z(n15438) );
  AND U15865 ( .A(n15439), .B(n15438), .Z(n15441) );
  NAND U15866 ( .A(n17308), .B(\stack[3][49] ), .Z(n15440) );
  NAND U15867 ( .A(n15441), .B(n15440), .Z(n2241) );
  NAND U15868 ( .A(n17311), .B(\stack[1][49] ), .Z(n15443) );
  NAND U15869 ( .A(n17305), .B(\stack[3][49] ), .Z(n15442) );
  AND U15870 ( .A(n15443), .B(n15442), .Z(n15445) );
  NAND U15871 ( .A(n17308), .B(\stack[2][49] ), .Z(n15444) );
  NAND U15872 ( .A(n15445), .B(n15444), .Z(n2242) );
  NAND U15873 ( .A(n17311), .B(o[49]), .Z(n15447) );
  NAND U15874 ( .A(n17305), .B(\stack[2][49] ), .Z(n15446) );
  AND U15875 ( .A(n15447), .B(n15446), .Z(n15449) );
  NAND U15876 ( .A(\stack[1][49] ), .B(n17308), .Z(n15448) );
  NAND U15877 ( .A(n15449), .B(n15448), .Z(n2243) );
  NAND U15878 ( .A(\stack[1][49] ), .B(n17313), .Z(n15450) );
  NAND U15879 ( .A(n17317), .B(n15450), .Z(n15451) );
  AND U15880 ( .A(o[49]), .B(n15451), .Z(n15460) );
  NAND U15881 ( .A(x[49]), .B(n17311), .Z(n15453) );
  NAND U15882 ( .A(\stack[1][49] ), .B(n17318), .Z(n15452) );
  AND U15883 ( .A(n15453), .B(n15452), .Z(n15458) );
  XNOR U15884 ( .A(n15455), .B(n15454), .Z(n15456) );
  NANDN U15885 ( .A(n17294), .B(n15456), .Z(n15457) );
  NAND U15886 ( .A(n15458), .B(n15457), .Z(n15459) );
  NOR U15887 ( .A(n15460), .B(n15459), .Z(n15461) );
  NAND U15888 ( .A(\stack[6][48] ), .B(n17311), .Z(n15463) );
  NANDN U15889 ( .A(n17311), .B(\stack[7][48] ), .Z(n15462) );
  NAND U15890 ( .A(n15463), .B(n15462), .Z(n2245) );
  NAND U15891 ( .A(\stack[5][48] ), .B(n17311), .Z(n15465) );
  NAND U15892 ( .A(n17305), .B(\stack[7][48] ), .Z(n15464) );
  AND U15893 ( .A(n15465), .B(n15464), .Z(n15467) );
  NAND U15894 ( .A(n17308), .B(\stack[6][48] ), .Z(n15466) );
  NAND U15895 ( .A(n15467), .B(n15466), .Z(n2246) );
  NAND U15896 ( .A(\stack[4][48] ), .B(n17311), .Z(n15469) );
  NAND U15897 ( .A(n17305), .B(\stack[6][48] ), .Z(n15468) );
  AND U15898 ( .A(n15469), .B(n15468), .Z(n15471) );
  NAND U15899 ( .A(n17308), .B(\stack[5][48] ), .Z(n15470) );
  NAND U15900 ( .A(n15471), .B(n15470), .Z(n2247) );
  NAND U15901 ( .A(\stack[3][48] ), .B(n17311), .Z(n15473) );
  NAND U15902 ( .A(n17305), .B(\stack[5][48] ), .Z(n15472) );
  AND U15903 ( .A(n15473), .B(n15472), .Z(n15475) );
  NAND U15904 ( .A(n17308), .B(\stack[4][48] ), .Z(n15474) );
  NAND U15905 ( .A(n15475), .B(n15474), .Z(n2248) );
  NAND U15906 ( .A(\stack[2][48] ), .B(n17311), .Z(n15477) );
  NAND U15907 ( .A(n17305), .B(\stack[4][48] ), .Z(n15476) );
  AND U15908 ( .A(n15477), .B(n15476), .Z(n15479) );
  NAND U15909 ( .A(n17308), .B(\stack[3][48] ), .Z(n15478) );
  NAND U15910 ( .A(n15479), .B(n15478), .Z(n2249) );
  NAND U15911 ( .A(n17311), .B(\stack[1][48] ), .Z(n15481) );
  NAND U15912 ( .A(n17305), .B(\stack[3][48] ), .Z(n15480) );
  AND U15913 ( .A(n15481), .B(n15480), .Z(n15483) );
  NAND U15914 ( .A(n17308), .B(\stack[2][48] ), .Z(n15482) );
  NAND U15915 ( .A(n15483), .B(n15482), .Z(n2250) );
  NAND U15916 ( .A(n17311), .B(o[48]), .Z(n15485) );
  NAND U15917 ( .A(n17305), .B(\stack[2][48] ), .Z(n15484) );
  AND U15918 ( .A(n15485), .B(n15484), .Z(n15487) );
  NAND U15919 ( .A(\stack[1][48] ), .B(n17308), .Z(n15486) );
  NAND U15920 ( .A(n15487), .B(n15486), .Z(n2251) );
  NAND U15921 ( .A(\stack[1][48] ), .B(n17313), .Z(n15488) );
  NAND U15922 ( .A(n17317), .B(n15488), .Z(n15489) );
  AND U15923 ( .A(o[48]), .B(n15489), .Z(n15498) );
  NAND U15924 ( .A(x[48]), .B(n17311), .Z(n15491) );
  NAND U15925 ( .A(\stack[1][48] ), .B(n17318), .Z(n15490) );
  AND U15926 ( .A(n15491), .B(n15490), .Z(n15496) );
  XNOR U15927 ( .A(n15493), .B(n15492), .Z(n15494) );
  NANDN U15928 ( .A(n17294), .B(n15494), .Z(n15495) );
  NAND U15929 ( .A(n15496), .B(n15495), .Z(n15497) );
  NOR U15930 ( .A(n15498), .B(n15497), .Z(n15499) );
  NAND U15931 ( .A(\stack[6][47] ), .B(n17311), .Z(n15501) );
  NANDN U15932 ( .A(n17311), .B(\stack[7][47] ), .Z(n15500) );
  NAND U15933 ( .A(n15501), .B(n15500), .Z(n2253) );
  NAND U15934 ( .A(\stack[5][47] ), .B(n17311), .Z(n15503) );
  NAND U15935 ( .A(n17305), .B(\stack[7][47] ), .Z(n15502) );
  AND U15936 ( .A(n15503), .B(n15502), .Z(n15505) );
  NAND U15937 ( .A(n17308), .B(\stack[6][47] ), .Z(n15504) );
  NAND U15938 ( .A(n15505), .B(n15504), .Z(n2254) );
  NAND U15939 ( .A(\stack[4][47] ), .B(n17311), .Z(n15507) );
  NAND U15940 ( .A(n17305), .B(\stack[6][47] ), .Z(n15506) );
  AND U15941 ( .A(n15507), .B(n15506), .Z(n15509) );
  NAND U15942 ( .A(n17308), .B(\stack[5][47] ), .Z(n15508) );
  NAND U15943 ( .A(n15509), .B(n15508), .Z(n2255) );
  NAND U15944 ( .A(\stack[3][47] ), .B(n17311), .Z(n15511) );
  NAND U15945 ( .A(n17305), .B(\stack[5][47] ), .Z(n15510) );
  AND U15946 ( .A(n15511), .B(n15510), .Z(n15513) );
  NAND U15947 ( .A(n17308), .B(\stack[4][47] ), .Z(n15512) );
  NAND U15948 ( .A(n15513), .B(n15512), .Z(n2256) );
  NAND U15949 ( .A(\stack[2][47] ), .B(n17311), .Z(n15515) );
  NAND U15950 ( .A(n17305), .B(\stack[4][47] ), .Z(n15514) );
  AND U15951 ( .A(n15515), .B(n15514), .Z(n15517) );
  NAND U15952 ( .A(n17308), .B(\stack[3][47] ), .Z(n15516) );
  NAND U15953 ( .A(n15517), .B(n15516), .Z(n2257) );
  NAND U15954 ( .A(n17311), .B(\stack[1][47] ), .Z(n15519) );
  NAND U15955 ( .A(n17305), .B(\stack[3][47] ), .Z(n15518) );
  AND U15956 ( .A(n15519), .B(n15518), .Z(n15521) );
  NAND U15957 ( .A(n17308), .B(\stack[2][47] ), .Z(n15520) );
  NAND U15958 ( .A(n15521), .B(n15520), .Z(n2258) );
  NAND U15959 ( .A(n17311), .B(o[47]), .Z(n15523) );
  NAND U15960 ( .A(n17305), .B(\stack[2][47] ), .Z(n15522) );
  AND U15961 ( .A(n15523), .B(n15522), .Z(n15525) );
  NAND U15962 ( .A(\stack[1][47] ), .B(n17308), .Z(n15524) );
  NAND U15963 ( .A(n15525), .B(n15524), .Z(n2259) );
  NAND U15964 ( .A(\stack[1][47] ), .B(n17313), .Z(n15526) );
  NAND U15965 ( .A(n17317), .B(n15526), .Z(n15527) );
  AND U15966 ( .A(o[47]), .B(n15527), .Z(n15536) );
  NAND U15967 ( .A(x[47]), .B(n17311), .Z(n15529) );
  NAND U15968 ( .A(\stack[1][47] ), .B(n17318), .Z(n15528) );
  AND U15969 ( .A(n15529), .B(n15528), .Z(n15534) );
  XNOR U15970 ( .A(n15531), .B(n15530), .Z(n15532) );
  NANDN U15971 ( .A(n17294), .B(n15532), .Z(n15533) );
  NAND U15972 ( .A(n15534), .B(n15533), .Z(n15535) );
  NOR U15973 ( .A(n15536), .B(n15535), .Z(n15537) );
  NAND U15974 ( .A(\stack[6][46] ), .B(n17311), .Z(n15539) );
  NANDN U15975 ( .A(n17311), .B(\stack[7][46] ), .Z(n15538) );
  NAND U15976 ( .A(n15539), .B(n15538), .Z(n2261) );
  NAND U15977 ( .A(\stack[5][46] ), .B(n17311), .Z(n15541) );
  NAND U15978 ( .A(n17305), .B(\stack[7][46] ), .Z(n15540) );
  AND U15979 ( .A(n15541), .B(n15540), .Z(n15543) );
  NAND U15980 ( .A(n17308), .B(\stack[6][46] ), .Z(n15542) );
  NAND U15981 ( .A(n15543), .B(n15542), .Z(n2262) );
  NAND U15982 ( .A(\stack[4][46] ), .B(n17311), .Z(n15545) );
  NAND U15983 ( .A(n17305), .B(\stack[6][46] ), .Z(n15544) );
  AND U15984 ( .A(n15545), .B(n15544), .Z(n15547) );
  NAND U15985 ( .A(n17308), .B(\stack[5][46] ), .Z(n15546) );
  NAND U15986 ( .A(n15547), .B(n15546), .Z(n2263) );
  NAND U15987 ( .A(\stack[3][46] ), .B(n17311), .Z(n15549) );
  NAND U15988 ( .A(n17305), .B(\stack[5][46] ), .Z(n15548) );
  AND U15989 ( .A(n15549), .B(n15548), .Z(n15551) );
  NAND U15990 ( .A(n17308), .B(\stack[4][46] ), .Z(n15550) );
  NAND U15991 ( .A(n15551), .B(n15550), .Z(n2264) );
  NAND U15992 ( .A(\stack[2][46] ), .B(n17311), .Z(n15553) );
  NAND U15993 ( .A(n17305), .B(\stack[4][46] ), .Z(n15552) );
  AND U15994 ( .A(n15553), .B(n15552), .Z(n15555) );
  NAND U15995 ( .A(n17308), .B(\stack[3][46] ), .Z(n15554) );
  NAND U15996 ( .A(n15555), .B(n15554), .Z(n2265) );
  NAND U15997 ( .A(n17311), .B(\stack[1][46] ), .Z(n15557) );
  NAND U15998 ( .A(n17305), .B(\stack[3][46] ), .Z(n15556) );
  AND U15999 ( .A(n15557), .B(n15556), .Z(n15559) );
  NAND U16000 ( .A(n17308), .B(\stack[2][46] ), .Z(n15558) );
  NAND U16001 ( .A(n15559), .B(n15558), .Z(n2266) );
  NAND U16002 ( .A(n17311), .B(o[46]), .Z(n15561) );
  NAND U16003 ( .A(n17305), .B(\stack[2][46] ), .Z(n15560) );
  AND U16004 ( .A(n15561), .B(n15560), .Z(n15563) );
  NAND U16005 ( .A(\stack[1][46] ), .B(n17308), .Z(n15562) );
  NAND U16006 ( .A(n15563), .B(n15562), .Z(n2267) );
  NAND U16007 ( .A(\stack[1][46] ), .B(n17313), .Z(n15564) );
  NAND U16008 ( .A(n17317), .B(n15564), .Z(n15565) );
  AND U16009 ( .A(o[46]), .B(n15565), .Z(n15574) );
  NAND U16010 ( .A(x[46]), .B(n17311), .Z(n15567) );
  NAND U16011 ( .A(\stack[1][46] ), .B(n17318), .Z(n15566) );
  AND U16012 ( .A(n15567), .B(n15566), .Z(n15572) );
  XNOR U16013 ( .A(n15569), .B(n15568), .Z(n15570) );
  NANDN U16014 ( .A(n17294), .B(n15570), .Z(n15571) );
  NAND U16015 ( .A(n15572), .B(n15571), .Z(n15573) );
  NOR U16016 ( .A(n15574), .B(n15573), .Z(n15575) );
  NAND U16017 ( .A(\stack[6][45] ), .B(n17311), .Z(n15577) );
  NANDN U16018 ( .A(n17311), .B(\stack[7][45] ), .Z(n15576) );
  NAND U16019 ( .A(n15577), .B(n15576), .Z(n2269) );
  NAND U16020 ( .A(\stack[5][45] ), .B(n17311), .Z(n15579) );
  NAND U16021 ( .A(n17305), .B(\stack[7][45] ), .Z(n15578) );
  AND U16022 ( .A(n15579), .B(n15578), .Z(n15581) );
  NAND U16023 ( .A(n17308), .B(\stack[6][45] ), .Z(n15580) );
  NAND U16024 ( .A(n15581), .B(n15580), .Z(n2270) );
  NAND U16025 ( .A(\stack[4][45] ), .B(n17311), .Z(n15583) );
  NAND U16026 ( .A(n17305), .B(\stack[6][45] ), .Z(n15582) );
  AND U16027 ( .A(n15583), .B(n15582), .Z(n15585) );
  NAND U16028 ( .A(n17308), .B(\stack[5][45] ), .Z(n15584) );
  NAND U16029 ( .A(n15585), .B(n15584), .Z(n2271) );
  NAND U16030 ( .A(\stack[3][45] ), .B(n17311), .Z(n15587) );
  NAND U16031 ( .A(n17305), .B(\stack[5][45] ), .Z(n15586) );
  AND U16032 ( .A(n15587), .B(n15586), .Z(n15589) );
  NAND U16033 ( .A(n17308), .B(\stack[4][45] ), .Z(n15588) );
  NAND U16034 ( .A(n15589), .B(n15588), .Z(n2272) );
  NAND U16035 ( .A(\stack[2][45] ), .B(n17311), .Z(n15591) );
  NAND U16036 ( .A(n17305), .B(\stack[4][45] ), .Z(n15590) );
  AND U16037 ( .A(n15591), .B(n15590), .Z(n15593) );
  NAND U16038 ( .A(n17308), .B(\stack[3][45] ), .Z(n15592) );
  NAND U16039 ( .A(n15593), .B(n15592), .Z(n2273) );
  NAND U16040 ( .A(n17311), .B(\stack[1][45] ), .Z(n15595) );
  NAND U16041 ( .A(n17305), .B(\stack[3][45] ), .Z(n15594) );
  AND U16042 ( .A(n15595), .B(n15594), .Z(n15597) );
  NAND U16043 ( .A(n17308), .B(\stack[2][45] ), .Z(n15596) );
  NAND U16044 ( .A(n15597), .B(n15596), .Z(n2274) );
  NAND U16045 ( .A(n17311), .B(o[45]), .Z(n15599) );
  NAND U16046 ( .A(n17305), .B(\stack[2][45] ), .Z(n15598) );
  AND U16047 ( .A(n15599), .B(n15598), .Z(n15601) );
  NAND U16048 ( .A(\stack[1][45] ), .B(n17308), .Z(n15600) );
  NAND U16049 ( .A(n15601), .B(n15600), .Z(n2275) );
  NAND U16050 ( .A(\stack[1][45] ), .B(n17313), .Z(n15602) );
  NAND U16051 ( .A(n17317), .B(n15602), .Z(n15603) );
  AND U16052 ( .A(o[45]), .B(n15603), .Z(n15612) );
  NAND U16053 ( .A(x[45]), .B(n17311), .Z(n15605) );
  NAND U16054 ( .A(\stack[1][45] ), .B(n17318), .Z(n15604) );
  AND U16055 ( .A(n15605), .B(n15604), .Z(n15610) );
  XNOR U16056 ( .A(n15607), .B(n15606), .Z(n15608) );
  NANDN U16057 ( .A(n17294), .B(n15608), .Z(n15609) );
  NAND U16058 ( .A(n15610), .B(n15609), .Z(n15611) );
  NOR U16059 ( .A(n15612), .B(n15611), .Z(n15613) );
  NAND U16060 ( .A(\stack[6][44] ), .B(n17311), .Z(n15615) );
  NANDN U16061 ( .A(n17311), .B(\stack[7][44] ), .Z(n15614) );
  NAND U16062 ( .A(n15615), .B(n15614), .Z(n2277) );
  NAND U16063 ( .A(\stack[5][44] ), .B(n17311), .Z(n15617) );
  NAND U16064 ( .A(n17305), .B(\stack[7][44] ), .Z(n15616) );
  AND U16065 ( .A(n15617), .B(n15616), .Z(n15619) );
  NAND U16066 ( .A(n17308), .B(\stack[6][44] ), .Z(n15618) );
  NAND U16067 ( .A(n15619), .B(n15618), .Z(n2278) );
  NAND U16068 ( .A(\stack[4][44] ), .B(n17311), .Z(n15621) );
  NAND U16069 ( .A(n17305), .B(\stack[6][44] ), .Z(n15620) );
  AND U16070 ( .A(n15621), .B(n15620), .Z(n15623) );
  NAND U16071 ( .A(n17308), .B(\stack[5][44] ), .Z(n15622) );
  NAND U16072 ( .A(n15623), .B(n15622), .Z(n2279) );
  NAND U16073 ( .A(\stack[3][44] ), .B(n17311), .Z(n15625) );
  NAND U16074 ( .A(n17305), .B(\stack[5][44] ), .Z(n15624) );
  AND U16075 ( .A(n15625), .B(n15624), .Z(n15627) );
  NAND U16076 ( .A(n17308), .B(\stack[4][44] ), .Z(n15626) );
  NAND U16077 ( .A(n15627), .B(n15626), .Z(n2280) );
  NAND U16078 ( .A(\stack[2][44] ), .B(n17311), .Z(n15629) );
  NAND U16079 ( .A(n17305), .B(\stack[4][44] ), .Z(n15628) );
  AND U16080 ( .A(n15629), .B(n15628), .Z(n15631) );
  NAND U16081 ( .A(n17308), .B(\stack[3][44] ), .Z(n15630) );
  NAND U16082 ( .A(n15631), .B(n15630), .Z(n2281) );
  NAND U16083 ( .A(n17311), .B(\stack[1][44] ), .Z(n15633) );
  NAND U16084 ( .A(n17305), .B(\stack[3][44] ), .Z(n15632) );
  AND U16085 ( .A(n15633), .B(n15632), .Z(n15635) );
  NAND U16086 ( .A(n17308), .B(\stack[2][44] ), .Z(n15634) );
  NAND U16087 ( .A(n15635), .B(n15634), .Z(n2282) );
  NAND U16088 ( .A(n17311), .B(o[44]), .Z(n15637) );
  NAND U16089 ( .A(n17305), .B(\stack[2][44] ), .Z(n15636) );
  AND U16090 ( .A(n15637), .B(n15636), .Z(n15639) );
  NAND U16091 ( .A(\stack[1][44] ), .B(n17308), .Z(n15638) );
  NAND U16092 ( .A(n15639), .B(n15638), .Z(n2283) );
  NAND U16093 ( .A(\stack[1][44] ), .B(n17313), .Z(n15640) );
  NAND U16094 ( .A(n17317), .B(n15640), .Z(n15641) );
  AND U16095 ( .A(o[44]), .B(n15641), .Z(n15650) );
  NAND U16096 ( .A(x[44]), .B(n17311), .Z(n15643) );
  NAND U16097 ( .A(\stack[1][44] ), .B(n17318), .Z(n15642) );
  AND U16098 ( .A(n15643), .B(n15642), .Z(n15648) );
  XNOR U16099 ( .A(n15645), .B(n15644), .Z(n15646) );
  NANDN U16100 ( .A(n17294), .B(n15646), .Z(n15647) );
  NAND U16101 ( .A(n15648), .B(n15647), .Z(n15649) );
  NOR U16102 ( .A(n15650), .B(n15649), .Z(n15651) );
  NAND U16103 ( .A(\stack[6][43] ), .B(n17311), .Z(n15653) );
  NANDN U16104 ( .A(n17311), .B(\stack[7][43] ), .Z(n15652) );
  NAND U16105 ( .A(n15653), .B(n15652), .Z(n2285) );
  NAND U16106 ( .A(\stack[5][43] ), .B(n17311), .Z(n15655) );
  NAND U16107 ( .A(n17305), .B(\stack[7][43] ), .Z(n15654) );
  AND U16108 ( .A(n15655), .B(n15654), .Z(n15657) );
  NAND U16109 ( .A(n17308), .B(\stack[6][43] ), .Z(n15656) );
  NAND U16110 ( .A(n15657), .B(n15656), .Z(n2286) );
  NAND U16111 ( .A(\stack[4][43] ), .B(n17311), .Z(n15659) );
  NAND U16112 ( .A(n17305), .B(\stack[6][43] ), .Z(n15658) );
  AND U16113 ( .A(n15659), .B(n15658), .Z(n15661) );
  NAND U16114 ( .A(n17308), .B(\stack[5][43] ), .Z(n15660) );
  NAND U16115 ( .A(n15661), .B(n15660), .Z(n2287) );
  NAND U16116 ( .A(\stack[3][43] ), .B(n17311), .Z(n15663) );
  NAND U16117 ( .A(n17305), .B(\stack[5][43] ), .Z(n15662) );
  AND U16118 ( .A(n15663), .B(n15662), .Z(n15665) );
  NAND U16119 ( .A(n17308), .B(\stack[4][43] ), .Z(n15664) );
  NAND U16120 ( .A(n15665), .B(n15664), .Z(n2288) );
  NAND U16121 ( .A(\stack[2][43] ), .B(n17311), .Z(n15667) );
  NAND U16122 ( .A(n17305), .B(\stack[4][43] ), .Z(n15666) );
  AND U16123 ( .A(n15667), .B(n15666), .Z(n15669) );
  NAND U16124 ( .A(n17308), .B(\stack[3][43] ), .Z(n15668) );
  NAND U16125 ( .A(n15669), .B(n15668), .Z(n2289) );
  NAND U16126 ( .A(n17311), .B(\stack[1][43] ), .Z(n15671) );
  NAND U16127 ( .A(n17305), .B(\stack[3][43] ), .Z(n15670) );
  AND U16128 ( .A(n15671), .B(n15670), .Z(n15673) );
  NAND U16129 ( .A(n17308), .B(\stack[2][43] ), .Z(n15672) );
  NAND U16130 ( .A(n15673), .B(n15672), .Z(n2290) );
  NAND U16131 ( .A(n17311), .B(o[43]), .Z(n15675) );
  NAND U16132 ( .A(n17305), .B(\stack[2][43] ), .Z(n15674) );
  AND U16133 ( .A(n15675), .B(n15674), .Z(n15677) );
  NAND U16134 ( .A(\stack[1][43] ), .B(n17308), .Z(n15676) );
  NAND U16135 ( .A(n15677), .B(n15676), .Z(n2291) );
  NAND U16136 ( .A(\stack[1][43] ), .B(n17313), .Z(n15678) );
  NAND U16137 ( .A(n17317), .B(n15678), .Z(n15679) );
  AND U16138 ( .A(o[43]), .B(n15679), .Z(n15688) );
  NAND U16139 ( .A(x[43]), .B(n17311), .Z(n15681) );
  NAND U16140 ( .A(\stack[1][43] ), .B(n17318), .Z(n15680) );
  AND U16141 ( .A(n15681), .B(n15680), .Z(n15686) );
  XNOR U16142 ( .A(n15683), .B(n15682), .Z(n15684) );
  NANDN U16143 ( .A(n17294), .B(n15684), .Z(n15685) );
  NAND U16144 ( .A(n15686), .B(n15685), .Z(n15687) );
  NOR U16145 ( .A(n15688), .B(n15687), .Z(n15689) );
  NAND U16146 ( .A(\stack[6][42] ), .B(n17311), .Z(n15691) );
  NANDN U16147 ( .A(n17311), .B(\stack[7][42] ), .Z(n15690) );
  NAND U16148 ( .A(n15691), .B(n15690), .Z(n2293) );
  NAND U16149 ( .A(\stack[5][42] ), .B(n17311), .Z(n15693) );
  NAND U16150 ( .A(n17305), .B(\stack[7][42] ), .Z(n15692) );
  AND U16151 ( .A(n15693), .B(n15692), .Z(n15695) );
  NAND U16152 ( .A(n17308), .B(\stack[6][42] ), .Z(n15694) );
  NAND U16153 ( .A(n15695), .B(n15694), .Z(n2294) );
  NAND U16154 ( .A(\stack[4][42] ), .B(n17311), .Z(n15697) );
  NAND U16155 ( .A(n17305), .B(\stack[6][42] ), .Z(n15696) );
  AND U16156 ( .A(n15697), .B(n15696), .Z(n15699) );
  NAND U16157 ( .A(n17308), .B(\stack[5][42] ), .Z(n15698) );
  NAND U16158 ( .A(n15699), .B(n15698), .Z(n2295) );
  NAND U16159 ( .A(\stack[3][42] ), .B(n17311), .Z(n15701) );
  NAND U16160 ( .A(n17305), .B(\stack[5][42] ), .Z(n15700) );
  AND U16161 ( .A(n15701), .B(n15700), .Z(n15703) );
  NAND U16162 ( .A(n17308), .B(\stack[4][42] ), .Z(n15702) );
  NAND U16163 ( .A(n15703), .B(n15702), .Z(n2296) );
  NAND U16164 ( .A(\stack[2][42] ), .B(n17311), .Z(n15705) );
  NAND U16165 ( .A(n17305), .B(\stack[4][42] ), .Z(n15704) );
  AND U16166 ( .A(n15705), .B(n15704), .Z(n15707) );
  NAND U16167 ( .A(n17308), .B(\stack[3][42] ), .Z(n15706) );
  NAND U16168 ( .A(n15707), .B(n15706), .Z(n2297) );
  NAND U16169 ( .A(n17311), .B(\stack[1][42] ), .Z(n15709) );
  NAND U16170 ( .A(n17305), .B(\stack[3][42] ), .Z(n15708) );
  AND U16171 ( .A(n15709), .B(n15708), .Z(n15711) );
  NAND U16172 ( .A(n17308), .B(\stack[2][42] ), .Z(n15710) );
  NAND U16173 ( .A(n15711), .B(n15710), .Z(n2298) );
  NAND U16174 ( .A(n17311), .B(o[42]), .Z(n15713) );
  NAND U16175 ( .A(n17305), .B(\stack[2][42] ), .Z(n15712) );
  AND U16176 ( .A(n15713), .B(n15712), .Z(n15715) );
  NAND U16177 ( .A(\stack[1][42] ), .B(n17308), .Z(n15714) );
  NAND U16178 ( .A(n15715), .B(n15714), .Z(n2299) );
  NAND U16179 ( .A(\stack[1][42] ), .B(n17313), .Z(n15716) );
  NAND U16180 ( .A(n17317), .B(n15716), .Z(n15717) );
  AND U16181 ( .A(o[42]), .B(n15717), .Z(n15726) );
  NAND U16182 ( .A(x[42]), .B(n17311), .Z(n15719) );
  NAND U16183 ( .A(\stack[1][42] ), .B(n17318), .Z(n15718) );
  AND U16184 ( .A(n15719), .B(n15718), .Z(n15724) );
  XNOR U16185 ( .A(n15721), .B(n15720), .Z(n15722) );
  NANDN U16186 ( .A(n17294), .B(n15722), .Z(n15723) );
  NAND U16187 ( .A(n15724), .B(n15723), .Z(n15725) );
  NOR U16188 ( .A(n15726), .B(n15725), .Z(n15727) );
  NAND U16189 ( .A(\stack[6][41] ), .B(n17311), .Z(n15729) );
  NANDN U16190 ( .A(n17311), .B(\stack[7][41] ), .Z(n15728) );
  NAND U16191 ( .A(n15729), .B(n15728), .Z(n2301) );
  NAND U16192 ( .A(\stack[5][41] ), .B(n17311), .Z(n15731) );
  NAND U16193 ( .A(n17305), .B(\stack[7][41] ), .Z(n15730) );
  AND U16194 ( .A(n15731), .B(n15730), .Z(n15733) );
  NAND U16195 ( .A(n17308), .B(\stack[6][41] ), .Z(n15732) );
  NAND U16196 ( .A(n15733), .B(n15732), .Z(n2302) );
  NAND U16197 ( .A(\stack[4][41] ), .B(n17311), .Z(n15735) );
  NAND U16198 ( .A(n17305), .B(\stack[6][41] ), .Z(n15734) );
  AND U16199 ( .A(n15735), .B(n15734), .Z(n15737) );
  NAND U16200 ( .A(n17308), .B(\stack[5][41] ), .Z(n15736) );
  NAND U16201 ( .A(n15737), .B(n15736), .Z(n2303) );
  NAND U16202 ( .A(\stack[3][41] ), .B(n17311), .Z(n15739) );
  NAND U16203 ( .A(n17305), .B(\stack[5][41] ), .Z(n15738) );
  AND U16204 ( .A(n15739), .B(n15738), .Z(n15741) );
  NAND U16205 ( .A(n17308), .B(\stack[4][41] ), .Z(n15740) );
  NAND U16206 ( .A(n15741), .B(n15740), .Z(n2304) );
  NAND U16207 ( .A(\stack[2][41] ), .B(n17311), .Z(n15743) );
  NAND U16208 ( .A(n17305), .B(\stack[4][41] ), .Z(n15742) );
  AND U16209 ( .A(n15743), .B(n15742), .Z(n15745) );
  NAND U16210 ( .A(n17308), .B(\stack[3][41] ), .Z(n15744) );
  NAND U16211 ( .A(n15745), .B(n15744), .Z(n2305) );
  NAND U16212 ( .A(n17311), .B(\stack[1][41] ), .Z(n15747) );
  NAND U16213 ( .A(n17305), .B(\stack[3][41] ), .Z(n15746) );
  AND U16214 ( .A(n15747), .B(n15746), .Z(n15749) );
  NAND U16215 ( .A(n17308), .B(\stack[2][41] ), .Z(n15748) );
  NAND U16216 ( .A(n15749), .B(n15748), .Z(n2306) );
  NAND U16217 ( .A(n17311), .B(o[41]), .Z(n15751) );
  NAND U16218 ( .A(n17305), .B(\stack[2][41] ), .Z(n15750) );
  AND U16219 ( .A(n15751), .B(n15750), .Z(n15753) );
  NAND U16220 ( .A(\stack[1][41] ), .B(n17308), .Z(n15752) );
  NAND U16221 ( .A(n15753), .B(n15752), .Z(n2307) );
  NAND U16222 ( .A(\stack[1][41] ), .B(n17313), .Z(n15754) );
  NAND U16223 ( .A(n17317), .B(n15754), .Z(n15755) );
  AND U16224 ( .A(o[41]), .B(n15755), .Z(n15764) );
  NAND U16225 ( .A(x[41]), .B(n17311), .Z(n15757) );
  NAND U16226 ( .A(\stack[1][41] ), .B(n17318), .Z(n15756) );
  AND U16227 ( .A(n15757), .B(n15756), .Z(n15762) );
  XNOR U16228 ( .A(n15759), .B(n15758), .Z(n15760) );
  NANDN U16229 ( .A(n17294), .B(n15760), .Z(n15761) );
  NAND U16230 ( .A(n15762), .B(n15761), .Z(n15763) );
  NOR U16231 ( .A(n15764), .B(n15763), .Z(n15765) );
  NAND U16232 ( .A(\stack[6][40] ), .B(n17311), .Z(n15767) );
  NANDN U16233 ( .A(n17311), .B(\stack[7][40] ), .Z(n15766) );
  NAND U16234 ( .A(n15767), .B(n15766), .Z(n2309) );
  NAND U16235 ( .A(\stack[5][40] ), .B(n17311), .Z(n15769) );
  NAND U16236 ( .A(n17305), .B(\stack[7][40] ), .Z(n15768) );
  AND U16237 ( .A(n15769), .B(n15768), .Z(n15771) );
  NAND U16238 ( .A(n17308), .B(\stack[6][40] ), .Z(n15770) );
  NAND U16239 ( .A(n15771), .B(n15770), .Z(n2310) );
  NAND U16240 ( .A(\stack[4][40] ), .B(n17311), .Z(n15773) );
  NAND U16241 ( .A(n17305), .B(\stack[6][40] ), .Z(n15772) );
  AND U16242 ( .A(n15773), .B(n15772), .Z(n15775) );
  NAND U16243 ( .A(n17308), .B(\stack[5][40] ), .Z(n15774) );
  NAND U16244 ( .A(n15775), .B(n15774), .Z(n2311) );
  NAND U16245 ( .A(\stack[3][40] ), .B(n17311), .Z(n15777) );
  NAND U16246 ( .A(n17305), .B(\stack[5][40] ), .Z(n15776) );
  AND U16247 ( .A(n15777), .B(n15776), .Z(n15779) );
  NAND U16248 ( .A(n17308), .B(\stack[4][40] ), .Z(n15778) );
  NAND U16249 ( .A(n15779), .B(n15778), .Z(n2312) );
  NAND U16250 ( .A(\stack[2][40] ), .B(n17311), .Z(n15781) );
  NAND U16251 ( .A(n17305), .B(\stack[4][40] ), .Z(n15780) );
  AND U16252 ( .A(n15781), .B(n15780), .Z(n15783) );
  NAND U16253 ( .A(n17308), .B(\stack[3][40] ), .Z(n15782) );
  NAND U16254 ( .A(n15783), .B(n15782), .Z(n2313) );
  NAND U16255 ( .A(n17311), .B(\stack[1][40] ), .Z(n15785) );
  NAND U16256 ( .A(n17305), .B(\stack[3][40] ), .Z(n15784) );
  AND U16257 ( .A(n15785), .B(n15784), .Z(n15787) );
  NAND U16258 ( .A(n17308), .B(\stack[2][40] ), .Z(n15786) );
  NAND U16259 ( .A(n15787), .B(n15786), .Z(n2314) );
  NAND U16260 ( .A(n17311), .B(o[40]), .Z(n15789) );
  NAND U16261 ( .A(n17305), .B(\stack[2][40] ), .Z(n15788) );
  AND U16262 ( .A(n15789), .B(n15788), .Z(n15791) );
  NAND U16263 ( .A(\stack[1][40] ), .B(n17308), .Z(n15790) );
  NAND U16264 ( .A(n15791), .B(n15790), .Z(n2315) );
  NAND U16265 ( .A(\stack[1][40] ), .B(n17313), .Z(n15792) );
  NAND U16266 ( .A(n17317), .B(n15792), .Z(n15793) );
  AND U16267 ( .A(o[40]), .B(n15793), .Z(n15802) );
  NAND U16268 ( .A(x[40]), .B(n17311), .Z(n15795) );
  NAND U16269 ( .A(\stack[1][40] ), .B(n17318), .Z(n15794) );
  AND U16270 ( .A(n15795), .B(n15794), .Z(n15800) );
  XNOR U16271 ( .A(n15797), .B(n15796), .Z(n15798) );
  NANDN U16272 ( .A(n17294), .B(n15798), .Z(n15799) );
  NAND U16273 ( .A(n15800), .B(n15799), .Z(n15801) );
  NOR U16274 ( .A(n15802), .B(n15801), .Z(n15803) );
  NAND U16275 ( .A(\stack[6][39] ), .B(n17311), .Z(n15805) );
  NANDN U16276 ( .A(n17311), .B(\stack[7][39] ), .Z(n15804) );
  NAND U16277 ( .A(n15805), .B(n15804), .Z(n2317) );
  NAND U16278 ( .A(\stack[5][39] ), .B(n17311), .Z(n15807) );
  NAND U16279 ( .A(n17305), .B(\stack[7][39] ), .Z(n15806) );
  AND U16280 ( .A(n15807), .B(n15806), .Z(n15809) );
  NAND U16281 ( .A(n17308), .B(\stack[6][39] ), .Z(n15808) );
  NAND U16282 ( .A(n15809), .B(n15808), .Z(n2318) );
  NAND U16283 ( .A(\stack[4][39] ), .B(n17311), .Z(n15811) );
  NAND U16284 ( .A(n17305), .B(\stack[6][39] ), .Z(n15810) );
  AND U16285 ( .A(n15811), .B(n15810), .Z(n15813) );
  NAND U16286 ( .A(n17308), .B(\stack[5][39] ), .Z(n15812) );
  NAND U16287 ( .A(n15813), .B(n15812), .Z(n2319) );
  NAND U16288 ( .A(\stack[3][39] ), .B(n17311), .Z(n15815) );
  NAND U16289 ( .A(n17305), .B(\stack[5][39] ), .Z(n15814) );
  AND U16290 ( .A(n15815), .B(n15814), .Z(n15817) );
  NAND U16291 ( .A(n17308), .B(\stack[4][39] ), .Z(n15816) );
  NAND U16292 ( .A(n15817), .B(n15816), .Z(n2320) );
  NAND U16293 ( .A(\stack[2][39] ), .B(n17311), .Z(n15819) );
  NAND U16294 ( .A(n17305), .B(\stack[4][39] ), .Z(n15818) );
  AND U16295 ( .A(n15819), .B(n15818), .Z(n15821) );
  NAND U16296 ( .A(n17308), .B(\stack[3][39] ), .Z(n15820) );
  NAND U16297 ( .A(n15821), .B(n15820), .Z(n2321) );
  NAND U16298 ( .A(n17311), .B(\stack[1][39] ), .Z(n15823) );
  NAND U16299 ( .A(n17305), .B(\stack[3][39] ), .Z(n15822) );
  AND U16300 ( .A(n15823), .B(n15822), .Z(n15825) );
  NAND U16301 ( .A(n17308), .B(\stack[2][39] ), .Z(n15824) );
  NAND U16302 ( .A(n15825), .B(n15824), .Z(n2322) );
  NAND U16303 ( .A(n17311), .B(o[39]), .Z(n15827) );
  NAND U16304 ( .A(n17305), .B(\stack[2][39] ), .Z(n15826) );
  AND U16305 ( .A(n15827), .B(n15826), .Z(n15829) );
  NAND U16306 ( .A(\stack[1][39] ), .B(n17308), .Z(n15828) );
  NAND U16307 ( .A(n15829), .B(n15828), .Z(n2323) );
  NAND U16308 ( .A(\stack[1][39] ), .B(n17313), .Z(n15830) );
  NAND U16309 ( .A(n17317), .B(n15830), .Z(n15831) );
  AND U16310 ( .A(o[39]), .B(n15831), .Z(n15840) );
  NAND U16311 ( .A(x[39]), .B(n17311), .Z(n15833) );
  NAND U16312 ( .A(\stack[1][39] ), .B(n17318), .Z(n15832) );
  AND U16313 ( .A(n15833), .B(n15832), .Z(n15838) );
  XNOR U16314 ( .A(n15835), .B(n15834), .Z(n15836) );
  NANDN U16315 ( .A(n17294), .B(n15836), .Z(n15837) );
  NAND U16316 ( .A(n15838), .B(n15837), .Z(n15839) );
  NOR U16317 ( .A(n15840), .B(n15839), .Z(n15841) );
  NAND U16318 ( .A(\stack[6][38] ), .B(n17311), .Z(n15843) );
  NANDN U16319 ( .A(n17311), .B(\stack[7][38] ), .Z(n15842) );
  NAND U16320 ( .A(n15843), .B(n15842), .Z(n2325) );
  NAND U16321 ( .A(\stack[5][38] ), .B(n17311), .Z(n15845) );
  NAND U16322 ( .A(n17305), .B(\stack[7][38] ), .Z(n15844) );
  AND U16323 ( .A(n15845), .B(n15844), .Z(n15847) );
  NAND U16324 ( .A(n17308), .B(\stack[6][38] ), .Z(n15846) );
  NAND U16325 ( .A(n15847), .B(n15846), .Z(n2326) );
  NAND U16326 ( .A(\stack[4][38] ), .B(n17311), .Z(n15849) );
  NAND U16327 ( .A(n17305), .B(\stack[6][38] ), .Z(n15848) );
  AND U16328 ( .A(n15849), .B(n15848), .Z(n15851) );
  NAND U16329 ( .A(n17308), .B(\stack[5][38] ), .Z(n15850) );
  NAND U16330 ( .A(n15851), .B(n15850), .Z(n2327) );
  NAND U16331 ( .A(\stack[3][38] ), .B(n17311), .Z(n15853) );
  NAND U16332 ( .A(n17305), .B(\stack[5][38] ), .Z(n15852) );
  AND U16333 ( .A(n15853), .B(n15852), .Z(n15855) );
  NAND U16334 ( .A(n17308), .B(\stack[4][38] ), .Z(n15854) );
  NAND U16335 ( .A(n15855), .B(n15854), .Z(n2328) );
  NAND U16336 ( .A(\stack[2][38] ), .B(n17311), .Z(n15857) );
  NAND U16337 ( .A(n17305), .B(\stack[4][38] ), .Z(n15856) );
  AND U16338 ( .A(n15857), .B(n15856), .Z(n15859) );
  NAND U16339 ( .A(n17308), .B(\stack[3][38] ), .Z(n15858) );
  NAND U16340 ( .A(n15859), .B(n15858), .Z(n2329) );
  NAND U16341 ( .A(n17311), .B(\stack[1][38] ), .Z(n15861) );
  NAND U16342 ( .A(n17305), .B(\stack[3][38] ), .Z(n15860) );
  AND U16343 ( .A(n15861), .B(n15860), .Z(n15863) );
  NAND U16344 ( .A(n17308), .B(\stack[2][38] ), .Z(n15862) );
  NAND U16345 ( .A(n15863), .B(n15862), .Z(n2330) );
  NAND U16346 ( .A(n17311), .B(o[38]), .Z(n15865) );
  NAND U16347 ( .A(n17305), .B(\stack[2][38] ), .Z(n15864) );
  AND U16348 ( .A(n15865), .B(n15864), .Z(n15867) );
  NAND U16349 ( .A(\stack[1][38] ), .B(n17308), .Z(n15866) );
  NAND U16350 ( .A(n15867), .B(n15866), .Z(n2331) );
  NAND U16351 ( .A(\stack[1][38] ), .B(n17313), .Z(n15868) );
  NAND U16352 ( .A(n17317), .B(n15868), .Z(n15869) );
  AND U16353 ( .A(o[38]), .B(n15869), .Z(n15878) );
  NAND U16354 ( .A(x[38]), .B(n17311), .Z(n15871) );
  NAND U16355 ( .A(\stack[1][38] ), .B(n17318), .Z(n15870) );
  AND U16356 ( .A(n15871), .B(n15870), .Z(n15876) );
  XNOR U16357 ( .A(n15873), .B(n15872), .Z(n15874) );
  NANDN U16358 ( .A(n17294), .B(n15874), .Z(n15875) );
  NAND U16359 ( .A(n15876), .B(n15875), .Z(n15877) );
  NOR U16360 ( .A(n15878), .B(n15877), .Z(n15879) );
  NAND U16361 ( .A(\stack[6][37] ), .B(n17311), .Z(n15881) );
  NANDN U16362 ( .A(n17311), .B(\stack[7][37] ), .Z(n15880) );
  NAND U16363 ( .A(n15881), .B(n15880), .Z(n2333) );
  NAND U16364 ( .A(\stack[5][37] ), .B(n17311), .Z(n15883) );
  NAND U16365 ( .A(n17305), .B(\stack[7][37] ), .Z(n15882) );
  AND U16366 ( .A(n15883), .B(n15882), .Z(n15885) );
  NAND U16367 ( .A(n17308), .B(\stack[6][37] ), .Z(n15884) );
  NAND U16368 ( .A(n15885), .B(n15884), .Z(n2334) );
  NAND U16369 ( .A(\stack[4][37] ), .B(n17311), .Z(n15887) );
  NAND U16370 ( .A(n17305), .B(\stack[6][37] ), .Z(n15886) );
  AND U16371 ( .A(n15887), .B(n15886), .Z(n15889) );
  NAND U16372 ( .A(n17308), .B(\stack[5][37] ), .Z(n15888) );
  NAND U16373 ( .A(n15889), .B(n15888), .Z(n2335) );
  NAND U16374 ( .A(\stack[3][37] ), .B(n17311), .Z(n15891) );
  NAND U16375 ( .A(n17305), .B(\stack[5][37] ), .Z(n15890) );
  AND U16376 ( .A(n15891), .B(n15890), .Z(n15893) );
  NAND U16377 ( .A(n17308), .B(\stack[4][37] ), .Z(n15892) );
  NAND U16378 ( .A(n15893), .B(n15892), .Z(n2336) );
  NAND U16379 ( .A(\stack[2][37] ), .B(n17311), .Z(n15895) );
  NAND U16380 ( .A(n17305), .B(\stack[4][37] ), .Z(n15894) );
  AND U16381 ( .A(n15895), .B(n15894), .Z(n15897) );
  NAND U16382 ( .A(n17308), .B(\stack[3][37] ), .Z(n15896) );
  NAND U16383 ( .A(n15897), .B(n15896), .Z(n2337) );
  NAND U16384 ( .A(n17311), .B(\stack[1][37] ), .Z(n15899) );
  NAND U16385 ( .A(n17305), .B(\stack[3][37] ), .Z(n15898) );
  AND U16386 ( .A(n15899), .B(n15898), .Z(n15901) );
  NAND U16387 ( .A(n17308), .B(\stack[2][37] ), .Z(n15900) );
  NAND U16388 ( .A(n15901), .B(n15900), .Z(n2338) );
  NAND U16389 ( .A(n17311), .B(o[37]), .Z(n15903) );
  NAND U16390 ( .A(n17305), .B(\stack[2][37] ), .Z(n15902) );
  AND U16391 ( .A(n15903), .B(n15902), .Z(n15905) );
  NAND U16392 ( .A(\stack[1][37] ), .B(n17308), .Z(n15904) );
  NAND U16393 ( .A(n15905), .B(n15904), .Z(n2339) );
  NAND U16394 ( .A(\stack[1][37] ), .B(n17313), .Z(n15906) );
  NAND U16395 ( .A(n17317), .B(n15906), .Z(n15907) );
  AND U16396 ( .A(o[37]), .B(n15907), .Z(n15916) );
  NAND U16397 ( .A(x[37]), .B(n17311), .Z(n15909) );
  NAND U16398 ( .A(\stack[1][37] ), .B(n17318), .Z(n15908) );
  AND U16399 ( .A(n15909), .B(n15908), .Z(n15914) );
  XNOR U16400 ( .A(n15911), .B(n15910), .Z(n15912) );
  NANDN U16401 ( .A(n17294), .B(n15912), .Z(n15913) );
  NAND U16402 ( .A(n15914), .B(n15913), .Z(n15915) );
  NOR U16403 ( .A(n15916), .B(n15915), .Z(n15917) );
  NAND U16404 ( .A(\stack[6][36] ), .B(n17311), .Z(n15919) );
  NANDN U16405 ( .A(n17311), .B(\stack[7][36] ), .Z(n15918) );
  NAND U16406 ( .A(n15919), .B(n15918), .Z(n2341) );
  NAND U16407 ( .A(\stack[5][36] ), .B(n17311), .Z(n15921) );
  NAND U16408 ( .A(n17305), .B(\stack[7][36] ), .Z(n15920) );
  AND U16409 ( .A(n15921), .B(n15920), .Z(n15923) );
  NAND U16410 ( .A(n17308), .B(\stack[6][36] ), .Z(n15922) );
  NAND U16411 ( .A(n15923), .B(n15922), .Z(n2342) );
  NAND U16412 ( .A(\stack[4][36] ), .B(n17311), .Z(n15925) );
  NAND U16413 ( .A(n17305), .B(\stack[6][36] ), .Z(n15924) );
  AND U16414 ( .A(n15925), .B(n15924), .Z(n15927) );
  NAND U16415 ( .A(n17308), .B(\stack[5][36] ), .Z(n15926) );
  NAND U16416 ( .A(n15927), .B(n15926), .Z(n2343) );
  NAND U16417 ( .A(\stack[3][36] ), .B(n17311), .Z(n15929) );
  NAND U16418 ( .A(n17305), .B(\stack[5][36] ), .Z(n15928) );
  AND U16419 ( .A(n15929), .B(n15928), .Z(n15931) );
  NAND U16420 ( .A(n17308), .B(\stack[4][36] ), .Z(n15930) );
  NAND U16421 ( .A(n15931), .B(n15930), .Z(n2344) );
  NAND U16422 ( .A(\stack[2][36] ), .B(n17311), .Z(n15933) );
  NAND U16423 ( .A(n17305), .B(\stack[4][36] ), .Z(n15932) );
  AND U16424 ( .A(n15933), .B(n15932), .Z(n15935) );
  NAND U16425 ( .A(n17308), .B(\stack[3][36] ), .Z(n15934) );
  NAND U16426 ( .A(n15935), .B(n15934), .Z(n2345) );
  NAND U16427 ( .A(n17311), .B(\stack[1][36] ), .Z(n15937) );
  NAND U16428 ( .A(n17305), .B(\stack[3][36] ), .Z(n15936) );
  AND U16429 ( .A(n15937), .B(n15936), .Z(n15939) );
  NAND U16430 ( .A(n17308), .B(\stack[2][36] ), .Z(n15938) );
  NAND U16431 ( .A(n15939), .B(n15938), .Z(n2346) );
  NAND U16432 ( .A(n17311), .B(o[36]), .Z(n15941) );
  NAND U16433 ( .A(n17305), .B(\stack[2][36] ), .Z(n15940) );
  AND U16434 ( .A(n15941), .B(n15940), .Z(n15943) );
  NAND U16435 ( .A(\stack[1][36] ), .B(n17308), .Z(n15942) );
  NAND U16436 ( .A(n15943), .B(n15942), .Z(n2347) );
  NAND U16437 ( .A(o[36]), .B(n17313), .Z(n15944) );
  NANDN U16438 ( .A(n17318), .B(n15944), .Z(n15945) );
  AND U16439 ( .A(\stack[1][36] ), .B(n15945), .Z(n15953) );
  NAND U16440 ( .A(x[36]), .B(n17311), .Z(n15946) );
  XNOR U16441 ( .A(n15948), .B(n15947), .Z(n15949) );
  NANDN U16442 ( .A(n17294), .B(n15949), .Z(n15950) );
  NAND U16443 ( .A(n15951), .B(n15950), .Z(n15952) );
  NOR U16444 ( .A(n15953), .B(n15952), .Z(n15955) );
  NANDN U16445 ( .A(n17317), .B(o[36]), .Z(n15954) );
  NAND U16446 ( .A(n15955), .B(n15954), .Z(n2348) );
  NAND U16447 ( .A(\stack[6][35] ), .B(n17311), .Z(n15957) );
  NANDN U16448 ( .A(n17311), .B(\stack[7][35] ), .Z(n15956) );
  NAND U16449 ( .A(n15957), .B(n15956), .Z(n2349) );
  NAND U16450 ( .A(\stack[5][35] ), .B(n17311), .Z(n15959) );
  NAND U16451 ( .A(n17305), .B(\stack[7][35] ), .Z(n15958) );
  AND U16452 ( .A(n15959), .B(n15958), .Z(n15961) );
  NAND U16453 ( .A(n17308), .B(\stack[6][35] ), .Z(n15960) );
  NAND U16454 ( .A(n15961), .B(n15960), .Z(n2350) );
  NAND U16455 ( .A(\stack[4][35] ), .B(n17311), .Z(n15963) );
  NAND U16456 ( .A(n17305), .B(\stack[6][35] ), .Z(n15962) );
  AND U16457 ( .A(n15963), .B(n15962), .Z(n15965) );
  NAND U16458 ( .A(n17308), .B(\stack[5][35] ), .Z(n15964) );
  NAND U16459 ( .A(n15965), .B(n15964), .Z(n2351) );
  NAND U16460 ( .A(\stack[3][35] ), .B(n17311), .Z(n15967) );
  NAND U16461 ( .A(n17305), .B(\stack[5][35] ), .Z(n15966) );
  AND U16462 ( .A(n15967), .B(n15966), .Z(n15969) );
  NAND U16463 ( .A(n17308), .B(\stack[4][35] ), .Z(n15968) );
  NAND U16464 ( .A(n15969), .B(n15968), .Z(n2352) );
  NAND U16465 ( .A(\stack[2][35] ), .B(n17311), .Z(n15971) );
  NAND U16466 ( .A(n17305), .B(\stack[4][35] ), .Z(n15970) );
  AND U16467 ( .A(n15971), .B(n15970), .Z(n15973) );
  NAND U16468 ( .A(n17308), .B(\stack[3][35] ), .Z(n15972) );
  NAND U16469 ( .A(n15973), .B(n15972), .Z(n2353) );
  NAND U16470 ( .A(n17311), .B(\stack[1][35] ), .Z(n15975) );
  NAND U16471 ( .A(n17305), .B(\stack[3][35] ), .Z(n15974) );
  AND U16472 ( .A(n15975), .B(n15974), .Z(n15977) );
  NAND U16473 ( .A(n17308), .B(\stack[2][35] ), .Z(n15976) );
  NAND U16474 ( .A(n15977), .B(n15976), .Z(n2354) );
  NAND U16475 ( .A(n17311), .B(o[35]), .Z(n15979) );
  NAND U16476 ( .A(n17305), .B(\stack[2][35] ), .Z(n15978) );
  AND U16477 ( .A(n15979), .B(n15978), .Z(n15981) );
  NAND U16478 ( .A(\stack[1][35] ), .B(n17308), .Z(n15980) );
  NAND U16479 ( .A(n15981), .B(n15980), .Z(n2355) );
  NAND U16480 ( .A(\stack[1][35] ), .B(n17313), .Z(n15982) );
  NAND U16481 ( .A(n17317), .B(n15982), .Z(n15983) );
  AND U16482 ( .A(o[35]), .B(n15983), .Z(n15992) );
  NAND U16483 ( .A(x[35]), .B(n17311), .Z(n15985) );
  NAND U16484 ( .A(\stack[1][35] ), .B(n17318), .Z(n15984) );
  AND U16485 ( .A(n15985), .B(n15984), .Z(n15990) );
  XNOR U16486 ( .A(n15987), .B(n15986), .Z(n15988) );
  NANDN U16487 ( .A(n17294), .B(n15988), .Z(n15989) );
  NAND U16488 ( .A(n15990), .B(n15989), .Z(n15991) );
  NOR U16489 ( .A(n15992), .B(n15991), .Z(n15993) );
  NAND U16490 ( .A(\stack[6][34] ), .B(n17311), .Z(n15995) );
  NANDN U16491 ( .A(n17311), .B(\stack[7][34] ), .Z(n15994) );
  NAND U16492 ( .A(n15995), .B(n15994), .Z(n2357) );
  NAND U16493 ( .A(\stack[5][34] ), .B(n17311), .Z(n15997) );
  NAND U16494 ( .A(n17305), .B(\stack[7][34] ), .Z(n15996) );
  AND U16495 ( .A(n15997), .B(n15996), .Z(n15999) );
  NAND U16496 ( .A(n17308), .B(\stack[6][34] ), .Z(n15998) );
  NAND U16497 ( .A(n15999), .B(n15998), .Z(n2358) );
  NAND U16498 ( .A(\stack[4][34] ), .B(n17311), .Z(n16001) );
  NAND U16499 ( .A(n17305), .B(\stack[6][34] ), .Z(n16000) );
  AND U16500 ( .A(n16001), .B(n16000), .Z(n16003) );
  NAND U16501 ( .A(n17308), .B(\stack[5][34] ), .Z(n16002) );
  NAND U16502 ( .A(n16003), .B(n16002), .Z(n2359) );
  NAND U16503 ( .A(\stack[3][34] ), .B(n17311), .Z(n16005) );
  NAND U16504 ( .A(n17305), .B(\stack[5][34] ), .Z(n16004) );
  AND U16505 ( .A(n16005), .B(n16004), .Z(n16007) );
  NAND U16506 ( .A(n17308), .B(\stack[4][34] ), .Z(n16006) );
  NAND U16507 ( .A(n16007), .B(n16006), .Z(n2360) );
  NAND U16508 ( .A(\stack[2][34] ), .B(n17311), .Z(n16009) );
  NAND U16509 ( .A(n17305), .B(\stack[4][34] ), .Z(n16008) );
  AND U16510 ( .A(n16009), .B(n16008), .Z(n16011) );
  NAND U16511 ( .A(n17308), .B(\stack[3][34] ), .Z(n16010) );
  NAND U16512 ( .A(n16011), .B(n16010), .Z(n2361) );
  NAND U16513 ( .A(n17311), .B(\stack[1][34] ), .Z(n16013) );
  NAND U16514 ( .A(n17305), .B(\stack[3][34] ), .Z(n16012) );
  AND U16515 ( .A(n16013), .B(n16012), .Z(n16015) );
  NAND U16516 ( .A(n17308), .B(\stack[2][34] ), .Z(n16014) );
  NAND U16517 ( .A(n16015), .B(n16014), .Z(n2362) );
  NAND U16518 ( .A(n17311), .B(o[34]), .Z(n16017) );
  NAND U16519 ( .A(n17305), .B(\stack[2][34] ), .Z(n16016) );
  AND U16520 ( .A(n16017), .B(n16016), .Z(n16019) );
  NAND U16521 ( .A(\stack[1][34] ), .B(n17308), .Z(n16018) );
  NAND U16522 ( .A(n16019), .B(n16018), .Z(n2363) );
  NAND U16523 ( .A(o[34]), .B(n17313), .Z(n16020) );
  NANDN U16524 ( .A(n17318), .B(n16020), .Z(n16021) );
  AND U16525 ( .A(\stack[1][34] ), .B(n16021), .Z(n16029) );
  NAND U16526 ( .A(x[34]), .B(n17311), .Z(n16022) );
  XNOR U16527 ( .A(n16024), .B(n16023), .Z(n16025) );
  NANDN U16528 ( .A(n17294), .B(n16025), .Z(n16026) );
  NAND U16529 ( .A(n16027), .B(n16026), .Z(n16028) );
  NOR U16530 ( .A(n16029), .B(n16028), .Z(n16031) );
  NANDN U16531 ( .A(n17317), .B(o[34]), .Z(n16030) );
  NAND U16532 ( .A(n16031), .B(n16030), .Z(n2364) );
  NAND U16533 ( .A(\stack[6][33] ), .B(n17311), .Z(n16033) );
  NANDN U16534 ( .A(n17311), .B(\stack[7][33] ), .Z(n16032) );
  NAND U16535 ( .A(n16033), .B(n16032), .Z(n2365) );
  NAND U16536 ( .A(\stack[5][33] ), .B(n17311), .Z(n16035) );
  NAND U16537 ( .A(n17305), .B(\stack[7][33] ), .Z(n16034) );
  AND U16538 ( .A(n16035), .B(n16034), .Z(n16037) );
  NAND U16539 ( .A(n17308), .B(\stack[6][33] ), .Z(n16036) );
  NAND U16540 ( .A(n16037), .B(n16036), .Z(n2366) );
  NAND U16541 ( .A(\stack[4][33] ), .B(n17311), .Z(n16039) );
  NAND U16542 ( .A(n17305), .B(\stack[6][33] ), .Z(n16038) );
  AND U16543 ( .A(n16039), .B(n16038), .Z(n16041) );
  NAND U16544 ( .A(n17308), .B(\stack[5][33] ), .Z(n16040) );
  NAND U16545 ( .A(n16041), .B(n16040), .Z(n2367) );
  NAND U16546 ( .A(\stack[3][33] ), .B(n17311), .Z(n16043) );
  NAND U16547 ( .A(n17305), .B(\stack[5][33] ), .Z(n16042) );
  AND U16548 ( .A(n16043), .B(n16042), .Z(n16045) );
  NAND U16549 ( .A(n17308), .B(\stack[4][33] ), .Z(n16044) );
  NAND U16550 ( .A(n16045), .B(n16044), .Z(n2368) );
  NAND U16551 ( .A(\stack[2][33] ), .B(n17311), .Z(n16047) );
  NAND U16552 ( .A(n17305), .B(\stack[4][33] ), .Z(n16046) );
  AND U16553 ( .A(n16047), .B(n16046), .Z(n16049) );
  NAND U16554 ( .A(n17308), .B(\stack[3][33] ), .Z(n16048) );
  NAND U16555 ( .A(n16049), .B(n16048), .Z(n2369) );
  NAND U16556 ( .A(n17311), .B(\stack[1][33] ), .Z(n16051) );
  NAND U16557 ( .A(n17305), .B(\stack[3][33] ), .Z(n16050) );
  AND U16558 ( .A(n16051), .B(n16050), .Z(n16053) );
  NAND U16559 ( .A(n17308), .B(\stack[2][33] ), .Z(n16052) );
  NAND U16560 ( .A(n16053), .B(n16052), .Z(n2370) );
  NAND U16561 ( .A(n17311), .B(o[33]), .Z(n16055) );
  NAND U16562 ( .A(n17305), .B(\stack[2][33] ), .Z(n16054) );
  AND U16563 ( .A(n16055), .B(n16054), .Z(n16057) );
  NAND U16564 ( .A(\stack[1][33] ), .B(n17308), .Z(n16056) );
  NAND U16565 ( .A(n16057), .B(n16056), .Z(n2371) );
  NAND U16566 ( .A(\stack[1][33] ), .B(n17313), .Z(n16058) );
  NAND U16567 ( .A(n17317), .B(n16058), .Z(n16059) );
  AND U16568 ( .A(o[33]), .B(n16059), .Z(n16068) );
  NAND U16569 ( .A(x[33]), .B(n17311), .Z(n16061) );
  NAND U16570 ( .A(\stack[1][33] ), .B(n17318), .Z(n16060) );
  AND U16571 ( .A(n16061), .B(n16060), .Z(n16066) );
  XNOR U16572 ( .A(n16063), .B(n16062), .Z(n16064) );
  NANDN U16573 ( .A(n17294), .B(n16064), .Z(n16065) );
  NAND U16574 ( .A(n16066), .B(n16065), .Z(n16067) );
  NOR U16575 ( .A(n16068), .B(n16067), .Z(n16069) );
  NAND U16576 ( .A(\stack[6][32] ), .B(n17311), .Z(n16071) );
  NANDN U16577 ( .A(n17311), .B(\stack[7][32] ), .Z(n16070) );
  NAND U16578 ( .A(n16071), .B(n16070), .Z(n2373) );
  NAND U16579 ( .A(\stack[5][32] ), .B(n17311), .Z(n16073) );
  NAND U16580 ( .A(n17305), .B(\stack[7][32] ), .Z(n16072) );
  AND U16581 ( .A(n16073), .B(n16072), .Z(n16075) );
  NAND U16582 ( .A(n17308), .B(\stack[6][32] ), .Z(n16074) );
  NAND U16583 ( .A(n16075), .B(n16074), .Z(n2374) );
  NAND U16584 ( .A(\stack[4][32] ), .B(n17311), .Z(n16077) );
  NAND U16585 ( .A(n17305), .B(\stack[6][32] ), .Z(n16076) );
  AND U16586 ( .A(n16077), .B(n16076), .Z(n16079) );
  NAND U16587 ( .A(n17308), .B(\stack[5][32] ), .Z(n16078) );
  NAND U16588 ( .A(n16079), .B(n16078), .Z(n2375) );
  NAND U16589 ( .A(\stack[3][32] ), .B(n17311), .Z(n16081) );
  NAND U16590 ( .A(n17305), .B(\stack[5][32] ), .Z(n16080) );
  AND U16591 ( .A(n16081), .B(n16080), .Z(n16083) );
  NAND U16592 ( .A(n17308), .B(\stack[4][32] ), .Z(n16082) );
  NAND U16593 ( .A(n16083), .B(n16082), .Z(n2376) );
  NAND U16594 ( .A(\stack[2][32] ), .B(n17311), .Z(n16085) );
  NAND U16595 ( .A(n17305), .B(\stack[4][32] ), .Z(n16084) );
  AND U16596 ( .A(n16085), .B(n16084), .Z(n16087) );
  NAND U16597 ( .A(n17308), .B(\stack[3][32] ), .Z(n16086) );
  NAND U16598 ( .A(n16087), .B(n16086), .Z(n2377) );
  NAND U16599 ( .A(n17311), .B(\stack[1][32] ), .Z(n16089) );
  NAND U16600 ( .A(n17305), .B(\stack[3][32] ), .Z(n16088) );
  AND U16601 ( .A(n16089), .B(n16088), .Z(n16091) );
  NAND U16602 ( .A(n17308), .B(\stack[2][32] ), .Z(n16090) );
  NAND U16603 ( .A(n16091), .B(n16090), .Z(n2378) );
  NAND U16604 ( .A(n17311), .B(o[32]), .Z(n16093) );
  NAND U16605 ( .A(n17305), .B(\stack[2][32] ), .Z(n16092) );
  AND U16606 ( .A(n16093), .B(n16092), .Z(n16095) );
  NAND U16607 ( .A(\stack[1][32] ), .B(n17308), .Z(n16094) );
  NAND U16608 ( .A(n16095), .B(n16094), .Z(n2379) );
  NAND U16609 ( .A(o[32]), .B(n17313), .Z(n16096) );
  NANDN U16610 ( .A(n17318), .B(n16096), .Z(n16097) );
  AND U16611 ( .A(\stack[1][32] ), .B(n16097), .Z(n16105) );
  NAND U16612 ( .A(x[32]), .B(n17311), .Z(n16098) );
  XNOR U16613 ( .A(n16100), .B(n16099), .Z(n16101) );
  NANDN U16614 ( .A(n17294), .B(n16101), .Z(n16102) );
  NAND U16615 ( .A(n16103), .B(n16102), .Z(n16104) );
  NOR U16616 ( .A(n16105), .B(n16104), .Z(n16107) );
  NANDN U16617 ( .A(n17317), .B(o[32]), .Z(n16106) );
  NAND U16618 ( .A(n16107), .B(n16106), .Z(n2380) );
  NAND U16619 ( .A(\stack[6][31] ), .B(n17311), .Z(n16109) );
  NANDN U16620 ( .A(n17311), .B(\stack[7][31] ), .Z(n16108) );
  NAND U16621 ( .A(n16109), .B(n16108), .Z(n2381) );
  NAND U16622 ( .A(\stack[5][31] ), .B(n17311), .Z(n16111) );
  NAND U16623 ( .A(n17305), .B(\stack[7][31] ), .Z(n16110) );
  AND U16624 ( .A(n16111), .B(n16110), .Z(n16113) );
  NAND U16625 ( .A(n17308), .B(\stack[6][31] ), .Z(n16112) );
  NAND U16626 ( .A(n16113), .B(n16112), .Z(n2382) );
  NAND U16627 ( .A(\stack[4][31] ), .B(n17311), .Z(n16115) );
  NAND U16628 ( .A(n17305), .B(\stack[6][31] ), .Z(n16114) );
  AND U16629 ( .A(n16115), .B(n16114), .Z(n16117) );
  NAND U16630 ( .A(n17308), .B(\stack[5][31] ), .Z(n16116) );
  NAND U16631 ( .A(n16117), .B(n16116), .Z(n2383) );
  NAND U16632 ( .A(\stack[3][31] ), .B(n17311), .Z(n16119) );
  NAND U16633 ( .A(n17305), .B(\stack[5][31] ), .Z(n16118) );
  AND U16634 ( .A(n16119), .B(n16118), .Z(n16121) );
  NAND U16635 ( .A(n17308), .B(\stack[4][31] ), .Z(n16120) );
  NAND U16636 ( .A(n16121), .B(n16120), .Z(n2384) );
  NAND U16637 ( .A(\stack[2][31] ), .B(n17311), .Z(n16123) );
  NAND U16638 ( .A(n17305), .B(\stack[4][31] ), .Z(n16122) );
  AND U16639 ( .A(n16123), .B(n16122), .Z(n16125) );
  NAND U16640 ( .A(n17308), .B(\stack[3][31] ), .Z(n16124) );
  NAND U16641 ( .A(n16125), .B(n16124), .Z(n2385) );
  NAND U16642 ( .A(n17311), .B(\stack[1][31] ), .Z(n16127) );
  NAND U16643 ( .A(n17305), .B(\stack[3][31] ), .Z(n16126) );
  AND U16644 ( .A(n16127), .B(n16126), .Z(n16129) );
  NAND U16645 ( .A(n17308), .B(\stack[2][31] ), .Z(n16128) );
  NAND U16646 ( .A(n16129), .B(n16128), .Z(n2386) );
  NAND U16647 ( .A(n17311), .B(o[31]), .Z(n16131) );
  NAND U16648 ( .A(n17305), .B(\stack[2][31] ), .Z(n16130) );
  AND U16649 ( .A(n16131), .B(n16130), .Z(n16133) );
  NAND U16650 ( .A(\stack[1][31] ), .B(n17308), .Z(n16132) );
  NAND U16651 ( .A(n16133), .B(n16132), .Z(n2387) );
  NAND U16652 ( .A(n17313), .B(o[31]), .Z(n16134) );
  NANDN U16653 ( .A(n17318), .B(n16134), .Z(n16135) );
  AND U16654 ( .A(\stack[1][31] ), .B(n16135), .Z(n16143) );
  NAND U16655 ( .A(x[31]), .B(n17311), .Z(n16136) );
  XNOR U16656 ( .A(n16138), .B(n16137), .Z(n16139) );
  NANDN U16657 ( .A(n17294), .B(n16139), .Z(n16140) );
  NAND U16658 ( .A(n16141), .B(n16140), .Z(n16142) );
  NOR U16659 ( .A(n16143), .B(n16142), .Z(n16145) );
  NANDN U16660 ( .A(n17317), .B(o[31]), .Z(n16144) );
  NAND U16661 ( .A(n16145), .B(n16144), .Z(n2388) );
  NAND U16662 ( .A(\stack[6][30] ), .B(n17311), .Z(n16147) );
  NANDN U16663 ( .A(n17311), .B(\stack[7][30] ), .Z(n16146) );
  NAND U16664 ( .A(n16147), .B(n16146), .Z(n2389) );
  NAND U16665 ( .A(\stack[5][30] ), .B(n17311), .Z(n16149) );
  NAND U16666 ( .A(n17305), .B(\stack[7][30] ), .Z(n16148) );
  AND U16667 ( .A(n16149), .B(n16148), .Z(n16151) );
  NAND U16668 ( .A(n17308), .B(\stack[6][30] ), .Z(n16150) );
  NAND U16669 ( .A(n16151), .B(n16150), .Z(n2390) );
  NAND U16670 ( .A(\stack[4][30] ), .B(n17311), .Z(n16153) );
  NAND U16671 ( .A(n17305), .B(\stack[6][30] ), .Z(n16152) );
  AND U16672 ( .A(n16153), .B(n16152), .Z(n16155) );
  NAND U16673 ( .A(n17308), .B(\stack[5][30] ), .Z(n16154) );
  NAND U16674 ( .A(n16155), .B(n16154), .Z(n2391) );
  NAND U16675 ( .A(\stack[3][30] ), .B(n17311), .Z(n16157) );
  NAND U16676 ( .A(n17305), .B(\stack[5][30] ), .Z(n16156) );
  AND U16677 ( .A(n16157), .B(n16156), .Z(n16159) );
  NAND U16678 ( .A(n17308), .B(\stack[4][30] ), .Z(n16158) );
  NAND U16679 ( .A(n16159), .B(n16158), .Z(n2392) );
  NAND U16680 ( .A(\stack[2][30] ), .B(n17311), .Z(n16161) );
  NAND U16681 ( .A(n17305), .B(\stack[4][30] ), .Z(n16160) );
  AND U16682 ( .A(n16161), .B(n16160), .Z(n16163) );
  NAND U16683 ( .A(n17308), .B(\stack[3][30] ), .Z(n16162) );
  NAND U16684 ( .A(n16163), .B(n16162), .Z(n2393) );
  NAND U16685 ( .A(n17311), .B(\stack[1][30] ), .Z(n16165) );
  NAND U16686 ( .A(n17305), .B(\stack[3][30] ), .Z(n16164) );
  AND U16687 ( .A(n16165), .B(n16164), .Z(n16167) );
  NAND U16688 ( .A(n17308), .B(\stack[2][30] ), .Z(n16166) );
  NAND U16689 ( .A(n16167), .B(n16166), .Z(n2394) );
  NAND U16690 ( .A(n17311), .B(o[30]), .Z(n16169) );
  NAND U16691 ( .A(n17305), .B(\stack[2][30] ), .Z(n16168) );
  AND U16692 ( .A(n16169), .B(n16168), .Z(n16171) );
  NAND U16693 ( .A(\stack[1][30] ), .B(n17308), .Z(n16170) );
  NAND U16694 ( .A(n16171), .B(n16170), .Z(n2395) );
  NAND U16695 ( .A(x[30]), .B(n17311), .Z(n16174) );
  NAND U16696 ( .A(n16172), .B(n17313), .Z(n16173) );
  NAND U16697 ( .A(n16174), .B(n16173), .Z(n16182) );
  NAND U16698 ( .A(n17318), .B(\stack[1][30] ), .Z(n16175) );
  XNOR U16699 ( .A(n16177), .B(n16176), .Z(n16178) );
  NANDN U16700 ( .A(n17294), .B(n16178), .Z(n16179) );
  NAND U16701 ( .A(n16180), .B(n16179), .Z(n16181) );
  NOR U16702 ( .A(n16182), .B(n16181), .Z(n16184) );
  NANDN U16703 ( .A(n17317), .B(o[30]), .Z(n16183) );
  NAND U16704 ( .A(n16184), .B(n16183), .Z(n2396) );
  NAND U16705 ( .A(\stack[6][29] ), .B(n17311), .Z(n16186) );
  NANDN U16706 ( .A(n17311), .B(\stack[7][29] ), .Z(n16185) );
  NAND U16707 ( .A(n16186), .B(n16185), .Z(n2397) );
  NAND U16708 ( .A(\stack[5][29] ), .B(n17311), .Z(n16188) );
  NAND U16709 ( .A(n17305), .B(\stack[7][29] ), .Z(n16187) );
  AND U16710 ( .A(n16188), .B(n16187), .Z(n16190) );
  NAND U16711 ( .A(n17308), .B(\stack[6][29] ), .Z(n16189) );
  NAND U16712 ( .A(n16190), .B(n16189), .Z(n2398) );
  NAND U16713 ( .A(\stack[4][29] ), .B(n17311), .Z(n16192) );
  NAND U16714 ( .A(n17305), .B(\stack[6][29] ), .Z(n16191) );
  AND U16715 ( .A(n16192), .B(n16191), .Z(n16194) );
  NAND U16716 ( .A(n17308), .B(\stack[5][29] ), .Z(n16193) );
  NAND U16717 ( .A(n16194), .B(n16193), .Z(n2399) );
  NAND U16718 ( .A(\stack[3][29] ), .B(n17311), .Z(n16196) );
  NAND U16719 ( .A(n17305), .B(\stack[5][29] ), .Z(n16195) );
  AND U16720 ( .A(n16196), .B(n16195), .Z(n16198) );
  NAND U16721 ( .A(n17308), .B(\stack[4][29] ), .Z(n16197) );
  NAND U16722 ( .A(n16198), .B(n16197), .Z(n2400) );
  NAND U16723 ( .A(\stack[2][29] ), .B(n17311), .Z(n16200) );
  NAND U16724 ( .A(n17305), .B(\stack[4][29] ), .Z(n16199) );
  AND U16725 ( .A(n16200), .B(n16199), .Z(n16202) );
  NAND U16726 ( .A(n17308), .B(\stack[3][29] ), .Z(n16201) );
  NAND U16727 ( .A(n16202), .B(n16201), .Z(n2401) );
  NAND U16728 ( .A(n17311), .B(\stack[1][29] ), .Z(n16204) );
  NAND U16729 ( .A(n17305), .B(\stack[3][29] ), .Z(n16203) );
  AND U16730 ( .A(n16204), .B(n16203), .Z(n16206) );
  NAND U16731 ( .A(n17308), .B(\stack[2][29] ), .Z(n16205) );
  NAND U16732 ( .A(n16206), .B(n16205), .Z(n2402) );
  NAND U16733 ( .A(n17311), .B(o[29]), .Z(n16208) );
  NAND U16734 ( .A(n17305), .B(\stack[2][29] ), .Z(n16207) );
  AND U16735 ( .A(n16208), .B(n16207), .Z(n16210) );
  NAND U16736 ( .A(\stack[1][29] ), .B(n17308), .Z(n16209) );
  NAND U16737 ( .A(n16210), .B(n16209), .Z(n2403) );
  NAND U16738 ( .A(n17313), .B(o[29]), .Z(n16211) );
  NANDN U16739 ( .A(n17318), .B(n16211), .Z(n16212) );
  AND U16740 ( .A(\stack[1][29] ), .B(n16212), .Z(n16220) );
  NAND U16741 ( .A(x[29]), .B(n17311), .Z(n16213) );
  XNOR U16742 ( .A(n16215), .B(n16214), .Z(n16216) );
  NANDN U16743 ( .A(n17294), .B(n16216), .Z(n16217) );
  NAND U16744 ( .A(n16218), .B(n16217), .Z(n16219) );
  NOR U16745 ( .A(n16220), .B(n16219), .Z(n16222) );
  NANDN U16746 ( .A(n17317), .B(o[29]), .Z(n16221) );
  NAND U16747 ( .A(n16222), .B(n16221), .Z(n2404) );
  NAND U16748 ( .A(\stack[6][28] ), .B(n17311), .Z(n16224) );
  NANDN U16749 ( .A(n17311), .B(\stack[7][28] ), .Z(n16223) );
  NAND U16750 ( .A(n16224), .B(n16223), .Z(n2405) );
  NAND U16751 ( .A(\stack[5][28] ), .B(n17311), .Z(n16226) );
  NAND U16752 ( .A(n17305), .B(\stack[7][28] ), .Z(n16225) );
  AND U16753 ( .A(n16226), .B(n16225), .Z(n16228) );
  NAND U16754 ( .A(n17308), .B(\stack[6][28] ), .Z(n16227) );
  NAND U16755 ( .A(n16228), .B(n16227), .Z(n2406) );
  NAND U16756 ( .A(\stack[4][28] ), .B(n17311), .Z(n16230) );
  NAND U16757 ( .A(n17305), .B(\stack[6][28] ), .Z(n16229) );
  AND U16758 ( .A(n16230), .B(n16229), .Z(n16232) );
  NAND U16759 ( .A(n17308), .B(\stack[5][28] ), .Z(n16231) );
  NAND U16760 ( .A(n16232), .B(n16231), .Z(n2407) );
  NAND U16761 ( .A(\stack[3][28] ), .B(n17311), .Z(n16234) );
  NAND U16762 ( .A(n17305), .B(\stack[5][28] ), .Z(n16233) );
  AND U16763 ( .A(n16234), .B(n16233), .Z(n16236) );
  NAND U16764 ( .A(n17308), .B(\stack[4][28] ), .Z(n16235) );
  NAND U16765 ( .A(n16236), .B(n16235), .Z(n2408) );
  NAND U16766 ( .A(\stack[2][28] ), .B(n17311), .Z(n16238) );
  NAND U16767 ( .A(n17305), .B(\stack[4][28] ), .Z(n16237) );
  AND U16768 ( .A(n16238), .B(n16237), .Z(n16240) );
  NAND U16769 ( .A(n17308), .B(\stack[3][28] ), .Z(n16239) );
  NAND U16770 ( .A(n16240), .B(n16239), .Z(n2409) );
  NAND U16771 ( .A(n17311), .B(\stack[1][28] ), .Z(n16242) );
  NAND U16772 ( .A(n17305), .B(\stack[3][28] ), .Z(n16241) );
  AND U16773 ( .A(n16242), .B(n16241), .Z(n16244) );
  NAND U16774 ( .A(n17308), .B(\stack[2][28] ), .Z(n16243) );
  NAND U16775 ( .A(n16244), .B(n16243), .Z(n2410) );
  NAND U16776 ( .A(n17311), .B(o[28]), .Z(n16246) );
  NAND U16777 ( .A(n17305), .B(\stack[2][28] ), .Z(n16245) );
  AND U16778 ( .A(n16246), .B(n16245), .Z(n16248) );
  NAND U16779 ( .A(\stack[1][28] ), .B(n17308), .Z(n16247) );
  NAND U16780 ( .A(n16248), .B(n16247), .Z(n2411) );
  NAND U16781 ( .A(x[28]), .B(n17311), .Z(n16250) );
  NAND U16782 ( .A(\stack[1][28] ), .B(n17318), .Z(n16249) );
  NAND U16783 ( .A(n16250), .B(n16249), .Z(n16259) );
  NAND U16784 ( .A(n17313), .B(n16251), .Z(n16252) );
  XNOR U16785 ( .A(n16254), .B(n16253), .Z(n16255) );
  NANDN U16786 ( .A(n17294), .B(n16255), .Z(n16256) );
  NAND U16787 ( .A(n16257), .B(n16256), .Z(n16258) );
  NOR U16788 ( .A(n16259), .B(n16258), .Z(n16261) );
  NANDN U16789 ( .A(n17317), .B(o[28]), .Z(n16260) );
  NAND U16790 ( .A(n16261), .B(n16260), .Z(n2412) );
  NAND U16791 ( .A(\stack[6][27] ), .B(n17311), .Z(n16263) );
  NANDN U16792 ( .A(n17311), .B(\stack[7][27] ), .Z(n16262) );
  NAND U16793 ( .A(n16263), .B(n16262), .Z(n2413) );
  NAND U16794 ( .A(\stack[5][27] ), .B(n17311), .Z(n16265) );
  NAND U16795 ( .A(n17305), .B(\stack[7][27] ), .Z(n16264) );
  AND U16796 ( .A(n16265), .B(n16264), .Z(n16267) );
  NAND U16797 ( .A(n17308), .B(\stack[6][27] ), .Z(n16266) );
  NAND U16798 ( .A(n16267), .B(n16266), .Z(n2414) );
  NAND U16799 ( .A(\stack[4][27] ), .B(n17311), .Z(n16269) );
  NAND U16800 ( .A(n17305), .B(\stack[6][27] ), .Z(n16268) );
  AND U16801 ( .A(n16269), .B(n16268), .Z(n16271) );
  NAND U16802 ( .A(n17308), .B(\stack[5][27] ), .Z(n16270) );
  NAND U16803 ( .A(n16271), .B(n16270), .Z(n2415) );
  NAND U16804 ( .A(\stack[3][27] ), .B(n17311), .Z(n16273) );
  NAND U16805 ( .A(n17305), .B(\stack[5][27] ), .Z(n16272) );
  AND U16806 ( .A(n16273), .B(n16272), .Z(n16275) );
  NAND U16807 ( .A(n17308), .B(\stack[4][27] ), .Z(n16274) );
  NAND U16808 ( .A(n16275), .B(n16274), .Z(n2416) );
  NAND U16809 ( .A(\stack[2][27] ), .B(n17311), .Z(n16277) );
  NAND U16810 ( .A(n17305), .B(\stack[4][27] ), .Z(n16276) );
  AND U16811 ( .A(n16277), .B(n16276), .Z(n16279) );
  NAND U16812 ( .A(n17308), .B(\stack[3][27] ), .Z(n16278) );
  NAND U16813 ( .A(n16279), .B(n16278), .Z(n2417) );
  NAND U16814 ( .A(n17311), .B(\stack[1][27] ), .Z(n16281) );
  NAND U16815 ( .A(n17305), .B(\stack[3][27] ), .Z(n16280) );
  AND U16816 ( .A(n16281), .B(n16280), .Z(n16283) );
  NAND U16817 ( .A(n17308), .B(\stack[2][27] ), .Z(n16282) );
  NAND U16818 ( .A(n16283), .B(n16282), .Z(n2418) );
  NAND U16819 ( .A(n17311), .B(o[27]), .Z(n16285) );
  NAND U16820 ( .A(n17305), .B(\stack[2][27] ), .Z(n16284) );
  AND U16821 ( .A(n16285), .B(n16284), .Z(n16287) );
  NAND U16822 ( .A(\stack[1][27] ), .B(n17308), .Z(n16286) );
  NAND U16823 ( .A(n16287), .B(n16286), .Z(n2419) );
  NAND U16824 ( .A(x[27]), .B(n17311), .Z(n16289) );
  NAND U16825 ( .A(\stack[1][27] ), .B(n17318), .Z(n16288) );
  NAND U16826 ( .A(n16289), .B(n16288), .Z(n16298) );
  NAND U16827 ( .A(n17313), .B(n16290), .Z(n16291) );
  XNOR U16828 ( .A(n16293), .B(n16292), .Z(n16294) );
  NANDN U16829 ( .A(n17294), .B(n16294), .Z(n16295) );
  NAND U16830 ( .A(n16296), .B(n16295), .Z(n16297) );
  NOR U16831 ( .A(n16298), .B(n16297), .Z(n16300) );
  NANDN U16832 ( .A(n17317), .B(o[27]), .Z(n16299) );
  NAND U16833 ( .A(n16300), .B(n16299), .Z(n2420) );
  NAND U16834 ( .A(\stack[6][26] ), .B(n17311), .Z(n16302) );
  NANDN U16835 ( .A(n17311), .B(\stack[7][26] ), .Z(n16301) );
  NAND U16836 ( .A(n16302), .B(n16301), .Z(n2421) );
  NAND U16837 ( .A(\stack[5][26] ), .B(n17311), .Z(n16304) );
  NAND U16838 ( .A(n17305), .B(\stack[7][26] ), .Z(n16303) );
  AND U16839 ( .A(n16304), .B(n16303), .Z(n16306) );
  NAND U16840 ( .A(n17308), .B(\stack[6][26] ), .Z(n16305) );
  NAND U16841 ( .A(n16306), .B(n16305), .Z(n2422) );
  NAND U16842 ( .A(\stack[4][26] ), .B(n17311), .Z(n16308) );
  NAND U16843 ( .A(n17305), .B(\stack[6][26] ), .Z(n16307) );
  AND U16844 ( .A(n16308), .B(n16307), .Z(n16310) );
  NAND U16845 ( .A(n17308), .B(\stack[5][26] ), .Z(n16309) );
  NAND U16846 ( .A(n16310), .B(n16309), .Z(n2423) );
  NAND U16847 ( .A(\stack[3][26] ), .B(n17311), .Z(n16312) );
  NAND U16848 ( .A(n17305), .B(\stack[5][26] ), .Z(n16311) );
  AND U16849 ( .A(n16312), .B(n16311), .Z(n16314) );
  NAND U16850 ( .A(n17308), .B(\stack[4][26] ), .Z(n16313) );
  NAND U16851 ( .A(n16314), .B(n16313), .Z(n2424) );
  NAND U16852 ( .A(\stack[2][26] ), .B(n17311), .Z(n16316) );
  NAND U16853 ( .A(n17305), .B(\stack[4][26] ), .Z(n16315) );
  AND U16854 ( .A(n16316), .B(n16315), .Z(n16318) );
  NAND U16855 ( .A(n17308), .B(\stack[3][26] ), .Z(n16317) );
  NAND U16856 ( .A(n16318), .B(n16317), .Z(n2425) );
  NAND U16857 ( .A(n17311), .B(\stack[1][26] ), .Z(n16320) );
  NAND U16858 ( .A(n17305), .B(\stack[3][26] ), .Z(n16319) );
  AND U16859 ( .A(n16320), .B(n16319), .Z(n16322) );
  NAND U16860 ( .A(n17308), .B(\stack[2][26] ), .Z(n16321) );
  NAND U16861 ( .A(n16322), .B(n16321), .Z(n2426) );
  NAND U16862 ( .A(n17311), .B(o[26]), .Z(n16324) );
  NAND U16863 ( .A(n17305), .B(\stack[2][26] ), .Z(n16323) );
  AND U16864 ( .A(n16324), .B(n16323), .Z(n16326) );
  NAND U16865 ( .A(\stack[1][26] ), .B(n17308), .Z(n16325) );
  NAND U16866 ( .A(n16326), .B(n16325), .Z(n2427) );
  NAND U16867 ( .A(x[26]), .B(n17311), .Z(n16329) );
  NAND U16868 ( .A(n16327), .B(n17313), .Z(n16328) );
  NAND U16869 ( .A(n16329), .B(n16328), .Z(n16337) );
  NAND U16870 ( .A(n17318), .B(\stack[1][26] ), .Z(n16330) );
  XNOR U16871 ( .A(n16332), .B(n16331), .Z(n16333) );
  NANDN U16872 ( .A(n17294), .B(n16333), .Z(n16334) );
  NAND U16873 ( .A(n16335), .B(n16334), .Z(n16336) );
  NOR U16874 ( .A(n16337), .B(n16336), .Z(n16339) );
  NANDN U16875 ( .A(n17317), .B(o[26]), .Z(n16338) );
  NAND U16876 ( .A(n16339), .B(n16338), .Z(n2428) );
  NAND U16877 ( .A(\stack[6][25] ), .B(n17311), .Z(n16341) );
  NANDN U16878 ( .A(n17311), .B(\stack[7][25] ), .Z(n16340) );
  NAND U16879 ( .A(n16341), .B(n16340), .Z(n2429) );
  NAND U16880 ( .A(\stack[5][25] ), .B(n17311), .Z(n16343) );
  NAND U16881 ( .A(n17305), .B(\stack[7][25] ), .Z(n16342) );
  AND U16882 ( .A(n16343), .B(n16342), .Z(n16345) );
  NAND U16883 ( .A(n17308), .B(\stack[6][25] ), .Z(n16344) );
  NAND U16884 ( .A(n16345), .B(n16344), .Z(n2430) );
  NAND U16885 ( .A(\stack[4][25] ), .B(n17311), .Z(n16347) );
  NAND U16886 ( .A(n17305), .B(\stack[6][25] ), .Z(n16346) );
  AND U16887 ( .A(n16347), .B(n16346), .Z(n16349) );
  NAND U16888 ( .A(n17308), .B(\stack[5][25] ), .Z(n16348) );
  NAND U16889 ( .A(n16349), .B(n16348), .Z(n2431) );
  NAND U16890 ( .A(\stack[3][25] ), .B(n17311), .Z(n16351) );
  NAND U16891 ( .A(n17305), .B(\stack[5][25] ), .Z(n16350) );
  AND U16892 ( .A(n16351), .B(n16350), .Z(n16353) );
  NAND U16893 ( .A(n17308), .B(\stack[4][25] ), .Z(n16352) );
  NAND U16894 ( .A(n16353), .B(n16352), .Z(n2432) );
  NAND U16895 ( .A(\stack[2][25] ), .B(n17311), .Z(n16355) );
  NAND U16896 ( .A(n17305), .B(\stack[4][25] ), .Z(n16354) );
  AND U16897 ( .A(n16355), .B(n16354), .Z(n16357) );
  NAND U16898 ( .A(n17308), .B(\stack[3][25] ), .Z(n16356) );
  NAND U16899 ( .A(n16357), .B(n16356), .Z(n2433) );
  NAND U16900 ( .A(n17311), .B(\stack[1][25] ), .Z(n16359) );
  NAND U16901 ( .A(n17305), .B(\stack[3][25] ), .Z(n16358) );
  AND U16902 ( .A(n16359), .B(n16358), .Z(n16361) );
  NAND U16903 ( .A(n17308), .B(\stack[2][25] ), .Z(n16360) );
  NAND U16904 ( .A(n16361), .B(n16360), .Z(n2434) );
  NAND U16905 ( .A(n17311), .B(o[25]), .Z(n16363) );
  NAND U16906 ( .A(n17305), .B(\stack[2][25] ), .Z(n16362) );
  AND U16907 ( .A(n16363), .B(n16362), .Z(n16365) );
  NAND U16908 ( .A(\stack[1][25] ), .B(n17308), .Z(n16364) );
  NAND U16909 ( .A(n16365), .B(n16364), .Z(n2435) );
  NAND U16910 ( .A(x[25]), .B(n17311), .Z(n16367) );
  NAND U16911 ( .A(\stack[1][25] ), .B(n17318), .Z(n16366) );
  NAND U16912 ( .A(n16367), .B(n16366), .Z(n16376) );
  NAND U16913 ( .A(n17313), .B(n16368), .Z(n16369) );
  XNOR U16914 ( .A(n16371), .B(n16370), .Z(n16372) );
  NANDN U16915 ( .A(n17294), .B(n16372), .Z(n16373) );
  NAND U16916 ( .A(n16374), .B(n16373), .Z(n16375) );
  NOR U16917 ( .A(n16376), .B(n16375), .Z(n16378) );
  NANDN U16918 ( .A(n17317), .B(o[25]), .Z(n16377) );
  NAND U16919 ( .A(n16378), .B(n16377), .Z(n2436) );
  NAND U16920 ( .A(\stack[6][24] ), .B(n17311), .Z(n16380) );
  NANDN U16921 ( .A(n17311), .B(\stack[7][24] ), .Z(n16379) );
  NAND U16922 ( .A(n16380), .B(n16379), .Z(n2437) );
  NAND U16923 ( .A(\stack[5][24] ), .B(n17311), .Z(n16382) );
  NAND U16924 ( .A(n17305), .B(\stack[7][24] ), .Z(n16381) );
  AND U16925 ( .A(n16382), .B(n16381), .Z(n16384) );
  NAND U16926 ( .A(n17308), .B(\stack[6][24] ), .Z(n16383) );
  NAND U16927 ( .A(n16384), .B(n16383), .Z(n2438) );
  NAND U16928 ( .A(\stack[4][24] ), .B(n17311), .Z(n16386) );
  NAND U16929 ( .A(n17305), .B(\stack[6][24] ), .Z(n16385) );
  AND U16930 ( .A(n16386), .B(n16385), .Z(n16388) );
  NAND U16931 ( .A(n17308), .B(\stack[5][24] ), .Z(n16387) );
  NAND U16932 ( .A(n16388), .B(n16387), .Z(n2439) );
  NAND U16933 ( .A(\stack[3][24] ), .B(n17311), .Z(n16390) );
  NAND U16934 ( .A(n17305), .B(\stack[5][24] ), .Z(n16389) );
  AND U16935 ( .A(n16390), .B(n16389), .Z(n16392) );
  NAND U16936 ( .A(n17308), .B(\stack[4][24] ), .Z(n16391) );
  NAND U16937 ( .A(n16392), .B(n16391), .Z(n2440) );
  NAND U16938 ( .A(\stack[2][24] ), .B(n17311), .Z(n16394) );
  NAND U16939 ( .A(n17305), .B(\stack[4][24] ), .Z(n16393) );
  AND U16940 ( .A(n16394), .B(n16393), .Z(n16396) );
  NAND U16941 ( .A(n17308), .B(\stack[3][24] ), .Z(n16395) );
  NAND U16942 ( .A(n16396), .B(n16395), .Z(n2441) );
  NAND U16943 ( .A(n17311), .B(\stack[1][24] ), .Z(n16398) );
  NAND U16944 ( .A(n17305), .B(\stack[3][24] ), .Z(n16397) );
  AND U16945 ( .A(n16398), .B(n16397), .Z(n16400) );
  NAND U16946 ( .A(n17308), .B(\stack[2][24] ), .Z(n16399) );
  NAND U16947 ( .A(n16400), .B(n16399), .Z(n2442) );
  NAND U16948 ( .A(n17311), .B(o[24]), .Z(n16402) );
  NAND U16949 ( .A(n17305), .B(\stack[2][24] ), .Z(n16401) );
  AND U16950 ( .A(n16402), .B(n16401), .Z(n16404) );
  NAND U16951 ( .A(\stack[1][24] ), .B(n17308), .Z(n16403) );
  NAND U16952 ( .A(n16404), .B(n16403), .Z(n2443) );
  NAND U16953 ( .A(n17313), .B(o[24]), .Z(n16405) );
  NANDN U16954 ( .A(n17318), .B(n16405), .Z(n16406) );
  AND U16955 ( .A(\stack[1][24] ), .B(n16406), .Z(n16414) );
  NAND U16956 ( .A(x[24]), .B(n17311), .Z(n16407) );
  XNOR U16957 ( .A(n16409), .B(n16408), .Z(n16410) );
  NANDN U16958 ( .A(n17294), .B(n16410), .Z(n16411) );
  NAND U16959 ( .A(n16412), .B(n16411), .Z(n16413) );
  NOR U16960 ( .A(n16414), .B(n16413), .Z(n16416) );
  NANDN U16961 ( .A(n17317), .B(o[24]), .Z(n16415) );
  NAND U16962 ( .A(n16416), .B(n16415), .Z(n2444) );
  NAND U16963 ( .A(\stack[6][23] ), .B(n17311), .Z(n16418) );
  NANDN U16964 ( .A(n17311), .B(\stack[7][23] ), .Z(n16417) );
  NAND U16965 ( .A(n16418), .B(n16417), .Z(n2445) );
  NAND U16966 ( .A(\stack[5][23] ), .B(n17311), .Z(n16420) );
  NAND U16967 ( .A(n17305), .B(\stack[7][23] ), .Z(n16419) );
  AND U16968 ( .A(n16420), .B(n16419), .Z(n16422) );
  NAND U16969 ( .A(n17308), .B(\stack[6][23] ), .Z(n16421) );
  NAND U16970 ( .A(n16422), .B(n16421), .Z(n2446) );
  NAND U16971 ( .A(\stack[4][23] ), .B(n17311), .Z(n16424) );
  NAND U16972 ( .A(n17305), .B(\stack[6][23] ), .Z(n16423) );
  AND U16973 ( .A(n16424), .B(n16423), .Z(n16426) );
  NAND U16974 ( .A(n17308), .B(\stack[5][23] ), .Z(n16425) );
  NAND U16975 ( .A(n16426), .B(n16425), .Z(n2447) );
  NAND U16976 ( .A(\stack[3][23] ), .B(n17311), .Z(n16428) );
  NAND U16977 ( .A(n17305), .B(\stack[5][23] ), .Z(n16427) );
  AND U16978 ( .A(n16428), .B(n16427), .Z(n16430) );
  NAND U16979 ( .A(n17308), .B(\stack[4][23] ), .Z(n16429) );
  NAND U16980 ( .A(n16430), .B(n16429), .Z(n2448) );
  NAND U16981 ( .A(\stack[2][23] ), .B(n17311), .Z(n16432) );
  NAND U16982 ( .A(n17305), .B(\stack[4][23] ), .Z(n16431) );
  AND U16983 ( .A(n16432), .B(n16431), .Z(n16434) );
  NAND U16984 ( .A(n17308), .B(\stack[3][23] ), .Z(n16433) );
  NAND U16985 ( .A(n16434), .B(n16433), .Z(n2449) );
  NAND U16986 ( .A(n17311), .B(\stack[1][23] ), .Z(n16436) );
  NAND U16987 ( .A(n17305), .B(\stack[3][23] ), .Z(n16435) );
  AND U16988 ( .A(n16436), .B(n16435), .Z(n16438) );
  NAND U16989 ( .A(n17308), .B(\stack[2][23] ), .Z(n16437) );
  NAND U16990 ( .A(n16438), .B(n16437), .Z(n2450) );
  NAND U16991 ( .A(n17311), .B(o[23]), .Z(n16440) );
  NAND U16992 ( .A(n17305), .B(\stack[2][23] ), .Z(n16439) );
  AND U16993 ( .A(n16440), .B(n16439), .Z(n16442) );
  NAND U16994 ( .A(\stack[1][23] ), .B(n17308), .Z(n16441) );
  NAND U16995 ( .A(n16442), .B(n16441), .Z(n2451) );
  NAND U16996 ( .A(n17313), .B(o[23]), .Z(n16443) );
  NANDN U16997 ( .A(n17318), .B(n16443), .Z(n16444) );
  AND U16998 ( .A(\stack[1][23] ), .B(n16444), .Z(n16452) );
  NAND U16999 ( .A(x[23]), .B(n17311), .Z(n16445) );
  XNOR U17000 ( .A(n16447), .B(n16446), .Z(n16448) );
  NANDN U17001 ( .A(n17294), .B(n16448), .Z(n16449) );
  NAND U17002 ( .A(n16450), .B(n16449), .Z(n16451) );
  NOR U17003 ( .A(n16452), .B(n16451), .Z(n16454) );
  NANDN U17004 ( .A(n17317), .B(o[23]), .Z(n16453) );
  NAND U17005 ( .A(n16454), .B(n16453), .Z(n2452) );
  NAND U17006 ( .A(\stack[6][22] ), .B(n17311), .Z(n16456) );
  NANDN U17007 ( .A(n17311), .B(\stack[7][22] ), .Z(n16455) );
  NAND U17008 ( .A(n16456), .B(n16455), .Z(n2453) );
  NAND U17009 ( .A(\stack[5][22] ), .B(n17311), .Z(n16458) );
  NAND U17010 ( .A(n17305), .B(\stack[7][22] ), .Z(n16457) );
  AND U17011 ( .A(n16458), .B(n16457), .Z(n16460) );
  NAND U17012 ( .A(n17308), .B(\stack[6][22] ), .Z(n16459) );
  NAND U17013 ( .A(n16460), .B(n16459), .Z(n2454) );
  NAND U17014 ( .A(\stack[4][22] ), .B(n17311), .Z(n16462) );
  NAND U17015 ( .A(n17305), .B(\stack[6][22] ), .Z(n16461) );
  AND U17016 ( .A(n16462), .B(n16461), .Z(n16464) );
  NAND U17017 ( .A(n17308), .B(\stack[5][22] ), .Z(n16463) );
  NAND U17018 ( .A(n16464), .B(n16463), .Z(n2455) );
  NAND U17019 ( .A(\stack[3][22] ), .B(n17311), .Z(n16466) );
  NAND U17020 ( .A(n17305), .B(\stack[5][22] ), .Z(n16465) );
  AND U17021 ( .A(n16466), .B(n16465), .Z(n16468) );
  NAND U17022 ( .A(n17308), .B(\stack[4][22] ), .Z(n16467) );
  NAND U17023 ( .A(n16468), .B(n16467), .Z(n2456) );
  NAND U17024 ( .A(\stack[2][22] ), .B(n17311), .Z(n16470) );
  NAND U17025 ( .A(n17305), .B(\stack[4][22] ), .Z(n16469) );
  AND U17026 ( .A(n16470), .B(n16469), .Z(n16472) );
  NAND U17027 ( .A(n17308), .B(\stack[3][22] ), .Z(n16471) );
  NAND U17028 ( .A(n16472), .B(n16471), .Z(n2457) );
  NAND U17029 ( .A(n17311), .B(\stack[1][22] ), .Z(n16474) );
  NAND U17030 ( .A(n17305), .B(\stack[3][22] ), .Z(n16473) );
  AND U17031 ( .A(n16474), .B(n16473), .Z(n16476) );
  NAND U17032 ( .A(n17308), .B(\stack[2][22] ), .Z(n16475) );
  NAND U17033 ( .A(n16476), .B(n16475), .Z(n2458) );
  NAND U17034 ( .A(n17311), .B(o[22]), .Z(n16478) );
  NAND U17035 ( .A(n17305), .B(\stack[2][22] ), .Z(n16477) );
  AND U17036 ( .A(n16478), .B(n16477), .Z(n16480) );
  NAND U17037 ( .A(\stack[1][22] ), .B(n17308), .Z(n16479) );
  NAND U17038 ( .A(n16480), .B(n16479), .Z(n2459) );
  NAND U17039 ( .A(o[22]), .B(n17313), .Z(n16481) );
  NANDN U17040 ( .A(n17318), .B(n16481), .Z(n16482) );
  AND U17041 ( .A(\stack[1][22] ), .B(n16482), .Z(n16490) );
  NAND U17042 ( .A(x[22]), .B(n17311), .Z(n16483) );
  XNOR U17043 ( .A(n16485), .B(n16484), .Z(n16486) );
  NANDN U17044 ( .A(n17294), .B(n16486), .Z(n16487) );
  NAND U17045 ( .A(n16488), .B(n16487), .Z(n16489) );
  NOR U17046 ( .A(n16490), .B(n16489), .Z(n16492) );
  NANDN U17047 ( .A(n17317), .B(o[22]), .Z(n16491) );
  NAND U17048 ( .A(n16492), .B(n16491), .Z(n2460) );
  NAND U17049 ( .A(\stack[6][21] ), .B(n17311), .Z(n16494) );
  NANDN U17050 ( .A(n17311), .B(\stack[7][21] ), .Z(n16493) );
  NAND U17051 ( .A(n16494), .B(n16493), .Z(n2461) );
  NAND U17052 ( .A(\stack[5][21] ), .B(n17311), .Z(n16496) );
  NAND U17053 ( .A(n17305), .B(\stack[7][21] ), .Z(n16495) );
  AND U17054 ( .A(n16496), .B(n16495), .Z(n16498) );
  NAND U17055 ( .A(n17308), .B(\stack[6][21] ), .Z(n16497) );
  NAND U17056 ( .A(n16498), .B(n16497), .Z(n2462) );
  NAND U17057 ( .A(\stack[4][21] ), .B(n17311), .Z(n16500) );
  NAND U17058 ( .A(n17305), .B(\stack[6][21] ), .Z(n16499) );
  AND U17059 ( .A(n16500), .B(n16499), .Z(n16502) );
  NAND U17060 ( .A(n17308), .B(\stack[5][21] ), .Z(n16501) );
  NAND U17061 ( .A(n16502), .B(n16501), .Z(n2463) );
  NAND U17062 ( .A(\stack[3][21] ), .B(n17311), .Z(n16504) );
  NAND U17063 ( .A(n17305), .B(\stack[5][21] ), .Z(n16503) );
  AND U17064 ( .A(n16504), .B(n16503), .Z(n16506) );
  NAND U17065 ( .A(n17308), .B(\stack[4][21] ), .Z(n16505) );
  NAND U17066 ( .A(n16506), .B(n16505), .Z(n2464) );
  NAND U17067 ( .A(\stack[2][21] ), .B(n17311), .Z(n16508) );
  NAND U17068 ( .A(n17305), .B(\stack[4][21] ), .Z(n16507) );
  AND U17069 ( .A(n16508), .B(n16507), .Z(n16510) );
  NAND U17070 ( .A(n17308), .B(\stack[3][21] ), .Z(n16509) );
  NAND U17071 ( .A(n16510), .B(n16509), .Z(n2465) );
  NAND U17072 ( .A(n17311), .B(\stack[1][21] ), .Z(n16512) );
  NAND U17073 ( .A(n17305), .B(\stack[3][21] ), .Z(n16511) );
  AND U17074 ( .A(n16512), .B(n16511), .Z(n16514) );
  NAND U17075 ( .A(n17308), .B(\stack[2][21] ), .Z(n16513) );
  NAND U17076 ( .A(n16514), .B(n16513), .Z(n2466) );
  NAND U17077 ( .A(n17311), .B(o[21]), .Z(n16516) );
  NAND U17078 ( .A(n17305), .B(\stack[2][21] ), .Z(n16515) );
  AND U17079 ( .A(n16516), .B(n16515), .Z(n16518) );
  NAND U17080 ( .A(\stack[1][21] ), .B(n17308), .Z(n16517) );
  NAND U17081 ( .A(n16518), .B(n16517), .Z(n2467) );
  NAND U17082 ( .A(x[21]), .B(n17311), .Z(n16520) );
  NAND U17083 ( .A(\stack[1][21] ), .B(n17318), .Z(n16519) );
  NAND U17084 ( .A(n16520), .B(n16519), .Z(n16529) );
  NAND U17085 ( .A(n17313), .B(n16521), .Z(n16522) );
  XNOR U17086 ( .A(n16524), .B(n16523), .Z(n16525) );
  NANDN U17087 ( .A(n17294), .B(n16525), .Z(n16526) );
  NAND U17088 ( .A(n16527), .B(n16526), .Z(n16528) );
  NOR U17089 ( .A(n16529), .B(n16528), .Z(n16531) );
  NANDN U17090 ( .A(n17317), .B(o[21]), .Z(n16530) );
  NAND U17091 ( .A(n16531), .B(n16530), .Z(n2468) );
  NAND U17092 ( .A(\stack[6][20] ), .B(n17311), .Z(n16533) );
  NANDN U17093 ( .A(n17311), .B(\stack[7][20] ), .Z(n16532) );
  NAND U17094 ( .A(n16533), .B(n16532), .Z(n2469) );
  NAND U17095 ( .A(\stack[5][20] ), .B(n17311), .Z(n16535) );
  NAND U17096 ( .A(n17305), .B(\stack[7][20] ), .Z(n16534) );
  AND U17097 ( .A(n16535), .B(n16534), .Z(n16537) );
  NAND U17098 ( .A(n17308), .B(\stack[6][20] ), .Z(n16536) );
  NAND U17099 ( .A(n16537), .B(n16536), .Z(n2470) );
  NAND U17100 ( .A(\stack[4][20] ), .B(n17311), .Z(n16539) );
  NAND U17101 ( .A(n17305), .B(\stack[6][20] ), .Z(n16538) );
  AND U17102 ( .A(n16539), .B(n16538), .Z(n16541) );
  NAND U17103 ( .A(n17308), .B(\stack[5][20] ), .Z(n16540) );
  NAND U17104 ( .A(n16541), .B(n16540), .Z(n2471) );
  NAND U17105 ( .A(\stack[3][20] ), .B(n17311), .Z(n16543) );
  NAND U17106 ( .A(n17305), .B(\stack[5][20] ), .Z(n16542) );
  AND U17107 ( .A(n16543), .B(n16542), .Z(n16545) );
  NAND U17108 ( .A(n17308), .B(\stack[4][20] ), .Z(n16544) );
  NAND U17109 ( .A(n16545), .B(n16544), .Z(n2472) );
  NAND U17110 ( .A(\stack[2][20] ), .B(n17311), .Z(n16547) );
  NAND U17111 ( .A(n17305), .B(\stack[4][20] ), .Z(n16546) );
  AND U17112 ( .A(n16547), .B(n16546), .Z(n16549) );
  NAND U17113 ( .A(n17308), .B(\stack[3][20] ), .Z(n16548) );
  NAND U17114 ( .A(n16549), .B(n16548), .Z(n2473) );
  NAND U17115 ( .A(n17311), .B(\stack[1][20] ), .Z(n16551) );
  NAND U17116 ( .A(n17305), .B(\stack[3][20] ), .Z(n16550) );
  AND U17117 ( .A(n16551), .B(n16550), .Z(n16553) );
  NAND U17118 ( .A(n17308), .B(\stack[2][20] ), .Z(n16552) );
  NAND U17119 ( .A(n16553), .B(n16552), .Z(n2474) );
  NAND U17120 ( .A(n17311), .B(o[20]), .Z(n16555) );
  NAND U17121 ( .A(n17305), .B(\stack[2][20] ), .Z(n16554) );
  AND U17122 ( .A(n16555), .B(n16554), .Z(n16557) );
  NAND U17123 ( .A(\stack[1][20] ), .B(n17308), .Z(n16556) );
  NAND U17124 ( .A(n16557), .B(n16556), .Z(n2475) );
  NAND U17125 ( .A(x[20]), .B(n17311), .Z(n16559) );
  NAND U17126 ( .A(\stack[1][20] ), .B(n17318), .Z(n16558) );
  NAND U17127 ( .A(n16559), .B(n16558), .Z(n16568) );
  NAND U17128 ( .A(n17313), .B(n16560), .Z(n16561) );
  XNOR U17129 ( .A(n16563), .B(n16562), .Z(n16564) );
  NANDN U17130 ( .A(n17294), .B(n16564), .Z(n16565) );
  NAND U17131 ( .A(n16566), .B(n16565), .Z(n16567) );
  NOR U17132 ( .A(n16568), .B(n16567), .Z(n16570) );
  NANDN U17133 ( .A(n17317), .B(o[20]), .Z(n16569) );
  NAND U17134 ( .A(n16570), .B(n16569), .Z(n2476) );
  NAND U17135 ( .A(\stack[6][19] ), .B(n17311), .Z(n16572) );
  NANDN U17136 ( .A(n17311), .B(\stack[7][19] ), .Z(n16571) );
  NAND U17137 ( .A(n16572), .B(n16571), .Z(n2477) );
  NAND U17138 ( .A(\stack[5][19] ), .B(n17311), .Z(n16574) );
  NAND U17139 ( .A(n17305), .B(\stack[7][19] ), .Z(n16573) );
  AND U17140 ( .A(n16574), .B(n16573), .Z(n16576) );
  NAND U17141 ( .A(n17308), .B(\stack[6][19] ), .Z(n16575) );
  NAND U17142 ( .A(n16576), .B(n16575), .Z(n2478) );
  NAND U17143 ( .A(\stack[4][19] ), .B(n17311), .Z(n16578) );
  NAND U17144 ( .A(n17305), .B(\stack[6][19] ), .Z(n16577) );
  AND U17145 ( .A(n16578), .B(n16577), .Z(n16580) );
  NAND U17146 ( .A(n17308), .B(\stack[5][19] ), .Z(n16579) );
  NAND U17147 ( .A(n16580), .B(n16579), .Z(n2479) );
  NAND U17148 ( .A(\stack[3][19] ), .B(n17311), .Z(n16582) );
  NAND U17149 ( .A(n17305), .B(\stack[5][19] ), .Z(n16581) );
  AND U17150 ( .A(n16582), .B(n16581), .Z(n16584) );
  NAND U17151 ( .A(n17308), .B(\stack[4][19] ), .Z(n16583) );
  NAND U17152 ( .A(n16584), .B(n16583), .Z(n2480) );
  NAND U17153 ( .A(\stack[2][19] ), .B(n17311), .Z(n16586) );
  NAND U17154 ( .A(n17305), .B(\stack[4][19] ), .Z(n16585) );
  AND U17155 ( .A(n16586), .B(n16585), .Z(n16588) );
  NAND U17156 ( .A(n17308), .B(\stack[3][19] ), .Z(n16587) );
  NAND U17157 ( .A(n16588), .B(n16587), .Z(n2481) );
  NAND U17158 ( .A(n17311), .B(\stack[1][19] ), .Z(n16590) );
  NAND U17159 ( .A(n17305), .B(\stack[3][19] ), .Z(n16589) );
  AND U17160 ( .A(n16590), .B(n16589), .Z(n16592) );
  NAND U17161 ( .A(n17308), .B(\stack[2][19] ), .Z(n16591) );
  NAND U17162 ( .A(n16592), .B(n16591), .Z(n2482) );
  NAND U17163 ( .A(n17311), .B(o[19]), .Z(n16594) );
  NAND U17164 ( .A(n17305), .B(\stack[2][19] ), .Z(n16593) );
  AND U17165 ( .A(n16594), .B(n16593), .Z(n16596) );
  NAND U17166 ( .A(\stack[1][19] ), .B(n17308), .Z(n16595) );
  NAND U17167 ( .A(n16596), .B(n16595), .Z(n2483) );
  NAND U17168 ( .A(n17313), .B(o[19]), .Z(n16597) );
  NANDN U17169 ( .A(n17318), .B(n16597), .Z(n16598) );
  AND U17170 ( .A(\stack[1][19] ), .B(n16598), .Z(n16606) );
  NAND U17171 ( .A(x[19]), .B(n17311), .Z(n16599) );
  XNOR U17172 ( .A(n16601), .B(n16600), .Z(n16602) );
  NANDN U17173 ( .A(n17294), .B(n16602), .Z(n16603) );
  NAND U17174 ( .A(n16604), .B(n16603), .Z(n16605) );
  NOR U17175 ( .A(n16606), .B(n16605), .Z(n16608) );
  NANDN U17176 ( .A(n17317), .B(o[19]), .Z(n16607) );
  NAND U17177 ( .A(n16608), .B(n16607), .Z(n2484) );
  NAND U17178 ( .A(\stack[6][18] ), .B(n17311), .Z(n16610) );
  NANDN U17179 ( .A(n17311), .B(\stack[7][18] ), .Z(n16609) );
  NAND U17180 ( .A(n16610), .B(n16609), .Z(n2485) );
  NAND U17181 ( .A(\stack[5][18] ), .B(n17311), .Z(n16612) );
  NAND U17182 ( .A(n17305), .B(\stack[7][18] ), .Z(n16611) );
  AND U17183 ( .A(n16612), .B(n16611), .Z(n16614) );
  NAND U17184 ( .A(n17308), .B(\stack[6][18] ), .Z(n16613) );
  NAND U17185 ( .A(n16614), .B(n16613), .Z(n2486) );
  NAND U17186 ( .A(\stack[4][18] ), .B(n17311), .Z(n16616) );
  NAND U17187 ( .A(n17305), .B(\stack[6][18] ), .Z(n16615) );
  AND U17188 ( .A(n16616), .B(n16615), .Z(n16618) );
  NAND U17189 ( .A(n17308), .B(\stack[5][18] ), .Z(n16617) );
  NAND U17190 ( .A(n16618), .B(n16617), .Z(n2487) );
  NAND U17191 ( .A(\stack[3][18] ), .B(n17311), .Z(n16620) );
  NAND U17192 ( .A(n17305), .B(\stack[5][18] ), .Z(n16619) );
  AND U17193 ( .A(n16620), .B(n16619), .Z(n16622) );
  NAND U17194 ( .A(n17308), .B(\stack[4][18] ), .Z(n16621) );
  NAND U17195 ( .A(n16622), .B(n16621), .Z(n2488) );
  NAND U17196 ( .A(\stack[2][18] ), .B(n17311), .Z(n16624) );
  NAND U17197 ( .A(n17305), .B(\stack[4][18] ), .Z(n16623) );
  AND U17198 ( .A(n16624), .B(n16623), .Z(n16626) );
  NAND U17199 ( .A(n17308), .B(\stack[3][18] ), .Z(n16625) );
  NAND U17200 ( .A(n16626), .B(n16625), .Z(n2489) );
  NAND U17201 ( .A(n17311), .B(\stack[1][18] ), .Z(n16628) );
  NAND U17202 ( .A(n17305), .B(\stack[3][18] ), .Z(n16627) );
  AND U17203 ( .A(n16628), .B(n16627), .Z(n16630) );
  NAND U17204 ( .A(n17308), .B(\stack[2][18] ), .Z(n16629) );
  NAND U17205 ( .A(n16630), .B(n16629), .Z(n2490) );
  NAND U17206 ( .A(n17311), .B(o[18]), .Z(n16632) );
  NAND U17207 ( .A(n17305), .B(\stack[2][18] ), .Z(n16631) );
  AND U17208 ( .A(n16632), .B(n16631), .Z(n16634) );
  NAND U17209 ( .A(\stack[1][18] ), .B(n17308), .Z(n16633) );
  NAND U17210 ( .A(n16634), .B(n16633), .Z(n2491) );
  NAND U17211 ( .A(x[18]), .B(n17311), .Z(n16636) );
  NAND U17212 ( .A(\stack[1][18] ), .B(n17318), .Z(n16635) );
  NAND U17213 ( .A(n16636), .B(n16635), .Z(n16645) );
  NAND U17214 ( .A(n17313), .B(n16637), .Z(n16638) );
  XNOR U17215 ( .A(n16640), .B(n16639), .Z(n16641) );
  NANDN U17216 ( .A(n17294), .B(n16641), .Z(n16642) );
  NAND U17217 ( .A(n16643), .B(n16642), .Z(n16644) );
  NOR U17218 ( .A(n16645), .B(n16644), .Z(n16647) );
  NANDN U17219 ( .A(n17317), .B(o[18]), .Z(n16646) );
  NAND U17220 ( .A(n16647), .B(n16646), .Z(n2492) );
  NAND U17221 ( .A(\stack[6][17] ), .B(n17311), .Z(n16649) );
  NANDN U17222 ( .A(n17311), .B(\stack[7][17] ), .Z(n16648) );
  NAND U17223 ( .A(n16649), .B(n16648), .Z(n2493) );
  NAND U17224 ( .A(\stack[5][17] ), .B(n17311), .Z(n16651) );
  NAND U17225 ( .A(n17305), .B(\stack[7][17] ), .Z(n16650) );
  AND U17226 ( .A(n16651), .B(n16650), .Z(n16653) );
  NAND U17227 ( .A(n17308), .B(\stack[6][17] ), .Z(n16652) );
  NAND U17228 ( .A(n16653), .B(n16652), .Z(n2494) );
  NAND U17229 ( .A(\stack[4][17] ), .B(n17311), .Z(n16655) );
  NAND U17230 ( .A(n17305), .B(\stack[6][17] ), .Z(n16654) );
  AND U17231 ( .A(n16655), .B(n16654), .Z(n16657) );
  NAND U17232 ( .A(n17308), .B(\stack[5][17] ), .Z(n16656) );
  NAND U17233 ( .A(n16657), .B(n16656), .Z(n2495) );
  NAND U17234 ( .A(\stack[3][17] ), .B(n17311), .Z(n16659) );
  NAND U17235 ( .A(n17305), .B(\stack[5][17] ), .Z(n16658) );
  AND U17236 ( .A(n16659), .B(n16658), .Z(n16661) );
  NAND U17237 ( .A(n17308), .B(\stack[4][17] ), .Z(n16660) );
  NAND U17238 ( .A(n16661), .B(n16660), .Z(n2496) );
  NAND U17239 ( .A(\stack[2][17] ), .B(n17311), .Z(n16663) );
  NAND U17240 ( .A(n17305), .B(\stack[4][17] ), .Z(n16662) );
  AND U17241 ( .A(n16663), .B(n16662), .Z(n16665) );
  NAND U17242 ( .A(n17308), .B(\stack[3][17] ), .Z(n16664) );
  NAND U17243 ( .A(n16665), .B(n16664), .Z(n2497) );
  NAND U17244 ( .A(n17311), .B(\stack[1][17] ), .Z(n16667) );
  NAND U17245 ( .A(n17305), .B(\stack[3][17] ), .Z(n16666) );
  AND U17246 ( .A(n16667), .B(n16666), .Z(n16669) );
  NAND U17247 ( .A(n17308), .B(\stack[2][17] ), .Z(n16668) );
  NAND U17248 ( .A(n16669), .B(n16668), .Z(n2498) );
  NAND U17249 ( .A(n17311), .B(o[17]), .Z(n16671) );
  NAND U17250 ( .A(n17305), .B(\stack[2][17] ), .Z(n16670) );
  AND U17251 ( .A(n16671), .B(n16670), .Z(n16673) );
  NAND U17252 ( .A(\stack[1][17] ), .B(n17308), .Z(n16672) );
  NAND U17253 ( .A(n16673), .B(n16672), .Z(n2499) );
  NAND U17254 ( .A(n17313), .B(o[17]), .Z(n16674) );
  NANDN U17255 ( .A(n17318), .B(n16674), .Z(n16675) );
  AND U17256 ( .A(\stack[1][17] ), .B(n16675), .Z(n16683) );
  NAND U17257 ( .A(x[17]), .B(n17311), .Z(n16676) );
  XNOR U17258 ( .A(n16678), .B(n16677), .Z(n16679) );
  NANDN U17259 ( .A(n17294), .B(n16679), .Z(n16680) );
  NAND U17260 ( .A(n16681), .B(n16680), .Z(n16682) );
  NOR U17261 ( .A(n16683), .B(n16682), .Z(n16685) );
  NANDN U17262 ( .A(n17317), .B(o[17]), .Z(n16684) );
  NAND U17263 ( .A(n16685), .B(n16684), .Z(n2500) );
  NAND U17264 ( .A(\stack[6][16] ), .B(n17311), .Z(n16687) );
  NANDN U17265 ( .A(n17311), .B(\stack[7][16] ), .Z(n16686) );
  NAND U17266 ( .A(n16687), .B(n16686), .Z(n2501) );
  NAND U17267 ( .A(\stack[5][16] ), .B(n17311), .Z(n16689) );
  NAND U17268 ( .A(n17305), .B(\stack[7][16] ), .Z(n16688) );
  AND U17269 ( .A(n16689), .B(n16688), .Z(n16691) );
  NAND U17270 ( .A(n17308), .B(\stack[6][16] ), .Z(n16690) );
  NAND U17271 ( .A(n16691), .B(n16690), .Z(n2502) );
  NAND U17272 ( .A(\stack[4][16] ), .B(n17311), .Z(n16693) );
  NAND U17273 ( .A(n17305), .B(\stack[6][16] ), .Z(n16692) );
  AND U17274 ( .A(n16693), .B(n16692), .Z(n16695) );
  NAND U17275 ( .A(n17308), .B(\stack[5][16] ), .Z(n16694) );
  NAND U17276 ( .A(n16695), .B(n16694), .Z(n2503) );
  NAND U17277 ( .A(\stack[3][16] ), .B(n17311), .Z(n16697) );
  NAND U17278 ( .A(n17305), .B(\stack[5][16] ), .Z(n16696) );
  AND U17279 ( .A(n16697), .B(n16696), .Z(n16699) );
  NAND U17280 ( .A(n17308), .B(\stack[4][16] ), .Z(n16698) );
  NAND U17281 ( .A(n16699), .B(n16698), .Z(n2504) );
  NAND U17282 ( .A(\stack[2][16] ), .B(n17311), .Z(n16701) );
  NAND U17283 ( .A(n17305), .B(\stack[4][16] ), .Z(n16700) );
  AND U17284 ( .A(n16701), .B(n16700), .Z(n16703) );
  NAND U17285 ( .A(n17308), .B(\stack[3][16] ), .Z(n16702) );
  NAND U17286 ( .A(n16703), .B(n16702), .Z(n2505) );
  NAND U17287 ( .A(n17311), .B(\stack[1][16] ), .Z(n16705) );
  NAND U17288 ( .A(n17305), .B(\stack[3][16] ), .Z(n16704) );
  AND U17289 ( .A(n16705), .B(n16704), .Z(n16707) );
  NAND U17290 ( .A(n17308), .B(\stack[2][16] ), .Z(n16706) );
  NAND U17291 ( .A(n16707), .B(n16706), .Z(n2506) );
  NAND U17292 ( .A(n17311), .B(o[16]), .Z(n16709) );
  NAND U17293 ( .A(n17305), .B(\stack[2][16] ), .Z(n16708) );
  AND U17294 ( .A(n16709), .B(n16708), .Z(n16711) );
  NAND U17295 ( .A(\stack[1][16] ), .B(n17308), .Z(n16710) );
  NAND U17296 ( .A(n16711), .B(n16710), .Z(n2507) );
  NAND U17297 ( .A(x[16]), .B(n17311), .Z(n16713) );
  NAND U17298 ( .A(\stack[1][16] ), .B(n17318), .Z(n16712) );
  NAND U17299 ( .A(n16713), .B(n16712), .Z(n16722) );
  NAND U17300 ( .A(n17313), .B(n16714), .Z(n16715) );
  XNOR U17301 ( .A(n16717), .B(n16716), .Z(n16718) );
  NANDN U17302 ( .A(n17294), .B(n16718), .Z(n16719) );
  NAND U17303 ( .A(n16720), .B(n16719), .Z(n16721) );
  NOR U17304 ( .A(n16722), .B(n16721), .Z(n16724) );
  NANDN U17305 ( .A(n17317), .B(o[16]), .Z(n16723) );
  NAND U17306 ( .A(n16724), .B(n16723), .Z(n2508) );
  NAND U17307 ( .A(\stack[6][15] ), .B(n17311), .Z(n16726) );
  NANDN U17308 ( .A(n17311), .B(\stack[7][15] ), .Z(n16725) );
  NAND U17309 ( .A(n16726), .B(n16725), .Z(n2509) );
  NAND U17310 ( .A(\stack[5][15] ), .B(n17311), .Z(n16728) );
  NAND U17311 ( .A(n17305), .B(\stack[7][15] ), .Z(n16727) );
  AND U17312 ( .A(n16728), .B(n16727), .Z(n16730) );
  NAND U17313 ( .A(n17308), .B(\stack[6][15] ), .Z(n16729) );
  NAND U17314 ( .A(n16730), .B(n16729), .Z(n2510) );
  NAND U17315 ( .A(\stack[4][15] ), .B(n17311), .Z(n16732) );
  NAND U17316 ( .A(n17305), .B(\stack[6][15] ), .Z(n16731) );
  AND U17317 ( .A(n16732), .B(n16731), .Z(n16734) );
  NAND U17318 ( .A(n17308), .B(\stack[5][15] ), .Z(n16733) );
  NAND U17319 ( .A(n16734), .B(n16733), .Z(n2511) );
  NAND U17320 ( .A(\stack[3][15] ), .B(n17311), .Z(n16736) );
  NAND U17321 ( .A(n17305), .B(\stack[5][15] ), .Z(n16735) );
  AND U17322 ( .A(n16736), .B(n16735), .Z(n16738) );
  NAND U17323 ( .A(n17308), .B(\stack[4][15] ), .Z(n16737) );
  NAND U17324 ( .A(n16738), .B(n16737), .Z(n2512) );
  NAND U17325 ( .A(\stack[2][15] ), .B(n17311), .Z(n16740) );
  NAND U17326 ( .A(n17305), .B(\stack[4][15] ), .Z(n16739) );
  AND U17327 ( .A(n16740), .B(n16739), .Z(n16742) );
  NAND U17328 ( .A(n17308), .B(\stack[3][15] ), .Z(n16741) );
  NAND U17329 ( .A(n16742), .B(n16741), .Z(n2513) );
  NAND U17330 ( .A(n17311), .B(\stack[1][15] ), .Z(n16744) );
  NAND U17331 ( .A(n17305), .B(\stack[3][15] ), .Z(n16743) );
  AND U17332 ( .A(n16744), .B(n16743), .Z(n16746) );
  NAND U17333 ( .A(n17308), .B(\stack[2][15] ), .Z(n16745) );
  NAND U17334 ( .A(n16746), .B(n16745), .Z(n2514) );
  NAND U17335 ( .A(n17311), .B(o[15]), .Z(n16748) );
  NAND U17336 ( .A(n17305), .B(\stack[2][15] ), .Z(n16747) );
  AND U17337 ( .A(n16748), .B(n16747), .Z(n16750) );
  NAND U17338 ( .A(\stack[1][15] ), .B(n17308), .Z(n16749) );
  NAND U17339 ( .A(n16750), .B(n16749), .Z(n2515) );
  NAND U17340 ( .A(o[15]), .B(n17313), .Z(n16751) );
  NANDN U17341 ( .A(n17318), .B(n16751), .Z(n16752) );
  AND U17342 ( .A(\stack[1][15] ), .B(n16752), .Z(n16760) );
  NAND U17343 ( .A(x[15]), .B(n17311), .Z(n16753) );
  XNOR U17344 ( .A(n16755), .B(n16754), .Z(n16756) );
  NANDN U17345 ( .A(n17294), .B(n16756), .Z(n16757) );
  NAND U17346 ( .A(n16758), .B(n16757), .Z(n16759) );
  NOR U17347 ( .A(n16760), .B(n16759), .Z(n16762) );
  NANDN U17348 ( .A(n17317), .B(o[15]), .Z(n16761) );
  NAND U17349 ( .A(n16762), .B(n16761), .Z(n2516) );
  NAND U17350 ( .A(\stack[6][14] ), .B(n17311), .Z(n16764) );
  NANDN U17351 ( .A(n17311), .B(\stack[7][14] ), .Z(n16763) );
  NAND U17352 ( .A(n16764), .B(n16763), .Z(n2517) );
  NAND U17353 ( .A(\stack[5][14] ), .B(n17311), .Z(n16766) );
  NAND U17354 ( .A(n17305), .B(\stack[7][14] ), .Z(n16765) );
  AND U17355 ( .A(n16766), .B(n16765), .Z(n16768) );
  NAND U17356 ( .A(n17308), .B(\stack[6][14] ), .Z(n16767) );
  NAND U17357 ( .A(n16768), .B(n16767), .Z(n2518) );
  NAND U17358 ( .A(\stack[4][14] ), .B(n17311), .Z(n16770) );
  NAND U17359 ( .A(n17305), .B(\stack[6][14] ), .Z(n16769) );
  AND U17360 ( .A(n16770), .B(n16769), .Z(n16772) );
  NAND U17361 ( .A(n17308), .B(\stack[5][14] ), .Z(n16771) );
  NAND U17362 ( .A(n16772), .B(n16771), .Z(n2519) );
  NAND U17363 ( .A(\stack[3][14] ), .B(n17311), .Z(n16774) );
  NAND U17364 ( .A(n17305), .B(\stack[5][14] ), .Z(n16773) );
  AND U17365 ( .A(n16774), .B(n16773), .Z(n16776) );
  NAND U17366 ( .A(n17308), .B(\stack[4][14] ), .Z(n16775) );
  NAND U17367 ( .A(n16776), .B(n16775), .Z(n2520) );
  NAND U17368 ( .A(\stack[2][14] ), .B(n17311), .Z(n16778) );
  NAND U17369 ( .A(n17305), .B(\stack[4][14] ), .Z(n16777) );
  AND U17370 ( .A(n16778), .B(n16777), .Z(n16780) );
  NAND U17371 ( .A(n17308), .B(\stack[3][14] ), .Z(n16779) );
  NAND U17372 ( .A(n16780), .B(n16779), .Z(n2521) );
  NAND U17373 ( .A(n17311), .B(\stack[1][14] ), .Z(n16782) );
  NAND U17374 ( .A(n17305), .B(\stack[3][14] ), .Z(n16781) );
  AND U17375 ( .A(n16782), .B(n16781), .Z(n16784) );
  NAND U17376 ( .A(n17308), .B(\stack[2][14] ), .Z(n16783) );
  NAND U17377 ( .A(n16784), .B(n16783), .Z(n2522) );
  NAND U17378 ( .A(n17311), .B(o[14]), .Z(n16786) );
  NAND U17379 ( .A(n17305), .B(\stack[2][14] ), .Z(n16785) );
  AND U17380 ( .A(n16786), .B(n16785), .Z(n16788) );
  NAND U17381 ( .A(\stack[1][14] ), .B(n17308), .Z(n16787) );
  NAND U17382 ( .A(n16788), .B(n16787), .Z(n2523) );
  NAND U17383 ( .A(n17313), .B(o[14]), .Z(n16789) );
  NANDN U17384 ( .A(n17318), .B(n16789), .Z(n16790) );
  AND U17385 ( .A(\stack[1][14] ), .B(n16790), .Z(n16798) );
  NAND U17386 ( .A(x[14]), .B(n17311), .Z(n16791) );
  XNOR U17387 ( .A(n16793), .B(n16792), .Z(n16794) );
  NANDN U17388 ( .A(n17294), .B(n16794), .Z(n16795) );
  NAND U17389 ( .A(n16796), .B(n16795), .Z(n16797) );
  NOR U17390 ( .A(n16798), .B(n16797), .Z(n16800) );
  NANDN U17391 ( .A(n17317), .B(o[14]), .Z(n16799) );
  NAND U17392 ( .A(n16800), .B(n16799), .Z(n2524) );
  NAND U17393 ( .A(\stack[6][13] ), .B(n17311), .Z(n16802) );
  NANDN U17394 ( .A(n17311), .B(\stack[7][13] ), .Z(n16801) );
  NAND U17395 ( .A(n16802), .B(n16801), .Z(n2525) );
  NAND U17396 ( .A(\stack[5][13] ), .B(n17311), .Z(n16804) );
  NAND U17397 ( .A(n17305), .B(\stack[7][13] ), .Z(n16803) );
  AND U17398 ( .A(n16804), .B(n16803), .Z(n16806) );
  NAND U17399 ( .A(n17308), .B(\stack[6][13] ), .Z(n16805) );
  NAND U17400 ( .A(n16806), .B(n16805), .Z(n2526) );
  NAND U17401 ( .A(\stack[4][13] ), .B(n17311), .Z(n16808) );
  NAND U17402 ( .A(n17305), .B(\stack[6][13] ), .Z(n16807) );
  AND U17403 ( .A(n16808), .B(n16807), .Z(n16810) );
  NAND U17404 ( .A(n17308), .B(\stack[5][13] ), .Z(n16809) );
  NAND U17405 ( .A(n16810), .B(n16809), .Z(n2527) );
  NAND U17406 ( .A(\stack[3][13] ), .B(n17311), .Z(n16812) );
  NAND U17407 ( .A(n17305), .B(\stack[5][13] ), .Z(n16811) );
  AND U17408 ( .A(n16812), .B(n16811), .Z(n16814) );
  NAND U17409 ( .A(n17308), .B(\stack[4][13] ), .Z(n16813) );
  NAND U17410 ( .A(n16814), .B(n16813), .Z(n2528) );
  NAND U17411 ( .A(\stack[2][13] ), .B(n17311), .Z(n16816) );
  NAND U17412 ( .A(n17305), .B(\stack[4][13] ), .Z(n16815) );
  AND U17413 ( .A(n16816), .B(n16815), .Z(n16818) );
  NAND U17414 ( .A(n17308), .B(\stack[3][13] ), .Z(n16817) );
  NAND U17415 ( .A(n16818), .B(n16817), .Z(n2529) );
  NAND U17416 ( .A(n17311), .B(\stack[1][13] ), .Z(n16820) );
  NAND U17417 ( .A(n17305), .B(\stack[3][13] ), .Z(n16819) );
  AND U17418 ( .A(n16820), .B(n16819), .Z(n16822) );
  NAND U17419 ( .A(n17308), .B(\stack[2][13] ), .Z(n16821) );
  NAND U17420 ( .A(n16822), .B(n16821), .Z(n2530) );
  NAND U17421 ( .A(n17311), .B(o[13]), .Z(n16824) );
  NAND U17422 ( .A(n17305), .B(\stack[2][13] ), .Z(n16823) );
  AND U17423 ( .A(n16824), .B(n16823), .Z(n16826) );
  NAND U17424 ( .A(\stack[1][13] ), .B(n17308), .Z(n16825) );
  NAND U17425 ( .A(n16826), .B(n16825), .Z(n2531) );
  NAND U17426 ( .A(x[13]), .B(n17311), .Z(n16828) );
  NAND U17427 ( .A(\stack[1][13] ), .B(n17318), .Z(n16827) );
  NAND U17428 ( .A(n16828), .B(n16827), .Z(n16837) );
  NAND U17429 ( .A(n17313), .B(n16829), .Z(n16830) );
  XNOR U17430 ( .A(n16832), .B(n16831), .Z(n16833) );
  NANDN U17431 ( .A(n17294), .B(n16833), .Z(n16834) );
  NAND U17432 ( .A(n16835), .B(n16834), .Z(n16836) );
  NOR U17433 ( .A(n16837), .B(n16836), .Z(n16839) );
  NANDN U17434 ( .A(n17317), .B(o[13]), .Z(n16838) );
  NAND U17435 ( .A(n16839), .B(n16838), .Z(n2532) );
  NAND U17436 ( .A(\stack[6][12] ), .B(n17311), .Z(n16841) );
  NANDN U17437 ( .A(n17311), .B(\stack[7][12] ), .Z(n16840) );
  NAND U17438 ( .A(n16841), .B(n16840), .Z(n2533) );
  NAND U17439 ( .A(\stack[5][12] ), .B(n17311), .Z(n16843) );
  NAND U17440 ( .A(n17305), .B(\stack[7][12] ), .Z(n16842) );
  AND U17441 ( .A(n16843), .B(n16842), .Z(n16845) );
  NAND U17442 ( .A(n17308), .B(\stack[6][12] ), .Z(n16844) );
  NAND U17443 ( .A(n16845), .B(n16844), .Z(n2534) );
  NAND U17444 ( .A(\stack[4][12] ), .B(n17311), .Z(n16847) );
  NAND U17445 ( .A(n17305), .B(\stack[6][12] ), .Z(n16846) );
  AND U17446 ( .A(n16847), .B(n16846), .Z(n16849) );
  NAND U17447 ( .A(n17308), .B(\stack[5][12] ), .Z(n16848) );
  NAND U17448 ( .A(n16849), .B(n16848), .Z(n2535) );
  NAND U17449 ( .A(\stack[3][12] ), .B(n17311), .Z(n16851) );
  NAND U17450 ( .A(n17305), .B(\stack[5][12] ), .Z(n16850) );
  AND U17451 ( .A(n16851), .B(n16850), .Z(n16853) );
  NAND U17452 ( .A(n17308), .B(\stack[4][12] ), .Z(n16852) );
  NAND U17453 ( .A(n16853), .B(n16852), .Z(n2536) );
  NAND U17454 ( .A(\stack[2][12] ), .B(n17311), .Z(n16855) );
  NAND U17455 ( .A(n17305), .B(\stack[4][12] ), .Z(n16854) );
  AND U17456 ( .A(n16855), .B(n16854), .Z(n16857) );
  NAND U17457 ( .A(n17308), .B(\stack[3][12] ), .Z(n16856) );
  NAND U17458 ( .A(n16857), .B(n16856), .Z(n2537) );
  NAND U17459 ( .A(n17311), .B(\stack[1][12] ), .Z(n16859) );
  NAND U17460 ( .A(n17305), .B(\stack[3][12] ), .Z(n16858) );
  AND U17461 ( .A(n16859), .B(n16858), .Z(n16861) );
  NAND U17462 ( .A(n17308), .B(\stack[2][12] ), .Z(n16860) );
  NAND U17463 ( .A(n16861), .B(n16860), .Z(n2538) );
  NAND U17464 ( .A(n17311), .B(o[12]), .Z(n16863) );
  NAND U17465 ( .A(n17305), .B(\stack[2][12] ), .Z(n16862) );
  AND U17466 ( .A(n16863), .B(n16862), .Z(n16865) );
  NAND U17467 ( .A(\stack[1][12] ), .B(n17308), .Z(n16864) );
  NAND U17468 ( .A(n16865), .B(n16864), .Z(n2539) );
  NAND U17469 ( .A(x[12]), .B(n17311), .Z(n16867) );
  NAND U17470 ( .A(\stack[1][12] ), .B(n17318), .Z(n16866) );
  NAND U17471 ( .A(n16867), .B(n16866), .Z(n16876) );
  NAND U17472 ( .A(n16868), .B(n17313), .Z(n16869) );
  XNOR U17473 ( .A(n16871), .B(n16870), .Z(n16872) );
  NANDN U17474 ( .A(n17294), .B(n16872), .Z(n16873) );
  NAND U17475 ( .A(n16874), .B(n16873), .Z(n16875) );
  NOR U17476 ( .A(n16876), .B(n16875), .Z(n16878) );
  NANDN U17477 ( .A(n17317), .B(o[12]), .Z(n16877) );
  NAND U17478 ( .A(n16878), .B(n16877), .Z(n2540) );
  NAND U17479 ( .A(\stack[6][11] ), .B(n17311), .Z(n16880) );
  NANDN U17480 ( .A(n17311), .B(\stack[7][11] ), .Z(n16879) );
  NAND U17481 ( .A(n16880), .B(n16879), .Z(n2541) );
  NAND U17482 ( .A(\stack[5][11] ), .B(n17311), .Z(n16882) );
  NAND U17483 ( .A(n17305), .B(\stack[7][11] ), .Z(n16881) );
  AND U17484 ( .A(n16882), .B(n16881), .Z(n16884) );
  NAND U17485 ( .A(n17308), .B(\stack[6][11] ), .Z(n16883) );
  NAND U17486 ( .A(n16884), .B(n16883), .Z(n2542) );
  NAND U17487 ( .A(\stack[4][11] ), .B(n17311), .Z(n16886) );
  NAND U17488 ( .A(n17305), .B(\stack[6][11] ), .Z(n16885) );
  AND U17489 ( .A(n16886), .B(n16885), .Z(n16888) );
  NAND U17490 ( .A(n17308), .B(\stack[5][11] ), .Z(n16887) );
  NAND U17491 ( .A(n16888), .B(n16887), .Z(n2543) );
  NAND U17492 ( .A(\stack[3][11] ), .B(n17311), .Z(n16890) );
  NAND U17493 ( .A(n17305), .B(\stack[5][11] ), .Z(n16889) );
  AND U17494 ( .A(n16890), .B(n16889), .Z(n16892) );
  NAND U17495 ( .A(n17308), .B(\stack[4][11] ), .Z(n16891) );
  NAND U17496 ( .A(n16892), .B(n16891), .Z(n2544) );
  NAND U17497 ( .A(\stack[2][11] ), .B(n17311), .Z(n16894) );
  NAND U17498 ( .A(n17305), .B(\stack[4][11] ), .Z(n16893) );
  AND U17499 ( .A(n16894), .B(n16893), .Z(n16896) );
  NAND U17500 ( .A(n17308), .B(\stack[3][11] ), .Z(n16895) );
  NAND U17501 ( .A(n16896), .B(n16895), .Z(n2545) );
  NAND U17502 ( .A(n17311), .B(\stack[1][11] ), .Z(n16898) );
  NAND U17503 ( .A(n17305), .B(\stack[3][11] ), .Z(n16897) );
  AND U17504 ( .A(n16898), .B(n16897), .Z(n16900) );
  NAND U17505 ( .A(n17308), .B(\stack[2][11] ), .Z(n16899) );
  NAND U17506 ( .A(n16900), .B(n16899), .Z(n2546) );
  NAND U17507 ( .A(n17311), .B(o[11]), .Z(n16902) );
  NAND U17508 ( .A(n17305), .B(\stack[2][11] ), .Z(n16901) );
  AND U17509 ( .A(n16902), .B(n16901), .Z(n16904) );
  NAND U17510 ( .A(\stack[1][11] ), .B(n17308), .Z(n16903) );
  NAND U17511 ( .A(n16904), .B(n16903), .Z(n2547) );
  NAND U17512 ( .A(\stack[1][11] ), .B(n17318), .Z(n16905) );
  NANDN U17513 ( .A(o[11]), .B(n16905), .Z(n16906) );
  ANDN U17514 ( .B(n16906), .A(n17317), .Z(n16916) );
  NAND U17515 ( .A(x[11]), .B(n17311), .Z(n16909) );
  NANDN U17516 ( .A(n16907), .B(n17313), .Z(n16908) );
  AND U17517 ( .A(n16909), .B(n16908), .Z(n16914) );
  XNOR U17518 ( .A(n16911), .B(n16910), .Z(n16912) );
  NANDN U17519 ( .A(n17294), .B(n16912), .Z(n16913) );
  NAND U17520 ( .A(n16914), .B(n16913), .Z(n16915) );
  NOR U17521 ( .A(n16916), .B(n16915), .Z(n16917) );
  NAND U17522 ( .A(\stack[6][10] ), .B(n17311), .Z(n16919) );
  NANDN U17523 ( .A(n17311), .B(\stack[7][10] ), .Z(n16918) );
  NAND U17524 ( .A(n16919), .B(n16918), .Z(n2549) );
  NAND U17525 ( .A(\stack[5][10] ), .B(n17311), .Z(n16921) );
  NAND U17526 ( .A(n17305), .B(\stack[7][10] ), .Z(n16920) );
  AND U17527 ( .A(n16921), .B(n16920), .Z(n16923) );
  NAND U17528 ( .A(n17308), .B(\stack[6][10] ), .Z(n16922) );
  NAND U17529 ( .A(n16923), .B(n16922), .Z(n2550) );
  NAND U17530 ( .A(\stack[4][10] ), .B(n17311), .Z(n16925) );
  NAND U17531 ( .A(n17305), .B(\stack[6][10] ), .Z(n16924) );
  AND U17532 ( .A(n16925), .B(n16924), .Z(n16927) );
  NAND U17533 ( .A(n17308), .B(\stack[5][10] ), .Z(n16926) );
  NAND U17534 ( .A(n16927), .B(n16926), .Z(n2551) );
  NAND U17535 ( .A(\stack[3][10] ), .B(n17311), .Z(n16929) );
  NAND U17536 ( .A(n17305), .B(\stack[5][10] ), .Z(n16928) );
  AND U17537 ( .A(n16929), .B(n16928), .Z(n16931) );
  NAND U17538 ( .A(n17308), .B(\stack[4][10] ), .Z(n16930) );
  NAND U17539 ( .A(n16931), .B(n16930), .Z(n2552) );
  NAND U17540 ( .A(\stack[2][10] ), .B(n17311), .Z(n16933) );
  NAND U17541 ( .A(n17305), .B(\stack[4][10] ), .Z(n16932) );
  AND U17542 ( .A(n16933), .B(n16932), .Z(n16935) );
  NAND U17543 ( .A(n17308), .B(\stack[3][10] ), .Z(n16934) );
  NAND U17544 ( .A(n16935), .B(n16934), .Z(n2553) );
  NAND U17545 ( .A(n17311), .B(\stack[1][10] ), .Z(n16937) );
  NAND U17546 ( .A(n17305), .B(\stack[3][10] ), .Z(n16936) );
  AND U17547 ( .A(n16937), .B(n16936), .Z(n16939) );
  NAND U17548 ( .A(n17308), .B(\stack[2][10] ), .Z(n16938) );
  NAND U17549 ( .A(n16939), .B(n16938), .Z(n2554) );
  NAND U17550 ( .A(n17311), .B(o[10]), .Z(n16941) );
  NAND U17551 ( .A(n17305), .B(\stack[2][10] ), .Z(n16940) );
  AND U17552 ( .A(n16941), .B(n16940), .Z(n16943) );
  NAND U17553 ( .A(\stack[1][10] ), .B(n17308), .Z(n16942) );
  NAND U17554 ( .A(n16943), .B(n16942), .Z(n2555) );
  NAND U17555 ( .A(n17313), .B(o[10]), .Z(n16944) );
  NANDN U17556 ( .A(n17318), .B(n16944), .Z(n16945) );
  AND U17557 ( .A(\stack[1][10] ), .B(n16945), .Z(n16953) );
  NAND U17558 ( .A(x[10]), .B(n17311), .Z(n16946) );
  XNOR U17559 ( .A(n16948), .B(n16947), .Z(n16949) );
  NANDN U17560 ( .A(n17294), .B(n16949), .Z(n16950) );
  NAND U17561 ( .A(n16951), .B(n16950), .Z(n16952) );
  NOR U17562 ( .A(n16953), .B(n16952), .Z(n16955) );
  NANDN U17563 ( .A(n17317), .B(o[10]), .Z(n16954) );
  NAND U17564 ( .A(n16955), .B(n16954), .Z(n2556) );
  NAND U17565 ( .A(\stack[6][9] ), .B(n17311), .Z(n16957) );
  NANDN U17566 ( .A(n17311), .B(\stack[7][9] ), .Z(n16956) );
  NAND U17567 ( .A(n16957), .B(n16956), .Z(n2557) );
  NAND U17568 ( .A(\stack[5][9] ), .B(n17311), .Z(n16959) );
  NAND U17569 ( .A(n17305), .B(\stack[7][9] ), .Z(n16958) );
  AND U17570 ( .A(n16959), .B(n16958), .Z(n16961) );
  NAND U17571 ( .A(n17308), .B(\stack[6][9] ), .Z(n16960) );
  NAND U17572 ( .A(n16961), .B(n16960), .Z(n2558) );
  NAND U17573 ( .A(\stack[4][9] ), .B(n17311), .Z(n16963) );
  NAND U17574 ( .A(n17305), .B(\stack[6][9] ), .Z(n16962) );
  AND U17575 ( .A(n16963), .B(n16962), .Z(n16965) );
  NAND U17576 ( .A(n17308), .B(\stack[5][9] ), .Z(n16964) );
  NAND U17577 ( .A(n16965), .B(n16964), .Z(n2559) );
  NAND U17578 ( .A(\stack[3][9] ), .B(n17311), .Z(n16967) );
  NAND U17579 ( .A(n17305), .B(\stack[5][9] ), .Z(n16966) );
  AND U17580 ( .A(n16967), .B(n16966), .Z(n16969) );
  NAND U17581 ( .A(n17308), .B(\stack[4][9] ), .Z(n16968) );
  NAND U17582 ( .A(n16969), .B(n16968), .Z(n2560) );
  NAND U17583 ( .A(\stack[2][9] ), .B(n17311), .Z(n16971) );
  NAND U17584 ( .A(n17305), .B(\stack[4][9] ), .Z(n16970) );
  AND U17585 ( .A(n16971), .B(n16970), .Z(n16973) );
  NAND U17586 ( .A(n17308), .B(\stack[3][9] ), .Z(n16972) );
  NAND U17587 ( .A(n16973), .B(n16972), .Z(n2561) );
  NAND U17588 ( .A(n17311), .B(\stack[1][9] ), .Z(n16975) );
  NAND U17589 ( .A(n17305), .B(\stack[3][9] ), .Z(n16974) );
  AND U17590 ( .A(n16975), .B(n16974), .Z(n16977) );
  NAND U17591 ( .A(n17308), .B(\stack[2][9] ), .Z(n16976) );
  NAND U17592 ( .A(n16977), .B(n16976), .Z(n2562) );
  NAND U17593 ( .A(n17311), .B(o[9]), .Z(n16979) );
  NAND U17594 ( .A(n17305), .B(\stack[2][9] ), .Z(n16978) );
  AND U17595 ( .A(n16979), .B(n16978), .Z(n16981) );
  NAND U17596 ( .A(\stack[1][9] ), .B(n17308), .Z(n16980) );
  NAND U17597 ( .A(n16981), .B(n16980), .Z(n2563) );
  NAND U17598 ( .A(n17313), .B(o[9]), .Z(n16982) );
  NANDN U17599 ( .A(n17318), .B(n16982), .Z(n16983) );
  AND U17600 ( .A(\stack[1][9] ), .B(n16983), .Z(n16991) );
  NAND U17601 ( .A(x[9]), .B(n17311), .Z(n16984) );
  XNOR U17602 ( .A(n16986), .B(n16985), .Z(n16987) );
  NANDN U17603 ( .A(n17294), .B(n16987), .Z(n16988) );
  NAND U17604 ( .A(n16989), .B(n16988), .Z(n16990) );
  NOR U17605 ( .A(n16991), .B(n16990), .Z(n16993) );
  NANDN U17606 ( .A(n17317), .B(o[9]), .Z(n16992) );
  NAND U17607 ( .A(n16993), .B(n16992), .Z(n2564) );
  NAND U17608 ( .A(\stack[6][8] ), .B(n17311), .Z(n16995) );
  NANDN U17609 ( .A(n17311), .B(\stack[7][8] ), .Z(n16994) );
  NAND U17610 ( .A(n16995), .B(n16994), .Z(n2565) );
  NAND U17611 ( .A(\stack[5][8] ), .B(n17311), .Z(n16997) );
  NAND U17612 ( .A(n17305), .B(\stack[7][8] ), .Z(n16996) );
  AND U17613 ( .A(n16997), .B(n16996), .Z(n16999) );
  NAND U17614 ( .A(n17308), .B(\stack[6][8] ), .Z(n16998) );
  NAND U17615 ( .A(n16999), .B(n16998), .Z(n2566) );
  NAND U17616 ( .A(\stack[4][8] ), .B(n17311), .Z(n17001) );
  NAND U17617 ( .A(n17305), .B(\stack[6][8] ), .Z(n17000) );
  AND U17618 ( .A(n17001), .B(n17000), .Z(n17003) );
  NAND U17619 ( .A(n17308), .B(\stack[5][8] ), .Z(n17002) );
  NAND U17620 ( .A(n17003), .B(n17002), .Z(n2567) );
  NAND U17621 ( .A(\stack[3][8] ), .B(n17311), .Z(n17005) );
  NAND U17622 ( .A(n17305), .B(\stack[5][8] ), .Z(n17004) );
  AND U17623 ( .A(n17005), .B(n17004), .Z(n17007) );
  NAND U17624 ( .A(n17308), .B(\stack[4][8] ), .Z(n17006) );
  NAND U17625 ( .A(n17007), .B(n17006), .Z(n2568) );
  NAND U17626 ( .A(\stack[2][8] ), .B(n17311), .Z(n17009) );
  NAND U17627 ( .A(n17305), .B(\stack[4][8] ), .Z(n17008) );
  AND U17628 ( .A(n17009), .B(n17008), .Z(n17011) );
  NAND U17629 ( .A(n17308), .B(\stack[3][8] ), .Z(n17010) );
  NAND U17630 ( .A(n17011), .B(n17010), .Z(n2569) );
  NAND U17631 ( .A(n17311), .B(\stack[1][8] ), .Z(n17013) );
  NAND U17632 ( .A(n17305), .B(\stack[3][8] ), .Z(n17012) );
  AND U17633 ( .A(n17013), .B(n17012), .Z(n17015) );
  NAND U17634 ( .A(n17308), .B(\stack[2][8] ), .Z(n17014) );
  NAND U17635 ( .A(n17015), .B(n17014), .Z(n2570) );
  NAND U17636 ( .A(n17311), .B(o[8]), .Z(n17017) );
  NAND U17637 ( .A(n17305), .B(\stack[2][8] ), .Z(n17016) );
  AND U17638 ( .A(n17017), .B(n17016), .Z(n17019) );
  NAND U17639 ( .A(\stack[1][8] ), .B(n17308), .Z(n17018) );
  NAND U17640 ( .A(n17019), .B(n17018), .Z(n2571) );
  NAND U17641 ( .A(x[8]), .B(n17311), .Z(n17022) );
  NAND U17642 ( .A(n17020), .B(n17313), .Z(n17021) );
  NAND U17643 ( .A(n17022), .B(n17021), .Z(n17030) );
  NAND U17644 ( .A(n17318), .B(\stack[1][8] ), .Z(n17023) );
  XNOR U17645 ( .A(n17025), .B(n17024), .Z(n17026) );
  NANDN U17646 ( .A(n17294), .B(n17026), .Z(n17027) );
  NAND U17647 ( .A(n17028), .B(n17027), .Z(n17029) );
  NOR U17648 ( .A(n17030), .B(n17029), .Z(n17032) );
  NANDN U17649 ( .A(n17317), .B(o[8]), .Z(n17031) );
  NAND U17650 ( .A(n17032), .B(n17031), .Z(n2572) );
  NAND U17651 ( .A(\stack[6][7] ), .B(n17311), .Z(n17034) );
  NANDN U17652 ( .A(n17311), .B(\stack[7][7] ), .Z(n17033) );
  NAND U17653 ( .A(n17034), .B(n17033), .Z(n2573) );
  NAND U17654 ( .A(\stack[5][7] ), .B(n17311), .Z(n17036) );
  NAND U17655 ( .A(n17305), .B(\stack[7][7] ), .Z(n17035) );
  AND U17656 ( .A(n17036), .B(n17035), .Z(n17038) );
  NAND U17657 ( .A(n17308), .B(\stack[6][7] ), .Z(n17037) );
  NAND U17658 ( .A(n17038), .B(n17037), .Z(n2574) );
  NAND U17659 ( .A(\stack[4][7] ), .B(n17311), .Z(n17040) );
  NAND U17660 ( .A(n17305), .B(\stack[6][7] ), .Z(n17039) );
  AND U17661 ( .A(n17040), .B(n17039), .Z(n17042) );
  NAND U17662 ( .A(n17308), .B(\stack[5][7] ), .Z(n17041) );
  NAND U17663 ( .A(n17042), .B(n17041), .Z(n2575) );
  NAND U17664 ( .A(\stack[3][7] ), .B(n17311), .Z(n17044) );
  NAND U17665 ( .A(n17305), .B(\stack[5][7] ), .Z(n17043) );
  AND U17666 ( .A(n17044), .B(n17043), .Z(n17046) );
  NAND U17667 ( .A(n17308), .B(\stack[4][7] ), .Z(n17045) );
  NAND U17668 ( .A(n17046), .B(n17045), .Z(n2576) );
  NAND U17669 ( .A(\stack[2][7] ), .B(n17311), .Z(n17048) );
  NAND U17670 ( .A(n17305), .B(\stack[4][7] ), .Z(n17047) );
  AND U17671 ( .A(n17048), .B(n17047), .Z(n17050) );
  NAND U17672 ( .A(n17308), .B(\stack[3][7] ), .Z(n17049) );
  NAND U17673 ( .A(n17050), .B(n17049), .Z(n2577) );
  NAND U17674 ( .A(n17311), .B(\stack[1][7] ), .Z(n17052) );
  NAND U17675 ( .A(n17305), .B(\stack[3][7] ), .Z(n17051) );
  AND U17676 ( .A(n17052), .B(n17051), .Z(n17054) );
  NAND U17677 ( .A(n17308), .B(\stack[2][7] ), .Z(n17053) );
  NAND U17678 ( .A(n17054), .B(n17053), .Z(n2578) );
  NAND U17679 ( .A(n17311), .B(o[7]), .Z(n17056) );
  NAND U17680 ( .A(n17305), .B(\stack[2][7] ), .Z(n17055) );
  AND U17681 ( .A(n17056), .B(n17055), .Z(n17058) );
  NAND U17682 ( .A(\stack[1][7] ), .B(n17308), .Z(n17057) );
  NAND U17683 ( .A(n17058), .B(n17057), .Z(n2579) );
  NAND U17684 ( .A(n17313), .B(o[7]), .Z(n17059) );
  NANDN U17685 ( .A(n17318), .B(n17059), .Z(n17060) );
  AND U17686 ( .A(\stack[1][7] ), .B(n17060), .Z(n17068) );
  NAND U17687 ( .A(x[7]), .B(n17311), .Z(n17061) );
  XNOR U17688 ( .A(n17063), .B(n17062), .Z(n17064) );
  NANDN U17689 ( .A(n17294), .B(n17064), .Z(n17065) );
  NAND U17690 ( .A(n17066), .B(n17065), .Z(n17067) );
  NOR U17691 ( .A(n17068), .B(n17067), .Z(n17070) );
  NANDN U17692 ( .A(n17317), .B(o[7]), .Z(n17069) );
  NAND U17693 ( .A(n17070), .B(n17069), .Z(n2580) );
  NAND U17694 ( .A(\stack[6][6] ), .B(n17311), .Z(n17072) );
  NANDN U17695 ( .A(n17311), .B(\stack[7][6] ), .Z(n17071) );
  NAND U17696 ( .A(n17072), .B(n17071), .Z(n2581) );
  NAND U17697 ( .A(\stack[5][6] ), .B(n17311), .Z(n17074) );
  NAND U17698 ( .A(n17305), .B(\stack[7][6] ), .Z(n17073) );
  AND U17699 ( .A(n17074), .B(n17073), .Z(n17076) );
  NAND U17700 ( .A(n17308), .B(\stack[6][6] ), .Z(n17075) );
  NAND U17701 ( .A(n17076), .B(n17075), .Z(n2582) );
  NAND U17702 ( .A(\stack[4][6] ), .B(n17311), .Z(n17078) );
  NAND U17703 ( .A(n17305), .B(\stack[6][6] ), .Z(n17077) );
  AND U17704 ( .A(n17078), .B(n17077), .Z(n17080) );
  NAND U17705 ( .A(n17308), .B(\stack[5][6] ), .Z(n17079) );
  NAND U17706 ( .A(n17080), .B(n17079), .Z(n2583) );
  NAND U17707 ( .A(\stack[3][6] ), .B(n17311), .Z(n17082) );
  NAND U17708 ( .A(n17305), .B(\stack[5][6] ), .Z(n17081) );
  AND U17709 ( .A(n17082), .B(n17081), .Z(n17084) );
  NAND U17710 ( .A(n17308), .B(\stack[4][6] ), .Z(n17083) );
  NAND U17711 ( .A(n17084), .B(n17083), .Z(n2584) );
  NAND U17712 ( .A(\stack[2][6] ), .B(n17311), .Z(n17086) );
  NAND U17713 ( .A(n17305), .B(\stack[4][6] ), .Z(n17085) );
  AND U17714 ( .A(n17086), .B(n17085), .Z(n17088) );
  NAND U17715 ( .A(n17308), .B(\stack[3][6] ), .Z(n17087) );
  NAND U17716 ( .A(n17088), .B(n17087), .Z(n2585) );
  NAND U17717 ( .A(n17311), .B(\stack[1][6] ), .Z(n17090) );
  NAND U17718 ( .A(n17305), .B(\stack[3][6] ), .Z(n17089) );
  AND U17719 ( .A(n17090), .B(n17089), .Z(n17092) );
  NAND U17720 ( .A(n17308), .B(\stack[2][6] ), .Z(n17091) );
  NAND U17721 ( .A(n17092), .B(n17091), .Z(n2586) );
  NAND U17722 ( .A(n17311), .B(o[6]), .Z(n17094) );
  NAND U17723 ( .A(n17305), .B(\stack[2][6] ), .Z(n17093) );
  AND U17724 ( .A(n17094), .B(n17093), .Z(n17096) );
  NAND U17725 ( .A(\stack[1][6] ), .B(n17308), .Z(n17095) );
  NAND U17726 ( .A(n17096), .B(n17095), .Z(n2587) );
  NAND U17727 ( .A(x[6]), .B(n17311), .Z(n17099) );
  NAND U17728 ( .A(n17097), .B(n17313), .Z(n17098) );
  NAND U17729 ( .A(n17099), .B(n17098), .Z(n17107) );
  NAND U17730 ( .A(n17318), .B(\stack[1][6] ), .Z(n17100) );
  XNOR U17731 ( .A(n17102), .B(n17101), .Z(n17103) );
  NANDN U17732 ( .A(n17294), .B(n17103), .Z(n17104) );
  NAND U17733 ( .A(n17105), .B(n17104), .Z(n17106) );
  NOR U17734 ( .A(n17107), .B(n17106), .Z(n17109) );
  NANDN U17735 ( .A(n17317), .B(o[6]), .Z(n17108) );
  NAND U17736 ( .A(n17109), .B(n17108), .Z(n2588) );
  NAND U17737 ( .A(\stack[6][5] ), .B(n17311), .Z(n17111) );
  NANDN U17738 ( .A(n17311), .B(\stack[7][5] ), .Z(n17110) );
  NAND U17739 ( .A(n17111), .B(n17110), .Z(n2589) );
  NAND U17740 ( .A(\stack[5][5] ), .B(n17311), .Z(n17113) );
  NAND U17741 ( .A(n17305), .B(\stack[7][5] ), .Z(n17112) );
  AND U17742 ( .A(n17113), .B(n17112), .Z(n17115) );
  NAND U17743 ( .A(n17308), .B(\stack[6][5] ), .Z(n17114) );
  NAND U17744 ( .A(n17115), .B(n17114), .Z(n2590) );
  NAND U17745 ( .A(\stack[4][5] ), .B(n17311), .Z(n17117) );
  NAND U17746 ( .A(n17305), .B(\stack[6][5] ), .Z(n17116) );
  AND U17747 ( .A(n17117), .B(n17116), .Z(n17119) );
  NAND U17748 ( .A(n17308), .B(\stack[5][5] ), .Z(n17118) );
  NAND U17749 ( .A(n17119), .B(n17118), .Z(n2591) );
  NAND U17750 ( .A(\stack[3][5] ), .B(n17311), .Z(n17121) );
  NAND U17751 ( .A(n17305), .B(\stack[5][5] ), .Z(n17120) );
  AND U17752 ( .A(n17121), .B(n17120), .Z(n17123) );
  NAND U17753 ( .A(n17308), .B(\stack[4][5] ), .Z(n17122) );
  NAND U17754 ( .A(n17123), .B(n17122), .Z(n2592) );
  NAND U17755 ( .A(\stack[2][5] ), .B(n17311), .Z(n17125) );
  NAND U17756 ( .A(n17305), .B(\stack[4][5] ), .Z(n17124) );
  AND U17757 ( .A(n17125), .B(n17124), .Z(n17127) );
  NAND U17758 ( .A(n17308), .B(\stack[3][5] ), .Z(n17126) );
  NAND U17759 ( .A(n17127), .B(n17126), .Z(n2593) );
  NAND U17760 ( .A(n17311), .B(\stack[1][5] ), .Z(n17129) );
  NAND U17761 ( .A(n17305), .B(\stack[3][5] ), .Z(n17128) );
  AND U17762 ( .A(n17129), .B(n17128), .Z(n17131) );
  NAND U17763 ( .A(n17308), .B(\stack[2][5] ), .Z(n17130) );
  NAND U17764 ( .A(n17131), .B(n17130), .Z(n2594) );
  NAND U17765 ( .A(n17311), .B(o[5]), .Z(n17133) );
  NAND U17766 ( .A(n17305), .B(\stack[2][5] ), .Z(n17132) );
  AND U17767 ( .A(n17133), .B(n17132), .Z(n17135) );
  NAND U17768 ( .A(\stack[1][5] ), .B(n17308), .Z(n17134) );
  NAND U17769 ( .A(n17135), .B(n17134), .Z(n2595) );
  NAND U17770 ( .A(x[5]), .B(n17311), .Z(n17138) );
  NAND U17771 ( .A(n17136), .B(n17313), .Z(n17137) );
  NAND U17772 ( .A(n17138), .B(n17137), .Z(n17146) );
  NAND U17773 ( .A(n17318), .B(\stack[1][5] ), .Z(n17139) );
  XNOR U17774 ( .A(n17141), .B(n17140), .Z(n17142) );
  NANDN U17775 ( .A(n17294), .B(n17142), .Z(n17143) );
  NAND U17776 ( .A(n17144), .B(n17143), .Z(n17145) );
  NOR U17777 ( .A(n17146), .B(n17145), .Z(n17148) );
  NANDN U17778 ( .A(n17317), .B(o[5]), .Z(n17147) );
  NAND U17779 ( .A(n17148), .B(n17147), .Z(n2596) );
  NAND U17780 ( .A(\stack[6][4] ), .B(n17311), .Z(n17150) );
  NANDN U17781 ( .A(n17311), .B(\stack[7][4] ), .Z(n17149) );
  NAND U17782 ( .A(n17150), .B(n17149), .Z(n2597) );
  NAND U17783 ( .A(\stack[5][4] ), .B(n17311), .Z(n17152) );
  NAND U17784 ( .A(n17305), .B(\stack[7][4] ), .Z(n17151) );
  AND U17785 ( .A(n17152), .B(n17151), .Z(n17154) );
  NAND U17786 ( .A(n17308), .B(\stack[6][4] ), .Z(n17153) );
  NAND U17787 ( .A(n17154), .B(n17153), .Z(n2598) );
  NAND U17788 ( .A(\stack[4][4] ), .B(n17311), .Z(n17156) );
  NAND U17789 ( .A(n17305), .B(\stack[6][4] ), .Z(n17155) );
  AND U17790 ( .A(n17156), .B(n17155), .Z(n17158) );
  NAND U17791 ( .A(n17308), .B(\stack[5][4] ), .Z(n17157) );
  NAND U17792 ( .A(n17158), .B(n17157), .Z(n2599) );
  NAND U17793 ( .A(\stack[3][4] ), .B(n17311), .Z(n17160) );
  NAND U17794 ( .A(n17305), .B(\stack[5][4] ), .Z(n17159) );
  AND U17795 ( .A(n17160), .B(n17159), .Z(n17162) );
  NAND U17796 ( .A(n17308), .B(\stack[4][4] ), .Z(n17161) );
  NAND U17797 ( .A(n17162), .B(n17161), .Z(n2600) );
  NAND U17798 ( .A(\stack[2][4] ), .B(n17311), .Z(n17164) );
  NAND U17799 ( .A(n17305), .B(\stack[4][4] ), .Z(n17163) );
  AND U17800 ( .A(n17164), .B(n17163), .Z(n17166) );
  NAND U17801 ( .A(n17308), .B(\stack[3][4] ), .Z(n17165) );
  NAND U17802 ( .A(n17166), .B(n17165), .Z(n2601) );
  NAND U17803 ( .A(n17311), .B(\stack[1][4] ), .Z(n17168) );
  NAND U17804 ( .A(n17305), .B(\stack[3][4] ), .Z(n17167) );
  AND U17805 ( .A(n17168), .B(n17167), .Z(n17170) );
  NAND U17806 ( .A(n17308), .B(\stack[2][4] ), .Z(n17169) );
  NAND U17807 ( .A(n17170), .B(n17169), .Z(n2602) );
  NAND U17808 ( .A(n17311), .B(o[4]), .Z(n17172) );
  NAND U17809 ( .A(n17305), .B(\stack[2][4] ), .Z(n17171) );
  AND U17810 ( .A(n17172), .B(n17171), .Z(n17174) );
  NAND U17811 ( .A(\stack[1][4] ), .B(n17308), .Z(n17173) );
  NAND U17812 ( .A(n17174), .B(n17173), .Z(n2603) );
  NAND U17813 ( .A(x[4]), .B(n17311), .Z(n17177) );
  NAND U17814 ( .A(n17175), .B(n17313), .Z(n17176) );
  NAND U17815 ( .A(n17177), .B(n17176), .Z(n17185) );
  NAND U17816 ( .A(n17318), .B(\stack[1][4] ), .Z(n17178) );
  XNOR U17817 ( .A(n17180), .B(n17179), .Z(n17181) );
  NANDN U17818 ( .A(n17294), .B(n17181), .Z(n17182) );
  NAND U17819 ( .A(n17183), .B(n17182), .Z(n17184) );
  NOR U17820 ( .A(n17185), .B(n17184), .Z(n17187) );
  NANDN U17821 ( .A(n17317), .B(o[4]), .Z(n17186) );
  NAND U17822 ( .A(n17187), .B(n17186), .Z(n2604) );
  NAND U17823 ( .A(\stack[6][3] ), .B(n17311), .Z(n17189) );
  NANDN U17824 ( .A(n17311), .B(\stack[7][3] ), .Z(n17188) );
  NAND U17825 ( .A(n17189), .B(n17188), .Z(n2605) );
  NAND U17826 ( .A(\stack[5][3] ), .B(n17311), .Z(n17191) );
  NAND U17827 ( .A(n17305), .B(\stack[7][3] ), .Z(n17190) );
  AND U17828 ( .A(n17191), .B(n17190), .Z(n17193) );
  NAND U17829 ( .A(n17308), .B(\stack[6][3] ), .Z(n17192) );
  NAND U17830 ( .A(n17193), .B(n17192), .Z(n2606) );
  NAND U17831 ( .A(\stack[4][3] ), .B(n17311), .Z(n17195) );
  NAND U17832 ( .A(n17305), .B(\stack[6][3] ), .Z(n17194) );
  AND U17833 ( .A(n17195), .B(n17194), .Z(n17197) );
  NAND U17834 ( .A(n17308), .B(\stack[5][3] ), .Z(n17196) );
  NAND U17835 ( .A(n17197), .B(n17196), .Z(n2607) );
  NAND U17836 ( .A(\stack[3][3] ), .B(n17311), .Z(n17199) );
  NAND U17837 ( .A(n17305), .B(\stack[5][3] ), .Z(n17198) );
  AND U17838 ( .A(n17199), .B(n17198), .Z(n17201) );
  NAND U17839 ( .A(n17308), .B(\stack[4][3] ), .Z(n17200) );
  NAND U17840 ( .A(n17201), .B(n17200), .Z(n2608) );
  NAND U17841 ( .A(\stack[2][3] ), .B(n17311), .Z(n17203) );
  NAND U17842 ( .A(n17305), .B(\stack[4][3] ), .Z(n17202) );
  AND U17843 ( .A(n17203), .B(n17202), .Z(n17205) );
  NAND U17844 ( .A(n17308), .B(\stack[3][3] ), .Z(n17204) );
  NAND U17845 ( .A(n17205), .B(n17204), .Z(n2609) );
  NAND U17846 ( .A(n17311), .B(\stack[1][3] ), .Z(n17207) );
  NAND U17847 ( .A(n17305), .B(\stack[3][3] ), .Z(n17206) );
  AND U17848 ( .A(n17207), .B(n17206), .Z(n17209) );
  NAND U17849 ( .A(n17308), .B(\stack[2][3] ), .Z(n17208) );
  NAND U17850 ( .A(n17209), .B(n17208), .Z(n2610) );
  NAND U17851 ( .A(n17311), .B(o[3]), .Z(n17211) );
  NAND U17852 ( .A(n17305), .B(\stack[2][3] ), .Z(n17210) );
  AND U17853 ( .A(n17211), .B(n17210), .Z(n17213) );
  NAND U17854 ( .A(\stack[1][3] ), .B(n17308), .Z(n17212) );
  NAND U17855 ( .A(n17213), .B(n17212), .Z(n2611) );
  NAND U17856 ( .A(x[3]), .B(n17311), .Z(n17216) );
  NAND U17857 ( .A(n17214), .B(n17313), .Z(n17215) );
  NAND U17858 ( .A(n17216), .B(n17215), .Z(n17224) );
  NAND U17859 ( .A(n17318), .B(\stack[1][3] ), .Z(n17217) );
  XNOR U17860 ( .A(n17219), .B(n17218), .Z(n17220) );
  NANDN U17861 ( .A(n17294), .B(n17220), .Z(n17221) );
  NAND U17862 ( .A(n17222), .B(n17221), .Z(n17223) );
  NOR U17863 ( .A(n17224), .B(n17223), .Z(n17226) );
  NANDN U17864 ( .A(n17317), .B(o[3]), .Z(n17225) );
  NAND U17865 ( .A(n17226), .B(n17225), .Z(n2612) );
  NAND U17866 ( .A(\stack[6][2] ), .B(n17311), .Z(n17228) );
  NANDN U17867 ( .A(n17311), .B(\stack[7][2] ), .Z(n17227) );
  NAND U17868 ( .A(n17228), .B(n17227), .Z(n2613) );
  NAND U17869 ( .A(\stack[5][2] ), .B(n17311), .Z(n17230) );
  NAND U17870 ( .A(n17305), .B(\stack[7][2] ), .Z(n17229) );
  AND U17871 ( .A(n17230), .B(n17229), .Z(n17232) );
  NAND U17872 ( .A(n17308), .B(\stack[6][2] ), .Z(n17231) );
  NAND U17873 ( .A(n17232), .B(n17231), .Z(n2614) );
  NAND U17874 ( .A(\stack[4][2] ), .B(n17311), .Z(n17234) );
  NAND U17875 ( .A(n17305), .B(\stack[6][2] ), .Z(n17233) );
  AND U17876 ( .A(n17234), .B(n17233), .Z(n17236) );
  NAND U17877 ( .A(n17308), .B(\stack[5][2] ), .Z(n17235) );
  NAND U17878 ( .A(n17236), .B(n17235), .Z(n2615) );
  NAND U17879 ( .A(\stack[3][2] ), .B(n17311), .Z(n17238) );
  NAND U17880 ( .A(n17305), .B(\stack[5][2] ), .Z(n17237) );
  AND U17881 ( .A(n17238), .B(n17237), .Z(n17240) );
  NAND U17882 ( .A(n17308), .B(\stack[4][2] ), .Z(n17239) );
  NAND U17883 ( .A(n17240), .B(n17239), .Z(n2616) );
  NAND U17884 ( .A(\stack[2][2] ), .B(n17311), .Z(n17242) );
  NAND U17885 ( .A(n17305), .B(\stack[4][2] ), .Z(n17241) );
  AND U17886 ( .A(n17242), .B(n17241), .Z(n17244) );
  NAND U17887 ( .A(n17308), .B(\stack[3][2] ), .Z(n17243) );
  NAND U17888 ( .A(n17244), .B(n17243), .Z(n2617) );
  NAND U17889 ( .A(n17311), .B(\stack[1][2] ), .Z(n17246) );
  NAND U17890 ( .A(n17305), .B(\stack[3][2] ), .Z(n17245) );
  AND U17891 ( .A(n17246), .B(n17245), .Z(n17248) );
  NAND U17892 ( .A(n17308), .B(\stack[2][2] ), .Z(n17247) );
  NAND U17893 ( .A(n17248), .B(n17247), .Z(n2618) );
  NAND U17894 ( .A(n17311), .B(o[2]), .Z(n17250) );
  NAND U17895 ( .A(n17305), .B(\stack[2][2] ), .Z(n17249) );
  AND U17896 ( .A(n17250), .B(n17249), .Z(n17252) );
  NAND U17897 ( .A(\stack[1][2] ), .B(n17308), .Z(n17251) );
  NAND U17898 ( .A(n17252), .B(n17251), .Z(n2619) );
  NAND U17899 ( .A(o[2]), .B(n17313), .Z(n17253) );
  NANDN U17900 ( .A(n17318), .B(n17253), .Z(n17254) );
  NAND U17901 ( .A(\stack[1][2] ), .B(n17254), .Z(n17257) );
  NAND U17902 ( .A(x[2]), .B(n17311), .Z(n17255) );
  AND U17903 ( .A(n17257), .B(n17256), .Z(n17259) );
  NANDN U17904 ( .A(n17317), .B(o[2]), .Z(n17258) );
  AND U17905 ( .A(n17259), .B(n17258), .Z(n17264) );
  XNOR U17906 ( .A(n17261), .B(n17260), .Z(n17262) );
  NANDN U17907 ( .A(n17294), .B(n17262), .Z(n17263) );
  NAND U17908 ( .A(n17264), .B(n17263), .Z(n2620) );
  NAND U17909 ( .A(\stack[6][1] ), .B(n17311), .Z(n17266) );
  NANDN U17910 ( .A(n17311), .B(\stack[7][1] ), .Z(n17265) );
  NAND U17911 ( .A(n17266), .B(n17265), .Z(n2621) );
  NAND U17912 ( .A(\stack[5][1] ), .B(n17311), .Z(n17268) );
  NAND U17913 ( .A(n17305), .B(\stack[7][1] ), .Z(n17267) );
  AND U17914 ( .A(n17268), .B(n17267), .Z(n17270) );
  NAND U17915 ( .A(n17308), .B(\stack[6][1] ), .Z(n17269) );
  NAND U17916 ( .A(n17270), .B(n17269), .Z(n2622) );
  NAND U17917 ( .A(\stack[4][1] ), .B(n17311), .Z(n17272) );
  NAND U17918 ( .A(n17305), .B(\stack[6][1] ), .Z(n17271) );
  AND U17919 ( .A(n17272), .B(n17271), .Z(n17274) );
  NAND U17920 ( .A(n17308), .B(\stack[5][1] ), .Z(n17273) );
  NAND U17921 ( .A(n17274), .B(n17273), .Z(n2623) );
  NAND U17922 ( .A(\stack[3][1] ), .B(n17311), .Z(n17276) );
  NAND U17923 ( .A(n17305), .B(\stack[5][1] ), .Z(n17275) );
  AND U17924 ( .A(n17276), .B(n17275), .Z(n17278) );
  NAND U17925 ( .A(n17308), .B(\stack[4][1] ), .Z(n17277) );
  NAND U17926 ( .A(n17278), .B(n17277), .Z(n2624) );
  NAND U17927 ( .A(\stack[2][1] ), .B(n17311), .Z(n17280) );
  NAND U17928 ( .A(n17305), .B(\stack[4][1] ), .Z(n17279) );
  AND U17929 ( .A(n17280), .B(n17279), .Z(n17282) );
  NAND U17930 ( .A(n17308), .B(\stack[3][1] ), .Z(n17281) );
  NAND U17931 ( .A(n17282), .B(n17281), .Z(n2625) );
  NAND U17932 ( .A(n17311), .B(\stack[1][1] ), .Z(n17284) );
  NAND U17933 ( .A(n17305), .B(\stack[3][1] ), .Z(n17283) );
  AND U17934 ( .A(n17284), .B(n17283), .Z(n17286) );
  NAND U17935 ( .A(n17308), .B(\stack[2][1] ), .Z(n17285) );
  NAND U17936 ( .A(n17286), .B(n17285), .Z(n2626) );
  NAND U17937 ( .A(n17311), .B(o[1]), .Z(n17288) );
  NAND U17938 ( .A(n17305), .B(\stack[2][1] ), .Z(n17287) );
  AND U17939 ( .A(n17288), .B(n17287), .Z(n17290) );
  NAND U17940 ( .A(\stack[1][1] ), .B(n17308), .Z(n17289) );
  NAND U17941 ( .A(n17290), .B(n17289), .Z(n2627) );
  XOR U17942 ( .A(n17292), .B(n17291), .Z(n17293) );
  NANDN U17943 ( .A(n17294), .B(n17293), .Z(n17299) );
  NAND U17944 ( .A(x[1]), .B(n17311), .Z(n17297) );
  NAND U17945 ( .A(o[1]), .B(\stack[1][1] ), .Z(n17295) );
  NANDN U17946 ( .A(n17295), .B(n17313), .Z(n17296) );
  AND U17947 ( .A(n17297), .B(n17296), .Z(n17298) );
  AND U17948 ( .A(n17299), .B(n17298), .Z(n17301) );
  NAND U17949 ( .A(\stack[1][1] ), .B(n17318), .Z(n17300) );
  AND U17950 ( .A(n17301), .B(n17300), .Z(n17304) );
  NANDN U17951 ( .A(n17317), .B(o[1]), .Z(n17302) );
  NAND U17952 ( .A(n17304), .B(n17303), .Z(n2628) );
  NAND U17953 ( .A(n17311), .B(o[0]), .Z(n17307) );
  NAND U17954 ( .A(n17305), .B(\stack[2][0] ), .Z(n17306) );
  AND U17955 ( .A(n17307), .B(n17306), .Z(n17310) );
  NAND U17956 ( .A(\stack[1][0] ), .B(n17308), .Z(n17309) );
  NAND U17957 ( .A(n17310), .B(n17309), .Z(n2629) );
  NAND U17958 ( .A(x[0]), .B(n17311), .Z(n17312) );
  OR U17959 ( .A(n17314), .B(n17313), .Z(n17315) );
  NAND U17960 ( .A(\stack[1][0] ), .B(n17315), .Z(n17316) );
  AND U17961 ( .A(n17317), .B(n17316), .Z(n17321) );
  NAND U17962 ( .A(\stack[1][0] ), .B(n17318), .Z(n17319) );
  NANDN U17963 ( .A(o[0]), .B(n17319), .Z(n17320) );
  NANDN U17964 ( .A(n17321), .B(n17320), .Z(n17322) );
  NAND U17965 ( .A(n17323), .B(n17322), .Z(n2630) );
endmodule

