
module first_nns_comb_W7_N512 ( q, DB, min_val_out );
  input [6:0] q;
  input [3583:0] DB;
  output [6:0] min_val_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001,
         n10002, n10003, n10004, n10005, n10006, n10007, n10008, n10009,
         n10010, n10011, n10012, n10013, n10014, n10015, n10016, n10017,
         n10018, n10019, n10020, n10021, n10022, n10023, n10024, n10025,
         n10026, n10027, n10028, n10029, n10030, n10031, n10032, n10033,
         n10034, n10035, n10036, n10037, n10038, n10039, n10040, n10041,
         n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049,
         n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057,
         n10058, n10059, n10060, n10061, n10062, n10063, n10064, n10065,
         n10066, n10067, n10068, n10069, n10070, n10071, n10072, n10073,
         n10074, n10075, n10076, n10077, n10078, n10079, n10080, n10081,
         n10082, n10083, n10084, n10085, n10086, n10087, n10088, n10089,
         n10090, n10091, n10092, n10093, n10094, n10095, n10096, n10097,
         n10098, n10099, n10100, n10101, n10102, n10103, n10104, n10105,
         n10106, n10107, n10108, n10109, n10110, n10111, n10112, n10113,
         n10114, n10115, n10116, n10117, n10118, n10119, n10120, n10121,
         n10122, n10123, n10124, n10125, n10126, n10127, n10128, n10129,
         n10130, n10131, n10132, n10133, n10134, n10135, n10136, n10137,
         n10138, n10139, n10140, n10141, n10142, n10143, n10144, n10145,
         n10146, n10147, n10148, n10149, n10150, n10151, n10152, n10153,
         n10154, n10155, n10156, n10157, n10158, n10159, n10160, n10161,
         n10162, n10163, n10164, n10165, n10166, n10167, n10168, n10169,
         n10170, n10171, n10172, n10173, n10174, n10175, n10176, n10177,
         n10178, n10179, n10180, n10181, n10182, n10183, n10184, n10185,
         n10186, n10187, n10188, n10189, n10190, n10191, n10192, n10193,
         n10194, n10195, n10196, n10197, n10198, n10199, n10200, n10201,
         n10202, n10203, n10204, n10205, n10206, n10207, n10208, n10209,
         n10210, n10211, n10212, n10213, n10214, n10215, n10216, n10217,
         n10218, n10219, n10220, n10221, n10222, n10223, n10224, n10225,
         n10226, n10227, n10228, n10229, n10230, n10231, n10232, n10233,
         n10234, n10235, n10236, n10237, n10238, n10239, n10240, n10241,
         n10242, n10243, n10244, n10245, n10246, n10247, n10248, n10249,
         n10250, n10251, n10252, n10253, n10254, n10255, n10256, n10257,
         n10258, n10259, n10260, n10261, n10262, n10263, n10264, n10265,
         n10266, n10267, n10268, n10269, n10270, n10271, n10272, n10273,
         n10274, n10275, n10276, n10277, n10278, n10279, n10280, n10281,
         n10282, n10283, n10284, n10285, n10286, n10287, n10288, n10289,
         n10290, n10291, n10292, n10293, n10294, n10295, n10296, n10297,
         n10298, n10299, n10300, n10301, n10302, n10303, n10304, n10305,
         n10306, n10307, n10308, n10309, n10310, n10311, n10312, n10313,
         n10314, n10315, n10316, n10317, n10318, n10319, n10320, n10321,
         n10322, n10323, n10324, n10325, n10326, n10327, n10328, n10329,
         n10330, n10331, n10332, n10333, n10334, n10335, n10336, n10337,
         n10338, n10339, n10340, n10341, n10342, n10343, n10344, n10345,
         n10346, n10347, n10348, n10349, n10350, n10351, n10352, n10353,
         n10354, n10355, n10356, n10357, n10358, n10359, n10360, n10361,
         n10362, n10363, n10364, n10365, n10366, n10367, n10368, n10369,
         n10370, n10371, n10372, n10373, n10374, n10375, n10376, n10377,
         n10378, n10379, n10380, n10381, n10382, n10383, n10384, n10385,
         n10386, n10387, n10388, n10389, n10390, n10391, n10392, n10393,
         n10394, n10395, n10396, n10397, n10398, n10399, n10400, n10401,
         n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409,
         n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417,
         n10418, n10419, n10420, n10421, n10422, n10423, n10424, n10425,
         n10426, n10427, n10428, n10429, n10430, n10431, n10432, n10433,
         n10434, n10435, n10436, n10437, n10438, n10439, n10440, n10441,
         n10442, n10443, n10444, n10445, n10446, n10447, n10448, n10449,
         n10450, n10451, n10452, n10453, n10454, n10455, n10456, n10457,
         n10458, n10459, n10460, n10461, n10462, n10463, n10464, n10465,
         n10466, n10467, n10468, n10469, n10470, n10471, n10472, n10473,
         n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481,
         n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489,
         n10490, n10491, n10492, n10493, n10494, n10495, n10496, n10497,
         n10498, n10499, n10500, n10501, n10502, n10503, n10504, n10505,
         n10506, n10507, n10508, n10509, n10510, n10511, n10512, n10513,
         n10514, n10515, n10516, n10517, n10518, n10519, n10520, n10521,
         n10522, n10523, n10524, n10525, n10526, n10527, n10528, n10529,
         n10530, n10531, n10532, n10533, n10534, n10535, n10536, n10537,
         n10538, n10539, n10540, n10541, n10542, n10543, n10544, n10545,
         n10546, n10547, n10548, n10549, n10550, n10551, n10552, n10553,
         n10554, n10555, n10556, n10557, n10558, n10559, n10560, n10561,
         n10562, n10563, n10564, n10565, n10566, n10567, n10568, n10569,
         n10570, n10571, n10572, n10573, n10574, n10575, n10576, n10577,
         n10578, n10579, n10580, n10581, n10582, n10583, n10584, n10585,
         n10586, n10587, n10588, n10589, n10590, n10591, n10592, n10593,
         n10594, n10595, n10596, n10597, n10598, n10599, n10600, n10601,
         n10602, n10603, n10604, n10605, n10606, n10607, n10608, n10609,
         n10610, n10611, n10612, n10613, n10614, n10615, n10616, n10617,
         n10618, n10619, n10620, n10621, n10622, n10623, n10624, n10625,
         n10626, n10627, n10628, n10629, n10630, n10631, n10632, n10633,
         n10634, n10635, n10636, n10637, n10638, n10639, n10640, n10641,
         n10642, n10643, n10644, n10645, n10646, n10647, n10648, n10649,
         n10650, n10651, n10652, n10653, n10654, n10655, n10656, n10657,
         n10658, n10659, n10660, n10661, n10662, n10663, n10664, n10665,
         n10666, n10667, n10668, n10669, n10670, n10671, n10672, n10673,
         n10674, n10675, n10676, n10677, n10678, n10679, n10680, n10681,
         n10682, n10683, n10684, n10685, n10686, n10687, n10688, n10689,
         n10690, n10691, n10692, n10693, n10694, n10695, n10696, n10697,
         n10698, n10699, n10700, n10701, n10702, n10703, n10704, n10705,
         n10706, n10707, n10708, n10709, n10710, n10711, n10712, n10713,
         n10714, n10715, n10716, n10717, n10718, n10719, n10720, n10721,
         n10722, n10723, n10724, n10725, n10726, n10727, n10728, n10729,
         n10730, n10731, n10732, n10733, n10734, n10735, n10736, n10737,
         n10738, n10739, n10740, n10741, n10742, n10743, n10744, n10745,
         n10746, n10747, n10748, n10749, n10750, n10751, n10752, n10753,
         n10754, n10755, n10756, n10757, n10758, n10759, n10760, n10761,
         n10762, n10763, n10764, n10765, n10766, n10767, n10768, n10769,
         n10770, n10771, n10772, n10773, n10774, n10775, n10776, n10777,
         n10778, n10779, n10780, n10781, n10782, n10783, n10784, n10785,
         n10786, n10787, n10788, n10789, n10790, n10791, n10792, n10793,
         n10794, n10795, n10796, n10797, n10798, n10799, n10800, n10801,
         n10802, n10803, n10804, n10805, n10806, n10807, n10808, n10809,
         n10810, n10811, n10812, n10813, n10814, n10815, n10816, n10817,
         n10818, n10819, n10820, n10821, n10822, n10823, n10824, n10825,
         n10826, n10827, n10828, n10829, n10830, n10831, n10832, n10833,
         n10834, n10835, n10836, n10837, n10838, n10839, n10840, n10841,
         n10842, n10843, n10844, n10845, n10846, n10847, n10848, n10849,
         n10850, n10851, n10852, n10853, n10854, n10855, n10856, n10857,
         n10858, n10859, n10860, n10861, n10862, n10863, n10864, n10865,
         n10866, n10867, n10868, n10869, n10870, n10871, n10872, n10873,
         n10874, n10875, n10876, n10877, n10878, n10879, n10880, n10881,
         n10882, n10883, n10884, n10885, n10886, n10887, n10888, n10889,
         n10890, n10891, n10892, n10893, n10894, n10895, n10896, n10897,
         n10898, n10899, n10900, n10901, n10902, n10903, n10904, n10905,
         n10906, n10907, n10908, n10909, n10910, n10911, n10912, n10913,
         n10914, n10915, n10916, n10917, n10918, n10919, n10920, n10921,
         n10922, n10923, n10924, n10925, n10926, n10927, n10928, n10929,
         n10930, n10931, n10932, n10933, n10934, n10935, n10936, n10937,
         n10938, n10939, n10940, n10941, n10942, n10943, n10944, n10945,
         n10946, n10947, n10948, n10949, n10950, n10951, n10952, n10953,
         n10954, n10955, n10956, n10957, n10958, n10959, n10960, n10961,
         n10962, n10963, n10964, n10965, n10966, n10967, n10968, n10969,
         n10970, n10971, n10972, n10973, n10974, n10975, n10976, n10977,
         n10978, n10979, n10980, n10981, n10982, n10983, n10984, n10985,
         n10986, n10987, n10988, n10989, n10990, n10991, n10992, n10993,
         n10994, n10995, n10996, n10997, n10998, n10999, n11000, n11001,
         n11002, n11003, n11004, n11005, n11006, n11007, n11008, n11009,
         n11010, n11011, n11012, n11013, n11014, n11015, n11016, n11017,
         n11018, n11019, n11020, n11021, n11022, n11023, n11024, n11025,
         n11026, n11027, n11028, n11029, n11030, n11031, n11032, n11033,
         n11034, n11035, n11036, n11037, n11038, n11039, n11040, n11041,
         n11042, n11043, n11044, n11045, n11046, n11047, n11048, n11049,
         n11050, n11051, n11052, n11053, n11054, n11055, n11056, n11057,
         n11058, n11059, n11060, n11061, n11062, n11063, n11064, n11065,
         n11066, n11067, n11068, n11069, n11070, n11071, n11072, n11073,
         n11074, n11075, n11076, n11077, n11078, n11079, n11080, n11081,
         n11082, n11083, n11084, n11085, n11086, n11087, n11088, n11089,
         n11090, n11091, n11092, n11093, n11094, n11095, n11096, n11097,
         n11098, n11099, n11100, n11101, n11102, n11103, n11104, n11105,
         n11106, n11107, n11108, n11109, n11110, n11111, n11112, n11113,
         n11114, n11115, n11116, n11117, n11118, n11119, n11120, n11121,
         n11122, n11123, n11124, n11125, n11126, n11127, n11128, n11129,
         n11130, n11131, n11132, n11133, n11134, n11135, n11136, n11137,
         n11138, n11139, n11140, n11141, n11142, n11143, n11144, n11145,
         n11146, n11147, n11148, n11149, n11150, n11151, n11152, n11153,
         n11154, n11155, n11156, n11157, n11158, n11159, n11160, n11161,
         n11162, n11163, n11164, n11165, n11166, n11167, n11168, n11169,
         n11170, n11171, n11172, n11173, n11174, n11175, n11176, n11177,
         n11178, n11179, n11180, n11181, n11182, n11183, n11184, n11185,
         n11186, n11187, n11188, n11189, n11190, n11191, n11192, n11193,
         n11194, n11195, n11196, n11197, n11198, n11199, n11200, n11201,
         n11202, n11203, n11204, n11205, n11206, n11207, n11208, n11209,
         n11210, n11211, n11212, n11213, n11214, n11215, n11216, n11217,
         n11218, n11219, n11220, n11221, n11222, n11223, n11224, n11225,
         n11226, n11227, n11228, n11229, n11230, n11231, n11232, n11233,
         n11234, n11235, n11236, n11237, n11238, n11239, n11240, n11241,
         n11242, n11243, n11244, n11245, n11246, n11247, n11248, n11249,
         n11250, n11251, n11252, n11253, n11254, n11255, n11256, n11257,
         n11258, n11259, n11260, n11261, n11262, n11263, n11264, n11265,
         n11266, n11267, n11268, n11269, n11270, n11271, n11272, n11273,
         n11274, n11275, n11276, n11277, n11278, n11279, n11280, n11281,
         n11282, n11283, n11284, n11285, n11286, n11287, n11288, n11289,
         n11290, n11291, n11292, n11293, n11294, n11295, n11296, n11297,
         n11298, n11299, n11300, n11301, n11302, n11303, n11304, n11305,
         n11306, n11307, n11308, n11309, n11310, n11311, n11312, n11313,
         n11314, n11315, n11316, n11317, n11318, n11319, n11320, n11321,
         n11322, n11323, n11324, n11325, n11326, n11327, n11328, n11329,
         n11330, n11331, n11332, n11333, n11334, n11335, n11336, n11337,
         n11338, n11339, n11340, n11341, n11342, n11343, n11344, n11345,
         n11346, n11347, n11348, n11349, n11350, n11351, n11352, n11353,
         n11354, n11355, n11356, n11357, n11358, n11359, n11360, n11361,
         n11362, n11363, n11364, n11365, n11366, n11367, n11368, n11369,
         n11370, n11371, n11372, n11373, n11374, n11375, n11376, n11377,
         n11378, n11379, n11380, n11381, n11382, n11383, n11384, n11385,
         n11386, n11387, n11388, n11389, n11390, n11391, n11392, n11393,
         n11394, n11395, n11396, n11397, n11398, n11399, n11400, n11401,
         n11402, n11403, n11404, n11405, n11406, n11407, n11408, n11409,
         n11410, n11411, n11412, n11413, n11414, n11415, n11416, n11417,
         n11418, n11419, n11420, n11421, n11422, n11423, n11424, n11425,
         n11426, n11427, n11428, n11429, n11430, n11431, n11432, n11433,
         n11434, n11435, n11436, n11437, n11438, n11439, n11440, n11441,
         n11442, n11443, n11444, n11445, n11446, n11447, n11448, n11449,
         n11450, n11451, n11452, n11453, n11454, n11455, n11456, n11457,
         n11458, n11459, n11460, n11461, n11462, n11463, n11464, n11465,
         n11466, n11467, n11468, n11469, n11470, n11471, n11472, n11473,
         n11474, n11475, n11476, n11477, n11478, n11479, n11480, n11481,
         n11482, n11483, n11484, n11485, n11486, n11487, n11488, n11489,
         n11490, n11491, n11492, n11493, n11494, n11495, n11496, n11497,
         n11498, n11499, n11500, n11501, n11502, n11503, n11504, n11505,
         n11506, n11507, n11508, n11509, n11510, n11511, n11512, n11513,
         n11514, n11515, n11516, n11517, n11518, n11519, n11520, n11521,
         n11522, n11523, n11524, n11525, n11526, n11527, n11528, n11529,
         n11530, n11531, n11532, n11533, n11534, n11535, n11536, n11537,
         n11538, n11539, n11540, n11541, n11542, n11543, n11544, n11545,
         n11546, n11547, n11548, n11549, n11550, n11551, n11552, n11553,
         n11554, n11555, n11556, n11557, n11558, n11559, n11560, n11561,
         n11562, n11563, n11564, n11565, n11566, n11567, n11568, n11569,
         n11570, n11571, n11572, n11573, n11574, n11575, n11576, n11577,
         n11578, n11579, n11580, n11581, n11582, n11583, n11584, n11585,
         n11586, n11587, n11588, n11589, n11590, n11591, n11592, n11593,
         n11594, n11595, n11596, n11597, n11598, n11599, n11600, n11601,
         n11602, n11603, n11604, n11605, n11606, n11607, n11608, n11609,
         n11610, n11611, n11612, n11613, n11614, n11615, n11616, n11617,
         n11618, n11619, n11620, n11621, n11622, n11623, n11624, n11625,
         n11626, n11627, n11628, n11629, n11630, n11631, n11632, n11633,
         n11634, n11635, n11636, n11637, n11638, n11639, n11640, n11641,
         n11642, n11643, n11644, n11645, n11646, n11647, n11648, n11649,
         n11650, n11651, n11652, n11653, n11654, n11655, n11656, n11657,
         n11658, n11659, n11660, n11661, n11662, n11663, n11664, n11665,
         n11666, n11667, n11668, n11669, n11670, n11671, n11672, n11673,
         n11674, n11675, n11676, n11677, n11678, n11679, n11680, n11681,
         n11682, n11683, n11684, n11685, n11686, n11687, n11688, n11689,
         n11690, n11691, n11692, n11693, n11694, n11695, n11696, n11697,
         n11698, n11699, n11700, n11701, n11702, n11703, n11704, n11705,
         n11706, n11707, n11708, n11709, n11710, n11711, n11712, n11713,
         n11714, n11715, n11716, n11717, n11718, n11719, n11720, n11721,
         n11722, n11723, n11724, n11725, n11726, n11727, n11728, n11729,
         n11730, n11731, n11732, n11733, n11734, n11735, n11736, n11737,
         n11738, n11739, n11740, n11741, n11742, n11743, n11744, n11745,
         n11746, n11747, n11748, n11749, n11750, n11751, n11752, n11753,
         n11754, n11755, n11756, n11757, n11758, n11759, n11760, n11761,
         n11762, n11763, n11764, n11765, n11766, n11767, n11768, n11769,
         n11770, n11771, n11772, n11773, n11774, n11775, n11776, n11777,
         n11778, n11779, n11780, n11781, n11782, n11783, n11784, n11785,
         n11786, n11787, n11788, n11789, n11790, n11791, n11792, n11793,
         n11794, n11795, n11796, n11797, n11798, n11799, n11800, n11801,
         n11802, n11803, n11804, n11805, n11806, n11807, n11808, n11809,
         n11810, n11811, n11812, n11813, n11814, n11815, n11816, n11817,
         n11818, n11819, n11820, n11821, n11822, n11823, n11824, n11825,
         n11826, n11827, n11828, n11829, n11830, n11831, n11832, n11833,
         n11834, n11835, n11836, n11837, n11838, n11839, n11840, n11841,
         n11842, n11843, n11844, n11845, n11846, n11847, n11848, n11849,
         n11850, n11851, n11852, n11853, n11854, n11855, n11856, n11857,
         n11858, n11859, n11860, n11861, n11862, n11863, n11864, n11865,
         n11866, n11867, n11868, n11869, n11870, n11871, n11872, n11873,
         n11874, n11875, n11876, n11877, n11878, n11879, n11880, n11881,
         n11882, n11883, n11884, n11885, n11886, n11887, n11888, n11889,
         n11890, n11891, n11892, n11893, n11894, n11895, n11896, n11897,
         n11898, n11899, n11900, n11901, n11902, n11903, n11904, n11905,
         n11906, n11907, n11908, n11909, n11910, n11911, n11912, n11913,
         n11914, n11915, n11916, n11917, n11918, n11919, n11920, n11921,
         n11922, n11923, n11924, n11925, n11926, n11927, n11928, n11929,
         n11930, n11931, n11932, n11933, n11934, n11935, n11936, n11937,
         n11938, n11939, n11940, n11941, n11942, n11943, n11944, n11945,
         n11946, n11947, n11948, n11949, n11950, n11951, n11952, n11953,
         n11954, n11955, n11956, n11957, n11958, n11959, n11960, n11961,
         n11962, n11963, n11964, n11965, n11966, n11967, n11968, n11969,
         n11970, n11971, n11972, n11973, n11974, n11975, n11976, n11977,
         n11978, n11979, n11980, n11981, n11982, n11983, n11984, n11985,
         n11986, n11987, n11988, n11989, n11990, n11991, n11992, n11993,
         n11994, n11995, n11996, n11997, n11998, n11999, n12000, n12001,
         n12002, n12003, n12004, n12005, n12006, n12007, n12008, n12009,
         n12010, n12011, n12012, n12013, n12014, n12015, n12016, n12017,
         n12018, n12019, n12020, n12021, n12022, n12023, n12024, n12025,
         n12026, n12027, n12028, n12029, n12030, n12031, n12032, n12033,
         n12034, n12035, n12036, n12037, n12038, n12039, n12040, n12041,
         n12042, n12043, n12044, n12045, n12046, n12047, n12048, n12049,
         n12050, n12051, n12052, n12053, n12054, n12055, n12056, n12057,
         n12058, n12059, n12060, n12061, n12062, n12063, n12064, n12065,
         n12066, n12067, n12068, n12069, n12070, n12071, n12072, n12073,
         n12074, n12075, n12076, n12077, n12078, n12079, n12080, n12081,
         n12082, n12083, n12084, n12085, n12086, n12087, n12088, n12089,
         n12090, n12091, n12092, n12093, n12094, n12095, n12096, n12097,
         n12098, n12099, n12100, n12101, n12102, n12103, n12104, n12105,
         n12106, n12107, n12108, n12109, n12110, n12111, n12112, n12113,
         n12114, n12115, n12116, n12117, n12118, n12119, n12120, n12121,
         n12122, n12123, n12124, n12125, n12126, n12127, n12128, n12129,
         n12130, n12131, n12132, n12133, n12134, n12135, n12136, n12137,
         n12138, n12139, n12140, n12141, n12142, n12143, n12144, n12145,
         n12146, n12147, n12148, n12149, n12150, n12151, n12152, n12153,
         n12154, n12155, n12156, n12157, n12158, n12159, n12160, n12161,
         n12162, n12163, n12164, n12165, n12166, n12167, n12168, n12169,
         n12170, n12171, n12172, n12173, n12174, n12175, n12176, n12177,
         n12178, n12179, n12180, n12181, n12182, n12183, n12184, n12185,
         n12186, n12187, n12188, n12189, n12190, n12191, n12192, n12193,
         n12194, n12195, n12196, n12197, n12198, n12199, n12200, n12201,
         n12202, n12203, n12204, n12205, n12206, n12207, n12208, n12209,
         n12210, n12211, n12212, n12213, n12214, n12215, n12216, n12217,
         n12218, n12219, n12220, n12221, n12222, n12223, n12224, n12225,
         n12226, n12227, n12228, n12229, n12230, n12231, n12232, n12233,
         n12234, n12235, n12236, n12237, n12238, n12239, n12240, n12241,
         n12242, n12243, n12244, n12245, n12246, n12247, n12248, n12249,
         n12250, n12251, n12252, n12253, n12254, n12255, n12256, n12257,
         n12258, n12259, n12260, n12261, n12262, n12263, n12264, n12265,
         n12266, n12267, n12268, n12269, n12270, n12271, n12272, n12273,
         n12274, n12275, n12276, n12277, n12278, n12279, n12280, n12281,
         n12282, n12283, n12284, n12285, n12286, n12287, n12288, n12289,
         n12290, n12291, n12292, n12293, n12294, n12295, n12296, n12297,
         n12298, n12299, n12300, n12301, n12302, n12303, n12304, n12305,
         n12306, n12307, n12308, n12309, n12310, n12311, n12312, n12313,
         n12314, n12315, n12316, n12317, n12318, n12319, n12320, n12321,
         n12322, n12323, n12324, n12325, n12326, n12327, n12328, n12329,
         n12330, n12331, n12332, n12333, n12334, n12335, n12336, n12337,
         n12338, n12339, n12340, n12341, n12342, n12343, n12344, n12345,
         n12346, n12347, n12348, n12349, n12350, n12351, n12352, n12353,
         n12354, n12355, n12356, n12357, n12358, n12359, n12360, n12361,
         n12362, n12363, n12364, n12365, n12366, n12367, n12368, n12369,
         n12370, n12371, n12372, n12373, n12374, n12375, n12376, n12377,
         n12378, n12379, n12380, n12381, n12382, n12383, n12384, n12385,
         n12386, n12387, n12388, n12389, n12390, n12391, n12392, n12393,
         n12394, n12395, n12396, n12397, n12398, n12399, n12400, n12401,
         n12402, n12403, n12404, n12405, n12406, n12407, n12408, n12409,
         n12410, n12411, n12412, n12413, n12414, n12415, n12416, n12417,
         n12418, n12419, n12420, n12421, n12422, n12423, n12424, n12425,
         n12426, n12427, n12428, n12429, n12430, n12431, n12432, n12433,
         n12434, n12435, n12436, n12437, n12438, n12439, n12440, n12441,
         n12442, n12443, n12444, n12445, n12446, n12447, n12448, n12449,
         n12450, n12451, n12452, n12453, n12454, n12455, n12456, n12457,
         n12458, n12459, n12460, n12461, n12462, n12463, n12464, n12465,
         n12466, n12467, n12468, n12469, n12470, n12471, n12472, n12473,
         n12474, n12475, n12476, n12477, n12478, n12479, n12480, n12481,
         n12482, n12483, n12484, n12485, n12486, n12487, n12488, n12489,
         n12490, n12491, n12492, n12493, n12494, n12495, n12496, n12497,
         n12498, n12499, n12500, n12501, n12502, n12503, n12504, n12505,
         n12506, n12507, n12508, n12509, n12510, n12511, n12512, n12513,
         n12514, n12515, n12516, n12517, n12518, n12519, n12520, n12521,
         n12522, n12523, n12524, n12525, n12526, n12527, n12528, n12529,
         n12530, n12531, n12532, n12533, n12534, n12535, n12536, n12537,
         n12538, n12539, n12540, n12541, n12542, n12543, n12544, n12545,
         n12546, n12547, n12548, n12549, n12550, n12551, n12552, n12553,
         n12554, n12555, n12556, n12557, n12558, n12559, n12560, n12561,
         n12562, n12563, n12564, n12565, n12566, n12567, n12568, n12569,
         n12570, n12571, n12572, n12573, n12574, n12575, n12576, n12577,
         n12578, n12579, n12580, n12581, n12582, n12583, n12584, n12585,
         n12586, n12587, n12588, n12589, n12590, n12591, n12592, n12593,
         n12594, n12595, n12596, n12597, n12598, n12599, n12600, n12601,
         n12602, n12603, n12604, n12605, n12606, n12607, n12608, n12609,
         n12610, n12611, n12612, n12613, n12614, n12615, n12616, n12617,
         n12618, n12619, n12620, n12621, n12622, n12623, n12624, n12625,
         n12626, n12627, n12628, n12629, n12630, n12631, n12632, n12633,
         n12634, n12635, n12636, n12637, n12638, n12639, n12640, n12641,
         n12642, n12643, n12644, n12645, n12646, n12647, n12648, n12649,
         n12650, n12651, n12652, n12653, n12654, n12655, n12656, n12657,
         n12658, n12659, n12660, n12661, n12662, n12663, n12664, n12665,
         n12666, n12667, n12668, n12669, n12670, n12671, n12672, n12673,
         n12674, n12675, n12676, n12677, n12678, n12679, n12680, n12681,
         n12682, n12683, n12684, n12685, n12686, n12687, n12688, n12689,
         n12690, n12691, n12692, n12693, n12694, n12695, n12696, n12697,
         n12698, n12699, n12700, n12701, n12702, n12703, n12704, n12705,
         n12706, n12707, n12708, n12709, n12710, n12711, n12712, n12713,
         n12714, n12715, n12716, n12717, n12718, n12719, n12720, n12721,
         n12722, n12723, n12724, n12725, n12726, n12727, n12728, n12729,
         n12730, n12731, n12732, n12733, n12734, n12735, n12736, n12737,
         n12738, n12739, n12740, n12741, n12742, n12743, n12744, n12745,
         n12746, n12747, n12748, n12749, n12750, n12751, n12752, n12753,
         n12754, n12755, n12756, n12757, n12758, n12759, n12760, n12761,
         n12762, n12763, n12764, n12765, n12766, n12767, n12768, n12769,
         n12770, n12771, n12772, n12773, n12774, n12775, n12776, n12777,
         n12778, n12779, n12780, n12781, n12782, n12783, n12784, n12785,
         n12786, n12787, n12788, n12789, n12790, n12791, n12792, n12793,
         n12794, n12795, n12796, n12797, n12798, n12799, n12800, n12801,
         n12802, n12803, n12804, n12805, n12806, n12807, n12808, n12809,
         n12810, n12811, n12812, n12813, n12814, n12815, n12816, n12817,
         n12818, n12819, n12820, n12821, n12822, n12823, n12824, n12825,
         n12826, n12827, n12828, n12829, n12830, n12831, n12832, n12833,
         n12834, n12835, n12836, n12837, n12838, n12839, n12840, n12841,
         n12842, n12843, n12844, n12845, n12846, n12847, n12848, n12849,
         n12850, n12851, n12852, n12853, n12854, n12855, n12856, n12857,
         n12858, n12859, n12860, n12861, n12862, n12863, n12864, n12865,
         n12866, n12867, n12868, n12869, n12870, n12871, n12872, n12873,
         n12874, n12875, n12876, n12877, n12878, n12879, n12880, n12881,
         n12882, n12883, n12884, n12885, n12886, n12887, n12888, n12889,
         n12890, n12891, n12892, n12893, n12894, n12895, n12896, n12897,
         n12898, n12899, n12900, n12901, n12902, n12903, n12904, n12905,
         n12906, n12907, n12908, n12909, n12910, n12911, n12912, n12913,
         n12914, n12915, n12916, n12917, n12918, n12919, n12920, n12921,
         n12922, n12923, n12924, n12925, n12926, n12927, n12928, n12929,
         n12930, n12931, n12932, n12933, n12934, n12935, n12936, n12937,
         n12938, n12939, n12940, n12941, n12942, n12943, n12944, n12945,
         n12946, n12947, n12948, n12949, n12950, n12951, n12952, n12953,
         n12954, n12955, n12956, n12957, n12958, n12959, n12960, n12961,
         n12962, n12963, n12964, n12965, n12966, n12967, n12968, n12969,
         n12970, n12971, n12972, n12973, n12974, n12975, n12976, n12977,
         n12978, n12979, n12980, n12981, n12982, n12983, n12984, n12985,
         n12986, n12987, n12988, n12989, n12990, n12991, n12992, n12993,
         n12994, n12995, n12996, n12997, n12998, n12999, n13000, n13001,
         n13002, n13003, n13004, n13005, n13006, n13007, n13008, n13009,
         n13010, n13011, n13012, n13013, n13014, n13015, n13016, n13017,
         n13018, n13019, n13020, n13021, n13022, n13023, n13024, n13025,
         n13026, n13027, n13028, n13029, n13030, n13031, n13032, n13033,
         n13034, n13035, n13036, n13037, n13038, n13039, n13040, n13041,
         n13042, n13043, n13044, n13045, n13046, n13047, n13048, n13049,
         n13050, n13051, n13052, n13053, n13054, n13055, n13056, n13057,
         n13058, n13059, n13060, n13061, n13062, n13063, n13064, n13065,
         n13066, n13067, n13068, n13069, n13070, n13071, n13072, n13073,
         n13074, n13075, n13076, n13077, n13078, n13079, n13080, n13081,
         n13082, n13083, n13084, n13085, n13086, n13087, n13088, n13089,
         n13090, n13091, n13092, n13093, n13094, n13095, n13096, n13097,
         n13098, n13099, n13100, n13101, n13102, n13103, n13104, n13105,
         n13106, n13107, n13108, n13109, n13110, n13111, n13112, n13113,
         n13114, n13115, n13116, n13117, n13118, n13119, n13120, n13121,
         n13122, n13123, n13124, n13125, n13126, n13127, n13128, n13129,
         n13130, n13131, n13132, n13133, n13134, n13135, n13136, n13137,
         n13138, n13139, n13140, n13141, n13142, n13143, n13144, n13145,
         n13146, n13147, n13148, n13149, n13150, n13151, n13152, n13153,
         n13154, n13155, n13156, n13157, n13158, n13159, n13160, n13161,
         n13162, n13163, n13164, n13165, n13166, n13167, n13168, n13169,
         n13170, n13171, n13172, n13173, n13174, n13175, n13176, n13177,
         n13178, n13179, n13180, n13181, n13182, n13183, n13184, n13185,
         n13186, n13187, n13188, n13189, n13190, n13191, n13192, n13193,
         n13194, n13195, n13196, n13197, n13198, n13199, n13200, n13201,
         n13202, n13203, n13204, n13205, n13206, n13207, n13208, n13209,
         n13210, n13211, n13212, n13213, n13214, n13215, n13216, n13217,
         n13218, n13219, n13220, n13221, n13222, n13223, n13224, n13225,
         n13226, n13227, n13228, n13229, n13230, n13231, n13232, n13233,
         n13234, n13235, n13236, n13237, n13238, n13239, n13240, n13241,
         n13242, n13243, n13244, n13245, n13246, n13247, n13248, n13249,
         n13250, n13251, n13252, n13253, n13254, n13255, n13256, n13257,
         n13258, n13259, n13260, n13261, n13262, n13263, n13264, n13265,
         n13266, n13267, n13268, n13269, n13270, n13271, n13272, n13273,
         n13274, n13275, n13276, n13277, n13278, n13279, n13280, n13281,
         n13282, n13283, n13284, n13285, n13286, n13287, n13288, n13289,
         n13290, n13291, n13292, n13293, n13294, n13295, n13296, n13297,
         n13298, n13299, n13300, n13301, n13302, n13303, n13304, n13305,
         n13306, n13307, n13308, n13309, n13310, n13311, n13312, n13313,
         n13314, n13315, n13316, n13317, n13318, n13319, n13320, n13321,
         n13322, n13323, n13324, n13325, n13326, n13327, n13328, n13329,
         n13330, n13331, n13332, n13333, n13334, n13335, n13336, n13337,
         n13338, n13339, n13340, n13341, n13342, n13343, n13344, n13345,
         n13346, n13347, n13348, n13349, n13350, n13351, n13352, n13353,
         n13354, n13355, n13356, n13357, n13358, n13359, n13360, n13361,
         n13362, n13363, n13364, n13365, n13366, n13367, n13368, n13369,
         n13370, n13371, n13372, n13373, n13374, n13375, n13376, n13377,
         n13378, n13379, n13380, n13381, n13382, n13383, n13384, n13385,
         n13386, n13387, n13388, n13389, n13390, n13391, n13392, n13393,
         n13394, n13395, n13396, n13397, n13398, n13399, n13400, n13401,
         n13402, n13403, n13404, n13405, n13406, n13407, n13408, n13409,
         n13410, n13411, n13412, n13413, n13414, n13415, n13416, n13417,
         n13418, n13419, n13420, n13421, n13422, n13423, n13424, n13425,
         n13426, n13427, n13428, n13429, n13430, n13431, n13432, n13433,
         n13434, n13435, n13436, n13437, n13438, n13439, n13440, n13441,
         n13442, n13443, n13444, n13445, n13446, n13447, n13448, n13449,
         n13450, n13451, n13452, n13453, n13454, n13455, n13456, n13457,
         n13458, n13459, n13460, n13461, n13462, n13463, n13464, n13465,
         n13466, n13467, n13468, n13469, n13470, n13471, n13472, n13473,
         n13474, n13475, n13476, n13477, n13478, n13479, n13480, n13481,
         n13482, n13483, n13484, n13485, n13486, n13487, n13488, n13489,
         n13490, n13491, n13492, n13493, n13494, n13495, n13496, n13497,
         n13498, n13499, n13500, n13501, n13502, n13503, n13504, n13505,
         n13506, n13507, n13508, n13509, n13510, n13511, n13512, n13513,
         n13514, n13515, n13516, n13517, n13518, n13519, n13520, n13521,
         n13522, n13523, n13524, n13525, n13526, n13527, n13528, n13529,
         n13530, n13531, n13532, n13533, n13534, n13535, n13536, n13537,
         n13538, n13539, n13540, n13541, n13542, n13543, n13544, n13545,
         n13546, n13547, n13548, n13549, n13550, n13551, n13552, n13553,
         n13554, n13555, n13556, n13557, n13558, n13559, n13560, n13561,
         n13562, n13563, n13564, n13565, n13566, n13567, n13568, n13569,
         n13570, n13571, n13572, n13573, n13574, n13575, n13576, n13577,
         n13578, n13579, n13580, n13581, n13582, n13583, n13584, n13585,
         n13586, n13587, n13588, n13589, n13590, n13591, n13592, n13593,
         n13594, n13595, n13596, n13597, n13598, n13599, n13600, n13601,
         n13602, n13603, n13604, n13605, n13606, n13607, n13608, n13609,
         n13610, n13611, n13612, n13613, n13614, n13615, n13616, n13617,
         n13618, n13619, n13620, n13621, n13622, n13623, n13624, n13625,
         n13626, n13627, n13628, n13629, n13630, n13631, n13632, n13633,
         n13634, n13635, n13636, n13637, n13638, n13639, n13640, n13641,
         n13642, n13643, n13644, n13645, n13646, n13647, n13648, n13649,
         n13650, n13651, n13652, n13653, n13654, n13655, n13656, n13657,
         n13658, n13659, n13660, n13661, n13662, n13663, n13664, n13665,
         n13666, n13667, n13668, n13669, n13670, n13671, n13672, n13673,
         n13674, n13675, n13676, n13677, n13678, n13679, n13680, n13681,
         n13682, n13683, n13684, n13685, n13686, n13687, n13688, n13689,
         n13690, n13691, n13692, n13693, n13694, n13695, n13696, n13697,
         n13698, n13699, n13700, n13701, n13702, n13703, n13704, n13705,
         n13706, n13707, n13708, n13709, n13710, n13711, n13712, n13713,
         n13714, n13715, n13716, n13717, n13718, n13719, n13720, n13721,
         n13722, n13723, n13724, n13725, n13726, n13727, n13728, n13729,
         n13730, n13731, n13732, n13733, n13734, n13735, n13736, n13737,
         n13738, n13739, n13740, n13741, n13742, n13743, n13744, n13745,
         n13746, n13747, n13748, n13749, n13750, n13751, n13752, n13753,
         n13754, n13755, n13756, n13757, n13758, n13759, n13760, n13761,
         n13762, n13763, n13764, n13765, n13766, n13767, n13768, n13769,
         n13770, n13771, n13772, n13773, n13774, n13775, n13776, n13777,
         n13778, n13779, n13780, n13781, n13782, n13783, n13784, n13785,
         n13786, n13787, n13788, n13789, n13790, n13791, n13792, n13793,
         n13794, n13795, n13796, n13797, n13798, n13799, n13800, n13801,
         n13802, n13803, n13804, n13805, n13806, n13807, n13808, n13809,
         n13810, n13811, n13812, n13813, n13814, n13815, n13816, n13817,
         n13818, n13819, n13820, n13821, n13822, n13823, n13824, n13825,
         n13826, n13827, n13828, n13829, n13830, n13831, n13832, n13833,
         n13834, n13835, n13836, n13837, n13838, n13839, n13840, n13841,
         n13842, n13843, n13844, n13845, n13846, n13847, n13848, n13849,
         n13850, n13851, n13852, n13853, n13854, n13855, n13856, n13857,
         n13858, n13859, n13860, n13861, n13862, n13863, n13864, n13865,
         n13866, n13867, n13868, n13869, n13870, n13871, n13872, n13873,
         n13874, n13875, n13876, n13877, n13878, n13879, n13880, n13881,
         n13882, n13883, n13884, n13885, n13886, n13887, n13888, n13889,
         n13890, n13891, n13892, n13893, n13894, n13895, n13896, n13897,
         n13898, n13899, n13900, n13901, n13902, n13903, n13904, n13905,
         n13906, n13907, n13908, n13909, n13910, n13911, n13912, n13913,
         n13914, n13915, n13916, n13917, n13918, n13919, n13920, n13921,
         n13922, n13923, n13924, n13925, n13926, n13927, n13928, n13929,
         n13930, n13931, n13932, n13933, n13934, n13935, n13936, n13937,
         n13938, n13939, n13940, n13941, n13942, n13943, n13944, n13945,
         n13946, n13947, n13948, n13949, n13950, n13951, n13952, n13953,
         n13954, n13955, n13956, n13957, n13958, n13959, n13960, n13961,
         n13962, n13963, n13964, n13965, n13966, n13967, n13968, n13969,
         n13970, n13971, n13972, n13973, n13974, n13975, n13976, n13977,
         n13978, n13979, n13980, n13981, n13982, n13983, n13984, n13985,
         n13986, n13987, n13988, n13989, n13990, n13991, n13992, n13993,
         n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001,
         n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009,
         n14010, n14011, n14012, n14013, n14014, n14015, n14016, n14017,
         n14018, n14019, n14020, n14021, n14022, n14023, n14024, n14025,
         n14026, n14027, n14028, n14029, n14030, n14031, n14032, n14033,
         n14034, n14035, n14036, n14037, n14038, n14039, n14040, n14041,
         n14042, n14043, n14044, n14045, n14046, n14047, n14048, n14049,
         n14050, n14051, n14052, n14053, n14054, n14055, n14056, n14057,
         n14058, n14059, n14060, n14061, n14062, n14063, n14064, n14065,
         n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073,
         n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081,
         n14082, n14083, n14084, n14085, n14086, n14087, n14088, n14089,
         n14090, n14091, n14092, n14093, n14094, n14095, n14096, n14097,
         n14098, n14099, n14100, n14101, n14102, n14103, n14104, n14105,
         n14106, n14107, n14108, n14109, n14110, n14111, n14112, n14113,
         n14114, n14115, n14116, n14117, n14118, n14119, n14120, n14121,
         n14122, n14123, n14124, n14125, n14126, n14127, n14128, n14129,
         n14130, n14131, n14132, n14133, n14134, n14135, n14136, n14137,
         n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145,
         n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153,
         n14154, n14155, n14156, n14157, n14158, n14159, n14160, n14161,
         n14162, n14163, n14164, n14165, n14166, n14167, n14168, n14169,
         n14170, n14171, n14172, n14173, n14174, n14175, n14176, n14177,
         n14178, n14179, n14180, n14181, n14182, n14183, n14184, n14185,
         n14186, n14187, n14188, n14189, n14190, n14191, n14192, n14193,
         n14194, n14195, n14196, n14197, n14198, n14199, n14200, n14201,
         n14202, n14203, n14204, n14205, n14206, n14207, n14208, n14209,
         n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217,
         n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225,
         n14226, n14227, n14228, n14229, n14230, n14231, n14232, n14233,
         n14234, n14235, n14236, n14237, n14238, n14239, n14240, n14241,
         n14242, n14243, n14244, n14245, n14246, n14247, n14248, n14249,
         n14250, n14251, n14252, n14253, n14254, n14255, n14256, n14257,
         n14258, n14259, n14260, n14261, n14262, n14263, n14264, n14265,
         n14266, n14267, n14268, n14269, n14270, n14271, n14272, n14273,
         n14274, n14275, n14276, n14277, n14278, n14279, n14280, n14281,
         n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289,
         n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297,
         n14298, n14299, n14300, n14301, n14302, n14303, n14304, n14305,
         n14306, n14307, n14308, n14309, n14310, n14311, n14312, n14313,
         n14314, n14315, n14316, n14317, n14318, n14319, n14320, n14321,
         n14322, n14323, n14324, n14325, n14326, n14327, n14328, n14329,
         n14330, n14331, n14332, n14333, n14334, n14335, n14336, n14337,
         n14338, n14339, n14340, n14341, n14342, n14343, n14344, n14345,
         n14346, n14347, n14348, n14349, n14350, n14351, n14352, n14353,
         n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361,
         n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369,
         n14370, n14371, n14372, n14373, n14374, n14375, n14376, n14377,
         n14378, n14379, n14380, n14381, n14382, n14383, n14384, n14385,
         n14386, n14387, n14388, n14389, n14390, n14391, n14392, n14393,
         n14394, n14395, n14396, n14397, n14398, n14399, n14400, n14401,
         n14402, n14403, n14404, n14405, n14406, n14407, n14408, n14409,
         n14410, n14411, n14412, n14413, n14414, n14415, n14416, n14417,
         n14418, n14419, n14420, n14421, n14422, n14423, n14424, n14425,
         n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433,
         n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441,
         n14442, n14443, n14444, n14445, n14446, n14447, n14448, n14449,
         n14450, n14451, n14452, n14453, n14454, n14455, n14456, n14457,
         n14458, n14459, n14460, n14461, n14462, n14463, n14464, n14465,
         n14466, n14467, n14468, n14469, n14470, n14471, n14472, n14473,
         n14474, n14475, n14476, n14477, n14478, n14479, n14480, n14481,
         n14482, n14483, n14484, n14485, n14486, n14487, n14488, n14489,
         n14490, n14491, n14492, n14493, n14494, n14495, n14496, n14497,
         n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505,
         n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513,
         n14514, n14515, n14516, n14517, n14518, n14519, n14520, n14521,
         n14522, n14523, n14524, n14525, n14526, n14527, n14528, n14529,
         n14530, n14531, n14532, n14533, n14534, n14535, n14536, n14537,
         n14538, n14539, n14540, n14541, n14542, n14543, n14544, n14545,
         n14546, n14547, n14548, n14549, n14550, n14551, n14552, n14553,
         n14554, n14555, n14556, n14557, n14558, n14559, n14560, n14561,
         n14562, n14563, n14564, n14565, n14566, n14567, n14568, n14569,
         n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577,
         n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585,
         n14586, n14587, n14588, n14589, n14590, n14591, n14592, n14593,
         n14594, n14595, n14596, n14597, n14598, n14599, n14600, n14601,
         n14602, n14603, n14604, n14605, n14606, n14607, n14608, n14609,
         n14610, n14611, n14612, n14613, n14614, n14615, n14616, n14617,
         n14618, n14619, n14620, n14621, n14622, n14623, n14624, n14625,
         n14626, n14627, n14628, n14629, n14630, n14631, n14632, n14633,
         n14634, n14635, n14636, n14637, n14638, n14639, n14640, n14641,
         n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649,
         n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657,
         n14658, n14659, n14660, n14661, n14662, n14663, n14664, n14665,
         n14666, n14667, n14668, n14669, n14670, n14671, n14672, n14673,
         n14674, n14675, n14676, n14677, n14678, n14679, n14680, n14681,
         n14682, n14683, n14684, n14685, n14686, n14687, n14688, n14689,
         n14690, n14691, n14692, n14693, n14694, n14695, n14696, n14697,
         n14698, n14699, n14700, n14701, n14702, n14703, n14704, n14705,
         n14706, n14707, n14708, n14709, n14710, n14711, n14712, n14713,
         n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721,
         n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729,
         n14730, n14731, n14732, n14733, n14734, n14735, n14736, n14737,
         n14738, n14739, n14740, n14741, n14742, n14743, n14744, n14745,
         n14746, n14747, n14748, n14749, n14750, n14751, n14752, n14753,
         n14754, n14755, n14756, n14757, n14758, n14759, n14760, n14761,
         n14762, n14763, n14764, n14765, n14766, n14767, n14768, n14769,
         n14770, n14771, n14772, n14773, n14774, n14775, n14776, n14777,
         n14778, n14779, n14780, n14781, n14782, n14783, n14784, n14785,
         n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793,
         n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801,
         n14802, n14803, n14804, n14805, n14806, n14807, n14808, n14809,
         n14810, n14811, n14812, n14813, n14814, n14815, n14816, n14817,
         n14818, n14819, n14820, n14821, n14822, n14823, n14824, n14825,
         n14826, n14827, n14828, n14829, n14830, n14831, n14832, n14833,
         n14834, n14835, n14836, n14837, n14838, n14839, n14840, n14841,
         n14842, n14843, n14844, n14845, n14846, n14847, n14848, n14849,
         n14850, n14851, n14852, n14853, n14854, n14855, n14856, n14857,
         n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865,
         n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873,
         n14874, n14875, n14876, n14877, n14878, n14879, n14880, n14881,
         n14882, n14883, n14884, n14885, n14886, n14887, n14888, n14889,
         n14890, n14891, n14892, n14893, n14894, n14895, n14896, n14897,
         n14898, n14899, n14900, n14901, n14902, n14903, n14904, n14905,
         n14906, n14907, n14908, n14909, n14910, n14911, n14912, n14913,
         n14914, n14915, n14916, n14917, n14918, n14919, n14920, n14921,
         n14922, n14923, n14924, n14925, n14926, n14927, n14928, n14929,
         n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937,
         n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945,
         n14946, n14947, n14948, n14949, n14950, n14951, n14952, n14953,
         n14954, n14955, n14956, n14957, n14958, n14959, n14960, n14961,
         n14962, n14963, n14964, n14965, n14966, n14967, n14968, n14969,
         n14970, n14971, n14972, n14973, n14974, n14975, n14976, n14977,
         n14978, n14979, n14980, n14981, n14982, n14983, n14984, n14985,
         n14986, n14987, n14988, n14989, n14990, n14991, n14992, n14993,
         n14994, n14995, n14996, n14997, n14998, n14999, n15000, n15001,
         n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009,
         n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017,
         n15018, n15019, n15020, n15021, n15022, n15023, n15024, n15025,
         n15026, n15027, n15028, n15029, n15030, n15031, n15032, n15033,
         n15034, n15035, n15036, n15037, n15038, n15039, n15040, n15041,
         n15042, n15043, n15044, n15045, n15046, n15047, n15048, n15049,
         n15050, n15051, n15052, n15053, n15054, n15055, n15056, n15057,
         n15058, n15059, n15060, n15061, n15062, n15063, n15064, n15065,
         n15066, n15067, n15068, n15069, n15070, n15071, n15072, n15073,
         n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081,
         n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089,
         n15090, n15091, n15092, n15093, n15094, n15095, n15096, n15097,
         n15098, n15099, n15100, n15101, n15102, n15103, n15104, n15105,
         n15106, n15107, n15108, n15109, n15110, n15111, n15112, n15113,
         n15114, n15115, n15116, n15117, n15118, n15119, n15120, n15121,
         n15122, n15123, n15124, n15125, n15126, n15127, n15128, n15129,
         n15130, n15131, n15132, n15133, n15134, n15135, n15136, n15137,
         n15138, n15139, n15140, n15141, n15142, n15143, n15144, n15145,
         n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153,
         n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161,
         n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169,
         n15170, n15171, n15172, n15173, n15174, n15175, n15176, n15177,
         n15178, n15179, n15180, n15181, n15182, n15183, n15184, n15185,
         n15186, n15187, n15188, n15189, n15190, n15191, n15192, n15193,
         n15194, n15195, n15196, n15197, n15198, n15199, n15200, n15201,
         n15202, n15203, n15204, n15205, n15206, n15207, n15208, n15209,
         n15210, n15211, n15212, n15213, n15214, n15215, n15216, n15217,
         n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225,
         n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233,
         n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241,
         n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249,
         n15250, n15251, n15252, n15253, n15254, n15255, n15256, n15257,
         n15258, n15259, n15260, n15261, n15262, n15263, n15264, n15265,
         n15266, n15267, n15268, n15269, n15270, n15271, n15272, n15273,
         n15274, n15275, n15276, n15277, n15278, n15279, n15280, n15281,
         n15282, n15283, n15284, n15285, n15286, n15287, n15288, n15289,
         n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297,
         n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305,
         n15306, n15307, n15308, n15309, n15310, n15311, n15312, n15313,
         n15314, n15315, n15316, n15317, n15318, n15319, n15320, n15321,
         n15322, n15323, n15324, n15325, n15326, n15327, n15328, n15329,
         n15330, n15331, n15332, n15333, n15334, n15335, n15336, n15337,
         n15338, n15339, n15340, n15341, n15342, n15343, n15344, n15345,
         n15346, n15347, n15348, n15349, n15350, n15351, n15352, n15353,
         n15354, n15355, n15356, n15357, n15358, n15359, n15360, n15361,
         n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369,
         n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377,
         n15378, n15379, n15380, n15381, n15382, n15383, n15384, n15385,
         n15386, n15387, n15388, n15389, n15390, n15391, n15392, n15393,
         n15394, n15395, n15396, n15397, n15398, n15399, n15400, n15401,
         n15402, n15403, n15404, n15405, n15406, n15407, n15408, n15409,
         n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417,
         n15418, n15419, n15420, n15421, n15422, n15423, n15424, n15425,
         n15426, n15427, n15428, n15429, n15430, n15431, n15432, n15433,
         n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441,
         n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449,
         n15450, n15451, n15452, n15453, n15454, n15455, n15456, n15457,
         n15458, n15459, n15460, n15461, n15462, n15463, n15464, n15465,
         n15466, n15467, n15468, n15469, n15470, n15471, n15472, n15473,
         n15474, n15475, n15476, n15477, n15478, n15479, n15480, n15481,
         n15482, n15483, n15484, n15485, n15486, n15487, n15488, n15489,
         n15490, n15491, n15492, n15493, n15494, n15495, n15496, n15497,
         n15498, n15499, n15500, n15501, n15502, n15503, n15504, n15505,
         n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513,
         n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521,
         n15522, n15523, n15524, n15525, n15526, n15527, n15528, n15529,
         n15530, n15531, n15532, n15533, n15534, n15535, n15536, n15537,
         n15538, n15539, n15540, n15541, n15542, n15543, n15544, n15545,
         n15546, n15547, n15548, n15549, n15550, n15551, n15552, n15553,
         n15554, n15555, n15556, n15557, n15558, n15559, n15560, n15561,
         n15562, n15563, n15564, n15565, n15566, n15567, n15568, n15569,
         n15570, n15571, n15572, n15573, n15574, n15575, n15576, n15577,
         n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585,
         n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593,
         n15594, n15595, n15596, n15597, n15598, n15599, n15600, n15601,
         n15602, n15603, n15604, n15605, n15606, n15607, n15608, n15609,
         n15610, n15611, n15612, n15613, n15614, n15615, n15616, n15617,
         n15618, n15619, n15620, n15621, n15622, n15623, n15624, n15625,
         n15626, n15627, n15628, n15629, n15630, n15631, n15632, n15633,
         n15634, n15635, n15636, n15637, n15638, n15639, n15640, n15641,
         n15642, n15643, n15644, n15645, n15646, n15647, n15648, n15649,
         n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657,
         n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665,
         n15666, n15667, n15668, n15669, n15670, n15671, n15672, n15673,
         n15674, n15675, n15676, n15677, n15678, n15679, n15680, n15681,
         n15682, n15683, n15684, n15685, n15686, n15687, n15688, n15689,
         n15690, n15691, n15692, n15693, n15694, n15695, n15696, n15697,
         n15698, n15699, n15700, n15701, n15702, n15703, n15704, n15705,
         n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713,
         n15714, n15715, n15716, n15717, n15718, n15719, n15720, n15721,
         n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729,
         n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737,
         n15738, n15739, n15740, n15741, n15742, n15743, n15744, n15745,
         n15746, n15747, n15748, n15749, n15750, n15751, n15752, n15753,
         n15754, n15755, n15756, n15757, n15758, n15759, n15760, n15761,
         n15762, n15763, n15764, n15765, n15766, n15767, n15768, n15769,
         n15770, n15771, n15772, n15773, n15774, n15775, n15776, n15777,
         n15778, n15779, n15780, n15781, n15782, n15783, n15784, n15785,
         n15786, n15787, n15788, n15789, n15790, n15791, n15792, n15793,
         n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801,
         n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809,
         n15810, n15811, n15812, n15813, n15814, n15815, n15816, n15817,
         n15818, n15819, n15820, n15821, n15822, n15823, n15824, n15825,
         n15826, n15827, n15828, n15829, n15830, n15831, n15832, n15833,
         n15834, n15835, n15836, n15837, n15838, n15839, n15840, n15841,
         n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849,
         n15850, n15851, n15852, n15853, n15854, n15855, n15856, n15857,
         n15858, n15859, n15860, n15861, n15862, n15863, n15864, n15865,
         n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873,
         n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881,
         n15882, n15883, n15884, n15885, n15886, n15887, n15888, n15889,
         n15890, n15891, n15892, n15893, n15894, n15895, n15896, n15897,
         n15898, n15899, n15900, n15901, n15902, n15903, n15904, n15905,
         n15906, n15907, n15908, n15909, n15910, n15911, n15912, n15913,
         n15914, n15915, n15916, n15917, n15918, n15919, n15920, n15921,
         n15922, n15923, n15924, n15925, n15926, n15927, n15928, n15929,
         n15930, n15931, n15932, n15933, n15934, n15935, n15936, n15937,
         n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945,
         n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953,
         n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961,
         n15962, n15963, n15964, n15965, n15966, n15967, n15968, n15969,
         n15970, n15971, n15972, n15973, n15974, n15975, n15976, n15977,
         n15978, n15979, n15980, n15981, n15982, n15983, n15984, n15985,
         n15986, n15987, n15988, n15989, n15990, n15991, n15992, n15993,
         n15994, n15995, n15996, n15997, n15998, n15999, n16000, n16001,
         n16002, n16003, n16004, n16005, n16006, n16007, n16008, n16009,
         n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017,
         n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025,
         n16026, n16027, n16028, n16029, n16030, n16031, n16032, n16033,
         n16034, n16035, n16036, n16037, n16038, n16039, n16040, n16041,
         n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049,
         n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057,
         n16058, n16059, n16060, n16061, n16062, n16063, n16064, n16065,
         n16066, n16067, n16068, n16069, n16070, n16071, n16072, n16073,
         n16074, n16075, n16076, n16077, n16078, n16079, n16080, n16081,
         n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089,
         n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097,
         n16098, n16099, n16100, n16101, n16102, n16103, n16104, n16105,
         n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113,
         n16114, n16115, n16116, n16117, n16118, n16119, n16120, n16121,
         n16122, n16123, n16124, n16125, n16126, n16127, n16128, n16129,
         n16130, n16131, n16132, n16133, n16134, n16135, n16136, n16137,
         n16138, n16139, n16140, n16141, n16142, n16143, n16144, n16145,
         n16146, n16147, n16148, n16149, n16150, n16151, n16152, n16153,
         n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161,
         n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169,
         n16170, n16171, n16172, n16173, n16174, n16175, n16176, n16177,
         n16178, n16179, n16180, n16181, n16182, n16183, n16184, n16185,
         n16186, n16187, n16188, n16189, n16190, n16191, n16192, n16193,
         n16194, n16195, n16196, n16197, n16198, n16199, n16200, n16201,
         n16202, n16203, n16204, n16205, n16206, n16207, n16208, n16209,
         n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217,
         n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225,
         n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233,
         n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241,
         n16242, n16243, n16244, n16245, n16246, n16247, n16248, n16249,
         n16250, n16251, n16252, n16253, n16254, n16255, n16256, n16257,
         n16258, n16259, n16260, n16261, n16262, n16263, n16264, n16265,
         n16266, n16267, n16268, n16269, n16270, n16271, n16272, n16273,
         n16274, n16275, n16276, n16277, n16278, n16279, n16280, n16281,
         n16282, n16283, n16284, n16285, n16286, n16287, n16288, n16289,
         n16290, n16291, n16292, n16293, n16294, n16295, n16296, n16297,
         n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305,
         n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313,
         n16314, n16315, n16316, n16317, n16318, n16319, n16320, n16321,
         n16322, n16323, n16324, n16325, n16326, n16327, n16328, n16329,
         n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337,
         n16338, n16339, n16340, n16341, n16342, n16343, n16344, n16345,
         n16346, n16347, n16348, n16349, n16350, n16351, n16352, n16353,
         n16354, n16355, n16356, n16357, n16358, n16359, n16360, n16361,
         n16362, n16363, n16364, n16365, n16366, n16367, n16368, n16369,
         n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377,
         n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385,
         n16386, n16387, n16388, n16389, n16390, n16391, n16392, n16393,
         n16394, n16395, n16396, n16397, n16398, n16399, n16400, n16401,
         n16402, n16403, n16404, n16405, n16406, n16407, n16408, n16409,
         n16410, n16411, n16412, n16413, n16414, n16415, n16416, n16417,
         n16418, n16419, n16420, n16421, n16422, n16423, n16424, n16425,
         n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433,
         n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441,
         n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449,
         n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457,
         n16458, n16459, n16460, n16461, n16462, n16463, n16464, n16465,
         n16466, n16467, n16468, n16469, n16470, n16471, n16472, n16473,
         n16474, n16475, n16476, n16477, n16478, n16479, n16480, n16481,
         n16482, n16483, n16484, n16485, n16486, n16487, n16488, n16489,
         n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497,
         n16498, n16499, n16500, n16501, n16502, n16503, n16504, n16505,
         n16506, n16507, n16508, n16509, n16510, n16511, n16512, n16513,
         n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521,
         n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529,
         n16530, n16531, n16532, n16533, n16534, n16535, n16536, n16537,
         n16538, n16539, n16540, n16541, n16542, n16543, n16544, n16545,
         n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553,
         n16554, n16555, n16556, n16557, n16558, n16559, n16560, n16561,
         n16562, n16563, n16564, n16565, n16566, n16567, n16568, n16569,
         n16570, n16571, n16572, n16573, n16574, n16575, n16576, n16577,
         n16578, n16579, n16580, n16581, n16582, n16583, n16584, n16585,
         n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593,
         n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601,
         n16602, n16603, n16604, n16605, n16606, n16607, n16608, n16609,
         n16610, n16611, n16612, n16613, n16614, n16615, n16616, n16617,
         n16618, n16619, n16620, n16621, n16622, n16623, n16624, n16625,
         n16626, n16627, n16628, n16629, n16630, n16631, n16632, n16633,
         n16634, n16635, n16636, n16637, n16638, n16639, n16640, n16641,
         n16642, n16643, n16644, n16645, n16646, n16647, n16648, n16649,
         n16650, n16651, n16652, n16653, n16654, n16655, n16656, n16657,
         n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665,
         n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673,
         n16674, n16675, n16676, n16677, n16678, n16679, n16680, n16681,
         n16682, n16683, n16684, n16685, n16686, n16687, n16688, n16689,
         n16690, n16691, n16692, n16693, n16694, n16695, n16696, n16697,
         n16698, n16699, n16700, n16701, n16702, n16703, n16704, n16705,
         n16706, n16707, n16708, n16709, n16710, n16711, n16712, n16713,
         n16714, n16715, n16716, n16717, n16718, n16719, n16720, n16721,
         n16722, n16723, n16724, n16725, n16726, n16727, n16728, n16729,
         n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737,
         n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745,
         n16746, n16747, n16748, n16749, n16750, n16751, n16752, n16753,
         n16754, n16755, n16756, n16757, n16758, n16759, n16760, n16761,
         n16762, n16763, n16764, n16765, n16766, n16767, n16768, n16769,
         n16770, n16771, n16772, n16773, n16774, n16775, n16776, n16777,
         n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785,
         n16786, n16787, n16788, n16789, n16790, n16791, n16792, n16793,
         n16794, n16795, n16796, n16797, n16798, n16799, n16800, n16801,
         n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809,
         n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817,
         n16818, n16819, n16820, n16821, n16822, n16823, n16824, n16825,
         n16826, n16827, n16828, n16829, n16830, n16831, n16832, n16833,
         n16834, n16835, n16836, n16837, n16838, n16839, n16840, n16841,
         n16842, n16843, n16844, n16845, n16846, n16847, n16848, n16849,
         n16850, n16851, n16852, n16853, n16854, n16855, n16856, n16857,
         n16858, n16859, n16860, n16861, n16862, n16863, n16864, n16865,
         n16866, n16867, n16868, n16869, n16870, n16871, n16872, n16873,
         n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881,
         n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889,
         n16890, n16891, n16892, n16893, n16894, n16895, n16896, n16897,
         n16898, n16899, n16900, n16901, n16902, n16903, n16904, n16905,
         n16906, n16907, n16908, n16909, n16910, n16911, n16912, n16913,
         n16914, n16915, n16916, n16917, n16918, n16919, n16920, n16921,
         n16922, n16923, n16924, n16925, n16926, n16927, n16928, n16929,
         n16930, n16931, n16932, n16933, n16934, n16935, n16936, n16937,
         n16938, n16939, n16940, n16941, n16942, n16943, n16944, n16945,
         n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953,
         n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961,
         n16962, n16963, n16964, n16965, n16966, n16967, n16968, n16969,
         n16970, n16971, n16972, n16973, n16974, n16975, n16976, n16977,
         n16978, n16979, n16980, n16981, n16982, n16983, n16984, n16985,
         n16986, n16987, n16988, n16989, n16990, n16991, n16992, n16993,
         n16994, n16995, n16996, n16997, n16998, n16999, n17000, n17001,
         n17002, n17003, n17004, n17005, n17006, n17007, n17008, n17009,
         n17010, n17011, n17012, n17013, n17014, n17015, n17016, n17017,
         n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025,
         n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033,
         n17034, n17035, n17036, n17037, n17038, n17039, n17040, n17041,
         n17042, n17043, n17044, n17045, n17046, n17047, n17048, n17049,
         n17050, n17051, n17052, n17053, n17054, n17055, n17056, n17057,
         n17058, n17059, n17060, n17061, n17062, n17063, n17064, n17065,
         n17066, n17067, n17068, n17069, n17070, n17071, n17072, n17073,
         n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17081,
         n17082, n17083, n17084, n17085, n17086, n17087, n17088, n17089,
         n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097,
         n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105,
         n17106, n17107, n17108, n17109, n17110, n17111, n17112, n17113,
         n17114, n17115, n17116, n17117, n17118, n17119, n17120, n17121,
         n17122, n17123, n17124, n17125, n17126, n17127, n17128, n17129,
         n17130, n17131, n17132, n17133, n17134, n17135, n17136, n17137,
         n17138, n17139, n17140, n17141, n17142, n17143, n17144, n17145,
         n17146, n17147, n17148, n17149, n17150, n17151, n17152, n17153,
         n17154, n17155, n17156, n17157, n17158, n17159, n17160, n17161,
         n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169,
         n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177,
         n17178, n17179, n17180, n17181, n17182, n17183, n17184, n17185,
         n17186, n17187, n17188, n17189, n17190, n17191, n17192, n17193,
         n17194, n17195, n17196, n17197, n17198, n17199, n17200, n17201,
         n17202, n17203, n17204, n17205, n17206, n17207, n17208, n17209,
         n17210, n17211, n17212, n17213, n17214, n17215, n17216, n17217,
         n17218, n17219, n17220, n17221, n17222, n17223, n17224, n17225,
         n17226, n17227, n17228, n17229, n17230, n17231, n17232, n17233,
         n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241,
         n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249,
         n17250, n17251, n17252, n17253, n17254, n17255, n17256, n17257,
         n17258, n17259, n17260, n17261, n17262, n17263, n17264, n17265,
         n17266, n17267, n17268, n17269, n17270, n17271, n17272, n17273,
         n17274, n17275, n17276, n17277, n17278, n17279, n17280, n17281,
         n17282, n17283, n17284, n17285, n17286, n17287, n17288, n17289,
         n17290, n17291, n17292, n17293, n17294, n17295, n17296, n17297,
         n17298, n17299, n17300, n17301, n17302, n17303, n17304, n17305,
         n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313,
         n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321,
         n17322, n17323, n17324, n17325, n17326, n17327, n17328, n17329,
         n17330, n17331, n17332, n17333, n17334, n17335, n17336, n17337,
         n17338, n17339, n17340, n17341, n17342, n17343, n17344, n17345,
         n17346, n17347, n17348, n17349, n17350, n17351, n17352, n17353,
         n17354, n17355, n17356, n17357, n17358, n17359, n17360, n17361,
         n17362, n17363, n17364, n17365, n17366, n17367, n17368, n17369,
         n17370, n17371, n17372, n17373, n17374, n17375, n17376, n17377,
         n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385,
         n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393,
         n17394, n17395, n17396, n17397, n17398, n17399, n17400, n17401,
         n17402, n17403, n17404, n17405, n17406, n17407, n17408, n17409,
         n17410, n17411, n17412, n17413, n17414, n17415, n17416, n17417,
         n17418, n17419, n17420, n17421, n17422, n17423, n17424, n17425,
         n17426, n17427, n17428, n17429, n17430, n17431, n17432, n17433,
         n17434, n17435, n17436, n17437, n17438, n17439, n17440, n17441,
         n17442, n17443, n17444, n17445, n17446, n17447, n17448, n17449,
         n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457,
         n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465,
         n17466, n17467, n17468, n17469, n17470, n17471, n17472, n17473,
         n17474, n17475, n17476, n17477, n17478, n17479, n17480, n17481,
         n17482, n17483, n17484, n17485, n17486, n17487, n17488, n17489,
         n17490, n17491, n17492, n17493, n17494, n17495, n17496, n17497,
         n17498, n17499, n17500, n17501, n17502, n17503, n17504, n17505,
         n17506, n17507, n17508, n17509, n17510, n17511, n17512, n17513,
         n17514, n17515, n17516, n17517, n17518, n17519, n17520, n17521,
         n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529,
         n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537,
         n17538, n17539, n17540, n17541, n17542, n17543, n17544, n17545,
         n17546, n17547, n17548, n17549, n17550, n17551, n17552, n17553,
         n17554, n17555, n17556, n17557, n17558, n17559, n17560, n17561,
         n17562, n17563, n17564, n17565, n17566, n17567, n17568, n17569,
         n17570, n17571, n17572, n17573, n17574, n17575, n17576, n17577,
         n17578, n17579, n17580, n17581, n17582, n17583, n17584, n17585,
         n17586, n17587, n17588, n17589, n17590, n17591, n17592, n17593,
         n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601,
         n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609,
         n17610, n17611, n17612, n17613, n17614, n17615, n17616, n17617,
         n17618, n17619, n17620, n17621, n17622, n17623, n17624, n17625,
         n17626, n17627, n17628, n17629, n17630, n17631, n17632, n17633,
         n17634, n17635, n17636, n17637, n17638, n17639, n17640, n17641,
         n17642, n17643, n17644, n17645, n17646, n17647, n17648, n17649,
         n17650, n17651, n17652, n17653, n17654, n17655, n17656, n17657,
         n17658, n17659, n17660, n17661, n17662, n17663, n17664, n17665,
         n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673,
         n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681,
         n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689,
         n17690, n17691, n17692, n17693, n17694, n17695, n17696, n17697,
         n17698, n17699, n17700, n17701, n17702, n17703, n17704, n17705,
         n17706, n17707, n17708, n17709, n17710, n17711, n17712, n17713,
         n17714, n17715, n17716, n17717, n17718, n17719, n17720, n17721,
         n17722, n17723, n17724, n17725, n17726, n17727, n17728, n17729,
         n17730, n17731, n17732, n17733, n17734, n17735, n17736, n17737,
         n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745,
         n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753,
         n17754, n17755, n17756, n17757, n17758, n17759, n17760, n17761,
         n17762, n17763, n17764, n17765, n17766, n17767, n17768, n17769,
         n17770, n17771, n17772, n17773, n17774, n17775, n17776, n17777,
         n17778, n17779, n17780, n17781, n17782, n17783, n17784, n17785,
         n17786, n17787, n17788, n17789, n17790, n17791, n17792, n17793,
         n17794, n17795, n17796, n17797, n17798, n17799, n17800, n17801,
         n17802, n17803, n17804, n17805, n17806, n17807, n17808, n17809,
         n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817,
         n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825,
         n17826, n17827, n17828, n17829, n17830, n17831, n17832, n17833,
         n17834, n17835, n17836, n17837, n17838, n17839, n17840, n17841,
         n17842, n17843, n17844, n17845, n17846, n17847, n17848, n17849,
         n17850, n17851, n17852, n17853, n17854, n17855, n17856, n17857,
         n17858, n17859, n17860, n17861, n17862, n17863, n17864, n17865,
         n17866, n17867, n17868, n17869, n17870, n17871, n17872, n17873,
         n17874, n17875, n17876, n17877, n17878, n17879, n17880, n17881,
         n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889,
         n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897,
         n17898, n17899, n17900, n17901, n17902, n17903, n17904, n17905,
         n17906, n17907, n17908, n17909, n17910, n17911, n17912, n17913,
         n17914, n17915, n17916, n17917, n17918, n17919, n17920, n17921,
         n17922, n17923, n17924, n17925, n17926, n17927, n17928, n17929,
         n17930, n17931, n17932, n17933, n17934, n17935, n17936, n17937,
         n17938, n17939, n17940, n17941, n17942, n17943, n17944, n17945,
         n17946, n17947, n17948, n17949, n17950, n17951, n17952, n17953,
         n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961,
         n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969,
         n17970, n17971, n17972, n17973, n17974, n17975, n17976, n17977,
         n17978, n17979, n17980, n17981, n17982, n17983, n17984, n17985,
         n17986, n17987, n17988, n17989, n17990, n17991, n17992, n17993,
         n17994, n17995, n17996, n17997, n17998, n17999, n18000, n18001,
         n18002, n18003, n18004, n18005, n18006, n18007, n18008, n18009,
         n18010, n18011, n18012, n18013, n18014, n18015, n18016, n18017,
         n18018, n18019, n18020, n18021, n18022, n18023, n18024, n18025,
         n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033,
         n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041,
         n18042, n18043, n18044, n18045, n18046, n18047, n18048, n18049,
         n18050, n18051, n18052, n18053, n18054, n18055, n18056, n18057,
         n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065,
         n18066, n18067, n18068, n18069, n18070, n18071, n18072, n18073,
         n18074, n18075, n18076, n18077, n18078, n18079, n18080, n18081,
         n18082, n18083, n18084, n18085, n18086, n18087, n18088, n18089,
         n18090, n18091, n18092, n18093, n18094, n18095, n18096, n18097,
         n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105,
         n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113,
         n18114, n18115, n18116, n18117, n18118, n18119, n18120, n18121,
         n18122, n18123, n18124, n18125, n18126, n18127, n18128, n18129,
         n18130, n18131, n18132, n18133, n18134, n18135, n18136, n18137,
         n18138, n18139, n18140, n18141, n18142, n18143, n18144, n18145,
         n18146, n18147, n18148, n18149, n18150, n18151, n18152, n18153,
         n18154, n18155, n18156, n18157, n18158, n18159, n18160, n18161,
         n18162, n18163, n18164, n18165, n18166, n18167, n18168, n18169,
         n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177,
         n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185,
         n18186, n18187, n18188, n18189, n18190, n18191, n18192, n18193,
         n18194, n18195, n18196, n18197, n18198, n18199, n18200, n18201,
         n18202, n18203, n18204, n18205, n18206, n18207, n18208, n18209,
         n18210, n18211, n18212, n18213, n18214, n18215, n18216, n18217,
         n18218, n18219, n18220, n18221, n18222, n18223, n18224, n18225,
         n18226, n18227, n18228, n18229, n18230, n18231, n18232, n18233,
         n18234, n18235, n18236, n18237, n18238, n18239, n18240, n18241,
         n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249,
         n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257,
         n18258, n18259, n18260, n18261, n18262, n18263, n18264, n18265,
         n18266, n18267, n18268, n18269, n18270, n18271, n18272, n18273,
         n18274, n18275, n18276, n18277, n18278, n18279, n18280, n18281,
         n18282, n18283, n18284, n18285, n18286, n18287, n18288, n18289,
         n18290, n18291, n18292, n18293, n18294, n18295, n18296, n18297,
         n18298, n18299, n18300, n18301, n18302, n18303, n18304, n18305,
         n18306, n18307, n18308, n18309, n18310, n18311, n18312, n18313,
         n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321,
         n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329,
         n18330, n18331, n18332, n18333, n18334, n18335, n18336, n18337,
         n18338, n18339, n18340, n18341, n18342, n18343, n18344, n18345,
         n18346, n18347, n18348, n18349, n18350, n18351, n18352, n18353,
         n18354, n18355, n18356, n18357, n18358, n18359, n18360, n18361,
         n18362, n18363, n18364, n18365, n18366, n18367, n18368, n18369,
         n18370, n18371, n18372, n18373, n18374, n18375, n18376, n18377,
         n18378, n18379, n18380, n18381, n18382, n18383, n18384, n18385,
         n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393,
         n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401,
         n18402, n18403, n18404, n18405, n18406, n18407, n18408, n18409,
         n18410, n18411, n18412, n18413, n18414, n18415, n18416, n18417,
         n18418, n18419, n18420, n18421, n18422, n18423, n18424, n18425,
         n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433,
         n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441,
         n18442, n18443, n18444, n18445, n18446, n18447, n18448, n18449,
         n18450, n18451, n18452, n18453, n18454, n18455, n18456, n18457,
         n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465,
         n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473,
         n18474, n18475, n18476, n18477, n18478, n18479, n18480, n18481,
         n18482, n18483, n18484, n18485, n18486, n18487, n18488, n18489,
         n18490, n18491, n18492, n18493, n18494, n18495, n18496, n18497,
         n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505,
         n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513,
         n18514, n18515, n18516, n18517, n18518, n18519, n18520, n18521,
         n18522, n18523, n18524, n18525, n18526, n18527, n18528, n18529,
         n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537,
         n18538, n18539, n18540, n18541, n18542, n18543, n18544, n18545,
         n18546, n18547, n18548, n18549, n18550, n18551, n18552, n18553,
         n18554, n18555, n18556, n18557, n18558, n18559, n18560, n18561,
         n18562, n18563, n18564, n18565, n18566, n18567, n18568, n18569,
         n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577,
         n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585,
         n18586, n18587, n18588, n18589, n18590, n18591, n18592, n18593,
         n18594, n18595, n18596, n18597, n18598, n18599, n18600, n18601,
         n18602, n18603, n18604, n18605, n18606, n18607, n18608, n18609,
         n18610, n18611, n18612, n18613, n18614, n18615, n18616, n18617,
         n18618, n18619, n18620, n18621, n18622, n18623, n18624, n18625,
         n18626, n18627, n18628, n18629, n18630, n18631, n18632, n18633,
         n18634, n18635, n18636, n18637, n18638, n18639, n18640, n18641,
         n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649,
         n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657,
         n18658, n18659, n18660, n18661, n18662, n18663, n18664, n18665,
         n18666, n18667, n18668, n18669, n18670, n18671, n18672, n18673,
         n18674, n18675, n18676, n18677, n18678, n18679, n18680, n18681,
         n18682, n18683, n18684, n18685, n18686, n18687, n18688, n18689,
         n18690, n18691, n18692, n18693, n18694, n18695, n18696, n18697,
         n18698, n18699, n18700, n18701, n18702, n18703, n18704, n18705,
         n18706, n18707, n18708, n18709, n18710, n18711, n18712, n18713,
         n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721,
         n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729,
         n18730, n18731, n18732, n18733, n18734, n18735, n18736, n18737,
         n18738, n18739, n18740, n18741, n18742, n18743, n18744, n18745,
         n18746, n18747, n18748, n18749, n18750, n18751, n18752, n18753,
         n18754, n18755, n18756, n18757, n18758, n18759, n18760, n18761,
         n18762, n18763, n18764, n18765, n18766, n18767, n18768, n18769,
         n18770, n18771, n18772, n18773, n18774, n18775, n18776, n18777,
         n18778, n18779, n18780, n18781, n18782, n18783, n18784, n18785,
         n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793,
         n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801,
         n18802, n18803, n18804, n18805, n18806, n18807, n18808, n18809,
         n18810, n18811, n18812, n18813, n18814, n18815, n18816, n18817,
         n18818, n18819, n18820, n18821, n18822, n18823, n18824, n18825,
         n18826, n18827, n18828, n18829, n18830, n18831, n18832, n18833,
         n18834, n18835, n18836, n18837, n18838, n18839, n18840, n18841,
         n18842, n18843, n18844, n18845, n18846, n18847, n18848, n18849,
         n18850, n18851, n18852, n18853, n18854, n18855, n18856, n18857,
         n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865,
         n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873,
         n18874, n18875, n18876, n18877, n18878, n18879, n18880, n18881,
         n18882, n18883, n18884, n18885, n18886, n18887, n18888, n18889,
         n18890, n18891, n18892, n18893, n18894, n18895, n18896, n18897,
         n18898, n18899, n18900, n18901, n18902, n18903, n18904, n18905,
         n18906, n18907, n18908, n18909, n18910, n18911, n18912, n18913,
         n18914, n18915, n18916, n18917, n18918, n18919, n18920, n18921,
         n18922, n18923, n18924, n18925, n18926, n18927, n18928, n18929,
         n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937,
         n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945,
         n18946, n18947, n18948, n18949, n18950, n18951, n18952, n18953,
         n18954, n18955, n18956, n18957, n18958, n18959, n18960, n18961,
         n18962, n18963, n18964, n18965, n18966, n18967, n18968, n18969,
         n18970, n18971, n18972, n18973, n18974, n18975, n18976, n18977,
         n18978, n18979, n18980, n18981, n18982, n18983, n18984, n18985,
         n18986, n18987, n18988, n18989, n18990, n18991, n18992, n18993,
         n18994, n18995, n18996, n18997, n18998, n18999, n19000, n19001,
         n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009,
         n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017,
         n19018, n19019, n19020, n19021, n19022, n19023, n19024, n19025,
         n19026, n19027, n19028, n19029, n19030, n19031, n19032, n19033,
         n19034, n19035, n19036, n19037, n19038, n19039, n19040, n19041,
         n19042, n19043, n19044, n19045, n19046, n19047, n19048, n19049,
         n19050, n19051, n19052, n19053, n19054, n19055, n19056, n19057,
         n19058, n19059, n19060, n19061, n19062, n19063, n19064, n19065,
         n19066, n19067, n19068, n19069, n19070, n19071, n19072, n19073,
         n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081,
         n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089,
         n19090, n19091, n19092, n19093, n19094, n19095, n19096, n19097,
         n19098, n19099, n19100, n19101, n19102, n19103, n19104, n19105,
         n19106, n19107, n19108, n19109, n19110, n19111, n19112, n19113,
         n19114, n19115, n19116, n19117, n19118, n19119, n19120, n19121,
         n19122, n19123, n19124, n19125, n19126, n19127, n19128, n19129,
         n19130, n19131, n19132, n19133, n19134, n19135, n19136, n19137,
         n19138, n19139, n19140, n19141, n19142, n19143, n19144, n19145,
         n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153,
         n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161,
         n19162, n19163, n19164, n19165, n19166, n19167, n19168, n19169,
         n19170, n19171, n19172, n19173, n19174, n19175, n19176, n19177,
         n19178, n19179, n19180, n19181, n19182, n19183, n19184, n19185,
         n19186, n19187, n19188, n19189, n19190, n19191, n19192, n19193,
         n19194, n19195, n19196, n19197, n19198, n19199, n19200, n19201,
         n19202, n19203, n19204, n19205, n19206, n19207, n19208, n19209,
         n19210, n19211, n19212, n19213, n19214, n19215, n19216, n19217,
         n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225,
         n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233,
         n19234, n19235, n19236, n19237, n19238, n19239, n19240, n19241,
         n19242, n19243, n19244, n19245, n19246, n19247, n19248, n19249,
         n19250, n19251, n19252, n19253, n19254, n19255, n19256, n19257,
         n19258, n19259, n19260, n19261, n19262, n19263, n19264, n19265,
         n19266, n19267, n19268, n19269, n19270, n19271, n19272, n19273,
         n19274, n19275, n19276, n19277, n19278, n19279, n19280, n19281,
         n19282, n19283, n19284, n19285, n19286, n19287, n19288, n19289,
         n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297,
         n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305,
         n19306, n19307, n19308, n19309, n19310, n19311, n19312, n19313,
         n19314, n19315, n19316, n19317, n19318, n19319, n19320, n19321,
         n19322, n19323, n19324, n19325, n19326, n19327, n19328, n19329,
         n19330, n19331, n19332, n19333, n19334, n19335, n19336, n19337,
         n19338, n19339, n19340, n19341, n19342, n19343, n19344, n19345,
         n19346, n19347, n19348, n19349, n19350, n19351, n19352, n19353,
         n19354, n19355, n19356, n19357, n19358, n19359, n19360, n19361,
         n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369,
         n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377,
         n19378, n19379, n19380, n19381, n19382, n19383, n19384, n19385,
         n19386, n19387, n19388, n19389, n19390, n19391, n19392, n19393,
         n19394, n19395, n19396, n19397, n19398, n19399, n19400, n19401,
         n19402, n19403, n19404, n19405, n19406, n19407, n19408, n19409,
         n19410, n19411, n19412, n19413, n19414, n19415, n19416, n19417,
         n19418, n19419, n19420, n19421, n19422, n19423, n19424, n19425,
         n19426, n19427, n19428, n19429, n19430, n19431, n19432, n19433,
         n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441,
         n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449,
         n19450, n19451, n19452, n19453, n19454, n19455, n19456, n19457,
         n19458, n19459, n19460, n19461, n19462, n19463, n19464, n19465,
         n19466, n19467, n19468, n19469, n19470, n19471, n19472, n19473,
         n19474, n19475, n19476, n19477, n19478, n19479, n19480, n19481,
         n19482, n19483, n19484, n19485, n19486, n19487, n19488, n19489,
         n19490, n19491, n19492, n19493, n19494, n19495, n19496, n19497,
         n19498, n19499, n19500, n19501, n19502, n19503, n19504, n19505,
         n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513,
         n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521,
         n19522, n19523, n19524, n19525, n19526, n19527, n19528, n19529,
         n19530, n19531, n19532, n19533, n19534, n19535, n19536, n19537,
         n19538, n19539, n19540, n19541, n19542, n19543, n19544, n19545,
         n19546, n19547, n19548, n19549, n19550, n19551, n19552, n19553,
         n19554, n19555, n19556, n19557, n19558, n19559, n19560, n19561,
         n19562, n19563, n19564, n19565, n19566, n19567, n19568, n19569,
         n19570, n19571, n19572, n19573, n19574, n19575, n19576, n19577,
         n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585,
         n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593,
         n19594, n19595, n19596, n19597, n19598, n19599, n19600, n19601,
         n19602, n19603, n19604, n19605, n19606, n19607, n19608, n19609,
         n19610, n19611, n19612, n19613, n19614, n19615, n19616, n19617,
         n19618, n19619, n19620, n19621, n19622, n19623, n19624, n19625,
         n19626, n19627, n19628, n19629, n19630, n19631, n19632, n19633,
         n19634, n19635, n19636, n19637, n19638, n19639, n19640, n19641,
         n19642, n19643, n19644, n19645, n19646, n19647, n19648, n19649,
         n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657,
         n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665,
         n19666, n19667, n19668, n19669, n19670, n19671, n19672, n19673,
         n19674, n19675, n19676, n19677, n19678, n19679, n19680, n19681,
         n19682, n19683, n19684, n19685, n19686, n19687, n19688, n19689,
         n19690, n19691, n19692, n19693, n19694, n19695, n19696, n19697,
         n19698, n19699, n19700, n19701, n19702, n19703, n19704, n19705,
         n19706, n19707, n19708, n19709, n19710, n19711, n19712, n19713,
         n19714, n19715, n19716, n19717, n19718, n19719, n19720, n19721,
         n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729,
         n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737,
         n19738, n19739, n19740, n19741, n19742, n19743, n19744, n19745,
         n19746, n19747, n19748, n19749, n19750, n19751, n19752, n19753,
         n19754, n19755, n19756, n19757, n19758, n19759, n19760, n19761,
         n19762, n19763, n19764, n19765, n19766, n19767, n19768, n19769,
         n19770, n19771, n19772, n19773, n19774, n19775, n19776, n19777,
         n19778, n19779, n19780, n19781, n19782, n19783, n19784, n19785,
         n19786, n19787, n19788, n19789, n19790, n19791, n19792, n19793,
         n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801,
         n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809,
         n19810, n19811, n19812, n19813, n19814, n19815, n19816, n19817,
         n19818, n19819, n19820, n19821, n19822, n19823, n19824, n19825,
         n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833,
         n19834, n19835, n19836, n19837, n19838, n19839, n19840, n19841,
         n19842, n19843, n19844, n19845, n19846, n19847, n19848, n19849,
         n19850, n19851, n19852, n19853, n19854, n19855, n19856, n19857,
         n19858, n19859, n19860, n19861, n19862, n19863, n19864, n19865,
         n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873,
         n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881,
         n19882, n19883, n19884, n19885, n19886, n19887, n19888, n19889,
         n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897,
         n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905,
         n19906, n19907, n19908, n19909, n19910, n19911, n19912, n19913,
         n19914, n19915, n19916, n19917, n19918, n19919, n19920, n19921,
         n19922, n19923, n19924, n19925, n19926, n19927, n19928, n19929,
         n19930, n19931, n19932, n19933, n19934, n19935, n19936, n19937,
         n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945,
         n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953,
         n19954, n19955, n19956, n19957, n19958, n19959, n19960, n19961,
         n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969,
         n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977,
         n19978, n19979, n19980, n19981, n19982, n19983, n19984, n19985,
         n19986, n19987, n19988, n19989, n19990, n19991, n19992, n19993,
         n19994, n19995, n19996, n19997, n19998, n19999, n20000, n20001,
         n20002, n20003, n20004, n20005, n20006, n20007, n20008, n20009,
         n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017,
         n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025,
         n20026, n20027, n20028, n20029, n20030, n20031, n20032, n20033,
         n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041,
         n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049,
         n20050, n20051, n20052, n20053, n20054, n20055, n20056, n20057,
         n20058, n20059, n20060, n20061, n20062, n20063, n20064, n20065,
         n20066, n20067, n20068, n20069, n20070, n20071, n20072, n20073,
         n20074, n20075, n20076, n20077, n20078, n20079, n20080, n20081,
         n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089,
         n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097,
         n20098, n20099, n20100, n20101, n20102, n20103, n20104, n20105,
         n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113,
         n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121,
         n20122, n20123, n20124, n20125, n20126, n20127, n20128, n20129,
         n20130, n20131, n20132, n20133, n20134, n20135, n20136, n20137,
         n20138, n20139, n20140, n20141, n20142, n20143, n20144, n20145,
         n20146, n20147, n20148, n20149, n20150, n20151, n20152, n20153,
         n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161,
         n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169,
         n20170, n20171, n20172, n20173, n20174, n20175, n20176, n20177,
         n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185,
         n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193,
         n20194, n20195, n20196, n20197, n20198, n20199, n20200, n20201,
         n20202, n20203, n20204, n20205, n20206, n20207, n20208, n20209,
         n20210, n20211, n20212, n20213, n20214, n20215, n20216, n20217,
         n20218, n20219, n20220, n20221, n20222, n20223, n20224, n20225,
         n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233,
         n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241,
         n20242, n20243, n20244, n20245, n20246, n20247, n20248, n20249,
         n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257,
         n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265,
         n20266, n20267, n20268, n20269, n20270, n20271, n20272, n20273,
         n20274, n20275, n20276, n20277, n20278, n20279, n20280, n20281,
         n20282, n20283, n20284, n20285, n20286, n20287, n20288, n20289,
         n20290, n20291, n20292, n20293, n20294, n20295, n20296, n20297,
         n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305,
         n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313,
         n20314, n20315, n20316, n20317, n20318, n20319, n20320, n20321,
         n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329,
         n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337,
         n20338, n20339, n20340, n20341, n20342, n20343, n20344, n20345,
         n20346, n20347, n20348, n20349, n20350, n20351, n20352, n20353,
         n20354, n20355, n20356, n20357, n20358, n20359, n20360, n20361,
         n20362, n20363, n20364, n20365, n20366, n20367, n20368, n20369,
         n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377,
         n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385,
         n20386, n20387, n20388, n20389, n20390, n20391, n20392, n20393,
         n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401,
         n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409,
         n20410, n20411, n20412, n20413, n20414, n20415, n20416, n20417,
         n20418, n20419, n20420, n20421, n20422, n20423, n20424, n20425,
         n20426, n20427, n20428, n20429, n20430, n20431, n20432, n20433,
         n20434, n20435, n20436, n20437, n20438, n20439, n20440, n20441,
         n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449,
         n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457,
         n20458, n20459, n20460, n20461, n20462, n20463, n20464, n20465,
         n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473,
         n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481,
         n20482, n20483, n20484, n20485, n20486, n20487, n20488, n20489,
         n20490, n20491, n20492, n20493, n20494, n20495, n20496, n20497,
         n20498, n20499, n20500, n20501, n20502, n20503, n20504, n20505,
         n20506, n20507, n20508, n20509, n20510, n20511, n20512, n20513,
         n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521,
         n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529,
         n20530, n20531, n20532, n20533, n20534, n20535, n20536, n20537,
         n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545,
         n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553,
         n20554, n20555, n20556, n20557, n20558, n20559, n20560, n20561,
         n20562, n20563, n20564, n20565, n20566, n20567, n20568, n20569,
         n20570, n20571, n20572, n20573, n20574, n20575, n20576, n20577,
         n20578, n20579, n20580, n20581, n20582, n20583, n20584, n20585,
         n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593,
         n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601,
         n20602, n20603, n20604, n20605, n20606, n20607, n20608, n20609,
         n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617,
         n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625,
         n20626, n20627, n20628, n20629, n20630, n20631, n20632, n20633,
         n20634, n20635, n20636, n20637, n20638, n20639, n20640, n20641,
         n20642, n20643, n20644, n20645, n20646, n20647, n20648, n20649,
         n20650, n20651, n20652, n20653, n20654, n20655, n20656, n20657,
         n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665,
         n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673,
         n20674, n20675, n20676, n20677, n20678, n20679, n20680, n20681,
         n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689,
         n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697,
         n20698, n20699, n20700, n20701, n20702, n20703, n20704, n20705,
         n20706, n20707, n20708, n20709, n20710, n20711, n20712, n20713,
         n20714, n20715, n20716, n20717, n20718, n20719, n20720, n20721,
         n20722, n20723, n20724, n20725, n20726, n20727, n20728, n20729,
         n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737,
         n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745,
         n20746, n20747, n20748, n20749, n20750, n20751, n20752, n20753,
         n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761,
         n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769,
         n20770, n20771, n20772, n20773, n20774, n20775, n20776, n20777,
         n20778, n20779, n20780, n20781, n20782, n20783, n20784, n20785,
         n20786, n20787, n20788, n20789, n20790, n20791, n20792, n20793,
         n20794, n20795, n20796, n20797, n20798, n20799, n20800, n20801,
         n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809,
         n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817,
         n20818, n20819, n20820, n20821, n20822, n20823, n20824, n20825,
         n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833,
         n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841,
         n20842, n20843, n20844, n20845, n20846, n20847, n20848, n20849,
         n20850, n20851, n20852, n20853, n20854, n20855, n20856, n20857,
         n20858, n20859, n20860, n20861, n20862, n20863, n20864, n20865,
         n20866, n20867, n20868, n20869, n20870, n20871, n20872, n20873,
         n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881,
         n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889,
         n20890, n20891, n20892, n20893, n20894, n20895, n20896, n20897,
         n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905,
         n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913,
         n20914, n20915, n20916, n20917, n20918, n20919, n20920, n20921,
         n20922, n20923, n20924, n20925, n20926, n20927, n20928, n20929,
         n20930, n20931, n20932, n20933, n20934, n20935, n20936, n20937,
         n20938, n20939, n20940, n20941, n20942, n20943, n20944, n20945,
         n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953,
         n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961,
         n20962, n20963, n20964, n20965, n20966, n20967, n20968, n20969,
         n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977,
         n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985,
         n20986, n20987, n20988, n20989, n20990, n20991, n20992, n20993,
         n20994, n20995, n20996, n20997, n20998, n20999, n21000, n21001,
         n21002, n21003, n21004, n21005, n21006, n21007, n21008, n21009,
         n21010, n21011, n21012, n21013, n21014, n21015, n21016, n21017,
         n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025,
         n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033,
         n21034, n21035, n21036, n21037, n21038, n21039, n21040, n21041,
         n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049,
         n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057,
         n21058, n21059, n21060, n21061, n21062, n21063, n21064, n21065,
         n21066, n21067, n21068, n21069, n21070, n21071, n21072, n21073,
         n21074, n21075, n21076, n21077, n21078, n21079, n21080, n21081,
         n21082, n21083, n21084, n21085, n21086, n21087, n21088, n21089,
         n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097,
         n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105,
         n21106, n21107, n21108, n21109, n21110, n21111, n21112, n21113,
         n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121,
         n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129,
         n21130, n21131, n21132, n21133, n21134, n21135, n21136, n21137,
         n21138, n21139, n21140, n21141, n21142, n21143, n21144, n21145,
         n21146, n21147, n21148, n21149, n21150, n21151, n21152, n21153,
         n21154, n21155, n21156, n21157, n21158, n21159, n21160, n21161,
         n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169,
         n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177,
         n21178, n21179, n21180, n21181, n21182, n21183, n21184, n21185,
         n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193,
         n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201,
         n21202, n21203, n21204, n21205, n21206, n21207, n21208, n21209,
         n21210, n21211, n21212, n21213, n21214, n21215, n21216, n21217,
         n21218, n21219, n21220, n21221, n21222, n21223, n21224, n21225,
         n21226, n21227, n21228, n21229, n21230, n21231, n21232, n21233,
         n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241,
         n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249,
         n21250, n21251, n21252, n21253, n21254, n21255, n21256, n21257,
         n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265,
         n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273,
         n21274, n21275, n21276, n21277, n21278, n21279, n21280, n21281,
         n21282, n21283, n21284, n21285, n21286, n21287, n21288, n21289,
         n21290, n21291, n21292, n21293, n21294, n21295, n21296, n21297,
         n21298, n21299, n21300, n21301, n21302, n21303, n21304, n21305,
         n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313,
         n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321,
         n21322, n21323, n21324, n21325, n21326, n21327, n21328, n21329,
         n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337,
         n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345,
         n21346, n21347, n21348, n21349, n21350, n21351, n21352, n21353,
         n21354, n21355, n21356, n21357, n21358, n21359, n21360, n21361,
         n21362, n21363, n21364, n21365, n21366, n21367, n21368, n21369,
         n21370, n21371, n21372, n21373, n21374, n21375, n21376, n21377,
         n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385,
         n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393,
         n21394, n21395, n21396, n21397, n21398, n21399, n21400, n21401,
         n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409,
         n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417,
         n21418, n21419, n21420, n21421, n21422, n21423, n21424, n21425,
         n21426, n21427, n21428, n21429, n21430, n21431, n21432, n21433,
         n21434, n21435, n21436, n21437, n21438, n21439, n21440, n21441,
         n21442, n21443, n21444, n21445, n21446, n21447, n21448, n21449,
         n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457,
         n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465,
         n21466, n21467, n21468, n21469, n21470, n21471, n21472, n21473,
         n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481,
         n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489,
         n21490, n21491, n21492, n21493, n21494, n21495, n21496, n21497,
         n21498, n21499, n21500, n21501, n21502, n21503, n21504, n21505,
         n21506, n21507, n21508, n21509, n21510, n21511, n21512, n21513,
         n21514, n21515, n21516, n21517, n21518, n21519, n21520, n21521,
         n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529,
         n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537,
         n21538, n21539, n21540, n21541, n21542, n21543, n21544, n21545,
         n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553,
         n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561,
         n21562, n21563, n21564, n21565, n21566, n21567, n21568, n21569,
         n21570, n21571, n21572, n21573, n21574, n21575, n21576, n21577,
         n21578, n21579, n21580, n21581, n21582, n21583, n21584, n21585,
         n21586, n21587, n21588, n21589, n21590, n21591, n21592, n21593,
         n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601,
         n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609,
         n21610, n21611, n21612, n21613, n21614, n21615, n21616, n21617,
         n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625,
         n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633,
         n21634, n21635, n21636, n21637, n21638, n21639, n21640, n21641,
         n21642, n21643, n21644, n21645, n21646, n21647, n21648, n21649,
         n21650, n21651, n21652, n21653, n21654, n21655, n21656, n21657,
         n21658, n21659, n21660, n21661, n21662, n21663, n21664, n21665,
         n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673,
         n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681,
         n21682, n21683, n21684, n21685, n21686, n21687, n21688, n21689,
         n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697,
         n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705,
         n21706, n21707, n21708, n21709, n21710, n21711, n21712, n21713,
         n21714, n21715, n21716, n21717, n21718, n21719, n21720, n21721,
         n21722, n21723, n21724, n21725, n21726, n21727, n21728, n21729,
         n21730, n21731, n21732, n21733, n21734, n21735, n21736, n21737,
         n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745,
         n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753,
         n21754, n21755, n21756, n21757, n21758, n21759, n21760, n21761,
         n21762, n21763, n21764, n21765, n21766, n21767, n21768, n21769,
         n21770, n21771, n21772, n21773, n21774, n21775, n21776, n21777,
         n21778, n21779, n21780, n21781, n21782, n21783, n21784, n21785,
         n21786, n21787, n21788, n21789, n21790, n21791, n21792, n21793,
         n21794, n21795, n21796, n21797, n21798, n21799, n21800, n21801,
         n21802, n21803, n21804, n21805, n21806, n21807, n21808, n21809,
         n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817,
         n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825,
         n21826, n21827, n21828, n21829, n21830, n21831, n21832, n21833,
         n21834, n21835, n21836, n21837, n21838, n21839, n21840, n21841,
         n21842, n21843, n21844, n21845, n21846, n21847, n21848, n21849,
         n21850, n21851, n21852, n21853, n21854, n21855, n21856, n21857,
         n21858, n21859, n21860, n21861, n21862, n21863, n21864, n21865,
         n21866, n21867, n21868, n21869, n21870, n21871, n21872, n21873,
         n21874, n21875, n21876, n21877, n21878, n21879, n21880, n21881,
         n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889,
         n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897,
         n21898, n21899, n21900, n21901, n21902, n21903, n21904, n21905,
         n21906, n21907, n21908, n21909, n21910, n21911, n21912, n21913,
         n21914, n21915, n21916, n21917, n21918, n21919, n21920, n21921,
         n21922, n21923, n21924, n21925, n21926, n21927, n21928, n21929,
         n21930, n21931, n21932, n21933, n21934, n21935, n21936, n21937,
         n21938, n21939, n21940, n21941, n21942, n21943, n21944, n21945,
         n21946, n21947, n21948, n21949, n21950, n21951, n21952, n21953,
         n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961,
         n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969,
         n21970, n21971, n21972, n21973, n21974, n21975, n21976, n21977,
         n21978, n21979, n21980, n21981, n21982, n21983, n21984, n21985,
         n21986, n21987, n21988, n21989, n21990, n21991, n21992, n21993,
         n21994, n21995, n21996, n21997, n21998, n21999, n22000, n22001,
         n22002, n22003, n22004, n22005, n22006, n22007, n22008, n22009,
         n22010, n22011, n22012, n22013, n22014, n22015, n22016, n22017,
         n22018, n22019, n22020, n22021, n22022, n22023, n22024, n22025,
         n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033,
         n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041,
         n22042, n22043, n22044, n22045, n22046, n22047, n22048, n22049,
         n22050, n22051, n22052, n22053, n22054, n22055, n22056, n22057,
         n22058, n22059, n22060, n22061, n22062, n22063, n22064, n22065,
         n22066, n22067, n22068, n22069, n22070, n22071, n22072, n22073,
         n22074, n22075, n22076, n22077, n22078, n22079, n22080, n22081,
         n22082, n22083, n22084, n22085, n22086, n22087, n22088, n22089,
         n22090, n22091, n22092, n22093, n22094, n22095, n22096, n22097,
         n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105,
         n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113,
         n22114, n22115, n22116, n22117, n22118, n22119, n22120, n22121,
         n22122, n22123, n22124, n22125, n22126, n22127, n22128, n22129,
         n22130, n22131, n22132, n22133, n22134, n22135, n22136, n22137,
         n22138, n22139, n22140, n22141, n22142, n22143, n22144, n22145,
         n22146, n22147, n22148, n22149, n22150, n22151, n22152, n22153,
         n22154, n22155, n22156, n22157, n22158, n22159, n22160, n22161,
         n22162, n22163, n22164, n22165, n22166, n22167, n22168, n22169,
         n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177,
         n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185,
         n22186, n22187, n22188, n22189, n22190, n22191, n22192, n22193,
         n22194, n22195, n22196, n22197, n22198, n22199, n22200, n22201,
         n22202, n22203, n22204, n22205, n22206, n22207, n22208, n22209,
         n22210, n22211, n22212, n22213, n22214, n22215, n22216, n22217,
         n22218, n22219, n22220, n22221, n22222, n22223, n22224, n22225,
         n22226, n22227, n22228, n22229, n22230, n22231, n22232, n22233,
         n22234, n22235, n22236, n22237, n22238, n22239, n22240, n22241,
         n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249,
         n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257,
         n22258, n22259, n22260, n22261, n22262, n22263, n22264, n22265,
         n22266, n22267, n22268, n22269, n22270, n22271, n22272, n22273,
         n22274, n22275, n22276, n22277, n22278, n22279, n22280, n22281,
         n22282, n22283, n22284, n22285, n22286, n22287, n22288, n22289,
         n22290, n22291, n22292, n22293, n22294, n22295, n22296, n22297,
         n22298, n22299, n22300, n22301, n22302, n22303, n22304, n22305,
         n22306, n22307, n22308, n22309, n22310, n22311, n22312, n22313,
         n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321,
         n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329,
         n22330, n22331, n22332, n22333, n22334, n22335, n22336, n22337,
         n22338, n22339, n22340, n22341, n22342, n22343, n22344, n22345,
         n22346, n22347, n22348, n22349, n22350, n22351, n22352, n22353,
         n22354, n22355, n22356, n22357, n22358, n22359, n22360, n22361,
         n22362, n22363, n22364, n22365, n22366, n22367, n22368, n22369,
         n22370, n22371, n22372, n22373, n22374, n22375, n22376, n22377,
         n22378, n22379, n22380, n22381, n22382, n22383, n22384, n22385,
         n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393,
         n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401,
         n22402, n22403, n22404, n22405, n22406, n22407, n22408, n22409,
         n22410, n22411, n22412, n22413, n22414, n22415, n22416, n22417,
         n22418, n22419, n22420, n22421, n22422, n22423, n22424, n22425,
         n22426, n22427, n22428, n22429, n22430, n22431, n22432, n22433,
         n22434, n22435, n22436, n22437, n22438, n22439, n22440, n22441,
         n22442, n22443, n22444, n22445, n22446, n22447, n22448, n22449,
         n22450, n22451, n22452, n22453, n22454, n22455, n22456, n22457,
         n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465,
         n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473,
         n22474, n22475, n22476, n22477, n22478, n22479, n22480, n22481,
         n22482, n22483, n22484, n22485, n22486, n22487, n22488, n22489,
         n22490, n22491, n22492, n22493, n22494, n22495, n22496, n22497,
         n22498, n22499, n22500, n22501, n22502, n22503, n22504, n22505,
         n22506, n22507, n22508, n22509, n22510, n22511, n22512, n22513,
         n22514, n22515, n22516, n22517, n22518, n22519, n22520, n22521,
         n22522, n22523, n22524, n22525, n22526, n22527, n22528, n22529,
         n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537,
         n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545,
         n22546, n22547, n22548, n22549, n22550, n22551, n22552, n22553,
         n22554, n22555, n22556, n22557, n22558, n22559, n22560, n22561,
         n22562, n22563, n22564, n22565, n22566, n22567, n22568, n22569,
         n22570, n22571, n22572, n22573, n22574, n22575, n22576, n22577,
         n22578, n22579, n22580, n22581, n22582, n22583, n22584, n22585,
         n22586, n22587, n22588, n22589, n22590, n22591, n22592, n22593,
         n22594, n22595, n22596, n22597, n22598, n22599, n22600, n22601,
         n22602, n22603, n22604, n22605, n22606, n22607, n22608, n22609,
         n22610, n22611, n22612, n22613, n22614, n22615, n22616, n22617,
         n22618, n22619, n22620, n22621, n22622, n22623, n22624, n22625,
         n22626, n22627, n22628, n22629, n22630, n22631, n22632, n22633,
         n22634, n22635, n22636, n22637, n22638, n22639, n22640, n22641,
         n22642, n22643, n22644, n22645, n22646, n22647, n22648, n22649,
         n22650, n22651, n22652, n22653, n22654, n22655, n22656, n22657,
         n22658, n22659, n22660, n22661, n22662, n22663, n22664, n22665,
         n22666, n22667, n22668, n22669, n22670, n22671, n22672, n22673,
         n22674, n22675, n22676, n22677, n22678, n22679, n22680, n22681,
         n22682, n22683, n22684, n22685, n22686, n22687, n22688, n22689,
         n22690, n22691, n22692, n22693, n22694, n22695, n22696, n22697,
         n22698, n22699, n22700, n22701, n22702, n22703, n22704, n22705,
         n22706, n22707, n22708, n22709, n22710, n22711, n22712, n22713,
         n22714, n22715, n22716, n22717, n22718, n22719, n22720, n22721,
         n22722, n22723, n22724, n22725, n22726, n22727, n22728, n22729,
         n22730, n22731, n22732, n22733, n22734, n22735, n22736, n22737,
         n22738, n22739, n22740, n22741, n22742, n22743, n22744, n22745,
         n22746, n22747, n22748, n22749, n22750, n22751, n22752, n22753,
         n22754, n22755, n22756, n22757, n22758, n22759, n22760, n22761,
         n22762, n22763, n22764, n22765, n22766, n22767, n22768, n22769,
         n22770, n22771, n22772, n22773, n22774, n22775, n22776, n22777,
         n22778, n22779, n22780, n22781, n22782, n22783, n22784, n22785,
         n22786, n22787, n22788, n22789, n22790, n22791, n22792, n22793,
         n22794, n22795, n22796, n22797, n22798, n22799, n22800, n22801,
         n22802, n22803, n22804, n22805, n22806, n22807, n22808, n22809,
         n22810, n22811, n22812, n22813, n22814, n22815, n22816, n22817,
         n22818, n22819, n22820, n22821, n22822, n22823, n22824, n22825,
         n22826, n22827, n22828, n22829, n22830, n22831, n22832, n22833,
         n22834, n22835, n22836, n22837, n22838, n22839, n22840, n22841,
         n22842, n22843, n22844, n22845, n22846, n22847, n22848, n22849,
         n22850, n22851, n22852, n22853, n22854, n22855, n22856, n22857,
         n22858, n22859, n22860, n22861, n22862, n22863, n22864, n22865,
         n22866, n22867, n22868, n22869, n22870, n22871, n22872, n22873,
         n22874, n22875, n22876, n22877, n22878, n22879, n22880, n22881,
         n22882, n22883, n22884, n22885, n22886, n22887, n22888, n22889,
         n22890, n22891, n22892, n22893, n22894, n22895, n22896, n22897,
         n22898, n22899, n22900, n22901, n22902, n22903, n22904, n22905,
         n22906, n22907, n22908, n22909, n22910, n22911, n22912, n22913,
         n22914, n22915, n22916, n22917, n22918, n22919, n22920, n22921,
         n22922, n22923, n22924, n22925, n22926, n22927, n22928, n22929,
         n22930, n22931, n22932, n22933, n22934, n22935, n22936, n22937,
         n22938, n22939, n22940, n22941, n22942, n22943, n22944, n22945,
         n22946, n22947, n22948, n22949, n22950, n22951, n22952, n22953,
         n22954, n22955, n22956, n22957, n22958, n22959, n22960, n22961,
         n22962, n22963, n22964, n22965, n22966, n22967, n22968, n22969,
         n22970, n22971, n22972, n22973, n22974, n22975, n22976, n22977,
         n22978, n22979, n22980, n22981, n22982, n22983, n22984, n22985,
         n22986, n22987, n22988, n22989, n22990, n22991, n22992, n22993,
         n22994, n22995, n22996, n22997, n22998, n22999, n23000, n23001,
         n23002, n23003, n23004, n23005, n23006, n23007, n23008, n23009,
         n23010, n23011, n23012, n23013, n23014, n23015, n23016, n23017,
         n23018, n23019, n23020, n23021, n23022, n23023, n23024, n23025,
         n23026, n23027, n23028, n23029, n23030, n23031, n23032, n23033,
         n23034, n23035, n23036, n23037, n23038, n23039, n23040, n23041,
         n23042, n23043, n23044, n23045, n23046, n23047, n23048, n23049,
         n23050, n23051, n23052, n23053, n23054, n23055, n23056, n23057,
         n23058, n23059, n23060, n23061, n23062, n23063, n23064, n23065,
         n23066, n23067, n23068, n23069, n23070, n23071, n23072, n23073,
         n23074, n23075, n23076, n23077, n23078, n23079, n23080, n23081,
         n23082, n23083, n23084, n23085, n23086, n23087, n23088, n23089,
         n23090, n23091, n23092, n23093, n23094, n23095, n23096, n23097,
         n23098, n23099, n23100, n23101, n23102, n23103, n23104, n23105,
         n23106, n23107, n23108, n23109, n23110, n23111, n23112, n23113,
         n23114, n23115, n23116, n23117, n23118, n23119, n23120, n23121,
         n23122, n23123, n23124, n23125, n23126, n23127, n23128, n23129,
         n23130, n23131, n23132, n23133, n23134, n23135, n23136, n23137,
         n23138, n23139, n23140, n23141, n23142, n23143, n23144, n23145,
         n23146, n23147, n23148, n23149, n23150, n23151, n23152, n23153,
         n23154, n23155, n23156, n23157, n23158, n23159, n23160, n23161,
         n23162, n23163, n23164, n23165, n23166, n23167, n23168, n23169,
         n23170, n23171, n23172, n23173, n23174, n23175, n23176, n23177,
         n23178, n23179, n23180, n23181, n23182, n23183, n23184, n23185,
         n23186, n23187, n23188, n23189, n23190, n23191, n23192, n23193,
         n23194, n23195, n23196, n23197, n23198, n23199, n23200, n23201,
         n23202, n23203, n23204, n23205, n23206, n23207, n23208, n23209,
         n23210, n23211, n23212, n23213, n23214, n23215, n23216, n23217,
         n23218, n23219, n23220, n23221, n23222, n23223, n23224, n23225,
         n23226, n23227, n23228, n23229, n23230, n23231, n23232, n23233,
         n23234, n23235, n23236, n23237, n23238, n23239, n23240, n23241,
         n23242, n23243, n23244, n23245, n23246, n23247, n23248, n23249,
         n23250, n23251, n23252, n23253, n23254, n23255, n23256, n23257,
         n23258, n23259, n23260, n23261, n23262, n23263, n23264, n23265,
         n23266, n23267, n23268, n23269, n23270, n23271, n23272, n23273,
         n23274, n23275, n23276, n23277, n23278, n23279, n23280, n23281,
         n23282, n23283, n23284, n23285, n23286, n23287, n23288, n23289,
         n23290, n23291, n23292, n23293, n23294, n23295, n23296, n23297,
         n23298, n23299, n23300, n23301, n23302, n23303, n23304, n23305,
         n23306, n23307, n23308, n23309, n23310, n23311, n23312, n23313,
         n23314, n23315, n23316, n23317, n23318, n23319, n23320, n23321,
         n23322, n23323, n23324, n23325, n23326, n23327, n23328, n23329,
         n23330, n23331, n23332, n23333, n23334, n23335, n23336, n23337,
         n23338, n23339, n23340, n23341, n23342, n23343, n23344, n23345,
         n23346, n23347, n23348, n23349, n23350, n23351, n23352, n23353,
         n23354, n23355, n23356, n23357, n23358, n23359, n23360, n23361,
         n23362, n23363, n23364, n23365, n23366, n23367, n23368, n23369,
         n23370, n23371, n23372, n23373, n23374, n23375, n23376, n23377,
         n23378, n23379, n23380, n23381, n23382, n23383, n23384, n23385,
         n23386, n23387, n23388, n23389, n23390, n23391, n23392, n23393,
         n23394, n23395, n23396, n23397, n23398, n23399, n23400, n23401,
         n23402, n23403, n23404, n23405, n23406, n23407, n23408, n23409,
         n23410, n23411, n23412, n23413, n23414, n23415, n23416, n23417,
         n23418, n23419, n23420, n23421, n23422, n23423, n23424, n23425,
         n23426, n23427, n23428, n23429, n23430, n23431, n23432, n23433,
         n23434, n23435, n23436, n23437, n23438, n23439, n23440, n23441,
         n23442, n23443, n23444, n23445, n23446, n23447, n23448, n23449,
         n23450, n23451, n23452, n23453, n23454, n23455, n23456, n23457,
         n23458, n23459, n23460, n23461, n23462, n23463, n23464, n23465,
         n23466, n23467, n23468, n23469, n23470, n23471, n23472, n23473,
         n23474, n23475, n23476, n23477, n23478, n23479, n23480, n23481,
         n23482, n23483, n23484, n23485, n23486, n23487, n23488, n23489,
         n23490, n23491, n23492, n23493, n23494, n23495, n23496, n23497,
         n23498, n23499, n23500, n23501, n23502, n23503, n23504, n23505,
         n23506, n23507, n23508, n23509, n23510, n23511, n23512, n23513,
         n23514, n23515, n23516, n23517, n23518, n23519, n23520, n23521,
         n23522, n23523, n23524, n23525, n23526, n23527, n23528, n23529,
         n23530, n23531, n23532, n23533, n23534, n23535, n23536, n23537,
         n23538, n23539, n23540, n23541, n23542, n23543, n23544, n23545,
         n23546, n23547, n23548, n23549, n23550, n23551, n23552, n23553,
         n23554, n23555, n23556, n23557, n23558, n23559, n23560, n23561,
         n23562, n23563, n23564, n23565, n23566, n23567, n23568, n23569,
         n23570, n23571, n23572, n23573, n23574, n23575, n23576, n23577,
         n23578, n23579, n23580, n23581, n23582, n23583, n23584, n23585,
         n23586, n23587, n23588, n23589, n23590, n23591, n23592, n23593,
         n23594, n23595, n23596, n23597, n23598, n23599, n23600, n23601,
         n23602, n23603, n23604, n23605, n23606, n23607, n23608, n23609,
         n23610, n23611, n23612, n23613, n23614, n23615, n23616, n23617,
         n23618, n23619, n23620, n23621, n23622, n23623, n23624, n23625,
         n23626, n23627, n23628, n23629, n23630, n23631, n23632, n23633,
         n23634, n23635, n23636, n23637, n23638, n23639, n23640, n23641,
         n23642, n23643, n23644, n23645, n23646, n23647, n23648, n23649,
         n23650, n23651, n23652, n23653, n23654, n23655, n23656, n23657,
         n23658, n23659, n23660, n23661, n23662, n23663, n23664, n23665,
         n23666, n23667, n23668, n23669, n23670, n23671, n23672, n23673,
         n23674, n23675, n23676, n23677, n23678, n23679, n23680, n23681,
         n23682, n23683, n23684, n23685, n23686, n23687, n23688, n23689,
         n23690, n23691, n23692, n23693, n23694, n23695, n23696, n23697,
         n23698, n23699, n23700, n23701, n23702, n23703, n23704, n23705,
         n23706, n23707, n23708, n23709, n23710, n23711, n23712, n23713,
         n23714, n23715, n23716, n23717, n23718, n23719, n23720, n23721,
         n23722, n23723, n23724, n23725, n23726, n23727, n23728, n23729,
         n23730, n23731, n23732, n23733, n23734, n23735, n23736, n23737,
         n23738, n23739, n23740, n23741, n23742, n23743, n23744, n23745,
         n23746, n23747, n23748, n23749, n23750, n23751, n23752, n23753,
         n23754, n23755, n23756, n23757, n23758, n23759, n23760, n23761,
         n23762, n23763, n23764, n23765, n23766, n23767, n23768, n23769,
         n23770, n23771, n23772, n23773, n23774, n23775, n23776, n23777,
         n23778, n23779, n23780, n23781, n23782, n23783, n23784, n23785,
         n23786, n23787, n23788, n23789, n23790, n23791, n23792, n23793,
         n23794, n23795, n23796, n23797, n23798, n23799, n23800, n23801,
         n23802, n23803, n23804, n23805, n23806, n23807, n23808, n23809,
         n23810, n23811, n23812, n23813, n23814, n23815, n23816, n23817,
         n23818, n23819, n23820, n23821, n23822, n23823, n23824, n23825,
         n23826, n23827, n23828, n23829, n23830, n23831, n23832, n23833,
         n23834, n23835, n23836, n23837, n23838, n23839, n23840, n23841,
         n23842, n23843, n23844, n23845, n23846, n23847, n23848, n23849,
         n23850, n23851, n23852, n23853, n23854, n23855, n23856, n23857,
         n23858, n23859, n23860, n23861, n23862, n23863, n23864, n23865,
         n23866, n23867, n23868, n23869, n23870, n23871, n23872, n23873,
         n23874, n23875, n23876, n23877, n23878, n23879, n23880, n23881,
         n23882, n23883, n23884, n23885, n23886, n23887, n23888, n23889,
         n23890, n23891, n23892, n23893, n23894, n23895, n23896, n23897,
         n23898, n23899, n23900, n23901, n23902, n23903, n23904, n23905,
         n23906, n23907, n23908, n23909, n23910, n23911, n23912, n23913,
         n23914, n23915, n23916, n23917, n23918, n23919, n23920, n23921,
         n23922, n23923, n23924, n23925, n23926, n23927, n23928, n23929,
         n23930, n23931, n23932, n23933, n23934, n23935, n23936, n23937,
         n23938, n23939, n23940, n23941, n23942, n23943, n23944, n23945,
         n23946, n23947, n23948, n23949, n23950, n23951, n23952, n23953,
         n23954, n23955, n23956, n23957, n23958, n23959, n23960, n23961,
         n23962, n23963, n23964, n23965, n23966, n23967, n23968, n23969,
         n23970, n23971, n23972, n23973, n23974, n23975, n23976, n23977,
         n23978, n23979, n23980, n23981, n23982, n23983, n23984, n23985,
         n23986, n23987, n23988, n23989, n23990, n23991, n23992, n23993,
         n23994, n23995, n23996, n23997, n23998, n23999, n24000, n24001,
         n24002, n24003, n24004, n24005, n24006, n24007, n24008, n24009,
         n24010, n24011, n24012, n24013, n24014, n24015, n24016, n24017,
         n24018, n24019, n24020, n24021, n24022, n24023, n24024, n24025,
         n24026, n24027, n24028, n24029, n24030, n24031, n24032, n24033,
         n24034, n24035, n24036, n24037, n24038, n24039, n24040, n24041,
         n24042, n24043, n24044, n24045, n24046, n24047, n24048, n24049,
         n24050, n24051, n24052, n24053, n24054, n24055, n24056, n24057,
         n24058, n24059, n24060, n24061, n24062, n24063, n24064, n24065,
         n24066, n24067, n24068, n24069, n24070, n24071, n24072, n24073,
         n24074, n24075, n24076, n24077, n24078, n24079, n24080, n24081,
         n24082, n24083, n24084, n24085, n24086, n24087, n24088, n24089,
         n24090, n24091, n24092, n24093, n24094, n24095, n24096, n24097,
         n24098, n24099, n24100, n24101, n24102, n24103, n24104, n24105,
         n24106, n24107, n24108, n24109, n24110, n24111, n24112, n24113,
         n24114, n24115, n24116, n24117, n24118, n24119, n24120, n24121,
         n24122, n24123, n24124, n24125, n24126, n24127, n24128, n24129,
         n24130, n24131, n24132, n24133, n24134, n24135, n24136, n24137,
         n24138, n24139, n24140, n24141, n24142, n24143, n24144, n24145,
         n24146, n24147, n24148, n24149, n24150, n24151, n24152, n24153,
         n24154, n24155, n24156, n24157, n24158, n24159, n24160, n24161,
         n24162, n24163, n24164, n24165, n24166, n24167, n24168, n24169,
         n24170, n24171, n24172, n24173, n24174, n24175, n24176, n24177,
         n24178, n24179, n24180, n24181, n24182, n24183, n24184, n24185,
         n24186, n24187, n24188, n24189, n24190, n24191, n24192, n24193,
         n24194, n24195, n24196, n24197, n24198, n24199, n24200, n24201,
         n24202, n24203, n24204, n24205, n24206, n24207, n24208, n24209,
         n24210, n24211, n24212, n24213, n24214, n24215, n24216, n24217,
         n24218, n24219, n24220, n24221, n24222, n24223, n24224, n24225,
         n24226, n24227, n24228, n24229, n24230, n24231, n24232, n24233,
         n24234, n24235, n24236, n24237, n24238, n24239, n24240, n24241,
         n24242, n24243, n24244, n24245, n24246, n24247, n24248, n24249,
         n24250, n24251, n24252, n24253, n24254, n24255, n24256, n24257,
         n24258, n24259, n24260, n24261, n24262, n24263, n24264, n24265,
         n24266, n24267, n24268, n24269, n24270, n24271, n24272, n24273,
         n24274, n24275, n24276, n24277, n24278, n24279, n24280, n24281,
         n24282, n24283, n24284, n24285, n24286, n24287, n24288, n24289,
         n24290, n24291, n24292, n24293, n24294, n24295, n24296, n24297,
         n24298, n24299, n24300, n24301, n24302, n24303, n24304, n24305,
         n24306, n24307, n24308, n24309, n24310, n24311, n24312, n24313,
         n24314, n24315, n24316, n24317, n24318, n24319, n24320, n24321,
         n24322, n24323, n24324, n24325, n24326, n24327, n24328, n24329,
         n24330, n24331, n24332, n24333, n24334, n24335, n24336, n24337,
         n24338, n24339, n24340, n24341, n24342, n24343, n24344, n24345,
         n24346, n24347, n24348, n24349, n24350, n24351, n24352, n24353,
         n24354, n24355, n24356, n24357, n24358, n24359, n24360, n24361,
         n24362, n24363, n24364, n24365, n24366, n24367, n24368, n24369,
         n24370, n24371, n24372, n24373, n24374, n24375, n24376, n24377,
         n24378, n24379, n24380, n24381, n24382, n24383, n24384, n24385,
         n24386, n24387, n24388, n24389, n24390, n24391, n24392, n24393,
         n24394, n24395, n24396, n24397, n24398, n24399, n24400, n24401,
         n24402, n24403, n24404, n24405, n24406, n24407, n24408, n24409,
         n24410, n24411, n24412, n24413, n24414, n24415, n24416, n24417,
         n24418, n24419, n24420, n24421, n24422, n24423, n24424, n24425,
         n24426, n24427, n24428, n24429, n24430, n24431, n24432, n24433,
         n24434, n24435, n24436, n24437, n24438, n24439, n24440, n24441,
         n24442, n24443, n24444, n24445, n24446, n24447, n24448, n24449,
         n24450, n24451, n24452, n24453, n24454, n24455, n24456, n24457,
         n24458, n24459, n24460, n24461, n24462, n24463, n24464, n24465,
         n24466, n24467, n24468, n24469, n24470, n24471, n24472, n24473,
         n24474, n24475, n24476, n24477, n24478, n24479, n24480, n24481,
         n24482, n24483, n24484, n24485, n24486, n24487, n24488, n24489,
         n24490, n24491, n24492, n24493, n24494, n24495, n24496, n24497,
         n24498, n24499, n24500, n24501, n24502, n24503, n24504, n24505,
         n24506, n24507, n24508, n24509, n24510, n24511, n24512, n24513,
         n24514, n24515, n24516, n24517, n24518, n24519, n24520, n24521,
         n24522, n24523, n24524, n24525, n24526, n24527, n24528, n24529,
         n24530, n24531, n24532, n24533, n24534, n24535, n24536, n24537,
         n24538, n24539, n24540, n24541, n24542, n24543, n24544, n24545,
         n24546, n24547, n24548, n24549, n24550, n24551, n24552, n24553,
         n24554, n24555, n24556, n24557, n24558, n24559, n24560, n24561,
         n24562, n24563, n24564, n24565, n24566, n24567, n24568, n24569,
         n24570, n24571, n24572, n24573, n24574, n24575, n24576, n24577,
         n24578, n24579, n24580, n24581, n24582, n24583, n24584, n24585,
         n24586, n24587, n24588, n24589, n24590, n24591, n24592, n24593,
         n24594, n24595, n24596, n24597, n24598, n24599, n24600, n24601,
         n24602, n24603, n24604, n24605, n24606, n24607, n24608, n24609,
         n24610, n24611, n24612, n24613, n24614, n24615, n24616, n24617,
         n24618, n24619, n24620, n24621, n24622, n24623, n24624, n24625,
         n24626, n24627, n24628, n24629, n24630, n24631, n24632, n24633,
         n24634, n24635, n24636, n24637, n24638, n24639, n24640, n24641,
         n24642, n24643, n24644, n24645, n24646, n24647, n24648, n24649,
         n24650, n24651, n24652, n24653, n24654, n24655, n24656, n24657,
         n24658, n24659, n24660, n24661, n24662, n24663, n24664, n24665,
         n24666, n24667, n24668, n24669, n24670, n24671, n24672, n24673,
         n24674, n24675, n24676, n24677, n24678, n24679, n24680, n24681,
         n24682, n24683, n24684, n24685, n24686, n24687, n24688, n24689,
         n24690, n24691, n24692, n24693, n24694, n24695, n24696, n24697,
         n24698, n24699, n24700, n24701, n24702, n24703, n24704, n24705,
         n24706, n24707, n24708, n24709, n24710, n24711, n24712, n24713,
         n24714, n24715, n24716, n24717, n24718, n24719, n24720, n24721,
         n24722, n24723, n24724, n24725, n24726, n24727, n24728, n24729,
         n24730, n24731, n24732, n24733, n24734, n24735, n24736, n24737,
         n24738, n24739, n24740, n24741, n24742, n24743, n24744, n24745,
         n24746, n24747, n24748, n24749, n24750, n24751, n24752, n24753,
         n24754, n24755, n24756, n24757, n24758, n24759, n24760, n24761,
         n24762, n24763, n24764, n24765, n24766, n24767, n24768, n24769,
         n24770, n24771, n24772, n24773, n24774, n24775, n24776, n24777,
         n24778, n24779, n24780, n24781, n24782, n24783, n24784, n24785,
         n24786, n24787, n24788, n24789, n24790, n24791, n24792, n24793,
         n24794, n24795, n24796, n24797, n24798, n24799, n24800, n24801,
         n24802, n24803, n24804, n24805, n24806, n24807, n24808, n24809,
         n24810, n24811, n24812, n24813, n24814, n24815, n24816, n24817,
         n24818, n24819, n24820, n24821, n24822, n24823, n24824, n24825,
         n24826, n24827, n24828, n24829, n24830, n24831, n24832, n24833,
         n24834, n24835, n24836, n24837, n24838, n24839, n24840, n24841,
         n24842, n24843, n24844, n24845, n24846, n24847, n24848, n24849,
         n24850, n24851, n24852, n24853, n24854, n24855, n24856, n24857,
         n24858, n24859, n24860, n24861, n24862, n24863, n24864, n24865,
         n24866, n24867, n24868, n24869, n24870, n24871, n24872, n24873,
         n24874, n24875, n24876, n24877, n24878, n24879, n24880, n24881,
         n24882, n24883, n24884, n24885, n24886, n24887, n24888, n24889,
         n24890, n24891, n24892, n24893, n24894, n24895, n24896, n24897,
         n24898, n24899, n24900, n24901, n24902, n24903, n24904, n24905,
         n24906, n24907, n24908, n24909, n24910, n24911, n24912, n24913,
         n24914, n24915, n24916, n24917, n24918, n24919, n24920, n24921,
         n24922, n24923, n24924, n24925, n24926, n24927, n24928, n24929,
         n24930, n24931, n24932, n24933, n24934, n24935, n24936, n24937,
         n24938, n24939, n24940, n24941, n24942, n24943, n24944, n24945,
         n24946, n24947, n24948, n24949, n24950, n24951, n24952, n24953,
         n24954, n24955, n24956, n24957, n24958, n24959, n24960, n24961,
         n24962, n24963, n24964, n24965, n24966, n24967, n24968, n24969,
         n24970, n24971, n24972, n24973, n24974, n24975, n24976, n24977,
         n24978, n24979, n24980, n24981, n24982, n24983, n24984, n24985,
         n24986, n24987, n24988, n24989, n24990, n24991, n24992, n24993,
         n24994, n24995, n24996, n24997, n24998, n24999, n25000, n25001,
         n25002, n25003, n25004, n25005, n25006, n25007, n25008, n25009,
         n25010, n25011, n25012, n25013, n25014, n25015, n25016, n25017,
         n25018, n25019, n25020, n25021, n25022, n25023, n25024, n25025,
         n25026, n25027, n25028, n25029, n25030, n25031, n25032, n25033,
         n25034, n25035, n25036, n25037, n25038, n25039, n25040, n25041,
         n25042, n25043, n25044, n25045, n25046, n25047, n25048, n25049,
         n25050, n25051, n25052, n25053, n25054, n25055, n25056, n25057,
         n25058, n25059, n25060, n25061, n25062, n25063, n25064, n25065,
         n25066, n25067, n25068, n25069, n25070, n25071, n25072, n25073,
         n25074, n25075, n25076, n25077, n25078, n25079, n25080, n25081,
         n25082, n25083, n25084, n25085, n25086, n25087, n25088, n25089,
         n25090, n25091, n25092, n25093, n25094, n25095, n25096, n25097,
         n25098, n25099, n25100, n25101, n25102, n25103, n25104, n25105,
         n25106, n25107, n25108, n25109, n25110, n25111, n25112, n25113,
         n25114, n25115, n25116, n25117, n25118, n25119, n25120, n25121,
         n25122, n25123, n25124, n25125, n25126, n25127, n25128, n25129,
         n25130, n25131, n25132, n25133, n25134, n25135, n25136, n25137,
         n25138, n25139, n25140, n25141, n25142, n25143, n25144, n25145,
         n25146, n25147, n25148, n25149, n25150, n25151, n25152, n25153,
         n25154, n25155, n25156, n25157, n25158, n25159, n25160, n25161,
         n25162, n25163, n25164, n25165, n25166, n25167, n25168, n25169,
         n25170, n25171, n25172, n25173, n25174, n25175, n25176, n25177,
         n25178, n25179, n25180, n25181, n25182, n25183, n25184, n25185,
         n25186, n25187, n25188, n25189, n25190, n25191, n25192, n25193,
         n25194, n25195, n25196, n25197, n25198, n25199, n25200, n25201,
         n25202, n25203, n25204, n25205, n25206, n25207, n25208, n25209,
         n25210, n25211, n25212, n25213, n25214, n25215, n25216, n25217,
         n25218, n25219, n25220, n25221, n25222, n25223, n25224, n25225,
         n25226, n25227, n25228, n25229, n25230, n25231, n25232, n25233,
         n25234, n25235, n25236, n25237, n25238, n25239, n25240, n25241,
         n25242, n25243, n25244, n25245, n25246, n25247, n25248, n25249,
         n25250, n25251, n25252, n25253, n25254, n25255, n25256, n25257,
         n25258, n25259, n25260, n25261, n25262, n25263, n25264, n25265,
         n25266, n25267, n25268, n25269, n25270, n25271, n25272, n25273,
         n25274, n25275, n25276, n25277, n25278, n25279, n25280, n25281,
         n25282, n25283, n25284, n25285, n25286, n25287, n25288, n25289,
         n25290, n25291, n25292, n25293, n25294, n25295, n25296, n25297,
         n25298, n25299, n25300, n25301, n25302, n25303, n25304, n25305,
         n25306, n25307, n25308, n25309, n25310, n25311, n25312, n25313,
         n25314, n25315, n25316, n25317, n25318, n25319, n25320, n25321,
         n25322, n25323, n25324, n25325, n25326, n25327, n25328, n25329,
         n25330, n25331, n25332, n25333, n25334, n25335, n25336, n25337,
         n25338, n25339, n25340, n25341, n25342, n25343, n25344, n25345,
         n25346, n25347, n25348, n25349, n25350, n25351, n25352, n25353,
         n25354, n25355, n25356, n25357, n25358, n25359, n25360, n25361,
         n25362, n25363, n25364, n25365, n25366, n25367, n25368, n25369,
         n25370, n25371, n25372, n25373, n25374, n25375, n25376, n25377,
         n25378, n25379, n25380, n25381, n25382, n25383, n25384, n25385,
         n25386, n25387, n25388, n25389, n25390, n25391, n25392, n25393,
         n25394, n25395, n25396, n25397, n25398, n25399, n25400, n25401,
         n25402, n25403, n25404, n25405, n25406, n25407, n25408, n25409,
         n25410, n25411, n25412, n25413, n25414, n25415, n25416, n25417,
         n25418, n25419, n25420, n25421, n25422, n25423, n25424, n25425,
         n25426, n25427, n25428, n25429, n25430, n25431, n25432, n25433,
         n25434, n25435, n25436, n25437, n25438, n25439, n25440, n25441,
         n25442, n25443, n25444, n25445, n25446, n25447, n25448, n25449,
         n25450, n25451, n25452, n25453, n25454, n25455, n25456, n25457,
         n25458, n25459, n25460, n25461, n25462, n25463, n25464, n25465,
         n25466, n25467, n25468, n25469, n25470, n25471, n25472, n25473,
         n25474, n25475, n25476, n25477, n25478, n25479, n25480, n25481,
         n25482, n25483, n25484, n25485, n25486, n25487, n25488, n25489,
         n25490, n25491, n25492, n25493, n25494, n25495, n25496, n25497,
         n25498, n25499, n25500, n25501, n25502, n25503, n25504, n25505,
         n25506, n25507, n25508, n25509, n25510, n25511, n25512, n25513,
         n25514, n25515, n25516, n25517, n25518, n25519, n25520, n25521,
         n25522, n25523, n25524, n25525, n25526, n25527, n25528, n25529,
         n25530, n25531, n25532, n25533, n25534, n25535, n25536, n25537,
         n25538, n25539, n25540, n25541, n25542, n25543, n25544, n25545,
         n25546, n25547, n25548, n25549, n25550, n25551, n25552, n25553,
         n25554, n25555, n25556, n25557, n25558, n25559, n25560, n25561,
         n25562, n25563, n25564, n25565, n25566, n25567, n25568, n25569,
         n25570, n25571, n25572, n25573, n25574, n25575, n25576, n25577,
         n25578, n25579, n25580, n25581, n25582, n25583, n25584, n25585,
         n25586, n25587, n25588, n25589, n25590, n25591, n25592, n25593,
         n25594, n25595, n25596, n25597, n25598, n25599, n25600, n25601,
         n25602, n25603, n25604, n25605, n25606, n25607, n25608, n25609,
         n25610, n25611, n25612, n25613, n25614, n25615, n25616, n25617,
         n25618, n25619, n25620, n25621, n25622, n25623, n25624, n25625,
         n25626, n25627, n25628, n25629, n25630, n25631, n25632, n25633,
         n25634, n25635, n25636, n25637, n25638, n25639, n25640, n25641,
         n25642, n25643, n25644, n25645, n25646, n25647, n25648, n25649,
         n25650, n25651, n25652, n25653, n25654, n25655, n25656, n25657,
         n25658, n25659, n25660, n25661, n25662, n25663, n25664, n25665,
         n25666, n25667, n25668, n25669, n25670, n25671, n25672, n25673,
         n25674, n25675, n25676, n25677, n25678, n25679, n25680, n25681,
         n25682, n25683, n25684, n25685, n25686, n25687, n25688, n25689,
         n25690, n25691, n25692, n25693, n25694, n25695, n25696, n25697,
         n25698, n25699, n25700, n25701, n25702, n25703, n25704, n25705,
         n25706, n25707, n25708, n25709, n25710, n25711, n25712, n25713,
         n25714, n25715, n25716, n25717, n25718, n25719, n25720, n25721,
         n25722, n25723, n25724, n25725, n25726, n25727, n25728, n25729,
         n25730, n25731, n25732, n25733, n25734, n25735, n25736, n25737,
         n25738, n25739, n25740, n25741, n25742, n25743, n25744, n25745,
         n25746, n25747, n25748, n25749, n25750, n25751, n25752, n25753,
         n25754, n25755, n25756, n25757, n25758, n25759, n25760, n25761,
         n25762, n25763, n25764, n25765, n25766, n25767, n25768, n25769,
         n25770, n25771, n25772, n25773, n25774, n25775, n25776, n25777,
         n25778, n25779, n25780, n25781, n25782, n25783, n25784, n25785,
         n25786, n25787, n25788, n25789, n25790, n25791, n25792, n25793,
         n25794, n25795, n25796, n25797, n25798, n25799, n25800, n25801,
         n25802, n25803, n25804, n25805, n25806, n25807, n25808, n25809,
         n25810, n25811, n25812, n25813, n25814, n25815, n25816, n25817,
         n25818, n25819, n25820, n25821, n25822, n25823, n25824, n25825,
         n25826, n25827, n25828, n25829, n25830, n25831, n25832, n25833,
         n25834, n25835, n25836, n25837, n25838, n25839, n25840, n25841,
         n25842, n25843, n25844, n25845, n25846, n25847, n25848, n25849,
         n25850, n25851, n25852, n25853, n25854, n25855, n25856, n25857,
         n25858, n25859, n25860, n25861, n25862, n25863, n25864, n25865,
         n25866, n25867, n25868, n25869, n25870, n25871, n25872, n25873,
         n25874, n25875, n25876, n25877, n25878, n25879, n25880, n25881,
         n25882, n25883, n25884, n25885, n25886, n25887, n25888, n25889,
         n25890, n25891, n25892, n25893, n25894, n25895, n25896, n25897,
         n25898, n25899, n25900, n25901, n25902, n25903, n25904, n25905,
         n25906, n25907, n25908, n25909, n25910, n25911, n25912, n25913,
         n25914, n25915, n25916, n25917, n25918, n25919, n25920, n25921,
         n25922, n25923, n25924, n25925, n25926, n25927, n25928, n25929,
         n25930, n25931, n25932, n25933, n25934, n25935, n25936, n25937,
         n25938, n25939, n25940, n25941, n25942, n25943, n25944, n25945,
         n25946, n25947, n25948, n25949, n25950, n25951, n25952, n25953,
         n25954, n25955, n25956, n25957, n25958, n25959, n25960, n25961,
         n25962, n25963, n25964, n25965, n25966, n25967, n25968, n25969,
         n25970, n25971, n25972, n25973, n25974, n25975, n25976, n25977,
         n25978, n25979, n25980, n25981, n25982, n25983, n25984, n25985,
         n25986, n25987, n25988, n25989, n25990, n25991, n25992, n25993,
         n25994, n25995, n25996, n25997, n25998, n25999, n26000, n26001,
         n26002, n26003, n26004, n26005, n26006, n26007, n26008, n26009,
         n26010, n26011, n26012, n26013, n26014, n26015, n26016, n26017,
         n26018, n26019, n26020, n26021, n26022, n26023, n26024, n26025,
         n26026, n26027, n26028, n26029, n26030, n26031, n26032, n26033,
         n26034, n26035, n26036, n26037, n26038, n26039, n26040, n26041,
         n26042, n26043, n26044, n26045, n26046, n26047, n26048, n26049,
         n26050, n26051, n26052, n26053, n26054, n26055, n26056, n26057,
         n26058, n26059, n26060, n26061, n26062, n26063, n26064, n26065,
         n26066, n26067, n26068, n26069, n26070, n26071, n26072, n26073,
         n26074, n26075, n26076, n26077, n26078, n26079, n26080, n26081,
         n26082, n26083, n26084, n26085, n26086, n26087, n26088, n26089,
         n26090, n26091, n26092, n26093, n26094, n26095, n26096, n26097,
         n26098, n26099, n26100, n26101, n26102, n26103, n26104, n26105,
         n26106, n26107, n26108, n26109, n26110, n26111, n26112, n26113,
         n26114, n26115, n26116, n26117, n26118, n26119, n26120, n26121,
         n26122, n26123, n26124, n26125, n26126, n26127, n26128, n26129,
         n26130, n26131, n26132, n26133, n26134, n26135, n26136, n26137,
         n26138, n26139, n26140, n26141, n26142, n26143, n26144, n26145,
         n26146, n26147, n26148, n26149, n26150, n26151, n26152, n26153,
         n26154, n26155, n26156, n26157, n26158, n26159, n26160, n26161,
         n26162, n26163, n26164, n26165, n26166, n26167, n26168, n26169,
         n26170, n26171, n26172, n26173, n26174, n26175, n26176, n26177,
         n26178, n26179, n26180, n26181, n26182, n26183, n26184, n26185,
         n26186, n26187, n26188, n26189, n26190, n26191, n26192, n26193,
         n26194, n26195, n26196, n26197, n26198, n26199, n26200, n26201,
         n26202, n26203, n26204, n26205, n26206, n26207, n26208, n26209,
         n26210, n26211, n26212, n26213, n26214, n26215, n26216, n26217,
         n26218, n26219, n26220, n26221, n26222, n26223, n26224, n26225,
         n26226, n26227, n26228, n26229, n26230, n26231, n26232, n26233,
         n26234, n26235, n26236, n26237, n26238, n26239, n26240, n26241,
         n26242, n26243, n26244, n26245, n26246, n26247, n26248, n26249,
         n26250, n26251, n26252, n26253, n26254, n26255, n26256, n26257,
         n26258, n26259, n26260, n26261, n26262, n26263, n26264, n26265,
         n26266, n26267, n26268, n26269, n26270, n26271, n26272, n26273,
         n26274, n26275, n26276, n26277, n26278, n26279, n26280, n26281,
         n26282, n26283, n26284, n26285, n26286, n26287, n26288, n26289,
         n26290, n26291, n26292, n26293, n26294, n26295, n26296, n26297,
         n26298, n26299, n26300, n26301, n26302, n26303, n26304, n26305,
         n26306, n26307, n26308, n26309, n26310, n26311, n26312, n26313,
         n26314, n26315, n26316, n26317, n26318, n26319, n26320, n26321,
         n26322, n26323, n26324, n26325, n26326, n26327, n26328, n26329,
         n26330, n26331, n26332, n26333, n26334, n26335, n26336, n26337,
         n26338, n26339, n26340, n26341, n26342, n26343, n26344, n26345,
         n26346, n26347, n26348, n26349, n26350, n26351, n26352, n26353,
         n26354, n26355, n26356, n26357, n26358, n26359, n26360, n26361,
         n26362, n26363, n26364, n26365, n26366, n26367, n26368, n26369,
         n26370, n26371, n26372, n26373, n26374, n26375, n26376, n26377,
         n26378, n26379, n26380, n26381, n26382, n26383, n26384, n26385,
         n26386, n26387, n26388, n26389, n26390, n26391, n26392, n26393,
         n26394, n26395, n26396, n26397, n26398, n26399, n26400, n26401,
         n26402, n26403, n26404, n26405, n26406, n26407, n26408, n26409,
         n26410, n26411, n26412, n26413, n26414, n26415, n26416, n26417,
         n26418, n26419, n26420, n26421, n26422, n26423, n26424, n26425,
         n26426, n26427, n26428, n26429, n26430, n26431, n26432, n26433,
         n26434, n26435, n26436, n26437, n26438, n26439, n26440, n26441,
         n26442, n26443, n26444, n26445, n26446, n26447, n26448, n26449,
         n26450, n26451, n26452, n26453, n26454, n26455, n26456, n26457,
         n26458, n26459, n26460, n26461, n26462, n26463, n26464, n26465,
         n26466, n26467, n26468, n26469, n26470, n26471, n26472, n26473,
         n26474, n26475, n26476, n26477, n26478, n26479, n26480, n26481,
         n26482, n26483, n26484, n26485, n26486, n26487, n26488, n26489,
         n26490, n26491, n26492, n26493, n26494, n26495, n26496, n26497,
         n26498, n26499, n26500, n26501, n26502, n26503, n26504, n26505,
         n26506, n26507, n26508, n26509, n26510, n26511, n26512, n26513,
         n26514, n26515, n26516, n26517, n26518, n26519, n26520, n26521,
         n26522, n26523, n26524, n26525, n26526, n26527, n26528, n26529,
         n26530, n26531, n26532, n26533, n26534, n26535, n26536, n26537,
         n26538, n26539, n26540, n26541, n26542, n26543, n26544, n26545,
         n26546, n26547, n26548, n26549, n26550, n26551, n26552, n26553,
         n26554, n26555, n26556, n26557, n26558, n26559, n26560, n26561,
         n26562, n26563, n26564, n26565, n26566, n26567, n26568, n26569,
         n26570, n26571, n26572, n26573, n26574, n26575, n26576, n26577,
         n26578, n26579, n26580, n26581, n26582, n26583, n26584, n26585,
         n26586, n26587, n26588, n26589, n26590, n26591, n26592, n26593,
         n26594, n26595, n26596, n26597, n26598, n26599, n26600, n26601,
         n26602, n26603, n26604, n26605, n26606, n26607, n26608, n26609,
         n26610, n26611, n26612, n26613, n26614, n26615, n26616, n26617,
         n26618, n26619, n26620, n26621, n26622, n26623, n26624, n26625,
         n26626, n26627, n26628, n26629, n26630, n26631, n26632, n26633,
         n26634, n26635, n26636, n26637, n26638, n26639, n26640, n26641,
         n26642, n26643, n26644, n26645, n26646, n26647, n26648, n26649,
         n26650, n26651, n26652, n26653, n26654, n26655, n26656, n26657,
         n26658, n26659, n26660, n26661, n26662, n26663, n26664, n26665,
         n26666, n26667, n26668, n26669, n26670, n26671, n26672, n26673,
         n26674, n26675, n26676, n26677, n26678, n26679, n26680, n26681,
         n26682, n26683, n26684, n26685, n26686, n26687, n26688, n26689,
         n26690, n26691, n26692, n26693, n26694, n26695, n26696, n26697,
         n26698, n26699, n26700, n26701, n26702, n26703, n26704, n26705,
         n26706, n26707, n26708, n26709, n26710, n26711, n26712, n26713,
         n26714, n26715, n26716, n26717, n26718, n26719, n26720, n26721,
         n26722, n26723, n26724, n26725, n26726, n26727, n26728, n26729,
         n26730, n26731, n26732, n26733, n26734, n26735, n26736, n26737,
         n26738, n26739, n26740, n26741, n26742, n26743, n26744, n26745,
         n26746, n26747, n26748, n26749, n26750, n26751, n26752, n26753,
         n26754, n26755, n26756, n26757, n26758, n26759, n26760, n26761,
         n26762, n26763, n26764, n26765, n26766, n26767, n26768, n26769,
         n26770, n26771, n26772, n26773, n26774, n26775, n26776, n26777,
         n26778, n26779, n26780, n26781, n26782, n26783, n26784, n26785,
         n26786, n26787, n26788, n26789, n26790, n26791, n26792, n26793,
         n26794, n26795, n26796, n26797, n26798, n26799, n26800, n26801,
         n26802, n26803, n26804, n26805, n26806, n26807, n26808, n26809,
         n26810, n26811, n26812, n26813, n26814, n26815, n26816, n26817,
         n26818, n26819, n26820, n26821, n26822, n26823, n26824, n26825,
         n26826, n26827, n26828, n26829, n26830, n26831, n26832, n26833,
         n26834, n26835, n26836, n26837, n26838, n26839, n26840, n26841,
         n26842, n26843, n26844, n26845, n26846, n26847, n26848, n26849,
         n26850, n26851, n26852, n26853, n26854, n26855, n26856, n26857,
         n26858, n26859, n26860, n26861, n26862, n26863, n26864, n26865,
         n26866, n26867, n26868, n26869, n26870, n26871, n26872, n26873,
         n26874, n26875, n26876, n26877, n26878, n26879, n26880, n26881,
         n26882, n26883, n26884, n26885, n26886, n26887, n26888, n26889,
         n26890, n26891, n26892, n26893, n26894, n26895, n26896, n26897,
         n26898, n26899, n26900, n26901, n26902, n26903, n26904, n26905,
         n26906, n26907, n26908, n26909, n26910, n26911, n26912, n26913,
         n26914, n26915, n26916, n26917, n26918, n26919, n26920, n26921,
         n26922, n26923, n26924, n26925, n26926, n26927, n26928, n26929,
         n26930, n26931, n26932, n26933, n26934, n26935, n26936, n26937,
         n26938, n26939, n26940, n26941, n26942, n26943, n26944, n26945,
         n26946, n26947, n26948, n26949, n26950, n26951, n26952, n26953,
         n26954, n26955, n26956, n26957, n26958, n26959, n26960, n26961,
         n26962, n26963, n26964, n26965, n26966, n26967, n26968, n26969,
         n26970, n26971, n26972, n26973, n26974, n26975, n26976, n26977,
         n26978, n26979, n26980, n26981, n26982, n26983, n26984, n26985,
         n26986, n26987, n26988, n26989, n26990, n26991, n26992, n26993,
         n26994, n26995, n26996, n26997, n26998, n26999, n27000, n27001,
         n27002, n27003, n27004, n27005, n27006, n27007, n27008, n27009,
         n27010, n27011, n27012, n27013, n27014, n27015, n27016, n27017,
         n27018, n27019, n27020, n27021, n27022, n27023, n27024, n27025,
         n27026, n27027, n27028, n27029, n27030, n27031, n27032, n27033,
         n27034, n27035, n27036, n27037, n27038, n27039, n27040, n27041,
         n27042, n27043, n27044, n27045, n27046, n27047, n27048, n27049,
         n27050, n27051, n27052, n27053, n27054, n27055, n27056, n27057,
         n27058, n27059, n27060, n27061, n27062, n27063, n27064, n27065,
         n27066, n27067, n27068, n27069, n27070, n27071, n27072, n27073,
         n27074, n27075, n27076, n27077, n27078, n27079, n27080, n27081,
         n27082, n27083, n27084, n27085, n27086, n27087, n27088, n27089,
         n27090, n27091, n27092, n27093, n27094, n27095, n27096, n27097,
         n27098, n27099, n27100, n27101, n27102, n27103, n27104, n27105,
         n27106, n27107, n27108, n27109, n27110, n27111, n27112, n27113,
         n27114, n27115, n27116, n27117, n27118, n27119, n27120, n27121,
         n27122, n27123, n27124, n27125, n27126, n27127, n27128, n27129,
         n27130, n27131, n27132, n27133, n27134, n27135, n27136, n27137,
         n27138, n27139, n27140, n27141, n27142, n27143, n27144, n27145,
         n27146, n27147, n27148, n27149, n27150, n27151, n27152, n27153,
         n27154, n27155, n27156, n27157, n27158, n27159, n27160, n27161,
         n27162, n27163, n27164, n27165, n27166, n27167, n27168, n27169,
         n27170, n27171, n27172, n27173, n27174, n27175, n27176, n27177,
         n27178, n27179, n27180, n27181, n27182, n27183, n27184, n27185,
         n27186, n27187, n27188, n27189, n27190, n27191, n27192, n27193,
         n27194, n27195, n27196, n27197, n27198, n27199, n27200, n27201,
         n27202, n27203, n27204, n27205, n27206, n27207, n27208, n27209,
         n27210, n27211, n27212, n27213, n27214, n27215, n27216, n27217,
         n27218, n27219, n27220, n27221, n27222, n27223, n27224, n27225,
         n27226, n27227, n27228, n27229, n27230, n27231, n27232, n27233,
         n27234, n27235, n27236, n27237, n27238, n27239, n27240, n27241,
         n27242, n27243, n27244, n27245, n27246, n27247, n27248, n27249,
         n27250, n27251, n27252, n27253, n27254, n27255, n27256, n27257,
         n27258, n27259, n27260, n27261, n27262, n27263, n27264, n27265,
         n27266, n27267, n27268, n27269, n27270, n27271, n27272, n27273,
         n27274, n27275, n27276, n27277, n27278, n27279, n27280, n27281,
         n27282, n27283, n27284, n27285, n27286, n27287, n27288, n27289,
         n27290, n27291, n27292, n27293, n27294, n27295, n27296, n27297,
         n27298, n27299, n27300, n27301, n27302, n27303, n27304, n27305,
         n27306, n27307, n27308, n27309, n27310, n27311, n27312, n27313,
         n27314, n27315, n27316, n27317, n27318, n27319, n27320, n27321,
         n27322, n27323, n27324, n27325, n27326, n27327, n27328, n27329,
         n27330, n27331, n27332, n27333, n27334, n27335, n27336, n27337,
         n27338, n27339, n27340, n27341, n27342, n27343, n27344, n27345,
         n27346, n27347, n27348, n27349, n27350, n27351, n27352, n27353,
         n27354, n27355, n27356, n27357, n27358, n27359, n27360, n27361,
         n27362, n27363, n27364, n27365, n27366, n27367, n27368, n27369,
         n27370, n27371, n27372, n27373, n27374, n27375, n27376, n27377,
         n27378, n27379, n27380, n27381, n27382, n27383, n27384, n27385,
         n27386, n27387, n27388, n27389, n27390, n27391, n27392, n27393,
         n27394, n27395, n27396, n27397, n27398, n27399, n27400, n27401,
         n27402, n27403, n27404, n27405, n27406, n27407, n27408, n27409,
         n27410, n27411, n27412, n27413, n27414, n27415, n27416, n27417,
         n27418, n27419, n27420, n27421, n27422, n27423, n27424, n27425,
         n27426, n27427, n27428, n27429, n27430, n27431, n27432, n27433,
         n27434, n27435, n27436, n27437, n27438, n27439, n27440, n27441,
         n27442, n27443, n27444, n27445, n27446, n27447, n27448, n27449,
         n27450, n27451, n27452, n27453, n27454, n27455, n27456, n27457,
         n27458, n27459, n27460, n27461, n27462, n27463, n27464, n27465,
         n27466, n27467, n27468, n27469, n27470, n27471, n27472, n27473,
         n27474, n27475, n27476, n27477, n27478, n27479, n27480, n27481,
         n27482, n27483, n27484, n27485, n27486, n27487, n27488, n27489,
         n27490, n27491, n27492, n27493, n27494, n27495, n27496, n27497,
         n27498, n27499, n27500, n27501, n27502, n27503, n27504, n27505,
         n27506, n27507, n27508, n27509, n27510, n27511, n27512, n27513,
         n27514, n27515, n27516, n27517, n27518, n27519, n27520, n27521,
         n27522, n27523, n27524, n27525, n27526, n27527, n27528, n27529,
         n27530, n27531, n27532, n27533, n27534, n27535, n27536, n27537,
         n27538, n27539, n27540, n27541, n27542, n27543, n27544, n27545,
         n27546, n27547, n27548, n27549, n27550, n27551, n27552, n27553,
         n27554, n27555, n27556, n27557, n27558, n27559, n27560, n27561,
         n27562, n27563, n27564, n27565, n27566, n27567, n27568, n27569,
         n27570, n27571, n27572, n27573, n27574, n27575, n27576, n27577,
         n27578, n27579, n27580, n27581, n27582, n27583, n27584, n27585,
         n27586, n27587, n27588, n27589, n27590, n27591, n27592, n27593,
         n27594, n27595, n27596, n27597, n27598, n27599, n27600, n27601,
         n27602, n27603, n27604, n27605, n27606, n27607, n27608, n27609,
         n27610, n27611, n27612, n27613, n27614, n27615, n27616, n27617,
         n27618, n27619, n27620, n27621, n27622, n27623, n27624, n27625,
         n27626, n27627, n27628, n27629, n27630, n27631, n27632, n27633,
         n27634, n27635, n27636, n27637, n27638, n27639, n27640, n27641,
         n27642, n27643, n27644, n27645, n27646, n27647, n27648, n27649,
         n27650, n27651, n27652, n27653, n27654, n27655, n27656, n27657,
         n27658, n27659, n27660, n27661, n27662, n27663, n27664, n27665,
         n27666, n27667, n27668, n27669, n27670, n27671, n27672, n27673,
         n27674, n27675, n27676, n27677, n27678, n27679, n27680, n27681,
         n27682, n27683, n27684, n27685, n27686, n27687, n27688, n27689,
         n27690, n27691, n27692, n27693, n27694, n27695, n27696, n27697,
         n27698, n27699, n27700, n27701, n27702, n27703, n27704, n27705,
         n27706, n27707, n27708, n27709, n27710, n27711, n27712, n27713,
         n27714, n27715, n27716, n27717, n27718, n27719, n27720, n27721,
         n27722, n27723, n27724, n27725, n27726, n27727, n27728, n27729,
         n27730, n27731, n27732, n27733, n27734, n27735, n27736, n27737,
         n27738, n27739, n27740, n27741, n27742, n27743, n27744, n27745,
         n27746, n27747, n27748, n27749, n27750, n27751, n27752, n27753,
         n27754, n27755, n27756, n27757, n27758, n27759, n27760, n27761,
         n27762, n27763, n27764, n27765, n27766, n27767, n27768, n27769,
         n27770, n27771, n27772, n27773, n27774, n27775, n27776, n27777,
         n27778, n27779, n27780, n27781, n27782, n27783, n27784, n27785,
         n27786, n27787, n27788, n27789, n27790, n27791, n27792, n27793,
         n27794, n27795, n27796, n27797, n27798, n27799, n27800, n27801,
         n27802, n27803, n27804, n27805, n27806, n27807, n27808, n27809,
         n27810, n27811, n27812, n27813, n27814, n27815, n27816, n27817,
         n27818, n27819, n27820, n27821, n27822, n27823, n27824, n27825,
         n27826, n27827, n27828, n27829, n27830, n27831, n27832, n27833,
         n27834, n27835, n27836, n27837, n27838, n27839, n27840, n27841,
         n27842, n27843, n27844, n27845, n27846, n27847, n27848, n27849,
         n27850, n27851, n27852, n27853, n27854, n27855, n27856, n27857,
         n27858, n27859, n27860, n27861, n27862, n27863, n27864, n27865,
         n27866, n27867, n27868, n27869, n27870, n27871, n27872, n27873,
         n27874, n27875, n27876, n27877, n27878, n27879, n27880, n27881,
         n27882, n27883, n27884, n27885, n27886, n27887, n27888, n27889,
         n27890, n27891, n27892, n27893, n27894, n27895, n27896, n27897,
         n27898, n27899, n27900, n27901, n27902, n27903, n27904, n27905,
         n27906, n27907, n27908, n27909, n27910, n27911, n27912, n27913,
         n27914, n27915, n27916, n27917, n27918, n27919, n27920, n27921,
         n27922, n27923, n27924, n27925, n27926, n27927, n27928, n27929,
         n27930, n27931, n27932, n27933, n27934, n27935, n27936, n27937,
         n27938, n27939, n27940, n27941, n27942, n27943, n27944, n27945,
         n27946, n27947, n27948, n27949, n27950, n27951, n27952, n27953,
         n27954, n27955, n27956, n27957, n27958, n27959, n27960, n27961,
         n27962, n27963, n27964, n27965, n27966, n27967, n27968, n27969,
         n27970, n27971, n27972, n27973, n27974, n27975, n27976, n27977,
         n27978, n27979, n27980, n27981, n27982, n27983, n27984, n27985,
         n27986, n27987, n27988, n27989, n27990, n27991, n27992, n27993,
         n27994, n27995, n27996, n27997, n27998, n27999, n28000, n28001,
         n28002, n28003, n28004, n28005, n28006, n28007, n28008, n28009,
         n28010, n28011, n28012, n28013, n28014, n28015, n28016, n28017,
         n28018, n28019, n28020, n28021, n28022, n28023, n28024, n28025,
         n28026, n28027, n28028, n28029, n28030, n28031, n28032, n28033,
         n28034, n28035, n28036, n28037, n28038, n28039, n28040, n28041,
         n28042, n28043, n28044, n28045, n28046, n28047, n28048, n28049,
         n28050, n28051, n28052, n28053, n28054, n28055, n28056, n28057,
         n28058, n28059, n28060, n28061, n28062, n28063, n28064, n28065,
         n28066, n28067, n28068, n28069, n28070, n28071, n28072, n28073,
         n28074, n28075, n28076, n28077, n28078, n28079, n28080, n28081,
         n28082, n28083, n28084, n28085, n28086, n28087, n28088, n28089,
         n28090, n28091, n28092, n28093, n28094, n28095, n28096, n28097,
         n28098, n28099, n28100, n28101, n28102, n28103, n28104, n28105,
         n28106, n28107, n28108, n28109, n28110, n28111, n28112, n28113,
         n28114, n28115, n28116, n28117, n28118, n28119, n28120, n28121,
         n28122, n28123, n28124, n28125, n28126, n28127, n28128, n28129,
         n28130, n28131, n28132, n28133, n28134, n28135, n28136, n28137,
         n28138, n28139, n28140, n28141, n28142, n28143, n28144, n28145,
         n28146, n28147, n28148, n28149, n28150, n28151, n28152, n28153,
         n28154, n28155, n28156, n28157, n28158, n28159, n28160, n28161,
         n28162, n28163, n28164, n28165, n28166, n28167, n28168, n28169,
         n28170, n28171, n28172, n28173, n28174, n28175, n28176, n28177,
         n28178, n28179, n28180, n28181, n28182, n28183, n28184, n28185,
         n28186, n28187, n28188, n28189, n28190, n28191, n28192, n28193,
         n28194, n28195, n28196, n28197, n28198, n28199, n28200, n28201,
         n28202, n28203, n28204, n28205, n28206, n28207, n28208, n28209,
         n28210, n28211, n28212, n28213, n28214, n28215, n28216, n28217,
         n28218, n28219, n28220, n28221, n28222, n28223, n28224, n28225,
         n28226, n28227, n28228, n28229, n28230, n28231, n28232, n28233,
         n28234, n28235, n28236, n28237, n28238, n28239, n28240, n28241,
         n28242, n28243, n28244, n28245, n28246, n28247, n28248, n28249,
         n28250, n28251, n28252, n28253, n28254, n28255, n28256, n28257,
         n28258, n28259, n28260, n28261, n28262, n28263, n28264, n28265,
         n28266, n28267, n28268, n28269, n28270, n28271, n28272, n28273,
         n28274, n28275, n28276, n28277, n28278, n28279, n28280, n28281,
         n28282, n28283, n28284, n28285, n28286, n28287, n28288, n28289,
         n28290, n28291, n28292, n28293, n28294, n28295, n28296, n28297,
         n28298, n28299, n28300, n28301, n28302, n28303, n28304, n28305,
         n28306, n28307, n28308, n28309, n28310, n28311, n28312, n28313,
         n28314, n28315, n28316, n28317, n28318, n28319, n28320, n28321,
         n28322, n28323, n28324, n28325, n28326, n28327, n28328, n28329,
         n28330, n28331, n28332, n28333, n28334, n28335, n28336, n28337,
         n28338, n28339, n28340, n28341, n28342, n28343, n28344, n28345,
         n28346, n28347, n28348, n28349, n28350, n28351, n28352, n28353,
         n28354, n28355, n28356, n28357, n28358, n28359, n28360, n28361,
         n28362, n28363, n28364, n28365, n28366, n28367, n28368, n28369,
         n28370, n28371, n28372, n28373, n28374, n28375, n28376, n28377,
         n28378, n28379, n28380, n28381, n28382, n28383, n28384, n28385,
         n28386, n28387, n28388, n28389, n28390, n28391, n28392, n28393,
         n28394, n28395, n28396, n28397, n28398, n28399, n28400, n28401,
         n28402, n28403, n28404, n28405, n28406, n28407, n28408, n28409,
         n28410, n28411, n28412, n28413, n28414, n28415, n28416, n28417,
         n28418, n28419, n28420, n28421, n28422, n28423, n28424, n28425,
         n28426, n28427, n28428, n28429, n28430, n28431, n28432, n28433,
         n28434, n28435, n28436, n28437, n28438, n28439, n28440, n28441,
         n28442, n28443, n28444, n28445, n28446, n28447, n28448, n28449,
         n28450, n28451, n28452, n28453, n28454, n28455, n28456, n28457,
         n28458, n28459, n28460, n28461, n28462, n28463, n28464, n28465,
         n28466, n28467, n28468, n28469, n28470, n28471, n28472, n28473,
         n28474, n28475, n28476, n28477, n28478, n28479, n28480, n28481,
         n28482, n28483, n28484, n28485, n28486, n28487, n28488, n28489,
         n28490, n28491, n28492, n28493, n28494, n28495, n28496, n28497,
         n28498, n28499, n28500, n28501, n28502, n28503, n28504, n28505,
         n28506, n28507, n28508, n28509, n28510, n28511, n28512, n28513,
         n28514, n28515, n28516, n28517, n28518, n28519, n28520, n28521,
         n28522, n28523, n28524, n28525, n28526, n28527, n28528, n28529,
         n28530, n28531, n28532, n28533, n28534, n28535, n28536, n28537,
         n28538, n28539, n28540, n28541, n28542, n28543, n28544, n28545,
         n28546, n28547, n28548, n28549, n28550, n28551, n28552, n28553,
         n28554, n28555, n28556, n28557, n28558, n28559, n28560, n28561,
         n28562, n28563, n28564, n28565, n28566, n28567, n28568, n28569,
         n28570, n28571, n28572, n28573, n28574, n28575, n28576, n28577,
         n28578, n28579, n28580, n28581, n28582, n28583, n28584, n28585,
         n28586, n28587, n28588, n28589, n28590, n28591, n28592, n28593,
         n28594, n28595, n28596, n28597, n28598, n28599, n28600, n28601,
         n28602, n28603, n28604, n28605, n28606, n28607, n28608, n28609,
         n28610, n28611, n28612, n28613, n28614, n28615, n28616, n28617,
         n28618, n28619, n28620, n28621, n28622, n28623, n28624, n28625,
         n28626, n28627, n28628, n28629, n28630, n28631, n28632, n28633,
         n28634, n28635, n28636, n28637, n28638, n28639, n28640, n28641,
         n28642, n28643, n28644, n28645, n28646, n28647, n28648, n28649,
         n28650, n28651, n28652, n28653, n28654, n28655, n28656, n28657,
         n28658, n28659, n28660, n28661, n28662, n28663, n28664, n28665,
         n28666, n28667, n28668, n28669, n28670, n28671, n28672, n28673,
         n28674, n28675, n28676, n28677, n28678, n28679, n28680, n28681,
         n28682, n28683, n28684, n28685, n28686, n28687, n28688, n28689,
         n28690, n28691, n28692, n28693, n28694, n28695, n28696, n28697,
         n28698, n28699, n28700, n28701, n28702, n28703, n28704, n28705,
         n28706, n28707, n28708, n28709, n28710, n28711, n28712, n28713,
         n28714, n28715, n28716, n28717, n28718, n28719, n28720, n28721,
         n28722, n28723, n28724, n28725, n28726, n28727, n28728, n28729,
         n28730, n28731, n28732, n28733, n28734, n28735, n28736, n28737,
         n28738, n28739, n28740, n28741, n28742, n28743, n28744, n28745,
         n28746, n28747, n28748, n28749, n28750, n28751, n28752, n28753,
         n28754, n28755, n28756, n28757, n28758, n28759, n28760, n28761,
         n28762, n28763, n28764, n28765, n28766, n28767, n28768, n28769,
         n28770, n28771, n28772, n28773, n28774, n28775, n28776, n28777,
         n28778, n28779, n28780, n28781, n28782, n28783, n28784, n28785,
         n28786, n28787, n28788, n28789, n28790, n28791, n28792, n28793,
         n28794, n28795, n28796, n28797, n28798, n28799, n28800, n28801,
         n28802, n28803, n28804, n28805, n28806, n28807, n28808, n28809,
         n28810, n28811, n28812, n28813, n28814, n28815, n28816, n28817,
         n28818, n28819, n28820, n28821, n28822, n28823, n28824, n28825,
         n28826, n28827, n28828, n28829, n28830, n28831, n28832, n28833,
         n28834, n28835, n28836, n28837, n28838, n28839, n28840, n28841,
         n28842, n28843, n28844, n28845, n28846, n28847, n28848, n28849,
         n28850, n28851, n28852, n28853, n28854, n28855, n28856, n28857,
         n28858, n28859, n28860, n28861, n28862, n28863, n28864, n28865,
         n28866, n28867, n28868, n28869, n28870, n28871, n28872, n28873,
         n28874, n28875, n28876, n28877, n28878, n28879, n28880, n28881,
         n28882, n28883, n28884, n28885, n28886, n28887, n28888, n28889,
         n28890, n28891, n28892, n28893, n28894, n28895, n28896, n28897,
         n28898, n28899, n28900, n28901, n28902, n28903, n28904, n28905,
         n28906, n28907, n28908, n28909, n28910, n28911, n28912, n28913,
         n28914, n28915, n28916, n28917, n28918, n28919, n28920, n28921,
         n28922, n28923, n28924, n28925, n28926, n28927, n28928, n28929,
         n28930, n28931, n28932, n28933, n28934, n28935, n28936, n28937,
         n28938, n28939, n28940, n28941, n28942, n28943, n28944, n28945,
         n28946, n28947, n28948, n28949, n28950, n28951, n28952, n28953,
         n28954, n28955, n28956, n28957, n28958, n28959, n28960, n28961,
         n28962, n28963, n28964, n28965, n28966, n28967, n28968, n28969,
         n28970, n28971, n28972, n28973, n28974, n28975, n28976, n28977,
         n28978, n28979, n28980, n28981, n28982, n28983, n28984, n28985,
         n28986, n28987, n28988, n28989, n28990, n28991, n28992, n28993,
         n28994, n28995, n28996, n28997, n28998, n28999, n29000, n29001,
         n29002, n29003, n29004, n29005, n29006, n29007, n29008, n29009,
         n29010, n29011, n29012, n29013, n29014, n29015, n29016, n29017,
         n29018, n29019, n29020, n29021, n29022, n29023, n29024, n29025,
         n29026, n29027, n29028, n29029, n29030, n29031, n29032, n29033,
         n29034, n29035, n29036, n29037, n29038, n29039, n29040, n29041,
         n29042, n29043, n29044, n29045, n29046, n29047, n29048, n29049,
         n29050, n29051, n29052, n29053, n29054, n29055, n29056, n29057,
         n29058, n29059, n29060, n29061, n29062, n29063, n29064, n29065,
         n29066, n29067, n29068, n29069, n29070, n29071, n29072, n29073,
         n29074, n29075, n29076, n29077, n29078, n29079, n29080, n29081,
         n29082, n29083, n29084, n29085, n29086, n29087, n29088, n29089,
         n29090, n29091, n29092, n29093, n29094, n29095, n29096, n29097,
         n29098, n29099, n29100, n29101, n29102, n29103, n29104, n29105,
         n29106, n29107, n29108, n29109, n29110, n29111, n29112, n29113,
         n29114, n29115, n29116, n29117, n29118, n29119, n29120, n29121,
         n29122, n29123, n29124, n29125, n29126, n29127, n29128, n29129,
         n29130, n29131, n29132, n29133, n29134, n29135, n29136, n29137,
         n29138, n29139, n29140, n29141, n29142, n29143, n29144, n29145,
         n29146, n29147, n29148, n29149, n29150, n29151, n29152, n29153,
         n29154, n29155, n29156, n29157, n29158, n29159, n29160, n29161,
         n29162, n29163, n29164, n29165, n29166, n29167, n29168, n29169,
         n29170, n29171, n29172, n29173, n29174, n29175, n29176, n29177,
         n29178, n29179, n29180, n29181, n29182, n29183, n29184, n29185,
         n29186, n29187, n29188, n29189, n29190, n29191, n29192, n29193,
         n29194, n29195, n29196, n29197, n29198, n29199, n29200, n29201,
         n29202, n29203, n29204, n29205, n29206, n29207, n29208, n29209,
         n29210, n29211, n29212, n29213, n29214, n29215, n29216, n29217,
         n29218, n29219, n29220, n29221, n29222, n29223, n29224, n29225,
         n29226, n29227, n29228, n29229, n29230, n29231, n29232, n29233,
         n29234, n29235, n29236, n29237, n29238, n29239, n29240, n29241,
         n29242, n29243, n29244, n29245, n29246, n29247, n29248, n29249,
         n29250, n29251, n29252, n29253, n29254, n29255, n29256, n29257,
         n29258, n29259, n29260, n29261, n29262, n29263, n29264, n29265,
         n29266, n29267, n29268, n29269, n29270, n29271, n29272, n29273,
         n29274, n29275, n29276, n29277, n29278, n29279, n29280, n29281,
         n29282, n29283, n29284, n29285, n29286, n29287, n29288, n29289,
         n29290, n29291, n29292, n29293, n29294, n29295, n29296, n29297,
         n29298, n29299, n29300, n29301, n29302, n29303, n29304, n29305,
         n29306, n29307, n29308, n29309, n29310, n29311, n29312, n29313,
         n29314, n29315, n29316, n29317, n29318, n29319, n29320, n29321,
         n29322, n29323, n29324, n29325, n29326, n29327, n29328, n29329,
         n29330, n29331, n29332, n29333, n29334, n29335, n29336, n29337,
         n29338, n29339, n29340, n29341, n29342, n29343, n29344, n29345,
         n29346, n29347, n29348, n29349, n29350, n29351, n29352, n29353,
         n29354, n29355, n29356, n29357, n29358, n29359, n29360, n29361,
         n29362, n29363, n29364, n29365, n29366, n29367, n29368, n29369,
         n29370, n29371, n29372, n29373, n29374, n29375, n29376, n29377,
         n29378, n29379, n29380, n29381, n29382, n29383, n29384, n29385,
         n29386, n29387, n29388, n29389, n29390, n29391, n29392, n29393,
         n29394, n29395, n29396, n29397, n29398, n29399, n29400, n29401,
         n29402, n29403, n29404, n29405, n29406, n29407, n29408, n29409,
         n29410, n29411, n29412, n29413, n29414, n29415, n29416, n29417,
         n29418, n29419, n29420, n29421, n29422, n29423, n29424, n29425,
         n29426, n29427, n29428, n29429, n29430, n29431, n29432, n29433,
         n29434, n29435, n29436, n29437, n29438, n29439, n29440, n29441,
         n29442, n29443, n29444, n29445, n29446, n29447, n29448, n29449,
         n29450, n29451, n29452, n29453, n29454, n29455, n29456, n29457,
         n29458, n29459, n29460, n29461, n29462, n29463, n29464, n29465,
         n29466, n29467, n29468, n29469, n29470, n29471, n29472, n29473,
         n29474, n29475, n29476, n29477, n29478, n29479, n29480, n29481,
         n29482, n29483, n29484, n29485, n29486, n29487, n29488, n29489,
         n29490, n29491, n29492, n29493, n29494, n29495, n29496, n29497,
         n29498, n29499, n29500, n29501, n29502, n29503, n29504, n29505,
         n29506, n29507, n29508, n29509, n29510, n29511, n29512, n29513,
         n29514, n29515, n29516, n29517, n29518, n29519, n29520, n29521,
         n29522, n29523, n29524, n29525, n29526, n29527, n29528, n29529,
         n29530, n29531, n29532, n29533, n29534, n29535, n29536, n29537,
         n29538, n29539, n29540, n29541, n29542, n29543, n29544, n29545,
         n29546, n29547, n29548, n29549, n29550, n29551, n29552, n29553,
         n29554, n29555, n29556, n29557, n29558, n29559, n29560, n29561,
         n29562, n29563, n29564, n29565, n29566, n29567, n29568, n29569,
         n29570, n29571, n29572, n29573, n29574, n29575, n29576, n29577,
         n29578, n29579, n29580, n29581, n29582, n29583, n29584, n29585,
         n29586, n29587, n29588, n29589, n29590, n29591, n29592, n29593,
         n29594, n29595, n29596, n29597, n29598, n29599, n29600, n29601,
         n29602, n29603, n29604, n29605, n29606, n29607, n29608, n29609,
         n29610, n29611, n29612, n29613, n29614, n29615, n29616, n29617,
         n29618, n29619, n29620, n29621, n29622, n29623, n29624, n29625,
         n29626, n29627, n29628, n29629, n29630, n29631, n29632, n29633,
         n29634, n29635, n29636, n29637, n29638, n29639, n29640, n29641,
         n29642, n29643, n29644, n29645, n29646, n29647, n29648, n29649,
         n29650, n29651, n29652, n29653, n29654, n29655, n29656, n29657,
         n29658, n29659, n29660, n29661, n29662, n29663, n29664, n29665,
         n29666, n29667, n29668, n29669, n29670, n29671, n29672, n29673,
         n29674, n29675, n29676, n29677, n29678, n29679, n29680, n29681,
         n29682, n29683, n29684, n29685, n29686, n29687, n29688, n29689,
         n29690, n29691, n29692, n29693, n29694, n29695, n29696, n29697,
         n29698, n29699, n29700, n29701, n29702, n29703, n29704, n29705,
         n29706, n29707, n29708, n29709, n29710, n29711, n29712, n29713,
         n29714, n29715, n29716, n29717, n29718, n29719, n29720, n29721,
         n29722, n29723, n29724, n29725, n29726, n29727, n29728, n29729,
         n29730, n29731, n29732, n29733, n29734, n29735, n29736, n29737,
         n29738, n29739, n29740, n29741, n29742, n29743, n29744, n29745,
         n29746, n29747, n29748, n29749, n29750, n29751, n29752, n29753,
         n29754, n29755, n29756, n29757, n29758, n29759, n29760, n29761,
         n29762, n29763, n29764, n29765, n29766, n29767, n29768, n29769,
         n29770, n29771, n29772, n29773, n29774, n29775, n29776, n29777,
         n29778, n29779, n29780, n29781, n29782, n29783, n29784, n29785,
         n29786, n29787, n29788, n29789, n29790, n29791, n29792, n29793,
         n29794, n29795, n29796, n29797, n29798, n29799, n29800, n29801,
         n29802, n29803, n29804, n29805, n29806, n29807, n29808, n29809,
         n29810, n29811, n29812, n29813, n29814, n29815, n29816, n29817,
         n29818, n29819, n29820, n29821, n29822, n29823, n29824, n29825,
         n29826, n29827, n29828, n29829, n29830, n29831, n29832, n29833,
         n29834, n29835, n29836, n29837, n29838, n29839, n29840, n29841,
         n29842, n29843, n29844, n29845, n29846, n29847, n29848, n29849,
         n29850, n29851, n29852, n29853, n29854, n29855, n29856, n29857,
         n29858, n29859, n29860, n29861, n29862, n29863, n29864, n29865,
         n29866, n29867, n29868, n29869, n29870, n29871, n29872, n29873,
         n29874, n29875, n29876, n29877, n29878, n29879, n29880, n29881,
         n29882, n29883, n29884, n29885, n29886, n29887, n29888, n29889,
         n29890, n29891, n29892, n29893, n29894, n29895, n29896, n29897,
         n29898, n29899, n29900, n29901, n29902, n29903, n29904, n29905,
         n29906, n29907, n29908, n29909, n29910, n29911, n29912, n29913,
         n29914, n29915, n29916, n29917, n29918, n29919, n29920, n29921,
         n29922, n29923, n29924, n29925, n29926, n29927, n29928, n29929,
         n29930, n29931, n29932, n29933, n29934, n29935, n29936, n29937,
         n29938, n29939, n29940, n29941, n29942, n29943, n29944, n29945,
         n29946, n29947, n29948, n29949, n29950, n29951, n29952, n29953,
         n29954, n29955, n29956, n29957, n29958, n29959, n29960, n29961,
         n29962, n29963, n29964, n29965, n29966, n29967, n29968, n29969,
         n29970, n29971, n29972, n29973, n29974, n29975, n29976, n29977,
         n29978, n29979, n29980, n29981, n29982, n29983, n29984, n29985,
         n29986, n29987, n29988, n29989, n29990, n29991, n29992, n29993,
         n29994, n29995, n29996, n29997, n29998, n29999, n30000, n30001,
         n30002, n30003, n30004, n30005, n30006, n30007, n30008, n30009,
         n30010, n30011, n30012, n30013, n30014, n30015, n30016, n30017,
         n30018, n30019, n30020, n30021, n30022, n30023, n30024, n30025,
         n30026, n30027, n30028, n30029, n30030, n30031, n30032, n30033,
         n30034, n30035, n30036, n30037, n30038, n30039, n30040, n30041,
         n30042, n30043, n30044, n30045, n30046, n30047, n30048, n30049,
         n30050, n30051, n30052, n30053, n30054, n30055, n30056, n30057,
         n30058, n30059, n30060, n30061, n30062, n30063, n30064, n30065,
         n30066, n30067, n30068, n30069, n30070, n30071, n30072, n30073,
         n30074, n30075, n30076, n30077, n30078, n30079, n30080, n30081,
         n30082, n30083, n30084, n30085, n30086, n30087, n30088, n30089,
         n30090, n30091, n30092, n30093, n30094, n30095, n30096, n30097,
         n30098, n30099, n30100, n30101, n30102, n30103, n30104, n30105,
         n30106, n30107, n30108, n30109, n30110, n30111, n30112, n30113,
         n30114, n30115, n30116, n30117, n30118, n30119, n30120, n30121,
         n30122, n30123, n30124, n30125, n30126, n30127, n30128, n30129,
         n30130, n30131, n30132, n30133, n30134, n30135, n30136, n30137,
         n30138, n30139, n30140, n30141, n30142, n30143, n30144, n30145,
         n30146, n30147, n30148, n30149, n30150, n30151, n30152, n30153,
         n30154, n30155, n30156, n30157, n30158, n30159, n30160, n30161,
         n30162, n30163, n30164, n30165, n30166, n30167, n30168, n30169,
         n30170, n30171, n30172, n30173, n30174, n30175, n30176, n30177,
         n30178, n30179, n30180, n30181, n30182, n30183, n30184, n30185,
         n30186, n30187, n30188, n30189, n30190, n30191, n30192, n30193,
         n30194, n30195, n30196, n30197, n30198, n30199, n30200, n30201,
         n30202, n30203, n30204, n30205, n30206, n30207, n30208, n30209,
         n30210, n30211, n30212, n30213, n30214, n30215, n30216, n30217,
         n30218, n30219, n30220, n30221, n30222, n30223, n30224, n30225,
         n30226, n30227, n30228, n30229, n30230, n30231, n30232, n30233,
         n30234, n30235, n30236, n30237, n30238, n30239, n30240, n30241,
         n30242, n30243, n30244, n30245, n30246, n30247, n30248, n30249,
         n30250, n30251, n30252, n30253, n30254, n30255, n30256, n30257,
         n30258, n30259, n30260, n30261, n30262, n30263, n30264, n30265,
         n30266, n30267, n30268, n30269, n30270, n30271, n30272, n30273,
         n30274, n30275, n30276, n30277, n30278, n30279, n30280, n30281,
         n30282, n30283, n30284, n30285, n30286, n30287, n30288, n30289,
         n30290, n30291, n30292, n30293, n30294, n30295, n30296, n30297,
         n30298, n30299, n30300, n30301, n30302, n30303, n30304, n30305,
         n30306, n30307, n30308, n30309, n30310, n30311, n30312, n30313,
         n30314, n30315, n30316, n30317, n30318, n30319, n30320, n30321,
         n30322, n30323, n30324, n30325, n30326, n30327, n30328, n30329,
         n30330, n30331, n30332, n30333, n30334, n30335, n30336, n30337,
         n30338, n30339, n30340, n30341, n30342, n30343, n30344, n30345,
         n30346, n30347, n30348, n30349, n30350, n30351, n30352, n30353,
         n30354, n30355, n30356, n30357, n30358, n30359, n30360, n30361,
         n30362, n30363, n30364, n30365, n30366, n30367, n30368, n30369,
         n30370, n30371, n30372, n30373, n30374, n30375, n30376, n30377,
         n30378, n30379, n30380, n30381, n30382, n30383, n30384, n30385,
         n30386, n30387, n30388, n30389, n30390, n30391, n30392, n30393,
         n30394, n30395, n30396, n30397, n30398, n30399, n30400, n30401,
         n30402, n30403, n30404, n30405, n30406, n30407, n30408, n30409,
         n30410, n30411, n30412, n30413, n30414, n30415, n30416, n30417,
         n30418, n30419, n30420, n30421, n30422, n30423, n30424, n30425,
         n30426, n30427, n30428, n30429, n30430, n30431, n30432, n30433,
         n30434, n30435, n30436, n30437, n30438, n30439, n30440, n30441,
         n30442, n30443, n30444, n30445, n30446, n30447, n30448, n30449,
         n30450, n30451, n30452, n30453, n30454, n30455, n30456, n30457,
         n30458, n30459, n30460, n30461, n30462, n30463, n30464, n30465,
         n30466, n30467, n30468, n30469, n30470, n30471, n30472, n30473,
         n30474, n30475, n30476, n30477, n30478, n30479, n30480, n30481,
         n30482, n30483, n30484, n30485, n30486, n30487, n30488, n30489,
         n30490, n30491, n30492, n30493, n30494, n30495, n30496, n30497,
         n30498, n30499, n30500, n30501, n30502, n30503, n30504, n30505,
         n30506, n30507, n30508, n30509, n30510, n30511, n30512, n30513,
         n30514, n30515, n30516, n30517, n30518, n30519, n30520, n30521,
         n30522, n30523, n30524, n30525, n30526, n30527, n30528, n30529,
         n30530, n30531, n30532, n30533, n30534, n30535, n30536, n30537,
         n30538, n30539, n30540, n30541, n30542, n30543, n30544, n30545,
         n30546, n30547, n30548, n30549, n30550, n30551, n30552, n30553,
         n30554, n30555, n30556, n30557, n30558, n30559, n30560, n30561,
         n30562, n30563, n30564, n30565, n30566, n30567, n30568, n30569,
         n30570, n30571, n30572, n30573, n30574, n30575, n30576, n30577,
         n30578, n30579, n30580, n30581, n30582, n30583, n30584, n30585,
         n30586, n30587, n30588, n30589, n30590, n30591, n30592, n30593,
         n30594, n30595, n30596, n30597, n30598, n30599, n30600, n30601,
         n30602, n30603, n30604, n30605, n30606, n30607, n30608, n30609,
         n30610, n30611, n30612, n30613, n30614, n30615, n30616, n30617,
         n30618, n30619, n30620, n30621, n30622, n30623, n30624, n30625,
         n30626, n30627, n30628, n30629, n30630, n30631, n30632, n30633,
         n30634, n30635, n30636, n30637, n30638, n30639, n30640, n30641,
         n30642, n30643, n30644, n30645, n30646, n30647, n30648, n30649,
         n30650, n30651, n30652, n30653, n30654, n30655, n30656, n30657,
         n30658, n30659, n30660, n30661, n30662, n30663, n30664, n30665,
         n30666, n30667, n30668, n30669, n30670, n30671, n30672, n30673,
         n30674, n30675, n30676, n30677, n30678, n30679, n30680, n30681,
         n30682, n30683, n30684, n30685, n30686, n30687, n30688, n30689,
         n30690, n30691, n30692, n30693, n30694, n30695, n30696, n30697,
         n30698, n30699, n30700, n30701, n30702, n30703, n30704, n30705,
         n30706, n30707, n30708, n30709, n30710, n30711, n30712, n30713,
         n30714, n30715, n30716, n30717, n30718, n30719, n30720, n30721,
         n30722, n30723, n30724, n30725, n30726, n30727, n30728, n30729,
         n30730, n30731, n30732, n30733, n30734, n30735, n30736, n30737,
         n30738, n30739, n30740, n30741, n30742, n30743, n30744, n30745,
         n30746, n30747, n30748, n30749, n30750, n30751, n30752, n30753,
         n30754, n30755, n30756, n30757, n30758, n30759, n30760, n30761,
         n30762, n30763, n30764, n30765, n30766, n30767, n30768, n30769,
         n30770, n30771, n30772, n30773, n30774, n30775, n30776, n30777,
         n30778, n30779, n30780, n30781, n30782, n30783, n30784, n30785,
         n30786, n30787, n30788, n30789, n30790, n30791, n30792, n30793,
         n30794, n30795, n30796, n30797, n30798, n30799, n30800, n30801,
         n30802, n30803, n30804, n30805, n30806, n30807, n30808, n30809,
         n30810, n30811, n30812, n30813, n30814, n30815, n30816, n30817,
         n30818, n30819, n30820, n30821, n30822, n30823, n30824, n30825,
         n30826, n30827, n30828, n30829, n30830, n30831, n30832, n30833,
         n30834, n30835, n30836, n30837, n30838, n30839, n30840, n30841,
         n30842, n30843, n30844, n30845, n30846, n30847, n30848, n30849,
         n30850, n30851, n30852, n30853, n30854, n30855, n30856, n30857,
         n30858, n30859, n30860, n30861, n30862, n30863, n30864, n30865,
         n30866, n30867, n30868, n30869, n30870, n30871, n30872, n30873,
         n30874, n30875, n30876, n30877, n30878, n30879, n30880, n30881,
         n30882, n30883, n30884, n30885, n30886, n30887, n30888, n30889,
         n30890, n30891, n30892, n30893, n30894, n30895, n30896, n30897,
         n30898, n30899, n30900, n30901, n30902, n30903, n30904, n30905,
         n30906, n30907, n30908, n30909, n30910, n30911, n30912, n30913,
         n30914, n30915, n30916, n30917, n30918, n30919, n30920, n30921,
         n30922, n30923, n30924, n30925, n30926, n30927, n30928, n30929,
         n30930, n30931, n30932, n30933, n30934, n30935, n30936, n30937,
         n30938, n30939, n30940, n30941, n30942, n30943, n30944, n30945,
         n30946, n30947, n30948, n30949, n30950, n30951, n30952, n30953,
         n30954, n30955, n30956, n30957, n30958, n30959, n30960, n30961,
         n30962, n30963, n30964, n30965, n30966, n30967, n30968, n30969,
         n30970, n30971, n30972, n30973, n30974, n30975, n30976, n30977,
         n30978, n30979, n30980, n30981, n30982, n30983, n30984, n30985,
         n30986, n30987, n30988, n30989, n30990, n30991, n30992, n30993,
         n30994, n30995, n30996, n30997, n30998, n30999, n31000, n31001,
         n31002, n31003, n31004, n31005, n31006, n31007, n31008, n31009,
         n31010, n31011, n31012, n31013, n31014, n31015, n31016, n31017,
         n31018, n31019, n31020, n31021, n31022, n31023, n31024, n31025,
         n31026, n31027, n31028, n31029, n31030, n31031, n31032, n31033,
         n31034, n31035, n31036, n31037, n31038, n31039, n31040, n31041,
         n31042, n31043, n31044, n31045, n31046, n31047, n31048, n31049,
         n31050, n31051, n31052, n31053, n31054, n31055, n31056, n31057,
         n31058, n31059, n31060, n31061, n31062, n31063, n31064, n31065,
         n31066, n31067, n31068, n31069, n31070, n31071, n31072, n31073,
         n31074, n31075, n31076, n31077, n31078, n31079, n31080, n31081,
         n31082, n31083, n31084, n31085, n31086, n31087, n31088, n31089,
         n31090, n31091, n31092, n31093, n31094, n31095, n31096, n31097,
         n31098, n31099, n31100, n31101, n31102, n31103, n31104, n31105,
         n31106, n31107, n31108, n31109, n31110, n31111, n31112, n31113,
         n31114, n31115, n31116, n31117, n31118, n31119, n31120, n31121,
         n31122, n31123, n31124, n31125, n31126, n31127, n31128, n31129,
         n31130, n31131, n31132, n31133, n31134, n31135, n31136, n31137,
         n31138, n31139, n31140, n31141, n31142, n31143, n31144, n31145,
         n31146, n31147, n31148, n31149, n31150, n31151, n31152, n31153,
         n31154, n31155, n31156, n31157, n31158, n31159, n31160, n31161,
         n31162, n31163, n31164, n31165, n31166, n31167, n31168, n31169,
         n31170, n31171, n31172, n31173, n31174, n31175, n31176, n31177,
         n31178, n31179, n31180, n31181, n31182, n31183, n31184, n31185,
         n31186, n31187, n31188, n31189, n31190, n31191, n31192, n31193,
         n31194, n31195, n31196, n31197, n31198, n31199, n31200, n31201,
         n31202, n31203, n31204, n31205, n31206, n31207, n31208, n31209,
         n31210, n31211, n31212, n31213, n31214, n31215, n31216, n31217,
         n31218, n31219, n31220, n31221, n31222, n31223, n31224, n31225,
         n31226, n31227, n31228, n31229, n31230, n31231, n31232, n31233,
         n31234, n31235, n31236, n31237, n31238, n31239, n31240, n31241,
         n31242, n31243, n31244, n31245, n31246, n31247, n31248, n31249,
         n31250, n31251, n31252, n31253, n31254, n31255, n31256, n31257,
         n31258, n31259, n31260, n31261, n31262, n31263, n31264, n31265,
         n31266, n31267, n31268, n31269, n31270, n31271, n31272, n31273,
         n31274, n31275, n31276, n31277, n31278, n31279, n31280, n31281,
         n31282, n31283, n31284, n31285, n31286, n31287, n31288, n31289,
         n31290, n31291, n31292, n31293, n31294, n31295, n31296, n31297,
         n31298, n31299, n31300, n31301, n31302, n31303, n31304, n31305,
         n31306, n31307, n31308, n31309, n31310, n31311, n31312, n31313,
         n31314, n31315, n31316, n31317, n31318, n31319, n31320, n31321,
         n31322, n31323, n31324, n31325, n31326, n31327, n31328, n31329,
         n31330, n31331, n31332, n31333, n31334, n31335, n31336, n31337,
         n31338, n31339, n31340, n31341, n31342, n31343, n31344, n31345,
         n31346, n31347, n31348, n31349, n31350, n31351, n31352, n31353,
         n31354, n31355, n31356, n31357, n31358, n31359, n31360, n31361,
         n31362, n31363, n31364, n31365, n31366, n31367, n31368, n31369,
         n31370, n31371, n31372, n31373, n31374, n31375, n31376, n31377,
         n31378, n31379, n31380, n31381, n31382, n31383, n31384, n31385,
         n31386, n31387, n31388, n31389, n31390, n31391, n31392, n31393,
         n31394, n31395, n31396, n31397, n31398, n31399, n31400, n31401,
         n31402, n31403, n31404, n31405, n31406, n31407, n31408, n31409,
         n31410, n31411, n31412, n31413, n31414, n31415, n31416, n31417,
         n31418, n31419, n31420, n31421, n31422, n31423, n31424, n31425,
         n31426, n31427, n31428, n31429, n31430, n31431, n31432, n31433,
         n31434, n31435, n31436, n31437, n31438, n31439, n31440, n31441,
         n31442, n31443, n31444, n31445, n31446, n31447, n31448, n31449,
         n31450, n31451, n31452, n31453, n31454, n31455, n31456, n31457,
         n31458, n31459, n31460, n31461, n31462, n31463, n31464, n31465,
         n31466, n31467, n31468, n31469, n31470, n31471, n31472, n31473,
         n31474, n31475, n31476, n31477, n31478, n31479, n31480, n31481,
         n31482, n31483, n31484, n31485, n31486, n31487, n31488, n31489,
         n31490, n31491, n31492, n31493, n31494, n31495, n31496, n31497,
         n31498, n31499, n31500, n31501, n31502, n31503, n31504, n31505,
         n31506, n31507, n31508, n31509, n31510, n31511, n31512, n31513,
         n31514, n31515, n31516, n31517, n31518, n31519, n31520, n31521,
         n31522, n31523, n31524, n31525, n31526, n31527, n31528, n31529,
         n31530, n31531, n31532, n31533, n31534, n31535, n31536, n31537,
         n31538, n31539, n31540, n31541, n31542, n31543, n31544, n31545,
         n31546, n31547, n31548, n31549, n31550, n31551, n31552, n31553,
         n31554, n31555, n31556, n31557, n31558, n31559, n31560, n31561,
         n31562, n31563, n31564, n31565, n31566, n31567, n31568, n31569,
         n31570, n31571, n31572, n31573, n31574, n31575, n31576, n31577,
         n31578, n31579, n31580, n31581, n31582, n31583, n31584, n31585,
         n31586, n31587, n31588, n31589, n31590, n31591, n31592, n31593,
         n31594, n31595, n31596, n31597, n31598, n31599, n31600, n31601,
         n31602, n31603, n31604, n31605, n31606, n31607, n31608, n31609,
         n31610, n31611, n31612, n31613, n31614, n31615, n31616, n31617,
         n31618, n31619, n31620, n31621, n31622, n31623, n31624, n31625,
         n31626, n31627, n31628, n31629, n31630, n31631, n31632, n31633,
         n31634, n31635, n31636, n31637, n31638, n31639, n31640, n31641,
         n31642, n31643, n31644, n31645, n31646, n31647, n31648, n31649,
         n31650, n31651, n31652, n31653, n31654, n31655, n31656, n31657,
         n31658, n31659, n31660, n31661, n31662, n31663, n31664, n31665,
         n31666, n31667, n31668, n31669, n31670, n31671, n31672, n31673,
         n31674, n31675, n31676, n31677, n31678, n31679, n31680, n31681,
         n31682, n31683, n31684, n31685, n31686, n31687, n31688, n31689,
         n31690, n31691, n31692, n31693, n31694, n31695, n31696, n31697,
         n31698, n31699, n31700, n31701, n31702, n31703, n31704, n31705,
         n31706, n31707, n31708, n31709, n31710, n31711, n31712, n31713,
         n31714, n31715, n31716, n31717, n31718, n31719, n31720, n31721,
         n31722, n31723, n31724, n31725, n31726, n31727, n31728, n31729,
         n31730, n31731, n31732, n31733, n31734, n31735, n31736, n31737,
         n31738, n31739, n31740, n31741, n31742, n31743, n31744, n31745,
         n31746, n31747, n31748, n31749, n31750, n31751, n31752, n31753,
         n31754, n31755, n31756, n31757, n31758, n31759, n31760, n31761,
         n31762, n31763, n31764, n31765, n31766, n31767, n31768, n31769,
         n31770, n31771, n31772, n31773, n31774, n31775, n31776, n31777,
         n31778, n31779, n31780, n31781, n31782, n31783, n31784, n31785,
         n31786, n31787, n31788, n31789, n31790, n31791, n31792, n31793,
         n31794, n31795, n31796, n31797, n31798, n31799, n31800, n31801,
         n31802, n31803, n31804, n31805, n31806, n31807, n31808, n31809,
         n31810, n31811, n31812, n31813, n31814, n31815, n31816, n31817,
         n31818, n31819, n31820, n31821, n31822, n31823, n31824, n31825,
         n31826, n31827, n31828, n31829, n31830, n31831, n31832, n31833,
         n31834, n31835, n31836, n31837, n31838, n31839, n31840, n31841,
         n31842, n31843, n31844, n31845, n31846, n31847, n31848, n31849,
         n31850, n31851, n31852, n31853, n31854, n31855, n31856, n31857,
         n31858, n31859, n31860, n31861, n31862, n31863, n31864, n31865,
         n31866, n31867, n31868, n31869, n31870, n31871, n31872, n31873,
         n31874, n31875, n31876, n31877, n31878, n31879, n31880, n31881,
         n31882, n31883, n31884, n31885, n31886, n31887, n31888, n31889,
         n31890, n31891, n31892, n31893, n31894, n31895, n31896, n31897,
         n31898, n31899, n31900, n31901, n31902, n31903, n31904, n31905,
         n31906, n31907, n31908, n31909, n31910, n31911, n31912, n31913,
         n31914, n31915, n31916, n31917, n31918, n31919, n31920, n31921,
         n31922, n31923, n31924, n31925, n31926, n31927, n31928, n31929,
         n31930, n31931, n31932, n31933, n31934, n31935, n31936, n31937,
         n31938, n31939, n31940, n31941, n31942, n31943, n31944, n31945,
         n31946, n31947, n31948, n31949, n31950, n31951, n31952, n31953,
         n31954, n31955, n31956, n31957, n31958, n31959, n31960, n31961,
         n31962, n31963, n31964, n31965, n31966, n31967, n31968, n31969,
         n31970, n31971, n31972, n31973, n31974, n31975, n31976, n31977,
         n31978, n31979, n31980, n31981, n31982, n31983, n31984, n31985,
         n31986, n31987, n31988, n31989, n31990, n31991, n31992, n31993,
         n31994, n31995, n31996, n31997, n31998, n31999, n32000, n32001,
         n32002, n32003, n32004, n32005, n32006, n32007, n32008, n32009,
         n32010, n32011, n32012, n32013, n32014, n32015, n32016, n32017,
         n32018, n32019, n32020, n32021, n32022, n32023, n32024, n32025,
         n32026, n32027, n32028, n32029, n32030, n32031, n32032, n32033,
         n32034, n32035, n32036, n32037, n32038, n32039, n32040, n32041,
         n32042, n32043, n32044, n32045, n32046, n32047, n32048, n32049,
         n32050, n32051, n32052, n32053, n32054, n32055, n32056, n32057,
         n32058, n32059, n32060, n32061, n32062, n32063, n32064, n32065,
         n32066, n32067, n32068, n32069, n32070, n32071, n32072, n32073,
         n32074, n32075, n32076, n32077, n32078, n32079, n32080, n32081,
         n32082, n32083, n32084, n32085, n32086, n32087, n32088, n32089,
         n32090, n32091, n32092, n32093, n32094, n32095, n32096, n32097,
         n32098, n32099, n32100, n32101, n32102, n32103, n32104, n32105,
         n32106, n32107, n32108, n32109, n32110, n32111, n32112, n32113,
         n32114, n32115, n32116, n32117, n32118, n32119, n32120, n32121,
         n32122, n32123, n32124, n32125, n32126, n32127, n32128, n32129,
         n32130, n32131, n32132, n32133, n32134, n32135, n32136, n32137,
         n32138, n32139, n32140, n32141, n32142, n32143, n32144, n32145,
         n32146, n32147, n32148, n32149, n32150, n32151, n32152, n32153,
         n32154, n32155, n32156, n32157, n32158, n32159, n32160, n32161,
         n32162, n32163, n32164, n32165, n32166, n32167, n32168, n32169,
         n32170, n32171, n32172, n32173, n32174, n32175, n32176, n32177,
         n32178, n32179, n32180, n32181, n32182, n32183, n32184, n32185,
         n32186, n32187, n32188, n32189, n32190, n32191, n32192, n32193,
         n32194, n32195, n32196, n32197, n32198, n32199, n32200, n32201,
         n32202, n32203, n32204, n32205, n32206, n32207, n32208, n32209,
         n32210, n32211, n32212, n32213, n32214, n32215, n32216, n32217,
         n32218, n32219, n32220, n32221, n32222, n32223, n32224, n32225,
         n32226, n32227, n32228, n32229, n32230, n32231, n32232, n32233,
         n32234, n32235, n32236, n32237, n32238, n32239, n32240, n32241,
         n32242, n32243, n32244, n32245, n32246, n32247, n32248, n32249,
         n32250, n32251, n32252, n32253, n32254, n32255, n32256, n32257,
         n32258, n32259, n32260, n32261, n32262, n32263, n32264, n32265,
         n32266, n32267, n32268, n32269, n32270, n32271, n32272, n32273,
         n32274, n32275, n32276, n32277, n32278, n32279, n32280, n32281,
         n32282, n32283, n32284, n32285, n32286, n32287, n32288, n32289,
         n32290, n32291, n32292, n32293, n32294, n32295, n32296, n32297,
         n32298, n32299, n32300, n32301, n32302, n32303, n32304, n32305,
         n32306, n32307, n32308, n32309, n32310, n32311, n32312, n32313,
         n32314, n32315, n32316, n32317, n32318, n32319, n32320, n32321,
         n32322, n32323, n32324, n32325, n32326, n32327, n32328, n32329,
         n32330, n32331, n32332, n32333, n32334, n32335, n32336, n32337,
         n32338, n32339, n32340, n32341, n32342, n32343, n32344, n32345,
         n32346, n32347, n32348, n32349, n32350, n32351, n32352, n32353,
         n32354, n32355, n32356, n32357, n32358, n32359, n32360, n32361,
         n32362, n32363, n32364, n32365, n32366, n32367, n32368, n32369,
         n32370, n32371, n32372, n32373, n32374, n32375, n32376, n32377,
         n32378, n32379, n32380, n32381, n32382, n32383, n32384, n32385,
         n32386, n32387, n32388, n32389, n32390, n32391, n32392, n32393,
         n32394, n32395, n32396, n32397, n32398, n32399, n32400, n32401,
         n32402, n32403, n32404, n32405, n32406, n32407, n32408, n32409,
         n32410, n32411, n32412, n32413, n32414, n32415, n32416, n32417,
         n32418, n32419, n32420, n32421, n32422, n32423, n32424, n32425,
         n32426, n32427, n32428, n32429, n32430, n32431, n32432, n32433,
         n32434, n32435, n32436, n32437, n32438, n32439, n32440, n32441,
         n32442, n32443, n32444, n32445, n32446, n32447, n32448, n32449,
         n32450, n32451, n32452, n32453, n32454, n32455, n32456, n32457,
         n32458, n32459, n32460, n32461, n32462, n32463, n32464, n32465,
         n32466, n32467, n32468, n32469, n32470, n32471, n32472, n32473,
         n32474, n32475, n32476, n32477, n32478, n32479, n32480, n32481,
         n32482, n32483, n32484, n32485, n32486, n32487, n32488, n32489,
         n32490, n32491, n32492, n32493, n32494, n32495, n32496, n32497,
         n32498, n32499, n32500, n32501, n32502, n32503, n32504, n32505,
         n32506, n32507, n32508, n32509, n32510, n32511, n32512, n32513,
         n32514, n32515, n32516, n32517, n32518, n32519, n32520, n32521,
         n32522, n32523, n32524, n32525, n32526, n32527, n32528, n32529,
         n32530, n32531, n32532, n32533, n32534, n32535, n32536, n32537,
         n32538, n32539, n32540, n32541, n32542, n32543, n32544, n32545,
         n32546, n32547, n32548, n32549, n32550, n32551, n32552, n32553,
         n32554, n32555, n32556, n32557, n32558, n32559, n32560, n32561,
         n32562, n32563, n32564, n32565, n32566, n32567, n32568, n32569,
         n32570, n32571, n32572, n32573, n32574, n32575, n32576, n32577,
         n32578, n32579, n32580, n32581, n32582, n32583, n32584, n32585,
         n32586, n32587, n32588, n32589, n32590, n32591, n32592, n32593,
         n32594, n32595, n32596, n32597, n32598, n32599, n32600, n32601,
         n32602, n32603, n32604, n32605, n32606, n32607, n32608, n32609,
         n32610, n32611, n32612, n32613, n32614, n32615, n32616, n32617,
         n32618, n32619, n32620, n32621, n32622, n32623, n32624, n32625,
         n32626, n32627, n32628, n32629, n32630, n32631, n32632, n32633,
         n32634, n32635, n32636, n32637, n32638, n32639, n32640, n32641,
         n32642, n32643, n32644, n32645, n32646, n32647, n32648, n32649,
         n32650, n32651, n32652, n32653, n32654, n32655, n32656, n32657,
         n32658, n32659, n32660, n32661, n32662, n32663, n32664, n32665,
         n32666, n32667, n32668, n32669, n32670, n32671, n32672, n32673,
         n32674, n32675, n32676, n32677, n32678, n32679, n32680, n32681,
         n32682, n32683, n32684, n32685, n32686, n32687, n32688, n32689,
         n32690, n32691, n32692, n32693, n32694, n32695, n32696, n32697,
         n32698, n32699, n32700, n32701, n32702, n32703, n32704, n32705,
         n32706, n32707, n32708, n32709, n32710, n32711, n32712, n32713,
         n32714, n32715, n32716, n32717, n32718, n32719, n32720, n32721,
         n32722, n32723, n32724, n32725, n32726, n32727, n32728, n32729,
         n32730, n32731, n32732, n32733, n32734, n32735, n32736, n32737,
         n32738, n32739, n32740, n32741, n32742, n32743, n32744, n32745,
         n32746, n32747, n32748, n32749, n32750, n32751, n32752, n32753,
         n32754, n32755, n32756, n32757, n32758, n32759, n32760, n32761,
         n32762, n32763, n32764, n32765, n32766, n32767, n32768, n32769,
         n32770, n32771, n32772, n32773, n32774, n32775, n32776, n32777,
         n32778, n32779, n32780, n32781, n32782, n32783, n32784, n32785,
         n32786, n32787, n32788, n32789, n32790, n32791, n32792, n32793,
         n32794, n32795, n32796, n32797, n32798, n32799, n32800, n32801,
         n32802, n32803, n32804, n32805, n32806, n32807, n32808, n32809,
         n32810, n32811, n32812, n32813, n32814, n32815, n32816, n32817,
         n32818, n32819, n32820, n32821, n32822, n32823, n32824, n32825,
         n32826, n32827, n32828, n32829, n32830, n32831, n32832, n32833,
         n32834, n32835, n32836, n32837, n32838, n32839, n32840, n32841,
         n32842, n32843, n32844, n32845, n32846, n32847, n32848, n32849,
         n32850, n32851, n32852, n32853, n32854, n32855, n32856, n32857,
         n32858, n32859, n32860, n32861, n32862, n32863, n32864, n32865,
         n32866, n32867, n32868, n32869, n32870, n32871, n32872, n32873,
         n32874, n32875, n32876, n32877, n32878, n32879, n32880, n32881,
         n32882, n32883, n32884, n32885, n32886, n32887, n32888, n32889,
         n32890, n32891, n32892, n32893, n32894, n32895, n32896, n32897,
         n32898, n32899, n32900, n32901, n32902, n32903, n32904, n32905,
         n32906, n32907, n32908, n32909, n32910, n32911, n32912, n32913,
         n32914, n32915, n32916, n32917, n32918, n32919, n32920, n32921,
         n32922, n32923, n32924, n32925, n32926, n32927, n32928, n32929,
         n32930, n32931, n32932, n32933, n32934, n32935, n32936, n32937,
         n32938, n32939, n32940, n32941, n32942, n32943, n32944, n32945,
         n32946, n32947, n32948, n32949, n32950, n32951, n32952, n32953,
         n32954, n32955, n32956, n32957, n32958, n32959, n32960, n32961,
         n32962, n32963, n32964, n32965, n32966, n32967, n32968, n32969,
         n32970, n32971, n32972, n32973, n32974, n32975, n32976, n32977,
         n32978, n32979, n32980, n32981, n32982, n32983, n32984, n32985,
         n32986, n32987, n32988, n32989, n32990, n32991, n32992, n32993,
         n32994, n32995, n32996, n32997, n32998, n32999, n33000, n33001,
         n33002, n33003, n33004, n33005, n33006, n33007, n33008, n33009,
         n33010, n33011, n33012, n33013, n33014, n33015, n33016, n33017,
         n33018, n33019, n33020, n33021, n33022, n33023, n33024, n33025,
         n33026, n33027, n33028, n33029, n33030, n33031, n33032, n33033,
         n33034, n33035, n33036, n33037, n33038, n33039, n33040, n33041,
         n33042, n33043, n33044, n33045, n33046, n33047, n33048, n33049,
         n33050, n33051, n33052, n33053, n33054, n33055, n33056, n33057,
         n33058, n33059, n33060, n33061, n33062, n33063, n33064, n33065,
         n33066, n33067, n33068, n33069, n33070, n33071, n33072, n33073,
         n33074, n33075, n33076, n33077, n33078, n33079, n33080, n33081,
         n33082, n33083, n33084, n33085, n33086, n33087, n33088, n33089,
         n33090, n33091, n33092, n33093, n33094, n33095, n33096, n33097,
         n33098, n33099, n33100, n33101, n33102, n33103, n33104, n33105,
         n33106, n33107, n33108, n33109, n33110, n33111, n33112, n33113,
         n33114, n33115, n33116, n33117, n33118, n33119, n33120, n33121,
         n33122, n33123, n33124, n33125, n33126, n33127, n33128, n33129,
         n33130, n33131, n33132, n33133, n33134, n33135, n33136, n33137,
         n33138, n33139, n33140, n33141, n33142, n33143, n33144, n33145,
         n33146, n33147, n33148, n33149, n33150, n33151, n33152, n33153,
         n33154, n33155, n33156, n33157, n33158, n33159, n33160, n33161,
         n33162, n33163, n33164, n33165, n33166, n33167, n33168, n33169,
         n33170, n33171, n33172, n33173, n33174, n33175, n33176, n33177,
         n33178, n33179, n33180, n33181, n33182, n33183, n33184, n33185,
         n33186, n33187, n33188, n33189, n33190, n33191, n33192, n33193,
         n33194, n33195, n33196, n33197, n33198, n33199, n33200, n33201,
         n33202, n33203, n33204, n33205, n33206, n33207, n33208, n33209,
         n33210, n33211, n33212, n33213, n33214, n33215, n33216, n33217,
         n33218, n33219, n33220, n33221, n33222, n33223, n33224, n33225,
         n33226, n33227, n33228, n33229, n33230, n33231, n33232, n33233,
         n33234, n33235, n33236, n33237, n33238, n33239, n33240, n33241,
         n33242, n33243, n33244, n33245, n33246, n33247, n33248, n33249,
         n33250, n33251, n33252, n33253, n33254, n33255, n33256, n33257,
         n33258, n33259, n33260, n33261, n33262, n33263, n33264, n33265,
         n33266, n33267, n33268, n33269, n33270, n33271, n33272, n33273,
         n33274, n33275, n33276, n33277, n33278, n33279, n33280, n33281,
         n33282, n33283, n33284, n33285, n33286, n33287, n33288, n33289,
         n33290, n33291, n33292, n33293, n33294, n33295, n33296, n33297,
         n33298, n33299, n33300, n33301, n33302, n33303, n33304, n33305,
         n33306, n33307, n33308, n33309, n33310, n33311, n33312, n33313,
         n33314, n33315, n33316, n33317, n33318, n33319, n33320, n33321,
         n33322, n33323, n33324, n33325, n33326, n33327, n33328, n33329,
         n33330, n33331, n33332, n33333, n33334, n33335, n33336, n33337,
         n33338, n33339, n33340, n33341, n33342, n33343, n33344, n33345,
         n33346, n33347, n33348, n33349, n33350, n33351, n33352, n33353,
         n33354, n33355, n33356, n33357, n33358, n33359, n33360, n33361,
         n33362, n33363, n33364, n33365, n33366, n33367, n33368, n33369,
         n33370, n33371, n33372, n33373, n33374, n33375, n33376, n33377,
         n33378, n33379, n33380, n33381, n33382, n33383, n33384, n33385,
         n33386, n33387, n33388, n33389, n33390, n33391, n33392, n33393,
         n33394, n33395, n33396, n33397, n33398, n33399, n33400, n33401,
         n33402, n33403, n33404, n33405, n33406, n33407, n33408, n33409,
         n33410, n33411, n33412, n33413, n33414, n33415, n33416, n33417,
         n33418, n33419, n33420, n33421, n33422, n33423, n33424, n33425,
         n33426, n33427, n33428, n33429, n33430, n33431, n33432, n33433,
         n33434, n33435, n33436, n33437, n33438, n33439, n33440, n33441,
         n33442, n33443, n33444, n33445, n33446, n33447, n33448, n33449,
         n33450, n33451, n33452, n33453, n33454, n33455, n33456, n33457,
         n33458, n33459, n33460, n33461, n33462, n33463, n33464, n33465,
         n33466, n33467, n33468, n33469, n33470, n33471, n33472, n33473,
         n33474, n33475, n33476, n33477, n33478, n33479, n33480, n33481,
         n33482, n33483, n33484, n33485, n33486, n33487, n33488, n33489,
         n33490, n33491, n33492, n33493, n33494, n33495, n33496, n33497,
         n33498, n33499, n33500, n33501, n33502, n33503, n33504, n33505,
         n33506, n33507, n33508, n33509, n33510, n33511, n33512, n33513,
         n33514, n33515, n33516, n33517, n33518, n33519, n33520, n33521,
         n33522, n33523, n33524, n33525, n33526, n33527, n33528, n33529,
         n33530, n33531, n33532, n33533, n33534, n33535, n33536, n33537,
         n33538, n33539, n33540, n33541, n33542, n33543, n33544, n33545,
         n33546, n33547, n33548, n33549, n33550, n33551, n33552, n33553,
         n33554, n33555, n33556, n33557, n33558, n33559, n33560, n33561,
         n33562, n33563, n33564, n33565, n33566, n33567, n33568, n33569,
         n33570, n33571, n33572, n33573, n33574, n33575, n33576, n33577,
         n33578, n33579, n33580, n33581, n33582, n33583, n33584, n33585,
         n33586, n33587, n33588, n33589, n33590, n33591, n33592, n33593,
         n33594, n33595, n33596, n33597, n33598, n33599, n33600, n33601,
         n33602, n33603, n33604, n33605, n33606, n33607, n33608, n33609,
         n33610, n33611, n33612, n33613, n33614, n33615, n33616, n33617,
         n33618, n33619, n33620, n33621, n33622, n33623, n33624, n33625,
         n33626, n33627, n33628, n33629, n33630, n33631, n33632, n33633,
         n33634, n33635, n33636, n33637, n33638, n33639, n33640, n33641,
         n33642, n33643, n33644, n33645, n33646, n33647, n33648, n33649,
         n33650, n33651, n33652, n33653, n33654, n33655, n33656, n33657,
         n33658, n33659, n33660, n33661, n33662, n33663, n33664, n33665,
         n33666, n33667, n33668, n33669, n33670, n33671, n33672, n33673,
         n33674, n33675, n33676, n33677, n33678, n33679, n33680, n33681,
         n33682, n33683, n33684, n33685, n33686, n33687, n33688, n33689,
         n33690, n33691, n33692, n33693, n33694, n33695, n33696, n33697,
         n33698, n33699, n33700, n33701, n33702, n33703, n33704, n33705,
         n33706, n33707, n33708, n33709, n33710, n33711, n33712, n33713,
         n33714, n33715, n33716, n33717, n33718, n33719, n33720, n33721,
         n33722, n33723, n33724, n33725, n33726, n33727, n33728, n33729,
         n33730, n33731, n33732, n33733, n33734, n33735, n33736, n33737,
         n33738, n33739, n33740, n33741, n33742, n33743, n33744, n33745,
         n33746, n33747, n33748, n33749, n33750, n33751, n33752, n33753,
         n33754, n33755, n33756, n33757, n33758, n33759, n33760, n33761,
         n33762, n33763, n33764, n33765, n33766, n33767, n33768, n33769,
         n33770, n33771, n33772, n33773, n33774, n33775, n33776, n33777,
         n33778, n33779, n33780, n33781, n33782, n33783, n33784, n33785,
         n33786, n33787, n33788, n33789, n33790, n33791, n33792, n33793,
         n33794, n33795, n33796, n33797, n33798, n33799, n33800, n33801,
         n33802, n33803, n33804, n33805, n33806, n33807, n33808, n33809,
         n33810, n33811, n33812, n33813, n33814, n33815, n33816, n33817,
         n33818, n33819, n33820, n33821, n33822, n33823, n33824, n33825,
         n33826, n33827, n33828, n33829, n33830, n33831, n33832, n33833,
         n33834, n33835, n33836, n33837, n33838, n33839, n33840, n33841,
         n33842, n33843, n33844, n33845, n33846, n33847, n33848, n33849,
         n33850, n33851, n33852, n33853, n33854, n33855, n33856, n33857,
         n33858, n33859, n33860, n33861, n33862, n33863, n33864, n33865,
         n33866, n33867, n33868, n33869, n33870, n33871, n33872, n33873,
         n33874, n33875, n33876, n33877, n33878, n33879, n33880, n33881,
         n33882, n33883, n33884, n33885, n33886, n33887, n33888, n33889,
         n33890, n33891, n33892, n33893, n33894, n33895, n33896, n33897,
         n33898, n33899, n33900, n33901, n33902, n33903, n33904, n33905,
         n33906, n33907, n33908, n33909, n33910, n33911, n33912, n33913,
         n33914, n33915, n33916, n33917, n33918, n33919, n33920, n33921,
         n33922, n33923, n33924, n33925, n33926, n33927, n33928, n33929,
         n33930, n33931, n33932, n33933, n33934, n33935, n33936, n33937,
         n33938, n33939, n33940, n33941, n33942, n33943, n33944, n33945,
         n33946, n33947, n33948, n33949, n33950, n33951, n33952, n33953,
         n33954, n33955, n33956, n33957, n33958, n33959, n33960, n33961,
         n33962, n33963, n33964, n33965, n33966, n33967, n33968, n33969,
         n33970, n33971, n33972, n33973, n33974, n33975, n33976, n33977,
         n33978, n33979, n33980, n33981, n33982, n33983, n33984, n33985,
         n33986, n33987, n33988, n33989, n33990, n33991, n33992, n33993,
         n33994, n33995, n33996, n33997, n33998, n33999, n34000, n34001,
         n34002, n34003, n34004, n34005, n34006, n34007, n34008, n34009,
         n34010, n34011, n34012, n34013, n34014, n34015, n34016, n34017,
         n34018, n34019, n34020, n34021, n34022, n34023, n34024, n34025,
         n34026, n34027, n34028, n34029, n34030, n34031, n34032, n34033,
         n34034, n34035, n34036, n34037, n34038, n34039, n34040, n34041,
         n34042, n34043, n34044, n34045, n34046, n34047, n34048, n34049,
         n34050, n34051, n34052, n34053, n34054, n34055, n34056, n34057,
         n34058, n34059, n34060, n34061, n34062, n34063, n34064, n34065,
         n34066, n34067, n34068, n34069, n34070, n34071, n34072, n34073,
         n34074, n34075, n34076, n34077, n34078, n34079, n34080, n34081,
         n34082, n34083, n34084, n34085, n34086, n34087, n34088, n34089,
         n34090, n34091, n34092, n34093, n34094, n34095, n34096, n34097,
         n34098, n34099, n34100, n34101, n34102, n34103, n34104, n34105,
         n34106, n34107, n34108, n34109, n34110, n34111, n34112, n34113,
         n34114, n34115, n34116, n34117, n34118, n34119, n34120, n34121,
         n34122, n34123, n34124, n34125, n34126, n34127, n34128, n34129,
         n34130, n34131, n34132, n34133, n34134, n34135, n34136, n34137,
         n34138, n34139, n34140, n34141, n34142, n34143, n34144, n34145,
         n34146, n34147, n34148, n34149, n34150, n34151, n34152, n34153,
         n34154, n34155, n34156, n34157, n34158, n34159, n34160, n34161,
         n34162, n34163, n34164, n34165, n34166, n34167, n34168, n34169,
         n34170, n34171, n34172, n34173, n34174, n34175, n34176, n34177,
         n34178, n34179, n34180, n34181, n34182, n34183, n34184, n34185,
         n34186, n34187, n34188, n34189, n34190, n34191, n34192, n34193,
         n34194, n34195, n34196, n34197, n34198, n34199, n34200, n34201,
         n34202, n34203, n34204, n34205, n34206, n34207, n34208, n34209,
         n34210, n34211, n34212, n34213, n34214, n34215, n34216, n34217,
         n34218, n34219, n34220, n34221, n34222, n34223, n34224, n34225,
         n34226, n34227, n34228, n34229, n34230, n34231, n34232, n34233,
         n34234, n34235, n34236, n34237, n34238, n34239, n34240, n34241,
         n34242, n34243, n34244, n34245, n34246, n34247, n34248, n34249,
         n34250, n34251, n34252, n34253, n34254, n34255, n34256, n34257,
         n34258, n34259, n34260, n34261, n34262, n34263, n34264, n34265,
         n34266, n34267, n34268, n34269, n34270, n34271, n34272, n34273,
         n34274, n34275, n34276, n34277, n34278, n34279, n34280, n34281,
         n34282, n34283, n34284, n34285, n34286, n34287, n34288, n34289,
         n34290, n34291, n34292, n34293, n34294, n34295, n34296, n34297,
         n34298, n34299, n34300, n34301, n34302, n34303, n34304, n34305,
         n34306, n34307, n34308, n34309, n34310, n34311, n34312, n34313,
         n34314, n34315, n34316, n34317, n34318, n34319, n34320, n34321,
         n34322, n34323, n34324, n34325, n34326, n34327, n34328, n34329,
         n34330, n34331, n34332, n34333, n34334, n34335, n34336, n34337,
         n34338, n34339, n34340, n34341, n34342, n34343, n34344, n34345,
         n34346, n34347, n34348, n34349, n34350, n34351, n34352, n34353,
         n34354, n34355, n34356, n34357, n34358, n34359, n34360, n34361,
         n34362, n34363, n34364, n34365, n34366, n34367, n34368, n34369,
         n34370, n34371, n34372, n34373, n34374, n34375, n34376, n34377,
         n34378, n34379, n34380, n34381, n34382, n34383, n34384, n34385,
         n34386, n34387, n34388, n34389, n34390, n34391, n34392, n34393,
         n34394, n34395, n34396, n34397, n34398, n34399, n34400, n34401,
         n34402, n34403, n34404, n34405, n34406, n34407, n34408, n34409,
         n34410, n34411, n34412, n34413, n34414, n34415, n34416, n34417,
         n34418, n34419, n34420, n34421, n34422, n34423, n34424, n34425,
         n34426, n34427, n34428, n34429, n34430, n34431, n34432, n34433,
         n34434, n34435, n34436, n34437, n34438, n34439, n34440, n34441,
         n34442, n34443, n34444, n34445, n34446, n34447, n34448, n34449,
         n34450, n34451, n34452, n34453, n34454, n34455, n34456, n34457,
         n34458, n34459, n34460, n34461, n34462, n34463, n34464, n34465,
         n34466, n34467, n34468, n34469, n34470, n34471, n34472, n34473,
         n34474, n34475, n34476, n34477, n34478, n34479, n34480, n34481,
         n34482, n34483, n34484, n34485, n34486, n34487, n34488, n34489,
         n34490, n34491, n34492, n34493, n34494, n34495, n34496, n34497,
         n34498, n34499, n34500, n34501, n34502, n34503, n34504, n34505,
         n34506, n34507, n34508, n34509, n34510, n34511, n34512, n34513,
         n34514, n34515, n34516, n34517, n34518, n34519, n34520, n34521,
         n34522, n34523, n34524, n34525, n34526, n34527, n34528, n34529,
         n34530, n34531, n34532, n34533, n34534, n34535, n34536, n34537,
         n34538, n34539, n34540, n34541, n34542, n34543, n34544, n34545,
         n34546, n34547, n34548, n34549, n34550, n34551, n34552, n34553,
         n34554, n34555, n34556, n34557, n34558, n34559, n34560, n34561,
         n34562, n34563, n34564, n34565, n34566, n34567, n34568, n34569,
         n34570, n34571, n34572, n34573, n34574, n34575, n34576, n34577,
         n34578, n34579, n34580, n34581, n34582, n34583, n34584, n34585,
         n34586, n34587, n34588, n34589, n34590, n34591, n34592, n34593,
         n34594, n34595, n34596, n34597, n34598, n34599, n34600, n34601,
         n34602, n34603, n34604, n34605, n34606, n34607, n34608, n34609,
         n34610, n34611, n34612, n34613, n34614, n34615, n34616, n34617,
         n34618, n34619, n34620, n34621, n34622, n34623, n34624, n34625,
         n34626, n34627, n34628, n34629, n34630, n34631, n34632, n34633,
         n34634, n34635, n34636, n34637, n34638, n34639, n34640, n34641,
         n34642, n34643, n34644, n34645, n34646, n34647, n34648, n34649,
         n34650, n34651, n34652, n34653, n34654, n34655, n34656, n34657,
         n34658, n34659, n34660, n34661, n34662, n34663, n34664, n34665,
         n34666, n34667, n34668, n34669, n34670, n34671, n34672, n34673,
         n34674, n34675, n34676, n34677, n34678, n34679, n34680, n34681,
         n34682, n34683, n34684, n34685, n34686, n34687, n34688, n34689,
         n34690, n34691, n34692, n34693, n34694, n34695, n34696, n34697,
         n34698, n34699, n34700, n34701, n34702, n34703, n34704, n34705,
         n34706, n34707, n34708, n34709, n34710, n34711, n34712, n34713,
         n34714, n34715, n34716, n34717, n34718, n34719, n34720, n34721,
         n34722, n34723, n34724, n34725, n34726, n34727, n34728, n34729,
         n34730, n34731, n34732, n34733, n34734, n34735, n34736, n34737,
         n34738, n34739, n34740, n34741, n34742, n34743, n34744, n34745,
         n34746, n34747, n34748, n34749, n34750, n34751, n34752, n34753,
         n34754, n34755, n34756, n34757, n34758, n34759, n34760, n34761,
         n34762, n34763, n34764, n34765, n34766, n34767, n34768, n34769,
         n34770, n34771, n34772, n34773, n34774, n34775, n34776, n34777,
         n34778, n34779, n34780, n34781, n34782, n34783, n34784, n34785,
         n34786, n34787, n34788, n34789, n34790, n34791, n34792, n34793,
         n34794, n34795, n34796, n34797, n34798, n34799, n34800, n34801,
         n34802, n34803, n34804, n34805, n34806, n34807, n34808, n34809,
         n34810, n34811, n34812, n34813, n34814, n34815, n34816, n34817,
         n34818, n34819, n34820, n34821, n34822, n34823, n34824, n34825,
         n34826, n34827, n34828, n34829, n34830, n34831, n34832, n34833,
         n34834, n34835, n34836, n34837, n34838, n34839, n34840, n34841,
         n34842, n34843, n34844, n34845, n34846, n34847, n34848, n34849,
         n34850, n34851, n34852, n34853, n34854, n34855, n34856, n34857,
         n34858, n34859, n34860, n34861, n34862, n34863, n34864, n34865,
         n34866, n34867, n34868, n34869, n34870, n34871, n34872, n34873,
         n34874, n34875, n34876, n34877, n34878, n34879, n34880, n34881,
         n34882, n34883, n34884, n34885, n34886, n34887, n34888, n34889,
         n34890, n34891, n34892, n34893, n34894, n34895, n34896, n34897,
         n34898, n34899, n34900, n34901, n34902, n34903, n34904, n34905,
         n34906, n34907, n34908, n34909, n34910, n34911, n34912, n34913,
         n34914, n34915, n34916, n34917, n34918, n34919, n34920, n34921,
         n34922, n34923, n34924, n34925, n34926, n34927, n34928, n34929,
         n34930, n34931, n34932, n34933, n34934, n34935, n34936, n34937,
         n34938, n34939, n34940, n34941, n34942, n34943, n34944, n34945,
         n34946, n34947, n34948, n34949, n34950, n34951, n34952, n34953,
         n34954, n34955, n34956, n34957, n34958, n34959, n34960, n34961,
         n34962, n34963, n34964, n34965, n34966, n34967, n34968, n34969,
         n34970, n34971, n34972, n34973, n34974, n34975, n34976, n34977,
         n34978, n34979, n34980, n34981, n34982, n34983, n34984, n34985,
         n34986, n34987, n34988, n34989, n34990, n34991, n34992, n34993,
         n34994, n34995, n34996, n34997, n34998, n34999, n35000, n35001,
         n35002, n35003, n35004, n35005, n35006, n35007, n35008, n35009,
         n35010, n35011, n35012, n35013, n35014, n35015, n35016, n35017,
         n35018, n35019, n35020, n35021, n35022, n35023, n35024, n35025,
         n35026, n35027, n35028, n35029, n35030, n35031, n35032, n35033,
         n35034, n35035, n35036, n35037, n35038, n35039, n35040, n35041,
         n35042, n35043, n35044, n35045, n35046, n35047, n35048, n35049,
         n35050, n35051, n35052, n35053, n35054, n35055, n35056, n35057,
         n35058, n35059, n35060, n35061, n35062, n35063, n35064, n35065,
         n35066, n35067, n35068, n35069, n35070, n35071, n35072, n35073,
         n35074, n35075, n35076, n35077, n35078, n35079, n35080, n35081,
         n35082, n35083, n35084, n35085, n35086, n35087, n35088, n35089,
         n35090, n35091, n35092, n35093, n35094, n35095, n35096, n35097,
         n35098, n35099, n35100, n35101, n35102, n35103, n35104, n35105,
         n35106, n35107, n35108, n35109, n35110, n35111, n35112, n35113,
         n35114, n35115, n35116, n35117, n35118, n35119, n35120, n35121,
         n35122, n35123, n35124, n35125, n35126, n35127, n35128, n35129,
         n35130, n35131, n35132, n35133, n35134, n35135, n35136, n35137,
         n35138, n35139, n35140, n35141, n35142, n35143, n35144, n35145,
         n35146, n35147, n35148, n35149, n35150, n35151, n35152, n35153,
         n35154, n35155, n35156, n35157, n35158, n35159, n35160, n35161,
         n35162, n35163, n35164, n35165, n35166, n35167, n35168, n35169,
         n35170, n35171, n35172, n35173, n35174, n35175, n35176, n35177,
         n35178, n35179, n35180, n35181, n35182, n35183, n35184, n35185,
         n35186, n35187, n35188, n35189, n35190, n35191, n35192, n35193,
         n35194, n35195, n35196, n35197, n35198, n35199, n35200, n35201,
         n35202, n35203, n35204, n35205, n35206, n35207, n35208, n35209,
         n35210, n35211, n35212, n35213, n35214, n35215, n35216, n35217,
         n35218, n35219, n35220, n35221, n35222, n35223, n35224, n35225,
         n35226, n35227, n35228, n35229, n35230, n35231, n35232, n35233,
         n35234, n35235, n35236, n35237, n35238, n35239, n35240, n35241,
         n35242, n35243, n35244, n35245, n35246, n35247, n35248, n35249,
         n35250, n35251, n35252, n35253, n35254, n35255, n35256, n35257,
         n35258, n35259, n35260, n35261, n35262, n35263, n35264, n35265,
         n35266, n35267, n35268, n35269, n35270, n35271, n35272, n35273,
         n35274, n35275, n35276, n35277, n35278, n35279, n35280, n35281,
         n35282, n35283, n35284, n35285, n35286, n35287, n35288, n35289,
         n35290, n35291, n35292, n35293, n35294, n35295, n35296, n35297,
         n35298, n35299, n35300, n35301, n35302, n35303, n35304, n35305,
         n35306, n35307, n35308, n35309, n35310, n35311, n35312, n35313,
         n35314, n35315, n35316, n35317, n35318, n35319, n35320, n35321,
         n35322, n35323, n35324, n35325, n35326, n35327, n35328, n35329,
         n35330, n35331, n35332, n35333, n35334, n35335, n35336, n35337,
         n35338, n35339, n35340, n35341, n35342, n35343, n35344, n35345,
         n35346, n35347, n35348, n35349, n35350, n35351, n35352, n35353,
         n35354, n35355, n35356, n35357, n35358, n35359, n35360, n35361,
         n35362, n35363, n35364, n35365, n35366, n35367, n35368, n35369,
         n35370, n35371, n35372, n35373, n35374, n35375, n35376, n35377,
         n35378, n35379, n35380, n35381, n35382, n35383, n35384, n35385,
         n35386, n35387, n35388, n35389, n35390, n35391, n35392, n35393,
         n35394, n35395, n35396, n35397, n35398, n35399, n35400, n35401,
         n35402, n35403, n35404, n35405, n35406, n35407, n35408, n35409,
         n35410, n35411, n35412, n35413, n35414, n35415, n35416, n35417,
         n35418, n35419, n35420, n35421, n35422, n35423, n35424, n35425,
         n35426, n35427, n35428, n35429, n35430, n35431, n35432, n35433,
         n35434, n35435, n35436, n35437, n35438, n35439, n35440, n35441,
         n35442, n35443, n35444, n35445, n35446, n35447, n35448, n35449,
         n35450, n35451, n35452, n35453, n35454, n35455, n35456, n35457,
         n35458, n35459, n35460, n35461, n35462, n35463, n35464, n35465,
         n35466, n35467, n35468, n35469, n35470, n35471, n35472, n35473,
         n35474, n35475, n35476, n35477, n35478, n35479, n35480, n35481,
         n35482, n35483, n35484, n35485, n35486, n35487, n35488, n35489,
         n35490, n35491, n35492, n35493, n35494, n35495, n35496, n35497,
         n35498, n35499, n35500, n35501, n35502, n35503, n35504, n35505,
         n35506, n35507, n35508, n35509, n35510, n35511, n35512, n35513,
         n35514, n35515, n35516, n35517, n35518, n35519, n35520, n35521,
         n35522, n35523, n35524, n35525, n35526, n35527, n35528, n35529,
         n35530, n35531, n35532, n35533, n35534, n35535, n35536, n35537,
         n35538, n35539, n35540, n35541, n35542, n35543, n35544, n35545,
         n35546, n35547, n35548, n35549, n35550, n35551, n35552, n35553,
         n35554, n35555, n35556, n35557, n35558, n35559, n35560, n35561,
         n35562, n35563, n35564, n35565, n35566, n35567, n35568, n35569,
         n35570, n35571, n35572, n35573, n35574, n35575, n35576, n35577,
         n35578, n35579, n35580, n35581, n35582, n35583, n35584, n35585,
         n35586, n35587, n35588, n35589, n35590, n35591, n35592, n35593,
         n35594, n35595, n35596, n35597, n35598, n35599, n35600, n35601,
         n35602, n35603, n35604, n35605, n35606, n35607, n35608, n35609,
         n35610, n35611, n35612, n35613, n35614, n35615, n35616, n35617,
         n35618, n35619, n35620, n35621, n35622, n35623, n35624, n35625,
         n35626, n35627, n35628, n35629, n35630, n35631, n35632, n35633,
         n35634, n35635, n35636, n35637, n35638, n35639, n35640, n35641,
         n35642, n35643, n35644, n35645, n35646, n35647, n35648, n35649,
         n35650, n35651, n35652, n35653, n35654, n35655, n35656, n35657,
         n35658, n35659, n35660, n35661, n35662, n35663, n35664, n35665,
         n35666, n35667, n35668, n35669, n35670, n35671, n35672, n35673,
         n35674, n35675, n35676, n35677, n35678, n35679, n35680, n35681,
         n35682, n35683, n35684, n35685, n35686, n35687, n35688, n35689,
         n35690, n35691, n35692, n35693, n35694, n35695, n35696, n35697,
         n35698, n35699, n35700, n35701, n35702, n35703, n35704, n35705,
         n35706, n35707, n35708, n35709, n35710, n35711, n35712, n35713,
         n35714, n35715, n35716, n35717, n35718, n35719, n35720, n35721,
         n35722, n35723, n35724, n35725, n35726, n35727, n35728, n35729,
         n35730, n35731, n35732, n35733, n35734, n35735, n35736, n35737,
         n35738, n35739, n35740, n35741, n35742, n35743, n35744, n35745,
         n35746, n35747, n35748, n35749, n35750, n35751, n35752, n35753,
         n35754, n35755, n35756, n35757, n35758, n35759, n35760, n35761,
         n35762, n35763, n35764, n35765, n35766, n35767, n35768, n35769,
         n35770, n35771, n35772, n35773, n35774, n35775, n35776, n35777,
         n35778, n35779, n35780, n35781, n35782, n35783, n35784, n35785,
         n35786, n35787, n35788, n35789, n35790, n35791, n35792, n35793,
         n35794, n35795, n35796, n35797, n35798, n35799, n35800, n35801,
         n35802, n35803, n35804, n35805, n35806, n35807, n35808, n35809,
         n35810, n35811, n35812, n35813, n35814, n35815, n35816, n35817,
         n35818, n35819, n35820, n35821, n35822, n35823, n35824, n35825,
         n35826, n35827, n35828, n35829, n35830, n35831, n35832, n35833,
         n35834, n35835, n35836, n35837, n35838, n35839, n35840, n35841,
         n35842, n35843, n35844, n35845, n35846, n35847, n35848, n35849,
         n35850, n35851, n35852, n35853, n35854, n35855, n35856, n35857,
         n35858, n35859, n35860, n35861, n35862, n35863, n35864, n35865,
         n35866, n35867, n35868, n35869, n35870, n35871, n35872, n35873,
         n35874, n35875, n35876, n35877, n35878, n35879, n35880, n35881,
         n35882, n35883, n35884, n35885, n35886, n35887, n35888, n35889,
         n35890, n35891, n35892, n35893, n35894, n35895, n35896, n35897,
         n35898, n35899, n35900, n35901, n35902, n35903, n35904, n35905,
         n35906, n35907, n35908, n35909, n35910, n35911, n35912, n35913,
         n35914, n35915, n35916, n35917, n35918, n35919, n35920, n35921,
         n35922, n35923, n35924, n35925, n35926, n35927, n35928, n35929,
         n35930, n35931, n35932, n35933, n35934, n35935, n35936, n35937,
         n35938, n35939, n35940, n35941, n35942, n35943, n35944, n35945,
         n35946, n35947, n35948, n35949, n35950, n35951, n35952, n35953,
         n35954, n35955, n35956, n35957, n35958, n35959, n35960, n35961,
         n35962, n35963, n35964, n35965, n35966, n35967, n35968, n35969,
         n35970, n35971, n35972, n35973, n35974, n35975, n35976, n35977,
         n35978, n35979, n35980, n35981, n35982, n35983, n35984, n35985,
         n35986, n35987, n35988, n35989, n35990, n35991, n35992, n35993,
         n35994, n35995, n35996, n35997, n35998, n35999, n36000, n36001,
         n36002, n36003, n36004, n36005, n36006, n36007, n36008, n36009,
         n36010, n36011, n36012, n36013, n36014, n36015, n36016, n36017,
         n36018, n36019, n36020, n36021, n36022, n36023, n36024, n36025,
         n36026, n36027, n36028, n36029, n36030, n36031, n36032, n36033,
         n36034, n36035, n36036, n36037, n36038, n36039, n36040, n36041,
         n36042, n36043, n36044, n36045, n36046, n36047, n36048, n36049,
         n36050, n36051, n36052, n36053, n36054, n36055, n36056, n36057,
         n36058, n36059, n36060, n36061, n36062, n36063, n36064, n36065,
         n36066, n36067, n36068, n36069, n36070, n36071, n36072, n36073,
         n36074, n36075, n36076, n36077, n36078, n36079, n36080, n36081,
         n36082, n36083, n36084, n36085, n36086, n36087, n36088, n36089,
         n36090, n36091, n36092, n36093, n36094, n36095, n36096, n36097,
         n36098, n36099, n36100, n36101, n36102, n36103, n36104, n36105,
         n36106, n36107, n36108, n36109, n36110, n36111, n36112, n36113,
         n36114, n36115, n36116, n36117, n36118, n36119, n36120, n36121,
         n36122, n36123, n36124, n36125, n36126, n36127, n36128, n36129,
         n36130, n36131, n36132, n36133, n36134, n36135, n36136, n36137,
         n36138, n36139, n36140, n36141, n36142, n36143, n36144, n36145,
         n36146, n36147, n36148, n36149, n36150, n36151, n36152, n36153,
         n36154, n36155, n36156, n36157, n36158, n36159, n36160, n36161,
         n36162, n36163, n36164, n36165, n36166, n36167, n36168, n36169,
         n36170, n36171, n36172, n36173, n36174, n36175, n36176, n36177,
         n36178, n36179, n36180, n36181, n36182, n36183, n36184, n36185,
         n36186, n36187, n36188, n36189, n36190, n36191, n36192, n36193,
         n36194, n36195, n36196, n36197, n36198, n36199, n36200, n36201,
         n36202, n36203, n36204, n36205, n36206, n36207, n36208, n36209,
         n36210, n36211, n36212, n36213, n36214, n36215, n36216, n36217,
         n36218, n36219, n36220, n36221, n36222, n36223, n36224, n36225,
         n36226, n36227, n36228, n36229, n36230, n36231, n36232, n36233,
         n36234, n36235, n36236, n36237, n36238, n36239, n36240, n36241,
         n36242, n36243, n36244, n36245, n36246, n36247, n36248, n36249,
         n36250, n36251, n36252, n36253, n36254, n36255, n36256, n36257,
         n36258, n36259, n36260, n36261, n36262, n36263, n36264, n36265,
         n36266, n36267, n36268, n36269, n36270, n36271, n36272, n36273,
         n36274, n36275, n36276, n36277, n36278, n36279, n36280, n36281,
         n36282, n36283, n36284, n36285, n36286, n36287, n36288, n36289,
         n36290, n36291, n36292, n36293, n36294, n36295, n36296, n36297;

  XOR U3585 ( .A(DB[3583]), .B(n1), .Z(min_val_out[6]) );
  AND U3586 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3587 ( .A(n4), .B(n5), .Z(n3) );
  XOR U3588 ( .A(DB[3583]), .B(DB[3576]), .Z(n5) );
  AND U3589 ( .A(n6), .B(n7), .Z(n4) );
  XOR U3590 ( .A(n8), .B(n9), .Z(n7) );
  XOR U3591 ( .A(DB[3576]), .B(DB[3569]), .Z(n9) );
  AND U3592 ( .A(n10), .B(n11), .Z(n8) );
  XOR U3593 ( .A(n12), .B(n13), .Z(n11) );
  XOR U3594 ( .A(DB[3569]), .B(DB[3562]), .Z(n13) );
  AND U3595 ( .A(n14), .B(n15), .Z(n12) );
  XOR U3596 ( .A(n16), .B(n17), .Z(n15) );
  XOR U3597 ( .A(DB[3562]), .B(DB[3555]), .Z(n17) );
  AND U3598 ( .A(n18), .B(n19), .Z(n16) );
  XOR U3599 ( .A(n20), .B(n21), .Z(n19) );
  XOR U3600 ( .A(DB[3555]), .B(DB[3548]), .Z(n21) );
  AND U3601 ( .A(n22), .B(n23), .Z(n20) );
  XOR U3602 ( .A(n24), .B(n25), .Z(n23) );
  XOR U3603 ( .A(DB[3548]), .B(DB[3541]), .Z(n25) );
  AND U3604 ( .A(n26), .B(n27), .Z(n24) );
  XOR U3605 ( .A(n28), .B(n29), .Z(n27) );
  XOR U3606 ( .A(DB[3541]), .B(DB[3534]), .Z(n29) );
  AND U3607 ( .A(n30), .B(n31), .Z(n28) );
  XOR U3608 ( .A(n32), .B(n33), .Z(n31) );
  XOR U3609 ( .A(DB[3534]), .B(DB[3527]), .Z(n33) );
  AND U3610 ( .A(n34), .B(n35), .Z(n32) );
  XOR U3611 ( .A(n36), .B(n37), .Z(n35) );
  XOR U3612 ( .A(DB[3527]), .B(DB[3520]), .Z(n37) );
  AND U3613 ( .A(n38), .B(n39), .Z(n36) );
  XOR U3614 ( .A(n40), .B(n41), .Z(n39) );
  XOR U3615 ( .A(DB[3520]), .B(DB[3513]), .Z(n41) );
  AND U3616 ( .A(n42), .B(n43), .Z(n40) );
  XOR U3617 ( .A(n44), .B(n45), .Z(n43) );
  XOR U3618 ( .A(DB[3513]), .B(DB[3506]), .Z(n45) );
  AND U3619 ( .A(n46), .B(n47), .Z(n44) );
  XOR U3620 ( .A(n48), .B(n49), .Z(n47) );
  XOR U3621 ( .A(DB[3506]), .B(DB[3499]), .Z(n49) );
  AND U3622 ( .A(n50), .B(n51), .Z(n48) );
  XOR U3623 ( .A(n52), .B(n53), .Z(n51) );
  XOR U3624 ( .A(DB[3499]), .B(DB[3492]), .Z(n53) );
  AND U3625 ( .A(n54), .B(n55), .Z(n52) );
  XOR U3626 ( .A(n56), .B(n57), .Z(n55) );
  XOR U3627 ( .A(DB[3492]), .B(DB[3485]), .Z(n57) );
  AND U3628 ( .A(n58), .B(n59), .Z(n56) );
  XOR U3629 ( .A(n60), .B(n61), .Z(n59) );
  XOR U3630 ( .A(DB[3485]), .B(DB[3478]), .Z(n61) );
  AND U3631 ( .A(n62), .B(n63), .Z(n60) );
  XOR U3632 ( .A(n64), .B(n65), .Z(n63) );
  XOR U3633 ( .A(DB[3478]), .B(DB[3471]), .Z(n65) );
  AND U3634 ( .A(n66), .B(n67), .Z(n64) );
  XOR U3635 ( .A(n68), .B(n69), .Z(n67) );
  XOR U3636 ( .A(DB[3471]), .B(DB[3464]), .Z(n69) );
  AND U3637 ( .A(n70), .B(n71), .Z(n68) );
  XOR U3638 ( .A(n72), .B(n73), .Z(n71) );
  XOR U3639 ( .A(DB[3464]), .B(DB[3457]), .Z(n73) );
  AND U3640 ( .A(n74), .B(n75), .Z(n72) );
  XOR U3641 ( .A(n76), .B(n77), .Z(n75) );
  XOR U3642 ( .A(DB[3457]), .B(DB[3450]), .Z(n77) );
  AND U3643 ( .A(n78), .B(n79), .Z(n76) );
  XOR U3644 ( .A(n80), .B(n81), .Z(n79) );
  XOR U3645 ( .A(DB[3450]), .B(DB[3443]), .Z(n81) );
  AND U3646 ( .A(n82), .B(n83), .Z(n80) );
  XOR U3647 ( .A(n84), .B(n85), .Z(n83) );
  XOR U3648 ( .A(DB[3443]), .B(DB[3436]), .Z(n85) );
  AND U3649 ( .A(n86), .B(n87), .Z(n84) );
  XOR U3650 ( .A(n88), .B(n89), .Z(n87) );
  XOR U3651 ( .A(DB[3436]), .B(DB[3429]), .Z(n89) );
  AND U3652 ( .A(n90), .B(n91), .Z(n88) );
  XOR U3653 ( .A(n92), .B(n93), .Z(n91) );
  XOR U3654 ( .A(DB[3429]), .B(DB[3422]), .Z(n93) );
  AND U3655 ( .A(n94), .B(n95), .Z(n92) );
  XOR U3656 ( .A(n96), .B(n97), .Z(n95) );
  XOR U3657 ( .A(DB[3422]), .B(DB[3415]), .Z(n97) );
  AND U3658 ( .A(n98), .B(n99), .Z(n96) );
  XOR U3659 ( .A(n100), .B(n101), .Z(n99) );
  XOR U3660 ( .A(DB[3415]), .B(DB[3408]), .Z(n101) );
  AND U3661 ( .A(n102), .B(n103), .Z(n100) );
  XOR U3662 ( .A(n104), .B(n105), .Z(n103) );
  XOR U3663 ( .A(DB[3408]), .B(DB[3401]), .Z(n105) );
  AND U3664 ( .A(n106), .B(n107), .Z(n104) );
  XOR U3665 ( .A(n108), .B(n109), .Z(n107) );
  XOR U3666 ( .A(DB[3401]), .B(DB[3394]), .Z(n109) );
  AND U3667 ( .A(n110), .B(n111), .Z(n108) );
  XOR U3668 ( .A(n112), .B(n113), .Z(n111) );
  XOR U3669 ( .A(DB[3394]), .B(DB[3387]), .Z(n113) );
  AND U3670 ( .A(n114), .B(n115), .Z(n112) );
  XOR U3671 ( .A(n116), .B(n117), .Z(n115) );
  XOR U3672 ( .A(DB[3387]), .B(DB[3380]), .Z(n117) );
  AND U3673 ( .A(n118), .B(n119), .Z(n116) );
  XOR U3674 ( .A(n120), .B(n121), .Z(n119) );
  XOR U3675 ( .A(DB[3380]), .B(DB[3373]), .Z(n121) );
  AND U3676 ( .A(n122), .B(n123), .Z(n120) );
  XOR U3677 ( .A(n124), .B(n125), .Z(n123) );
  XOR U3678 ( .A(DB[3373]), .B(DB[3366]), .Z(n125) );
  AND U3679 ( .A(n126), .B(n127), .Z(n124) );
  XOR U3680 ( .A(n128), .B(n129), .Z(n127) );
  XOR U3681 ( .A(DB[3366]), .B(DB[3359]), .Z(n129) );
  AND U3682 ( .A(n130), .B(n131), .Z(n128) );
  XOR U3683 ( .A(n132), .B(n133), .Z(n131) );
  XOR U3684 ( .A(DB[3359]), .B(DB[3352]), .Z(n133) );
  AND U3685 ( .A(n134), .B(n135), .Z(n132) );
  XOR U3686 ( .A(n136), .B(n137), .Z(n135) );
  XOR U3687 ( .A(DB[3352]), .B(DB[3345]), .Z(n137) );
  AND U3688 ( .A(n138), .B(n139), .Z(n136) );
  XOR U3689 ( .A(n140), .B(n141), .Z(n139) );
  XOR U3690 ( .A(DB[3345]), .B(DB[3338]), .Z(n141) );
  AND U3691 ( .A(n142), .B(n143), .Z(n140) );
  XOR U3692 ( .A(n144), .B(n145), .Z(n143) );
  XOR U3693 ( .A(DB[3338]), .B(DB[3331]), .Z(n145) );
  AND U3694 ( .A(n146), .B(n147), .Z(n144) );
  XOR U3695 ( .A(n148), .B(n149), .Z(n147) );
  XOR U3696 ( .A(DB[3331]), .B(DB[3324]), .Z(n149) );
  AND U3697 ( .A(n150), .B(n151), .Z(n148) );
  XOR U3698 ( .A(n152), .B(n153), .Z(n151) );
  XOR U3699 ( .A(DB[3324]), .B(DB[3317]), .Z(n153) );
  AND U3700 ( .A(n154), .B(n155), .Z(n152) );
  XOR U3701 ( .A(n156), .B(n157), .Z(n155) );
  XOR U3702 ( .A(DB[3317]), .B(DB[3310]), .Z(n157) );
  AND U3703 ( .A(n158), .B(n159), .Z(n156) );
  XOR U3704 ( .A(n160), .B(n161), .Z(n159) );
  XOR U3705 ( .A(DB[3310]), .B(DB[3303]), .Z(n161) );
  AND U3706 ( .A(n162), .B(n163), .Z(n160) );
  XOR U3707 ( .A(n164), .B(n165), .Z(n163) );
  XOR U3708 ( .A(DB[3303]), .B(DB[3296]), .Z(n165) );
  AND U3709 ( .A(n166), .B(n167), .Z(n164) );
  XOR U3710 ( .A(n168), .B(n169), .Z(n167) );
  XOR U3711 ( .A(DB[3296]), .B(DB[3289]), .Z(n169) );
  AND U3712 ( .A(n170), .B(n171), .Z(n168) );
  XOR U3713 ( .A(n172), .B(n173), .Z(n171) );
  XOR U3714 ( .A(DB[3289]), .B(DB[3282]), .Z(n173) );
  AND U3715 ( .A(n174), .B(n175), .Z(n172) );
  XOR U3716 ( .A(n176), .B(n177), .Z(n175) );
  XOR U3717 ( .A(DB[3282]), .B(DB[3275]), .Z(n177) );
  AND U3718 ( .A(n178), .B(n179), .Z(n176) );
  XOR U3719 ( .A(n180), .B(n181), .Z(n179) );
  XOR U3720 ( .A(DB[3275]), .B(DB[3268]), .Z(n181) );
  AND U3721 ( .A(n182), .B(n183), .Z(n180) );
  XOR U3722 ( .A(n184), .B(n185), .Z(n183) );
  XOR U3723 ( .A(DB[3268]), .B(DB[3261]), .Z(n185) );
  AND U3724 ( .A(n186), .B(n187), .Z(n184) );
  XOR U3725 ( .A(n188), .B(n189), .Z(n187) );
  XOR U3726 ( .A(DB[3261]), .B(DB[3254]), .Z(n189) );
  AND U3727 ( .A(n190), .B(n191), .Z(n188) );
  XOR U3728 ( .A(n192), .B(n193), .Z(n191) );
  XOR U3729 ( .A(DB[3254]), .B(DB[3247]), .Z(n193) );
  AND U3730 ( .A(n194), .B(n195), .Z(n192) );
  XOR U3731 ( .A(n196), .B(n197), .Z(n195) );
  XOR U3732 ( .A(DB[3247]), .B(DB[3240]), .Z(n197) );
  AND U3733 ( .A(n198), .B(n199), .Z(n196) );
  XOR U3734 ( .A(n200), .B(n201), .Z(n199) );
  XOR U3735 ( .A(DB[3240]), .B(DB[3233]), .Z(n201) );
  AND U3736 ( .A(n202), .B(n203), .Z(n200) );
  XOR U3737 ( .A(n204), .B(n205), .Z(n203) );
  XOR U3738 ( .A(DB[3233]), .B(DB[3226]), .Z(n205) );
  AND U3739 ( .A(n206), .B(n207), .Z(n204) );
  XOR U3740 ( .A(n208), .B(n209), .Z(n207) );
  XOR U3741 ( .A(DB[3226]), .B(DB[3219]), .Z(n209) );
  AND U3742 ( .A(n210), .B(n211), .Z(n208) );
  XOR U3743 ( .A(n212), .B(n213), .Z(n211) );
  XOR U3744 ( .A(DB[3219]), .B(DB[3212]), .Z(n213) );
  AND U3745 ( .A(n214), .B(n215), .Z(n212) );
  XOR U3746 ( .A(n216), .B(n217), .Z(n215) );
  XOR U3747 ( .A(DB[3212]), .B(DB[3205]), .Z(n217) );
  AND U3748 ( .A(n218), .B(n219), .Z(n216) );
  XOR U3749 ( .A(n220), .B(n221), .Z(n219) );
  XOR U3750 ( .A(DB[3205]), .B(DB[3198]), .Z(n221) );
  AND U3751 ( .A(n222), .B(n223), .Z(n220) );
  XOR U3752 ( .A(n224), .B(n225), .Z(n223) );
  XOR U3753 ( .A(DB[3198]), .B(DB[3191]), .Z(n225) );
  AND U3754 ( .A(n226), .B(n227), .Z(n224) );
  XOR U3755 ( .A(n228), .B(n229), .Z(n227) );
  XOR U3756 ( .A(DB[3191]), .B(DB[3184]), .Z(n229) );
  AND U3757 ( .A(n230), .B(n231), .Z(n228) );
  XOR U3758 ( .A(n232), .B(n233), .Z(n231) );
  XOR U3759 ( .A(DB[3184]), .B(DB[3177]), .Z(n233) );
  AND U3760 ( .A(n234), .B(n235), .Z(n232) );
  XOR U3761 ( .A(n236), .B(n237), .Z(n235) );
  XOR U3762 ( .A(DB[3177]), .B(DB[3170]), .Z(n237) );
  AND U3763 ( .A(n238), .B(n239), .Z(n236) );
  XOR U3764 ( .A(n240), .B(n241), .Z(n239) );
  XOR U3765 ( .A(DB[3170]), .B(DB[3163]), .Z(n241) );
  AND U3766 ( .A(n242), .B(n243), .Z(n240) );
  XOR U3767 ( .A(n244), .B(n245), .Z(n243) );
  XOR U3768 ( .A(DB[3163]), .B(DB[3156]), .Z(n245) );
  AND U3769 ( .A(n246), .B(n247), .Z(n244) );
  XOR U3770 ( .A(n248), .B(n249), .Z(n247) );
  XOR U3771 ( .A(DB[3156]), .B(DB[3149]), .Z(n249) );
  AND U3772 ( .A(n250), .B(n251), .Z(n248) );
  XOR U3773 ( .A(n252), .B(n253), .Z(n251) );
  XOR U3774 ( .A(DB[3149]), .B(DB[3142]), .Z(n253) );
  AND U3775 ( .A(n254), .B(n255), .Z(n252) );
  XOR U3776 ( .A(n256), .B(n257), .Z(n255) );
  XOR U3777 ( .A(DB[3142]), .B(DB[3135]), .Z(n257) );
  AND U3778 ( .A(n258), .B(n259), .Z(n256) );
  XOR U3779 ( .A(n260), .B(n261), .Z(n259) );
  XOR U3780 ( .A(DB[3135]), .B(DB[3128]), .Z(n261) );
  AND U3781 ( .A(n262), .B(n263), .Z(n260) );
  XOR U3782 ( .A(n264), .B(n265), .Z(n263) );
  XOR U3783 ( .A(DB[3128]), .B(DB[3121]), .Z(n265) );
  AND U3784 ( .A(n266), .B(n267), .Z(n264) );
  XOR U3785 ( .A(n268), .B(n269), .Z(n267) );
  XOR U3786 ( .A(DB[3121]), .B(DB[3114]), .Z(n269) );
  AND U3787 ( .A(n270), .B(n271), .Z(n268) );
  XOR U3788 ( .A(n272), .B(n273), .Z(n271) );
  XOR U3789 ( .A(DB[3114]), .B(DB[3107]), .Z(n273) );
  AND U3790 ( .A(n274), .B(n275), .Z(n272) );
  XOR U3791 ( .A(n276), .B(n277), .Z(n275) );
  XOR U3792 ( .A(DB[3107]), .B(DB[3100]), .Z(n277) );
  AND U3793 ( .A(n278), .B(n279), .Z(n276) );
  XOR U3794 ( .A(n280), .B(n281), .Z(n279) );
  XOR U3795 ( .A(DB[3100]), .B(DB[3093]), .Z(n281) );
  AND U3796 ( .A(n282), .B(n283), .Z(n280) );
  XOR U3797 ( .A(n284), .B(n285), .Z(n283) );
  XOR U3798 ( .A(DB[3093]), .B(DB[3086]), .Z(n285) );
  AND U3799 ( .A(n286), .B(n287), .Z(n284) );
  XOR U3800 ( .A(n288), .B(n289), .Z(n287) );
  XOR U3801 ( .A(DB[3086]), .B(DB[3079]), .Z(n289) );
  AND U3802 ( .A(n290), .B(n291), .Z(n288) );
  XOR U3803 ( .A(n292), .B(n293), .Z(n291) );
  XOR U3804 ( .A(DB[3079]), .B(DB[3072]), .Z(n293) );
  AND U3805 ( .A(n294), .B(n295), .Z(n292) );
  XOR U3806 ( .A(n296), .B(n297), .Z(n295) );
  XOR U3807 ( .A(DB[3072]), .B(DB[3065]), .Z(n297) );
  AND U3808 ( .A(n298), .B(n299), .Z(n296) );
  XOR U3809 ( .A(n300), .B(n301), .Z(n299) );
  XOR U3810 ( .A(DB[3065]), .B(DB[3058]), .Z(n301) );
  AND U3811 ( .A(n302), .B(n303), .Z(n300) );
  XOR U3812 ( .A(n304), .B(n305), .Z(n303) );
  XOR U3813 ( .A(DB[3058]), .B(DB[3051]), .Z(n305) );
  AND U3814 ( .A(n306), .B(n307), .Z(n304) );
  XOR U3815 ( .A(n308), .B(n309), .Z(n307) );
  XOR U3816 ( .A(DB[3051]), .B(DB[3044]), .Z(n309) );
  AND U3817 ( .A(n310), .B(n311), .Z(n308) );
  XOR U3818 ( .A(n312), .B(n313), .Z(n311) );
  XOR U3819 ( .A(DB[3044]), .B(DB[3037]), .Z(n313) );
  AND U3820 ( .A(n314), .B(n315), .Z(n312) );
  XOR U3821 ( .A(n316), .B(n317), .Z(n315) );
  XOR U3822 ( .A(DB[3037]), .B(DB[3030]), .Z(n317) );
  AND U3823 ( .A(n318), .B(n319), .Z(n316) );
  XOR U3824 ( .A(n320), .B(n321), .Z(n319) );
  XOR U3825 ( .A(DB[3030]), .B(DB[3023]), .Z(n321) );
  AND U3826 ( .A(n322), .B(n323), .Z(n320) );
  XOR U3827 ( .A(n324), .B(n325), .Z(n323) );
  XOR U3828 ( .A(DB[3023]), .B(DB[3016]), .Z(n325) );
  AND U3829 ( .A(n326), .B(n327), .Z(n324) );
  XOR U3830 ( .A(n328), .B(n329), .Z(n327) );
  XOR U3831 ( .A(DB[3016]), .B(DB[3009]), .Z(n329) );
  AND U3832 ( .A(n330), .B(n331), .Z(n328) );
  XOR U3833 ( .A(n332), .B(n333), .Z(n331) );
  XOR U3834 ( .A(DB[3009]), .B(DB[3002]), .Z(n333) );
  AND U3835 ( .A(n334), .B(n335), .Z(n332) );
  XOR U3836 ( .A(n336), .B(n337), .Z(n335) );
  XOR U3837 ( .A(DB[3002]), .B(DB[2995]), .Z(n337) );
  AND U3838 ( .A(n338), .B(n339), .Z(n336) );
  XOR U3839 ( .A(n340), .B(n341), .Z(n339) );
  XOR U3840 ( .A(DB[2995]), .B(DB[2988]), .Z(n341) );
  AND U3841 ( .A(n342), .B(n343), .Z(n340) );
  XOR U3842 ( .A(n344), .B(n345), .Z(n343) );
  XOR U3843 ( .A(DB[2988]), .B(DB[2981]), .Z(n345) );
  AND U3844 ( .A(n346), .B(n347), .Z(n344) );
  XOR U3845 ( .A(n348), .B(n349), .Z(n347) );
  XOR U3846 ( .A(DB[2981]), .B(DB[2974]), .Z(n349) );
  AND U3847 ( .A(n350), .B(n351), .Z(n348) );
  XOR U3848 ( .A(n352), .B(n353), .Z(n351) );
  XOR U3849 ( .A(DB[2974]), .B(DB[2967]), .Z(n353) );
  AND U3850 ( .A(n354), .B(n355), .Z(n352) );
  XOR U3851 ( .A(n356), .B(n357), .Z(n355) );
  XOR U3852 ( .A(DB[2967]), .B(DB[2960]), .Z(n357) );
  AND U3853 ( .A(n358), .B(n359), .Z(n356) );
  XOR U3854 ( .A(n360), .B(n361), .Z(n359) );
  XOR U3855 ( .A(DB[2960]), .B(DB[2953]), .Z(n361) );
  AND U3856 ( .A(n362), .B(n363), .Z(n360) );
  XOR U3857 ( .A(n364), .B(n365), .Z(n363) );
  XOR U3858 ( .A(DB[2953]), .B(DB[2946]), .Z(n365) );
  AND U3859 ( .A(n366), .B(n367), .Z(n364) );
  XOR U3860 ( .A(n368), .B(n369), .Z(n367) );
  XOR U3861 ( .A(DB[2946]), .B(DB[2939]), .Z(n369) );
  AND U3862 ( .A(n370), .B(n371), .Z(n368) );
  XOR U3863 ( .A(n372), .B(n373), .Z(n371) );
  XOR U3864 ( .A(DB[2939]), .B(DB[2932]), .Z(n373) );
  AND U3865 ( .A(n374), .B(n375), .Z(n372) );
  XOR U3866 ( .A(n376), .B(n377), .Z(n375) );
  XOR U3867 ( .A(DB[2932]), .B(DB[2925]), .Z(n377) );
  AND U3868 ( .A(n378), .B(n379), .Z(n376) );
  XOR U3869 ( .A(n380), .B(n381), .Z(n379) );
  XOR U3870 ( .A(DB[2925]), .B(DB[2918]), .Z(n381) );
  AND U3871 ( .A(n382), .B(n383), .Z(n380) );
  XOR U3872 ( .A(n384), .B(n385), .Z(n383) );
  XOR U3873 ( .A(DB[2918]), .B(DB[2911]), .Z(n385) );
  AND U3874 ( .A(n386), .B(n387), .Z(n384) );
  XOR U3875 ( .A(n388), .B(n389), .Z(n387) );
  XOR U3876 ( .A(DB[2911]), .B(DB[2904]), .Z(n389) );
  AND U3877 ( .A(n390), .B(n391), .Z(n388) );
  XOR U3878 ( .A(n392), .B(n393), .Z(n391) );
  XOR U3879 ( .A(DB[2904]), .B(DB[2897]), .Z(n393) );
  AND U3880 ( .A(n394), .B(n395), .Z(n392) );
  XOR U3881 ( .A(n396), .B(n397), .Z(n395) );
  XOR U3882 ( .A(DB[2897]), .B(DB[2890]), .Z(n397) );
  AND U3883 ( .A(n398), .B(n399), .Z(n396) );
  XOR U3884 ( .A(n400), .B(n401), .Z(n399) );
  XOR U3885 ( .A(DB[2890]), .B(DB[2883]), .Z(n401) );
  AND U3886 ( .A(n402), .B(n403), .Z(n400) );
  XOR U3887 ( .A(n404), .B(n405), .Z(n403) );
  XOR U3888 ( .A(DB[2883]), .B(DB[2876]), .Z(n405) );
  AND U3889 ( .A(n406), .B(n407), .Z(n404) );
  XOR U3890 ( .A(n408), .B(n409), .Z(n407) );
  XOR U3891 ( .A(DB[2876]), .B(DB[2869]), .Z(n409) );
  AND U3892 ( .A(n410), .B(n411), .Z(n408) );
  XOR U3893 ( .A(n412), .B(n413), .Z(n411) );
  XOR U3894 ( .A(DB[2869]), .B(DB[2862]), .Z(n413) );
  AND U3895 ( .A(n414), .B(n415), .Z(n412) );
  XOR U3896 ( .A(n416), .B(n417), .Z(n415) );
  XOR U3897 ( .A(DB[2862]), .B(DB[2855]), .Z(n417) );
  AND U3898 ( .A(n418), .B(n419), .Z(n416) );
  XOR U3899 ( .A(n420), .B(n421), .Z(n419) );
  XOR U3900 ( .A(DB[2855]), .B(DB[2848]), .Z(n421) );
  AND U3901 ( .A(n422), .B(n423), .Z(n420) );
  XOR U3902 ( .A(n424), .B(n425), .Z(n423) );
  XOR U3903 ( .A(DB[2848]), .B(DB[2841]), .Z(n425) );
  AND U3904 ( .A(n426), .B(n427), .Z(n424) );
  XOR U3905 ( .A(n428), .B(n429), .Z(n427) );
  XOR U3906 ( .A(DB[2841]), .B(DB[2834]), .Z(n429) );
  AND U3907 ( .A(n430), .B(n431), .Z(n428) );
  XOR U3908 ( .A(n432), .B(n433), .Z(n431) );
  XOR U3909 ( .A(DB[2834]), .B(DB[2827]), .Z(n433) );
  AND U3910 ( .A(n434), .B(n435), .Z(n432) );
  XOR U3911 ( .A(n436), .B(n437), .Z(n435) );
  XOR U3912 ( .A(DB[2827]), .B(DB[2820]), .Z(n437) );
  AND U3913 ( .A(n438), .B(n439), .Z(n436) );
  XOR U3914 ( .A(n440), .B(n441), .Z(n439) );
  XOR U3915 ( .A(DB[2820]), .B(DB[2813]), .Z(n441) );
  AND U3916 ( .A(n442), .B(n443), .Z(n440) );
  XOR U3917 ( .A(n444), .B(n445), .Z(n443) );
  XOR U3918 ( .A(DB[2813]), .B(DB[2806]), .Z(n445) );
  AND U3919 ( .A(n446), .B(n447), .Z(n444) );
  XOR U3920 ( .A(n448), .B(n449), .Z(n447) );
  XOR U3921 ( .A(DB[2806]), .B(DB[2799]), .Z(n449) );
  AND U3922 ( .A(n450), .B(n451), .Z(n448) );
  XOR U3923 ( .A(n452), .B(n453), .Z(n451) );
  XOR U3924 ( .A(DB[2799]), .B(DB[2792]), .Z(n453) );
  AND U3925 ( .A(n454), .B(n455), .Z(n452) );
  XOR U3926 ( .A(n456), .B(n457), .Z(n455) );
  XOR U3927 ( .A(DB[2792]), .B(DB[2785]), .Z(n457) );
  AND U3928 ( .A(n458), .B(n459), .Z(n456) );
  XOR U3929 ( .A(n460), .B(n461), .Z(n459) );
  XOR U3930 ( .A(DB[2785]), .B(DB[2778]), .Z(n461) );
  AND U3931 ( .A(n462), .B(n463), .Z(n460) );
  XOR U3932 ( .A(n464), .B(n465), .Z(n463) );
  XOR U3933 ( .A(DB[2778]), .B(DB[2771]), .Z(n465) );
  AND U3934 ( .A(n466), .B(n467), .Z(n464) );
  XOR U3935 ( .A(n468), .B(n469), .Z(n467) );
  XOR U3936 ( .A(DB[2771]), .B(DB[2764]), .Z(n469) );
  AND U3937 ( .A(n470), .B(n471), .Z(n468) );
  XOR U3938 ( .A(n472), .B(n473), .Z(n471) );
  XOR U3939 ( .A(DB[2764]), .B(DB[2757]), .Z(n473) );
  AND U3940 ( .A(n474), .B(n475), .Z(n472) );
  XOR U3941 ( .A(n476), .B(n477), .Z(n475) );
  XOR U3942 ( .A(DB[2757]), .B(DB[2750]), .Z(n477) );
  AND U3943 ( .A(n478), .B(n479), .Z(n476) );
  XOR U3944 ( .A(n480), .B(n481), .Z(n479) );
  XOR U3945 ( .A(DB[2750]), .B(DB[2743]), .Z(n481) );
  AND U3946 ( .A(n482), .B(n483), .Z(n480) );
  XOR U3947 ( .A(n484), .B(n485), .Z(n483) );
  XOR U3948 ( .A(DB[2743]), .B(DB[2736]), .Z(n485) );
  AND U3949 ( .A(n486), .B(n487), .Z(n484) );
  XOR U3950 ( .A(n488), .B(n489), .Z(n487) );
  XOR U3951 ( .A(DB[2736]), .B(DB[2729]), .Z(n489) );
  AND U3952 ( .A(n490), .B(n491), .Z(n488) );
  XOR U3953 ( .A(n492), .B(n493), .Z(n491) );
  XOR U3954 ( .A(DB[2729]), .B(DB[2722]), .Z(n493) );
  AND U3955 ( .A(n494), .B(n495), .Z(n492) );
  XOR U3956 ( .A(n496), .B(n497), .Z(n495) );
  XOR U3957 ( .A(DB[2722]), .B(DB[2715]), .Z(n497) );
  AND U3958 ( .A(n498), .B(n499), .Z(n496) );
  XOR U3959 ( .A(n500), .B(n501), .Z(n499) );
  XOR U3960 ( .A(DB[2715]), .B(DB[2708]), .Z(n501) );
  AND U3961 ( .A(n502), .B(n503), .Z(n500) );
  XOR U3962 ( .A(n504), .B(n505), .Z(n503) );
  XOR U3963 ( .A(DB[2708]), .B(DB[2701]), .Z(n505) );
  AND U3964 ( .A(n506), .B(n507), .Z(n504) );
  XOR U3965 ( .A(n508), .B(n509), .Z(n507) );
  XOR U3966 ( .A(DB[2701]), .B(DB[2694]), .Z(n509) );
  AND U3967 ( .A(n510), .B(n511), .Z(n508) );
  XOR U3968 ( .A(n512), .B(n513), .Z(n511) );
  XOR U3969 ( .A(DB[2694]), .B(DB[2687]), .Z(n513) );
  AND U3970 ( .A(n514), .B(n515), .Z(n512) );
  XOR U3971 ( .A(n516), .B(n517), .Z(n515) );
  XOR U3972 ( .A(DB[2687]), .B(DB[2680]), .Z(n517) );
  AND U3973 ( .A(n518), .B(n519), .Z(n516) );
  XOR U3974 ( .A(n520), .B(n521), .Z(n519) );
  XOR U3975 ( .A(DB[2680]), .B(DB[2673]), .Z(n521) );
  AND U3976 ( .A(n522), .B(n523), .Z(n520) );
  XOR U3977 ( .A(n524), .B(n525), .Z(n523) );
  XOR U3978 ( .A(DB[2673]), .B(DB[2666]), .Z(n525) );
  AND U3979 ( .A(n526), .B(n527), .Z(n524) );
  XOR U3980 ( .A(n528), .B(n529), .Z(n527) );
  XOR U3981 ( .A(DB[2666]), .B(DB[2659]), .Z(n529) );
  AND U3982 ( .A(n530), .B(n531), .Z(n528) );
  XOR U3983 ( .A(n532), .B(n533), .Z(n531) );
  XOR U3984 ( .A(DB[2659]), .B(DB[2652]), .Z(n533) );
  AND U3985 ( .A(n534), .B(n535), .Z(n532) );
  XOR U3986 ( .A(n536), .B(n537), .Z(n535) );
  XOR U3987 ( .A(DB[2652]), .B(DB[2645]), .Z(n537) );
  AND U3988 ( .A(n538), .B(n539), .Z(n536) );
  XOR U3989 ( .A(n540), .B(n541), .Z(n539) );
  XOR U3990 ( .A(DB[2645]), .B(DB[2638]), .Z(n541) );
  AND U3991 ( .A(n542), .B(n543), .Z(n540) );
  XOR U3992 ( .A(n544), .B(n545), .Z(n543) );
  XOR U3993 ( .A(DB[2638]), .B(DB[2631]), .Z(n545) );
  AND U3994 ( .A(n546), .B(n547), .Z(n544) );
  XOR U3995 ( .A(n548), .B(n549), .Z(n547) );
  XOR U3996 ( .A(DB[2631]), .B(DB[2624]), .Z(n549) );
  AND U3997 ( .A(n550), .B(n551), .Z(n548) );
  XOR U3998 ( .A(n552), .B(n553), .Z(n551) );
  XOR U3999 ( .A(DB[2624]), .B(DB[2617]), .Z(n553) );
  AND U4000 ( .A(n554), .B(n555), .Z(n552) );
  XOR U4001 ( .A(n556), .B(n557), .Z(n555) );
  XOR U4002 ( .A(DB[2617]), .B(DB[2610]), .Z(n557) );
  AND U4003 ( .A(n558), .B(n559), .Z(n556) );
  XOR U4004 ( .A(n560), .B(n561), .Z(n559) );
  XOR U4005 ( .A(DB[2610]), .B(DB[2603]), .Z(n561) );
  AND U4006 ( .A(n562), .B(n563), .Z(n560) );
  XOR U4007 ( .A(n564), .B(n565), .Z(n563) );
  XOR U4008 ( .A(DB[2603]), .B(DB[2596]), .Z(n565) );
  AND U4009 ( .A(n566), .B(n567), .Z(n564) );
  XOR U4010 ( .A(n568), .B(n569), .Z(n567) );
  XOR U4011 ( .A(DB[2596]), .B(DB[2589]), .Z(n569) );
  AND U4012 ( .A(n570), .B(n571), .Z(n568) );
  XOR U4013 ( .A(n572), .B(n573), .Z(n571) );
  XOR U4014 ( .A(DB[2589]), .B(DB[2582]), .Z(n573) );
  AND U4015 ( .A(n574), .B(n575), .Z(n572) );
  XOR U4016 ( .A(n576), .B(n577), .Z(n575) );
  XOR U4017 ( .A(DB[2582]), .B(DB[2575]), .Z(n577) );
  AND U4018 ( .A(n578), .B(n579), .Z(n576) );
  XOR U4019 ( .A(n580), .B(n581), .Z(n579) );
  XOR U4020 ( .A(DB[2575]), .B(DB[2568]), .Z(n581) );
  AND U4021 ( .A(n582), .B(n583), .Z(n580) );
  XOR U4022 ( .A(n584), .B(n585), .Z(n583) );
  XOR U4023 ( .A(DB[2568]), .B(DB[2561]), .Z(n585) );
  AND U4024 ( .A(n586), .B(n587), .Z(n584) );
  XOR U4025 ( .A(n588), .B(n589), .Z(n587) );
  XOR U4026 ( .A(DB[2561]), .B(DB[2554]), .Z(n589) );
  AND U4027 ( .A(n590), .B(n591), .Z(n588) );
  XOR U4028 ( .A(n592), .B(n593), .Z(n591) );
  XOR U4029 ( .A(DB[2554]), .B(DB[2547]), .Z(n593) );
  AND U4030 ( .A(n594), .B(n595), .Z(n592) );
  XOR U4031 ( .A(n596), .B(n597), .Z(n595) );
  XOR U4032 ( .A(DB[2547]), .B(DB[2540]), .Z(n597) );
  AND U4033 ( .A(n598), .B(n599), .Z(n596) );
  XOR U4034 ( .A(n600), .B(n601), .Z(n599) );
  XOR U4035 ( .A(DB[2540]), .B(DB[2533]), .Z(n601) );
  AND U4036 ( .A(n602), .B(n603), .Z(n600) );
  XOR U4037 ( .A(n604), .B(n605), .Z(n603) );
  XOR U4038 ( .A(DB[2533]), .B(DB[2526]), .Z(n605) );
  AND U4039 ( .A(n606), .B(n607), .Z(n604) );
  XOR U4040 ( .A(n608), .B(n609), .Z(n607) );
  XOR U4041 ( .A(DB[2526]), .B(DB[2519]), .Z(n609) );
  AND U4042 ( .A(n610), .B(n611), .Z(n608) );
  XOR U4043 ( .A(n612), .B(n613), .Z(n611) );
  XOR U4044 ( .A(DB[2519]), .B(DB[2512]), .Z(n613) );
  AND U4045 ( .A(n614), .B(n615), .Z(n612) );
  XOR U4046 ( .A(n616), .B(n617), .Z(n615) );
  XOR U4047 ( .A(DB[2512]), .B(DB[2505]), .Z(n617) );
  AND U4048 ( .A(n618), .B(n619), .Z(n616) );
  XOR U4049 ( .A(n620), .B(n621), .Z(n619) );
  XOR U4050 ( .A(DB[2505]), .B(DB[2498]), .Z(n621) );
  AND U4051 ( .A(n622), .B(n623), .Z(n620) );
  XOR U4052 ( .A(n624), .B(n625), .Z(n623) );
  XOR U4053 ( .A(DB[2498]), .B(DB[2491]), .Z(n625) );
  AND U4054 ( .A(n626), .B(n627), .Z(n624) );
  XOR U4055 ( .A(n628), .B(n629), .Z(n627) );
  XOR U4056 ( .A(DB[2491]), .B(DB[2484]), .Z(n629) );
  AND U4057 ( .A(n630), .B(n631), .Z(n628) );
  XOR U4058 ( .A(n632), .B(n633), .Z(n631) );
  XOR U4059 ( .A(DB[2484]), .B(DB[2477]), .Z(n633) );
  AND U4060 ( .A(n634), .B(n635), .Z(n632) );
  XOR U4061 ( .A(n636), .B(n637), .Z(n635) );
  XOR U4062 ( .A(DB[2477]), .B(DB[2470]), .Z(n637) );
  AND U4063 ( .A(n638), .B(n639), .Z(n636) );
  XOR U4064 ( .A(n640), .B(n641), .Z(n639) );
  XOR U4065 ( .A(DB[2470]), .B(DB[2463]), .Z(n641) );
  AND U4066 ( .A(n642), .B(n643), .Z(n640) );
  XOR U4067 ( .A(n644), .B(n645), .Z(n643) );
  XOR U4068 ( .A(DB[2463]), .B(DB[2456]), .Z(n645) );
  AND U4069 ( .A(n646), .B(n647), .Z(n644) );
  XOR U4070 ( .A(n648), .B(n649), .Z(n647) );
  XOR U4071 ( .A(DB[2456]), .B(DB[2449]), .Z(n649) );
  AND U4072 ( .A(n650), .B(n651), .Z(n648) );
  XOR U4073 ( .A(n652), .B(n653), .Z(n651) );
  XOR U4074 ( .A(DB[2449]), .B(DB[2442]), .Z(n653) );
  AND U4075 ( .A(n654), .B(n655), .Z(n652) );
  XOR U4076 ( .A(n656), .B(n657), .Z(n655) );
  XOR U4077 ( .A(DB[2442]), .B(DB[2435]), .Z(n657) );
  AND U4078 ( .A(n658), .B(n659), .Z(n656) );
  XOR U4079 ( .A(n660), .B(n661), .Z(n659) );
  XOR U4080 ( .A(DB[2435]), .B(DB[2428]), .Z(n661) );
  AND U4081 ( .A(n662), .B(n663), .Z(n660) );
  XOR U4082 ( .A(n664), .B(n665), .Z(n663) );
  XOR U4083 ( .A(DB[2428]), .B(DB[2421]), .Z(n665) );
  AND U4084 ( .A(n666), .B(n667), .Z(n664) );
  XOR U4085 ( .A(n668), .B(n669), .Z(n667) );
  XOR U4086 ( .A(DB[2421]), .B(DB[2414]), .Z(n669) );
  AND U4087 ( .A(n670), .B(n671), .Z(n668) );
  XOR U4088 ( .A(n672), .B(n673), .Z(n671) );
  XOR U4089 ( .A(DB[2414]), .B(DB[2407]), .Z(n673) );
  AND U4090 ( .A(n674), .B(n675), .Z(n672) );
  XOR U4091 ( .A(n676), .B(n677), .Z(n675) );
  XOR U4092 ( .A(DB[2407]), .B(DB[2400]), .Z(n677) );
  AND U4093 ( .A(n678), .B(n679), .Z(n676) );
  XOR U4094 ( .A(n680), .B(n681), .Z(n679) );
  XOR U4095 ( .A(DB[2400]), .B(DB[2393]), .Z(n681) );
  AND U4096 ( .A(n682), .B(n683), .Z(n680) );
  XOR U4097 ( .A(n684), .B(n685), .Z(n683) );
  XOR U4098 ( .A(DB[2393]), .B(DB[2386]), .Z(n685) );
  AND U4099 ( .A(n686), .B(n687), .Z(n684) );
  XOR U4100 ( .A(n688), .B(n689), .Z(n687) );
  XOR U4101 ( .A(DB[2386]), .B(DB[2379]), .Z(n689) );
  AND U4102 ( .A(n690), .B(n691), .Z(n688) );
  XOR U4103 ( .A(n692), .B(n693), .Z(n691) );
  XOR U4104 ( .A(DB[2379]), .B(DB[2372]), .Z(n693) );
  AND U4105 ( .A(n694), .B(n695), .Z(n692) );
  XOR U4106 ( .A(n696), .B(n697), .Z(n695) );
  XOR U4107 ( .A(DB[2372]), .B(DB[2365]), .Z(n697) );
  AND U4108 ( .A(n698), .B(n699), .Z(n696) );
  XOR U4109 ( .A(n700), .B(n701), .Z(n699) );
  XOR U4110 ( .A(DB[2365]), .B(DB[2358]), .Z(n701) );
  AND U4111 ( .A(n702), .B(n703), .Z(n700) );
  XOR U4112 ( .A(n704), .B(n705), .Z(n703) );
  XOR U4113 ( .A(DB[2358]), .B(DB[2351]), .Z(n705) );
  AND U4114 ( .A(n706), .B(n707), .Z(n704) );
  XOR U4115 ( .A(n708), .B(n709), .Z(n707) );
  XOR U4116 ( .A(DB[2351]), .B(DB[2344]), .Z(n709) );
  AND U4117 ( .A(n710), .B(n711), .Z(n708) );
  XOR U4118 ( .A(n712), .B(n713), .Z(n711) );
  XOR U4119 ( .A(DB[2344]), .B(DB[2337]), .Z(n713) );
  AND U4120 ( .A(n714), .B(n715), .Z(n712) );
  XOR U4121 ( .A(n716), .B(n717), .Z(n715) );
  XOR U4122 ( .A(DB[2337]), .B(DB[2330]), .Z(n717) );
  AND U4123 ( .A(n718), .B(n719), .Z(n716) );
  XOR U4124 ( .A(n720), .B(n721), .Z(n719) );
  XOR U4125 ( .A(DB[2330]), .B(DB[2323]), .Z(n721) );
  AND U4126 ( .A(n722), .B(n723), .Z(n720) );
  XOR U4127 ( .A(n724), .B(n725), .Z(n723) );
  XOR U4128 ( .A(DB[2323]), .B(DB[2316]), .Z(n725) );
  AND U4129 ( .A(n726), .B(n727), .Z(n724) );
  XOR U4130 ( .A(n728), .B(n729), .Z(n727) );
  XOR U4131 ( .A(DB[2316]), .B(DB[2309]), .Z(n729) );
  AND U4132 ( .A(n730), .B(n731), .Z(n728) );
  XOR U4133 ( .A(n732), .B(n733), .Z(n731) );
  XOR U4134 ( .A(DB[2309]), .B(DB[2302]), .Z(n733) );
  AND U4135 ( .A(n734), .B(n735), .Z(n732) );
  XOR U4136 ( .A(n736), .B(n737), .Z(n735) );
  XOR U4137 ( .A(DB[2302]), .B(DB[2295]), .Z(n737) );
  AND U4138 ( .A(n738), .B(n739), .Z(n736) );
  XOR U4139 ( .A(n740), .B(n741), .Z(n739) );
  XOR U4140 ( .A(DB[2295]), .B(DB[2288]), .Z(n741) );
  AND U4141 ( .A(n742), .B(n743), .Z(n740) );
  XOR U4142 ( .A(n744), .B(n745), .Z(n743) );
  XOR U4143 ( .A(DB[2288]), .B(DB[2281]), .Z(n745) );
  AND U4144 ( .A(n746), .B(n747), .Z(n744) );
  XOR U4145 ( .A(n748), .B(n749), .Z(n747) );
  XOR U4146 ( .A(DB[2281]), .B(DB[2274]), .Z(n749) );
  AND U4147 ( .A(n750), .B(n751), .Z(n748) );
  XOR U4148 ( .A(n752), .B(n753), .Z(n751) );
  XOR U4149 ( .A(DB[2274]), .B(DB[2267]), .Z(n753) );
  AND U4150 ( .A(n754), .B(n755), .Z(n752) );
  XOR U4151 ( .A(n756), .B(n757), .Z(n755) );
  XOR U4152 ( .A(DB[2267]), .B(DB[2260]), .Z(n757) );
  AND U4153 ( .A(n758), .B(n759), .Z(n756) );
  XOR U4154 ( .A(n760), .B(n761), .Z(n759) );
  XOR U4155 ( .A(DB[2260]), .B(DB[2253]), .Z(n761) );
  AND U4156 ( .A(n762), .B(n763), .Z(n760) );
  XOR U4157 ( .A(n764), .B(n765), .Z(n763) );
  XOR U4158 ( .A(DB[2253]), .B(DB[2246]), .Z(n765) );
  AND U4159 ( .A(n766), .B(n767), .Z(n764) );
  XOR U4160 ( .A(n768), .B(n769), .Z(n767) );
  XOR U4161 ( .A(DB[2246]), .B(DB[2239]), .Z(n769) );
  AND U4162 ( .A(n770), .B(n771), .Z(n768) );
  XOR U4163 ( .A(n772), .B(n773), .Z(n771) );
  XOR U4164 ( .A(DB[2239]), .B(DB[2232]), .Z(n773) );
  AND U4165 ( .A(n774), .B(n775), .Z(n772) );
  XOR U4166 ( .A(n776), .B(n777), .Z(n775) );
  XOR U4167 ( .A(DB[2232]), .B(DB[2225]), .Z(n777) );
  AND U4168 ( .A(n778), .B(n779), .Z(n776) );
  XOR U4169 ( .A(n780), .B(n781), .Z(n779) );
  XOR U4170 ( .A(DB[2225]), .B(DB[2218]), .Z(n781) );
  AND U4171 ( .A(n782), .B(n783), .Z(n780) );
  XOR U4172 ( .A(n784), .B(n785), .Z(n783) );
  XOR U4173 ( .A(DB[2218]), .B(DB[2211]), .Z(n785) );
  AND U4174 ( .A(n786), .B(n787), .Z(n784) );
  XOR U4175 ( .A(n788), .B(n789), .Z(n787) );
  XOR U4176 ( .A(DB[2211]), .B(DB[2204]), .Z(n789) );
  AND U4177 ( .A(n790), .B(n791), .Z(n788) );
  XOR U4178 ( .A(n792), .B(n793), .Z(n791) );
  XOR U4179 ( .A(DB[2204]), .B(DB[2197]), .Z(n793) );
  AND U4180 ( .A(n794), .B(n795), .Z(n792) );
  XOR U4181 ( .A(n796), .B(n797), .Z(n795) );
  XOR U4182 ( .A(DB[2197]), .B(DB[2190]), .Z(n797) );
  AND U4183 ( .A(n798), .B(n799), .Z(n796) );
  XOR U4184 ( .A(n800), .B(n801), .Z(n799) );
  XOR U4185 ( .A(DB[2190]), .B(DB[2183]), .Z(n801) );
  AND U4186 ( .A(n802), .B(n803), .Z(n800) );
  XOR U4187 ( .A(n804), .B(n805), .Z(n803) );
  XOR U4188 ( .A(DB[2183]), .B(DB[2176]), .Z(n805) );
  AND U4189 ( .A(n806), .B(n807), .Z(n804) );
  XOR U4190 ( .A(n808), .B(n809), .Z(n807) );
  XOR U4191 ( .A(DB[2176]), .B(DB[2169]), .Z(n809) );
  AND U4192 ( .A(n810), .B(n811), .Z(n808) );
  XOR U4193 ( .A(n812), .B(n813), .Z(n811) );
  XOR U4194 ( .A(DB[2169]), .B(DB[2162]), .Z(n813) );
  AND U4195 ( .A(n814), .B(n815), .Z(n812) );
  XOR U4196 ( .A(n816), .B(n817), .Z(n815) );
  XOR U4197 ( .A(DB[2162]), .B(DB[2155]), .Z(n817) );
  AND U4198 ( .A(n818), .B(n819), .Z(n816) );
  XOR U4199 ( .A(n820), .B(n821), .Z(n819) );
  XOR U4200 ( .A(DB[2155]), .B(DB[2148]), .Z(n821) );
  AND U4201 ( .A(n822), .B(n823), .Z(n820) );
  XOR U4202 ( .A(n824), .B(n825), .Z(n823) );
  XOR U4203 ( .A(DB[2148]), .B(DB[2141]), .Z(n825) );
  AND U4204 ( .A(n826), .B(n827), .Z(n824) );
  XOR U4205 ( .A(n828), .B(n829), .Z(n827) );
  XOR U4206 ( .A(DB[2141]), .B(DB[2134]), .Z(n829) );
  AND U4207 ( .A(n830), .B(n831), .Z(n828) );
  XOR U4208 ( .A(n832), .B(n833), .Z(n831) );
  XOR U4209 ( .A(DB[2134]), .B(DB[2127]), .Z(n833) );
  AND U4210 ( .A(n834), .B(n835), .Z(n832) );
  XOR U4211 ( .A(n836), .B(n837), .Z(n835) );
  XOR U4212 ( .A(DB[2127]), .B(DB[2120]), .Z(n837) );
  AND U4213 ( .A(n838), .B(n839), .Z(n836) );
  XOR U4214 ( .A(n840), .B(n841), .Z(n839) );
  XOR U4215 ( .A(DB[2120]), .B(DB[2113]), .Z(n841) );
  AND U4216 ( .A(n842), .B(n843), .Z(n840) );
  XOR U4217 ( .A(n844), .B(n845), .Z(n843) );
  XOR U4218 ( .A(DB[2113]), .B(DB[2106]), .Z(n845) );
  AND U4219 ( .A(n846), .B(n847), .Z(n844) );
  XOR U4220 ( .A(n848), .B(n849), .Z(n847) );
  XOR U4221 ( .A(DB[2106]), .B(DB[2099]), .Z(n849) );
  AND U4222 ( .A(n850), .B(n851), .Z(n848) );
  XOR U4223 ( .A(n852), .B(n853), .Z(n851) );
  XOR U4224 ( .A(DB[2099]), .B(DB[2092]), .Z(n853) );
  AND U4225 ( .A(n854), .B(n855), .Z(n852) );
  XOR U4226 ( .A(n856), .B(n857), .Z(n855) );
  XOR U4227 ( .A(DB[2092]), .B(DB[2085]), .Z(n857) );
  AND U4228 ( .A(n858), .B(n859), .Z(n856) );
  XOR U4229 ( .A(n860), .B(n861), .Z(n859) );
  XOR U4230 ( .A(DB[2085]), .B(DB[2078]), .Z(n861) );
  AND U4231 ( .A(n862), .B(n863), .Z(n860) );
  XOR U4232 ( .A(n864), .B(n865), .Z(n863) );
  XOR U4233 ( .A(DB[2078]), .B(DB[2071]), .Z(n865) );
  AND U4234 ( .A(n866), .B(n867), .Z(n864) );
  XOR U4235 ( .A(n868), .B(n869), .Z(n867) );
  XOR U4236 ( .A(DB[2071]), .B(DB[2064]), .Z(n869) );
  AND U4237 ( .A(n870), .B(n871), .Z(n868) );
  XOR U4238 ( .A(n872), .B(n873), .Z(n871) );
  XOR U4239 ( .A(DB[2064]), .B(DB[2057]), .Z(n873) );
  AND U4240 ( .A(n874), .B(n875), .Z(n872) );
  XOR U4241 ( .A(n876), .B(n877), .Z(n875) );
  XOR U4242 ( .A(DB[2057]), .B(DB[2050]), .Z(n877) );
  AND U4243 ( .A(n878), .B(n879), .Z(n876) );
  XOR U4244 ( .A(n880), .B(n881), .Z(n879) );
  XOR U4245 ( .A(DB[2050]), .B(DB[2043]), .Z(n881) );
  AND U4246 ( .A(n882), .B(n883), .Z(n880) );
  XOR U4247 ( .A(n884), .B(n885), .Z(n883) );
  XOR U4248 ( .A(DB[2043]), .B(DB[2036]), .Z(n885) );
  AND U4249 ( .A(n886), .B(n887), .Z(n884) );
  XOR U4250 ( .A(n888), .B(n889), .Z(n887) );
  XOR U4251 ( .A(DB[2036]), .B(DB[2029]), .Z(n889) );
  AND U4252 ( .A(n890), .B(n891), .Z(n888) );
  XOR U4253 ( .A(n892), .B(n893), .Z(n891) );
  XOR U4254 ( .A(DB[2029]), .B(DB[2022]), .Z(n893) );
  AND U4255 ( .A(n894), .B(n895), .Z(n892) );
  XOR U4256 ( .A(n896), .B(n897), .Z(n895) );
  XOR U4257 ( .A(DB[2022]), .B(DB[2015]), .Z(n897) );
  AND U4258 ( .A(n898), .B(n899), .Z(n896) );
  XOR U4259 ( .A(n900), .B(n901), .Z(n899) );
  XOR U4260 ( .A(DB[2015]), .B(DB[2008]), .Z(n901) );
  AND U4261 ( .A(n902), .B(n903), .Z(n900) );
  XOR U4262 ( .A(n904), .B(n905), .Z(n903) );
  XOR U4263 ( .A(DB[2008]), .B(DB[2001]), .Z(n905) );
  AND U4264 ( .A(n906), .B(n907), .Z(n904) );
  XOR U4265 ( .A(n908), .B(n909), .Z(n907) );
  XOR U4266 ( .A(DB[2001]), .B(DB[1994]), .Z(n909) );
  AND U4267 ( .A(n910), .B(n911), .Z(n908) );
  XOR U4268 ( .A(n912), .B(n913), .Z(n911) );
  XOR U4269 ( .A(DB[1994]), .B(DB[1987]), .Z(n913) );
  AND U4270 ( .A(n914), .B(n915), .Z(n912) );
  XOR U4271 ( .A(n916), .B(n917), .Z(n915) );
  XOR U4272 ( .A(DB[1987]), .B(DB[1980]), .Z(n917) );
  AND U4273 ( .A(n918), .B(n919), .Z(n916) );
  XOR U4274 ( .A(n920), .B(n921), .Z(n919) );
  XOR U4275 ( .A(DB[1980]), .B(DB[1973]), .Z(n921) );
  AND U4276 ( .A(n922), .B(n923), .Z(n920) );
  XOR U4277 ( .A(n924), .B(n925), .Z(n923) );
  XOR U4278 ( .A(DB[1973]), .B(DB[1966]), .Z(n925) );
  AND U4279 ( .A(n926), .B(n927), .Z(n924) );
  XOR U4280 ( .A(n928), .B(n929), .Z(n927) );
  XOR U4281 ( .A(DB[1966]), .B(DB[1959]), .Z(n929) );
  AND U4282 ( .A(n930), .B(n931), .Z(n928) );
  XOR U4283 ( .A(n932), .B(n933), .Z(n931) );
  XOR U4284 ( .A(DB[1959]), .B(DB[1952]), .Z(n933) );
  AND U4285 ( .A(n934), .B(n935), .Z(n932) );
  XOR U4286 ( .A(n936), .B(n937), .Z(n935) );
  XOR U4287 ( .A(DB[1952]), .B(DB[1945]), .Z(n937) );
  AND U4288 ( .A(n938), .B(n939), .Z(n936) );
  XOR U4289 ( .A(n940), .B(n941), .Z(n939) );
  XOR U4290 ( .A(DB[1945]), .B(DB[1938]), .Z(n941) );
  AND U4291 ( .A(n942), .B(n943), .Z(n940) );
  XOR U4292 ( .A(n944), .B(n945), .Z(n943) );
  XOR U4293 ( .A(DB[1938]), .B(DB[1931]), .Z(n945) );
  AND U4294 ( .A(n946), .B(n947), .Z(n944) );
  XOR U4295 ( .A(n948), .B(n949), .Z(n947) );
  XOR U4296 ( .A(DB[1931]), .B(DB[1924]), .Z(n949) );
  AND U4297 ( .A(n950), .B(n951), .Z(n948) );
  XOR U4298 ( .A(n952), .B(n953), .Z(n951) );
  XOR U4299 ( .A(DB[1924]), .B(DB[1917]), .Z(n953) );
  AND U4300 ( .A(n954), .B(n955), .Z(n952) );
  XOR U4301 ( .A(n956), .B(n957), .Z(n955) );
  XOR U4302 ( .A(DB[1917]), .B(DB[1910]), .Z(n957) );
  AND U4303 ( .A(n958), .B(n959), .Z(n956) );
  XOR U4304 ( .A(n960), .B(n961), .Z(n959) );
  XOR U4305 ( .A(DB[1910]), .B(DB[1903]), .Z(n961) );
  AND U4306 ( .A(n962), .B(n963), .Z(n960) );
  XOR U4307 ( .A(n964), .B(n965), .Z(n963) );
  XOR U4308 ( .A(DB[1903]), .B(DB[1896]), .Z(n965) );
  AND U4309 ( .A(n966), .B(n967), .Z(n964) );
  XOR U4310 ( .A(n968), .B(n969), .Z(n967) );
  XOR U4311 ( .A(DB[1896]), .B(DB[1889]), .Z(n969) );
  AND U4312 ( .A(n970), .B(n971), .Z(n968) );
  XOR U4313 ( .A(n972), .B(n973), .Z(n971) );
  XOR U4314 ( .A(DB[1889]), .B(DB[1882]), .Z(n973) );
  AND U4315 ( .A(n974), .B(n975), .Z(n972) );
  XOR U4316 ( .A(n976), .B(n977), .Z(n975) );
  XOR U4317 ( .A(DB[1882]), .B(DB[1875]), .Z(n977) );
  AND U4318 ( .A(n978), .B(n979), .Z(n976) );
  XOR U4319 ( .A(n980), .B(n981), .Z(n979) );
  XOR U4320 ( .A(DB[1875]), .B(DB[1868]), .Z(n981) );
  AND U4321 ( .A(n982), .B(n983), .Z(n980) );
  XOR U4322 ( .A(n984), .B(n985), .Z(n983) );
  XOR U4323 ( .A(DB[1868]), .B(DB[1861]), .Z(n985) );
  AND U4324 ( .A(n986), .B(n987), .Z(n984) );
  XOR U4325 ( .A(n988), .B(n989), .Z(n987) );
  XOR U4326 ( .A(DB[1861]), .B(DB[1854]), .Z(n989) );
  AND U4327 ( .A(n990), .B(n991), .Z(n988) );
  XOR U4328 ( .A(n992), .B(n993), .Z(n991) );
  XOR U4329 ( .A(DB[1854]), .B(DB[1847]), .Z(n993) );
  AND U4330 ( .A(n994), .B(n995), .Z(n992) );
  XOR U4331 ( .A(n996), .B(n997), .Z(n995) );
  XOR U4332 ( .A(DB[1847]), .B(DB[1840]), .Z(n997) );
  AND U4333 ( .A(n998), .B(n999), .Z(n996) );
  XOR U4334 ( .A(n1000), .B(n1001), .Z(n999) );
  XOR U4335 ( .A(DB[1840]), .B(DB[1833]), .Z(n1001) );
  AND U4336 ( .A(n1002), .B(n1003), .Z(n1000) );
  XOR U4337 ( .A(n1004), .B(n1005), .Z(n1003) );
  XOR U4338 ( .A(DB[1833]), .B(DB[1826]), .Z(n1005) );
  AND U4339 ( .A(n1006), .B(n1007), .Z(n1004) );
  XOR U4340 ( .A(n1008), .B(n1009), .Z(n1007) );
  XOR U4341 ( .A(DB[1826]), .B(DB[1819]), .Z(n1009) );
  AND U4342 ( .A(n1010), .B(n1011), .Z(n1008) );
  XOR U4343 ( .A(n1012), .B(n1013), .Z(n1011) );
  XOR U4344 ( .A(DB[1819]), .B(DB[1812]), .Z(n1013) );
  AND U4345 ( .A(n1014), .B(n1015), .Z(n1012) );
  XOR U4346 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR U4347 ( .A(DB[1812]), .B(DB[1805]), .Z(n1017) );
  AND U4348 ( .A(n1018), .B(n1019), .Z(n1016) );
  XOR U4349 ( .A(n1020), .B(n1021), .Z(n1019) );
  XOR U4350 ( .A(DB[1805]), .B(DB[1798]), .Z(n1021) );
  AND U4351 ( .A(n1022), .B(n1023), .Z(n1020) );
  XOR U4352 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U4353 ( .A(DB[1798]), .B(DB[1791]), .Z(n1025) );
  AND U4354 ( .A(n1026), .B(n1027), .Z(n1024) );
  XOR U4355 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U4356 ( .A(DB[1791]), .B(DB[1784]), .Z(n1029) );
  AND U4357 ( .A(n1030), .B(n1031), .Z(n1028) );
  XOR U4358 ( .A(n1032), .B(n1033), .Z(n1031) );
  XOR U4359 ( .A(DB[1784]), .B(DB[1777]), .Z(n1033) );
  AND U4360 ( .A(n1034), .B(n1035), .Z(n1032) );
  XOR U4361 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR U4362 ( .A(DB[1777]), .B(DB[1770]), .Z(n1037) );
  AND U4363 ( .A(n1038), .B(n1039), .Z(n1036) );
  XOR U4364 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U4365 ( .A(DB[1770]), .B(DB[1763]), .Z(n1041) );
  AND U4366 ( .A(n1042), .B(n1043), .Z(n1040) );
  XOR U4367 ( .A(n1044), .B(n1045), .Z(n1043) );
  XOR U4368 ( .A(DB[1763]), .B(DB[1756]), .Z(n1045) );
  AND U4369 ( .A(n1046), .B(n1047), .Z(n1044) );
  XOR U4370 ( .A(n1048), .B(n1049), .Z(n1047) );
  XOR U4371 ( .A(DB[1756]), .B(DB[1749]), .Z(n1049) );
  AND U4372 ( .A(n1050), .B(n1051), .Z(n1048) );
  XOR U4373 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR U4374 ( .A(DB[1749]), .B(DB[1742]), .Z(n1053) );
  AND U4375 ( .A(n1054), .B(n1055), .Z(n1052) );
  XOR U4376 ( .A(n1056), .B(n1057), .Z(n1055) );
  XOR U4377 ( .A(DB[1742]), .B(DB[1735]), .Z(n1057) );
  AND U4378 ( .A(n1058), .B(n1059), .Z(n1056) );
  XOR U4379 ( .A(n1060), .B(n1061), .Z(n1059) );
  XOR U4380 ( .A(DB[1735]), .B(DB[1728]), .Z(n1061) );
  AND U4381 ( .A(n1062), .B(n1063), .Z(n1060) );
  XOR U4382 ( .A(n1064), .B(n1065), .Z(n1063) );
  XOR U4383 ( .A(DB[1728]), .B(DB[1721]), .Z(n1065) );
  AND U4384 ( .A(n1066), .B(n1067), .Z(n1064) );
  XOR U4385 ( .A(n1068), .B(n1069), .Z(n1067) );
  XOR U4386 ( .A(DB[1721]), .B(DB[1714]), .Z(n1069) );
  AND U4387 ( .A(n1070), .B(n1071), .Z(n1068) );
  XOR U4388 ( .A(n1072), .B(n1073), .Z(n1071) );
  XOR U4389 ( .A(DB[1714]), .B(DB[1707]), .Z(n1073) );
  AND U4390 ( .A(n1074), .B(n1075), .Z(n1072) );
  XOR U4391 ( .A(n1076), .B(n1077), .Z(n1075) );
  XOR U4392 ( .A(DB[1707]), .B(DB[1700]), .Z(n1077) );
  AND U4393 ( .A(n1078), .B(n1079), .Z(n1076) );
  XOR U4394 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR U4395 ( .A(DB[1700]), .B(DB[1693]), .Z(n1081) );
  AND U4396 ( .A(n1082), .B(n1083), .Z(n1080) );
  XOR U4397 ( .A(n1084), .B(n1085), .Z(n1083) );
  XOR U4398 ( .A(DB[1693]), .B(DB[1686]), .Z(n1085) );
  AND U4399 ( .A(n1086), .B(n1087), .Z(n1084) );
  XOR U4400 ( .A(n1088), .B(n1089), .Z(n1087) );
  XOR U4401 ( .A(DB[1686]), .B(DB[1679]), .Z(n1089) );
  AND U4402 ( .A(n1090), .B(n1091), .Z(n1088) );
  XOR U4403 ( .A(n1092), .B(n1093), .Z(n1091) );
  XOR U4404 ( .A(DB[1679]), .B(DB[1672]), .Z(n1093) );
  AND U4405 ( .A(n1094), .B(n1095), .Z(n1092) );
  XOR U4406 ( .A(n1096), .B(n1097), .Z(n1095) );
  XOR U4407 ( .A(DB[1672]), .B(DB[1665]), .Z(n1097) );
  AND U4408 ( .A(n1098), .B(n1099), .Z(n1096) );
  XOR U4409 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U4410 ( .A(DB[1665]), .B(DB[1658]), .Z(n1101) );
  AND U4411 ( .A(n1102), .B(n1103), .Z(n1100) );
  XOR U4412 ( .A(n1104), .B(n1105), .Z(n1103) );
  XOR U4413 ( .A(DB[1658]), .B(DB[1651]), .Z(n1105) );
  AND U4414 ( .A(n1106), .B(n1107), .Z(n1104) );
  XOR U4415 ( .A(n1108), .B(n1109), .Z(n1107) );
  XOR U4416 ( .A(DB[1651]), .B(DB[1644]), .Z(n1109) );
  AND U4417 ( .A(n1110), .B(n1111), .Z(n1108) );
  XOR U4418 ( .A(n1112), .B(n1113), .Z(n1111) );
  XOR U4419 ( .A(DB[1644]), .B(DB[1637]), .Z(n1113) );
  AND U4420 ( .A(n1114), .B(n1115), .Z(n1112) );
  XOR U4421 ( .A(n1116), .B(n1117), .Z(n1115) );
  XOR U4422 ( .A(DB[1637]), .B(DB[1630]), .Z(n1117) );
  AND U4423 ( .A(n1118), .B(n1119), .Z(n1116) );
  XOR U4424 ( .A(n1120), .B(n1121), .Z(n1119) );
  XOR U4425 ( .A(DB[1630]), .B(DB[1623]), .Z(n1121) );
  AND U4426 ( .A(n1122), .B(n1123), .Z(n1120) );
  XOR U4427 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U4428 ( .A(DB[1623]), .B(DB[1616]), .Z(n1125) );
  AND U4429 ( .A(n1126), .B(n1127), .Z(n1124) );
  XOR U4430 ( .A(n1128), .B(n1129), .Z(n1127) );
  XOR U4431 ( .A(DB[1616]), .B(DB[1609]), .Z(n1129) );
  AND U4432 ( .A(n1130), .B(n1131), .Z(n1128) );
  XOR U4433 ( .A(n1132), .B(n1133), .Z(n1131) );
  XOR U4434 ( .A(DB[1609]), .B(DB[1602]), .Z(n1133) );
  AND U4435 ( .A(n1134), .B(n1135), .Z(n1132) );
  XOR U4436 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U4437 ( .A(DB[1602]), .B(DB[1595]), .Z(n1137) );
  AND U4438 ( .A(n1138), .B(n1139), .Z(n1136) );
  XOR U4439 ( .A(n1140), .B(n1141), .Z(n1139) );
  XOR U4440 ( .A(DB[1595]), .B(DB[1588]), .Z(n1141) );
  AND U4441 ( .A(n1142), .B(n1143), .Z(n1140) );
  XOR U4442 ( .A(n1144), .B(n1145), .Z(n1143) );
  XOR U4443 ( .A(DB[1588]), .B(DB[1581]), .Z(n1145) );
  AND U4444 ( .A(n1146), .B(n1147), .Z(n1144) );
  XOR U4445 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U4446 ( .A(DB[1581]), .B(DB[1574]), .Z(n1149) );
  AND U4447 ( .A(n1150), .B(n1151), .Z(n1148) );
  XOR U4448 ( .A(n1152), .B(n1153), .Z(n1151) );
  XOR U4449 ( .A(DB[1574]), .B(DB[1567]), .Z(n1153) );
  AND U4450 ( .A(n1154), .B(n1155), .Z(n1152) );
  XOR U4451 ( .A(n1156), .B(n1157), .Z(n1155) );
  XOR U4452 ( .A(DB[1567]), .B(DB[1560]), .Z(n1157) );
  AND U4453 ( .A(n1158), .B(n1159), .Z(n1156) );
  XOR U4454 ( .A(n1160), .B(n1161), .Z(n1159) );
  XOR U4455 ( .A(DB[1560]), .B(DB[1553]), .Z(n1161) );
  AND U4456 ( .A(n1162), .B(n1163), .Z(n1160) );
  XOR U4457 ( .A(n1164), .B(n1165), .Z(n1163) );
  XOR U4458 ( .A(DB[1553]), .B(DB[1546]), .Z(n1165) );
  AND U4459 ( .A(n1166), .B(n1167), .Z(n1164) );
  XOR U4460 ( .A(n1168), .B(n1169), .Z(n1167) );
  XOR U4461 ( .A(DB[1546]), .B(DB[1539]), .Z(n1169) );
  AND U4462 ( .A(n1170), .B(n1171), .Z(n1168) );
  XOR U4463 ( .A(n1172), .B(n1173), .Z(n1171) );
  XOR U4464 ( .A(DB[1539]), .B(DB[1532]), .Z(n1173) );
  AND U4465 ( .A(n1174), .B(n1175), .Z(n1172) );
  XOR U4466 ( .A(n1176), .B(n1177), .Z(n1175) );
  XOR U4467 ( .A(DB[1532]), .B(DB[1525]), .Z(n1177) );
  AND U4468 ( .A(n1178), .B(n1179), .Z(n1176) );
  XOR U4469 ( .A(n1180), .B(n1181), .Z(n1179) );
  XOR U4470 ( .A(DB[1525]), .B(DB[1518]), .Z(n1181) );
  AND U4471 ( .A(n1182), .B(n1183), .Z(n1180) );
  XOR U4472 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U4473 ( .A(DB[1518]), .B(DB[1511]), .Z(n1185) );
  AND U4474 ( .A(n1186), .B(n1187), .Z(n1184) );
  XOR U4475 ( .A(n1188), .B(n1189), .Z(n1187) );
  XOR U4476 ( .A(DB[1511]), .B(DB[1504]), .Z(n1189) );
  AND U4477 ( .A(n1190), .B(n1191), .Z(n1188) );
  XOR U4478 ( .A(n1192), .B(n1193), .Z(n1191) );
  XOR U4479 ( .A(DB[1504]), .B(DB[1497]), .Z(n1193) );
  AND U4480 ( .A(n1194), .B(n1195), .Z(n1192) );
  XOR U4481 ( .A(n1196), .B(n1197), .Z(n1195) );
  XOR U4482 ( .A(DB[1497]), .B(DB[1490]), .Z(n1197) );
  AND U4483 ( .A(n1198), .B(n1199), .Z(n1196) );
  XOR U4484 ( .A(n1200), .B(n1201), .Z(n1199) );
  XOR U4485 ( .A(DB[1490]), .B(DB[1483]), .Z(n1201) );
  AND U4486 ( .A(n1202), .B(n1203), .Z(n1200) );
  XOR U4487 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U4488 ( .A(DB[1483]), .B(DB[1476]), .Z(n1205) );
  AND U4489 ( .A(n1206), .B(n1207), .Z(n1204) );
  XOR U4490 ( .A(n1208), .B(n1209), .Z(n1207) );
  XOR U4491 ( .A(DB[1476]), .B(DB[1469]), .Z(n1209) );
  AND U4492 ( .A(n1210), .B(n1211), .Z(n1208) );
  XOR U4493 ( .A(n1212), .B(n1213), .Z(n1211) );
  XOR U4494 ( .A(DB[1469]), .B(DB[1462]), .Z(n1213) );
  AND U4495 ( .A(n1214), .B(n1215), .Z(n1212) );
  XOR U4496 ( .A(n1216), .B(n1217), .Z(n1215) );
  XOR U4497 ( .A(DB[1462]), .B(DB[1455]), .Z(n1217) );
  AND U4498 ( .A(n1218), .B(n1219), .Z(n1216) );
  XOR U4499 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U4500 ( .A(DB[1455]), .B(DB[1448]), .Z(n1221) );
  AND U4501 ( .A(n1222), .B(n1223), .Z(n1220) );
  XOR U4502 ( .A(n1224), .B(n1225), .Z(n1223) );
  XOR U4503 ( .A(DB[1448]), .B(DB[1441]), .Z(n1225) );
  AND U4504 ( .A(n1226), .B(n1227), .Z(n1224) );
  XOR U4505 ( .A(n1228), .B(n1229), .Z(n1227) );
  XOR U4506 ( .A(DB[1441]), .B(DB[1434]), .Z(n1229) );
  AND U4507 ( .A(n1230), .B(n1231), .Z(n1228) );
  XOR U4508 ( .A(n1232), .B(n1233), .Z(n1231) );
  XOR U4509 ( .A(DB[1434]), .B(DB[1427]), .Z(n1233) );
  AND U4510 ( .A(n1234), .B(n1235), .Z(n1232) );
  XOR U4511 ( .A(n1236), .B(n1237), .Z(n1235) );
  XOR U4512 ( .A(DB[1427]), .B(DB[1420]), .Z(n1237) );
  AND U4513 ( .A(n1238), .B(n1239), .Z(n1236) );
  XOR U4514 ( .A(n1240), .B(n1241), .Z(n1239) );
  XOR U4515 ( .A(DB[1420]), .B(DB[1413]), .Z(n1241) );
  AND U4516 ( .A(n1242), .B(n1243), .Z(n1240) );
  XOR U4517 ( .A(n1244), .B(n1245), .Z(n1243) );
  XOR U4518 ( .A(DB[1413]), .B(DB[1406]), .Z(n1245) );
  AND U4519 ( .A(n1246), .B(n1247), .Z(n1244) );
  XOR U4520 ( .A(n1248), .B(n1249), .Z(n1247) );
  XOR U4521 ( .A(DB[1406]), .B(DB[1399]), .Z(n1249) );
  AND U4522 ( .A(n1250), .B(n1251), .Z(n1248) );
  XOR U4523 ( .A(n1252), .B(n1253), .Z(n1251) );
  XOR U4524 ( .A(DB[1399]), .B(DB[1392]), .Z(n1253) );
  AND U4525 ( .A(n1254), .B(n1255), .Z(n1252) );
  XOR U4526 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U4527 ( .A(DB[1392]), .B(DB[1385]), .Z(n1257) );
  AND U4528 ( .A(n1258), .B(n1259), .Z(n1256) );
  XOR U4529 ( .A(n1260), .B(n1261), .Z(n1259) );
  XOR U4530 ( .A(DB[1385]), .B(DB[1378]), .Z(n1261) );
  AND U4531 ( .A(n1262), .B(n1263), .Z(n1260) );
  XOR U4532 ( .A(n1264), .B(n1265), .Z(n1263) );
  XOR U4533 ( .A(DB[1378]), .B(DB[1371]), .Z(n1265) );
  AND U4534 ( .A(n1266), .B(n1267), .Z(n1264) );
  XOR U4535 ( .A(n1268), .B(n1269), .Z(n1267) );
  XOR U4536 ( .A(DB[1371]), .B(DB[1364]), .Z(n1269) );
  AND U4537 ( .A(n1270), .B(n1271), .Z(n1268) );
  XOR U4538 ( .A(n1272), .B(n1273), .Z(n1271) );
  XOR U4539 ( .A(DB[1364]), .B(DB[1357]), .Z(n1273) );
  AND U4540 ( .A(n1274), .B(n1275), .Z(n1272) );
  XOR U4541 ( .A(n1276), .B(n1277), .Z(n1275) );
  XOR U4542 ( .A(DB[1357]), .B(DB[1350]), .Z(n1277) );
  AND U4543 ( .A(n1278), .B(n1279), .Z(n1276) );
  XOR U4544 ( .A(n1280), .B(n1281), .Z(n1279) );
  XOR U4545 ( .A(DB[1350]), .B(DB[1343]), .Z(n1281) );
  AND U4546 ( .A(n1282), .B(n1283), .Z(n1280) );
  XOR U4547 ( .A(n1284), .B(n1285), .Z(n1283) );
  XOR U4548 ( .A(DB[1343]), .B(DB[1336]), .Z(n1285) );
  AND U4549 ( .A(n1286), .B(n1287), .Z(n1284) );
  XOR U4550 ( .A(n1288), .B(n1289), .Z(n1287) );
  XOR U4551 ( .A(DB[1336]), .B(DB[1329]), .Z(n1289) );
  AND U4552 ( .A(n1290), .B(n1291), .Z(n1288) );
  XOR U4553 ( .A(n1292), .B(n1293), .Z(n1291) );
  XOR U4554 ( .A(DB[1329]), .B(DB[1322]), .Z(n1293) );
  AND U4555 ( .A(n1294), .B(n1295), .Z(n1292) );
  XOR U4556 ( .A(n1296), .B(n1297), .Z(n1295) );
  XOR U4557 ( .A(DB[1322]), .B(DB[1315]), .Z(n1297) );
  AND U4558 ( .A(n1298), .B(n1299), .Z(n1296) );
  XOR U4559 ( .A(n1300), .B(n1301), .Z(n1299) );
  XOR U4560 ( .A(DB[1315]), .B(DB[1308]), .Z(n1301) );
  AND U4561 ( .A(n1302), .B(n1303), .Z(n1300) );
  XOR U4562 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U4563 ( .A(DB[1308]), .B(DB[1301]), .Z(n1305) );
  AND U4564 ( .A(n1306), .B(n1307), .Z(n1304) );
  XOR U4565 ( .A(n1308), .B(n1309), .Z(n1307) );
  XOR U4566 ( .A(DB[1301]), .B(DB[1294]), .Z(n1309) );
  AND U4567 ( .A(n1310), .B(n1311), .Z(n1308) );
  XOR U4568 ( .A(n1312), .B(n1313), .Z(n1311) );
  XOR U4569 ( .A(DB[1294]), .B(DB[1287]), .Z(n1313) );
  AND U4570 ( .A(n1314), .B(n1315), .Z(n1312) );
  XOR U4571 ( .A(n1316), .B(n1317), .Z(n1315) );
  XOR U4572 ( .A(DB[1287]), .B(DB[1280]), .Z(n1317) );
  AND U4573 ( .A(n1318), .B(n1319), .Z(n1316) );
  XOR U4574 ( .A(n1320), .B(n1321), .Z(n1319) );
  XOR U4575 ( .A(DB[1280]), .B(DB[1273]), .Z(n1321) );
  AND U4576 ( .A(n1322), .B(n1323), .Z(n1320) );
  XOR U4577 ( .A(n1324), .B(n1325), .Z(n1323) );
  XOR U4578 ( .A(DB[1273]), .B(DB[1266]), .Z(n1325) );
  AND U4579 ( .A(n1326), .B(n1327), .Z(n1324) );
  XOR U4580 ( .A(n1328), .B(n1329), .Z(n1327) );
  XOR U4581 ( .A(DB[1266]), .B(DB[1259]), .Z(n1329) );
  AND U4582 ( .A(n1330), .B(n1331), .Z(n1328) );
  XOR U4583 ( .A(n1332), .B(n1333), .Z(n1331) );
  XOR U4584 ( .A(DB[1259]), .B(DB[1252]), .Z(n1333) );
  AND U4585 ( .A(n1334), .B(n1335), .Z(n1332) );
  XOR U4586 ( .A(n1336), .B(n1337), .Z(n1335) );
  XOR U4587 ( .A(DB[1252]), .B(DB[1245]), .Z(n1337) );
  AND U4588 ( .A(n1338), .B(n1339), .Z(n1336) );
  XOR U4589 ( .A(n1340), .B(n1341), .Z(n1339) );
  XOR U4590 ( .A(DB[1245]), .B(DB[1238]), .Z(n1341) );
  AND U4591 ( .A(n1342), .B(n1343), .Z(n1340) );
  XOR U4592 ( .A(n1344), .B(n1345), .Z(n1343) );
  XOR U4593 ( .A(DB[1238]), .B(DB[1231]), .Z(n1345) );
  AND U4594 ( .A(n1346), .B(n1347), .Z(n1344) );
  XOR U4595 ( .A(n1348), .B(n1349), .Z(n1347) );
  XOR U4596 ( .A(DB[1231]), .B(DB[1224]), .Z(n1349) );
  AND U4597 ( .A(n1350), .B(n1351), .Z(n1348) );
  XOR U4598 ( .A(n1352), .B(n1353), .Z(n1351) );
  XOR U4599 ( .A(DB[1224]), .B(DB[1217]), .Z(n1353) );
  AND U4600 ( .A(n1354), .B(n1355), .Z(n1352) );
  XOR U4601 ( .A(n1356), .B(n1357), .Z(n1355) );
  XOR U4602 ( .A(DB[1217]), .B(DB[1210]), .Z(n1357) );
  AND U4603 ( .A(n1358), .B(n1359), .Z(n1356) );
  XOR U4604 ( .A(n1360), .B(n1361), .Z(n1359) );
  XOR U4605 ( .A(DB[1210]), .B(DB[1203]), .Z(n1361) );
  AND U4606 ( .A(n1362), .B(n1363), .Z(n1360) );
  XOR U4607 ( .A(n1364), .B(n1365), .Z(n1363) );
  XOR U4608 ( .A(DB[1203]), .B(DB[1196]), .Z(n1365) );
  AND U4609 ( .A(n1366), .B(n1367), .Z(n1364) );
  XOR U4610 ( .A(n1368), .B(n1369), .Z(n1367) );
  XOR U4611 ( .A(DB[1196]), .B(DB[1189]), .Z(n1369) );
  AND U4612 ( .A(n1370), .B(n1371), .Z(n1368) );
  XOR U4613 ( .A(n1372), .B(n1373), .Z(n1371) );
  XOR U4614 ( .A(DB[1189]), .B(DB[1182]), .Z(n1373) );
  AND U4615 ( .A(n1374), .B(n1375), .Z(n1372) );
  XOR U4616 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR U4617 ( .A(DB[1182]), .B(DB[1175]), .Z(n1377) );
  AND U4618 ( .A(n1378), .B(n1379), .Z(n1376) );
  XOR U4619 ( .A(n1380), .B(n1381), .Z(n1379) );
  XOR U4620 ( .A(DB[1175]), .B(DB[1168]), .Z(n1381) );
  AND U4621 ( .A(n1382), .B(n1383), .Z(n1380) );
  XOR U4622 ( .A(n1384), .B(n1385), .Z(n1383) );
  XOR U4623 ( .A(DB[1168]), .B(DB[1161]), .Z(n1385) );
  AND U4624 ( .A(n1386), .B(n1387), .Z(n1384) );
  XOR U4625 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR U4626 ( .A(DB[1161]), .B(DB[1154]), .Z(n1389) );
  AND U4627 ( .A(n1390), .B(n1391), .Z(n1388) );
  XOR U4628 ( .A(n1392), .B(n1393), .Z(n1391) );
  XOR U4629 ( .A(DB[1154]), .B(DB[1147]), .Z(n1393) );
  AND U4630 ( .A(n1394), .B(n1395), .Z(n1392) );
  XOR U4631 ( .A(n1396), .B(n1397), .Z(n1395) );
  XOR U4632 ( .A(DB[1147]), .B(DB[1140]), .Z(n1397) );
  AND U4633 ( .A(n1398), .B(n1399), .Z(n1396) );
  XOR U4634 ( .A(n1400), .B(n1401), .Z(n1399) );
  XOR U4635 ( .A(DB[1140]), .B(DB[1133]), .Z(n1401) );
  AND U4636 ( .A(n1402), .B(n1403), .Z(n1400) );
  XOR U4637 ( .A(n1404), .B(n1405), .Z(n1403) );
  XOR U4638 ( .A(DB[1133]), .B(DB[1126]), .Z(n1405) );
  AND U4639 ( .A(n1406), .B(n1407), .Z(n1404) );
  XOR U4640 ( .A(n1408), .B(n1409), .Z(n1407) );
  XOR U4641 ( .A(DB[1126]), .B(DB[1119]), .Z(n1409) );
  AND U4642 ( .A(n1410), .B(n1411), .Z(n1408) );
  XOR U4643 ( .A(n1412), .B(n1413), .Z(n1411) );
  XOR U4644 ( .A(DB[1119]), .B(DB[1112]), .Z(n1413) );
  AND U4645 ( .A(n1414), .B(n1415), .Z(n1412) );
  XOR U4646 ( .A(n1416), .B(n1417), .Z(n1415) );
  XOR U4647 ( .A(DB[1112]), .B(DB[1105]), .Z(n1417) );
  AND U4648 ( .A(n1418), .B(n1419), .Z(n1416) );
  XOR U4649 ( .A(n1420), .B(n1421), .Z(n1419) );
  XOR U4650 ( .A(DB[1105]), .B(DB[1098]), .Z(n1421) );
  AND U4651 ( .A(n1422), .B(n1423), .Z(n1420) );
  XOR U4652 ( .A(n1424), .B(n1425), .Z(n1423) );
  XOR U4653 ( .A(DB[1098]), .B(DB[1091]), .Z(n1425) );
  AND U4654 ( .A(n1426), .B(n1427), .Z(n1424) );
  XOR U4655 ( .A(n1428), .B(n1429), .Z(n1427) );
  XOR U4656 ( .A(DB[1091]), .B(DB[1084]), .Z(n1429) );
  AND U4657 ( .A(n1430), .B(n1431), .Z(n1428) );
  XOR U4658 ( .A(n1432), .B(n1433), .Z(n1431) );
  XOR U4659 ( .A(DB[1084]), .B(DB[1077]), .Z(n1433) );
  AND U4660 ( .A(n1434), .B(n1435), .Z(n1432) );
  XOR U4661 ( .A(n1436), .B(n1437), .Z(n1435) );
  XOR U4662 ( .A(DB[1077]), .B(DB[1070]), .Z(n1437) );
  AND U4663 ( .A(n1438), .B(n1439), .Z(n1436) );
  XOR U4664 ( .A(n1440), .B(n1441), .Z(n1439) );
  XOR U4665 ( .A(DB[1070]), .B(DB[1063]), .Z(n1441) );
  AND U4666 ( .A(n1442), .B(n1443), .Z(n1440) );
  XOR U4667 ( .A(n1444), .B(n1445), .Z(n1443) );
  XOR U4668 ( .A(DB[1063]), .B(DB[1056]), .Z(n1445) );
  AND U4669 ( .A(n1446), .B(n1447), .Z(n1444) );
  XOR U4670 ( .A(n1448), .B(n1449), .Z(n1447) );
  XOR U4671 ( .A(DB[1056]), .B(DB[1049]), .Z(n1449) );
  AND U4672 ( .A(n1450), .B(n1451), .Z(n1448) );
  XOR U4673 ( .A(n1452), .B(n1453), .Z(n1451) );
  XOR U4674 ( .A(DB[1049]), .B(DB[1042]), .Z(n1453) );
  AND U4675 ( .A(n1454), .B(n1455), .Z(n1452) );
  XOR U4676 ( .A(n1456), .B(n1457), .Z(n1455) );
  XOR U4677 ( .A(DB[1042]), .B(DB[1035]), .Z(n1457) );
  AND U4678 ( .A(n1458), .B(n1459), .Z(n1456) );
  XOR U4679 ( .A(n1460), .B(n1461), .Z(n1459) );
  XOR U4680 ( .A(DB[1035]), .B(DB[1028]), .Z(n1461) );
  AND U4681 ( .A(n1462), .B(n1463), .Z(n1460) );
  XOR U4682 ( .A(n1464), .B(n1465), .Z(n1463) );
  XOR U4683 ( .A(DB[1028]), .B(DB[1021]), .Z(n1465) );
  AND U4684 ( .A(n1466), .B(n1467), .Z(n1464) );
  XOR U4685 ( .A(n1468), .B(n1469), .Z(n1467) );
  XOR U4686 ( .A(DB[1021]), .B(DB[1014]), .Z(n1469) );
  AND U4687 ( .A(n1470), .B(n1471), .Z(n1468) );
  XOR U4688 ( .A(n1472), .B(n1473), .Z(n1471) );
  XOR U4689 ( .A(DB[1014]), .B(DB[1007]), .Z(n1473) );
  AND U4690 ( .A(n1474), .B(n1475), .Z(n1472) );
  XOR U4691 ( .A(n1476), .B(n1477), .Z(n1475) );
  XOR U4692 ( .A(DB[1007]), .B(DB[1000]), .Z(n1477) );
  AND U4693 ( .A(n1478), .B(n1479), .Z(n1476) );
  XOR U4694 ( .A(n1480), .B(n1481), .Z(n1479) );
  XOR U4695 ( .A(DB[993]), .B(DB[1000]), .Z(n1481) );
  AND U4696 ( .A(n1482), .B(n1483), .Z(n1480) );
  XOR U4697 ( .A(n1484), .B(n1485), .Z(n1483) );
  XOR U4698 ( .A(DB[993]), .B(DB[986]), .Z(n1485) );
  AND U4699 ( .A(n1486), .B(n1487), .Z(n1484) );
  XOR U4700 ( .A(n1488), .B(n1489), .Z(n1487) );
  XOR U4701 ( .A(DB[986]), .B(DB[979]), .Z(n1489) );
  AND U4702 ( .A(n1490), .B(n1491), .Z(n1488) );
  XOR U4703 ( .A(n1492), .B(n1493), .Z(n1491) );
  XOR U4704 ( .A(DB[979]), .B(DB[972]), .Z(n1493) );
  AND U4705 ( .A(n1494), .B(n1495), .Z(n1492) );
  XOR U4706 ( .A(n1496), .B(n1497), .Z(n1495) );
  XOR U4707 ( .A(DB[972]), .B(DB[965]), .Z(n1497) );
  AND U4708 ( .A(n1498), .B(n1499), .Z(n1496) );
  XOR U4709 ( .A(n1500), .B(n1501), .Z(n1499) );
  XOR U4710 ( .A(DB[965]), .B(DB[958]), .Z(n1501) );
  AND U4711 ( .A(n1502), .B(n1503), .Z(n1500) );
  XOR U4712 ( .A(n1504), .B(n1505), .Z(n1503) );
  XOR U4713 ( .A(DB[958]), .B(DB[951]), .Z(n1505) );
  AND U4714 ( .A(n1506), .B(n1507), .Z(n1504) );
  XOR U4715 ( .A(n1508), .B(n1509), .Z(n1507) );
  XOR U4716 ( .A(DB[951]), .B(DB[944]), .Z(n1509) );
  AND U4717 ( .A(n1510), .B(n1511), .Z(n1508) );
  XOR U4718 ( .A(n1512), .B(n1513), .Z(n1511) );
  XOR U4719 ( .A(DB[944]), .B(DB[937]), .Z(n1513) );
  AND U4720 ( .A(n1514), .B(n1515), .Z(n1512) );
  XOR U4721 ( .A(n1516), .B(n1517), .Z(n1515) );
  XOR U4722 ( .A(DB[937]), .B(DB[930]), .Z(n1517) );
  AND U4723 ( .A(n1518), .B(n1519), .Z(n1516) );
  XOR U4724 ( .A(n1520), .B(n1521), .Z(n1519) );
  XOR U4725 ( .A(DB[930]), .B(DB[923]), .Z(n1521) );
  AND U4726 ( .A(n1522), .B(n1523), .Z(n1520) );
  XOR U4727 ( .A(n1524), .B(n1525), .Z(n1523) );
  XOR U4728 ( .A(DB[923]), .B(DB[916]), .Z(n1525) );
  AND U4729 ( .A(n1526), .B(n1527), .Z(n1524) );
  XOR U4730 ( .A(n1528), .B(n1529), .Z(n1527) );
  XOR U4731 ( .A(DB[916]), .B(DB[909]), .Z(n1529) );
  AND U4732 ( .A(n1530), .B(n1531), .Z(n1528) );
  XOR U4733 ( .A(n1532), .B(n1533), .Z(n1531) );
  XOR U4734 ( .A(DB[909]), .B(DB[902]), .Z(n1533) );
  AND U4735 ( .A(n1534), .B(n1535), .Z(n1532) );
  XOR U4736 ( .A(n1536), .B(n1537), .Z(n1535) );
  XOR U4737 ( .A(DB[902]), .B(DB[895]), .Z(n1537) );
  AND U4738 ( .A(n1538), .B(n1539), .Z(n1536) );
  XOR U4739 ( .A(n1540), .B(n1541), .Z(n1539) );
  XOR U4740 ( .A(DB[895]), .B(DB[888]), .Z(n1541) );
  AND U4741 ( .A(n1542), .B(n1543), .Z(n1540) );
  XOR U4742 ( .A(n1544), .B(n1545), .Z(n1543) );
  XOR U4743 ( .A(DB[888]), .B(DB[881]), .Z(n1545) );
  AND U4744 ( .A(n1546), .B(n1547), .Z(n1544) );
  XOR U4745 ( .A(n1548), .B(n1549), .Z(n1547) );
  XOR U4746 ( .A(DB[881]), .B(DB[874]), .Z(n1549) );
  AND U4747 ( .A(n1550), .B(n1551), .Z(n1548) );
  XOR U4748 ( .A(n1552), .B(n1553), .Z(n1551) );
  XOR U4749 ( .A(DB[874]), .B(DB[867]), .Z(n1553) );
  AND U4750 ( .A(n1554), .B(n1555), .Z(n1552) );
  XOR U4751 ( .A(n1556), .B(n1557), .Z(n1555) );
  XOR U4752 ( .A(DB[867]), .B(DB[860]), .Z(n1557) );
  AND U4753 ( .A(n1558), .B(n1559), .Z(n1556) );
  XOR U4754 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U4755 ( .A(DB[860]), .B(DB[853]), .Z(n1561) );
  AND U4756 ( .A(n1562), .B(n1563), .Z(n1560) );
  XOR U4757 ( .A(n1564), .B(n1565), .Z(n1563) );
  XOR U4758 ( .A(DB[853]), .B(DB[846]), .Z(n1565) );
  AND U4759 ( .A(n1566), .B(n1567), .Z(n1564) );
  XOR U4760 ( .A(n1568), .B(n1569), .Z(n1567) );
  XOR U4761 ( .A(DB[846]), .B(DB[839]), .Z(n1569) );
  AND U4762 ( .A(n1570), .B(n1571), .Z(n1568) );
  XOR U4763 ( .A(n1572), .B(n1573), .Z(n1571) );
  XOR U4764 ( .A(DB[839]), .B(DB[832]), .Z(n1573) );
  AND U4765 ( .A(n1574), .B(n1575), .Z(n1572) );
  XOR U4766 ( .A(n1576), .B(n1577), .Z(n1575) );
  XOR U4767 ( .A(DB[832]), .B(DB[825]), .Z(n1577) );
  AND U4768 ( .A(n1578), .B(n1579), .Z(n1576) );
  XOR U4769 ( .A(n1580), .B(n1581), .Z(n1579) );
  XOR U4770 ( .A(DB[825]), .B(DB[818]), .Z(n1581) );
  AND U4771 ( .A(n1582), .B(n1583), .Z(n1580) );
  XOR U4772 ( .A(n1584), .B(n1585), .Z(n1583) );
  XOR U4773 ( .A(DB[818]), .B(DB[811]), .Z(n1585) );
  AND U4774 ( .A(n1586), .B(n1587), .Z(n1584) );
  XOR U4775 ( .A(n1588), .B(n1589), .Z(n1587) );
  XOR U4776 ( .A(DB[811]), .B(DB[804]), .Z(n1589) );
  AND U4777 ( .A(n1590), .B(n1591), .Z(n1588) );
  XOR U4778 ( .A(n1592), .B(n1593), .Z(n1591) );
  XOR U4779 ( .A(DB[804]), .B(DB[797]), .Z(n1593) );
  AND U4780 ( .A(n1594), .B(n1595), .Z(n1592) );
  XOR U4781 ( .A(n1596), .B(n1597), .Z(n1595) );
  XOR U4782 ( .A(DB[797]), .B(DB[790]), .Z(n1597) );
  AND U4783 ( .A(n1598), .B(n1599), .Z(n1596) );
  XOR U4784 ( .A(n1600), .B(n1601), .Z(n1599) );
  XOR U4785 ( .A(DB[790]), .B(DB[783]), .Z(n1601) );
  AND U4786 ( .A(n1602), .B(n1603), .Z(n1600) );
  XOR U4787 ( .A(n1604), .B(n1605), .Z(n1603) );
  XOR U4788 ( .A(DB[783]), .B(DB[776]), .Z(n1605) );
  AND U4789 ( .A(n1606), .B(n1607), .Z(n1604) );
  XOR U4790 ( .A(n1608), .B(n1609), .Z(n1607) );
  XOR U4791 ( .A(DB[776]), .B(DB[769]), .Z(n1609) );
  AND U4792 ( .A(n1610), .B(n1611), .Z(n1608) );
  XOR U4793 ( .A(n1612), .B(n1613), .Z(n1611) );
  XOR U4794 ( .A(DB[769]), .B(DB[762]), .Z(n1613) );
  AND U4795 ( .A(n1614), .B(n1615), .Z(n1612) );
  XOR U4796 ( .A(n1616), .B(n1617), .Z(n1615) );
  XOR U4797 ( .A(DB[762]), .B(DB[755]), .Z(n1617) );
  AND U4798 ( .A(n1618), .B(n1619), .Z(n1616) );
  XOR U4799 ( .A(n1620), .B(n1621), .Z(n1619) );
  XOR U4800 ( .A(DB[755]), .B(DB[748]), .Z(n1621) );
  AND U4801 ( .A(n1622), .B(n1623), .Z(n1620) );
  XOR U4802 ( .A(n1624), .B(n1625), .Z(n1623) );
  XOR U4803 ( .A(DB[748]), .B(DB[741]), .Z(n1625) );
  AND U4804 ( .A(n1626), .B(n1627), .Z(n1624) );
  XOR U4805 ( .A(n1628), .B(n1629), .Z(n1627) );
  XOR U4806 ( .A(DB[741]), .B(DB[734]), .Z(n1629) );
  AND U4807 ( .A(n1630), .B(n1631), .Z(n1628) );
  XOR U4808 ( .A(n1632), .B(n1633), .Z(n1631) );
  XOR U4809 ( .A(DB[734]), .B(DB[727]), .Z(n1633) );
  AND U4810 ( .A(n1634), .B(n1635), .Z(n1632) );
  XOR U4811 ( .A(n1636), .B(n1637), .Z(n1635) );
  XOR U4812 ( .A(DB[727]), .B(DB[720]), .Z(n1637) );
  AND U4813 ( .A(n1638), .B(n1639), .Z(n1636) );
  XOR U4814 ( .A(n1640), .B(n1641), .Z(n1639) );
  XOR U4815 ( .A(DB[720]), .B(DB[713]), .Z(n1641) );
  AND U4816 ( .A(n1642), .B(n1643), .Z(n1640) );
  XOR U4817 ( .A(n1644), .B(n1645), .Z(n1643) );
  XOR U4818 ( .A(DB[713]), .B(DB[706]), .Z(n1645) );
  AND U4819 ( .A(n1646), .B(n1647), .Z(n1644) );
  XOR U4820 ( .A(n1648), .B(n1649), .Z(n1647) );
  XOR U4821 ( .A(DB[706]), .B(DB[699]), .Z(n1649) );
  AND U4822 ( .A(n1650), .B(n1651), .Z(n1648) );
  XOR U4823 ( .A(n1652), .B(n1653), .Z(n1651) );
  XOR U4824 ( .A(DB[699]), .B(DB[692]), .Z(n1653) );
  AND U4825 ( .A(n1654), .B(n1655), .Z(n1652) );
  XOR U4826 ( .A(n1656), .B(n1657), .Z(n1655) );
  XOR U4827 ( .A(DB[692]), .B(DB[685]), .Z(n1657) );
  AND U4828 ( .A(n1658), .B(n1659), .Z(n1656) );
  XOR U4829 ( .A(n1660), .B(n1661), .Z(n1659) );
  XOR U4830 ( .A(DB[685]), .B(DB[678]), .Z(n1661) );
  AND U4831 ( .A(n1662), .B(n1663), .Z(n1660) );
  XOR U4832 ( .A(n1664), .B(n1665), .Z(n1663) );
  XOR U4833 ( .A(DB[678]), .B(DB[671]), .Z(n1665) );
  AND U4834 ( .A(n1666), .B(n1667), .Z(n1664) );
  XOR U4835 ( .A(n1668), .B(n1669), .Z(n1667) );
  XOR U4836 ( .A(DB[671]), .B(DB[664]), .Z(n1669) );
  AND U4837 ( .A(n1670), .B(n1671), .Z(n1668) );
  XOR U4838 ( .A(n1672), .B(n1673), .Z(n1671) );
  XOR U4839 ( .A(DB[664]), .B(DB[657]), .Z(n1673) );
  AND U4840 ( .A(n1674), .B(n1675), .Z(n1672) );
  XOR U4841 ( .A(n1676), .B(n1677), .Z(n1675) );
  XOR U4842 ( .A(DB[657]), .B(DB[650]), .Z(n1677) );
  AND U4843 ( .A(n1678), .B(n1679), .Z(n1676) );
  XOR U4844 ( .A(n1680), .B(n1681), .Z(n1679) );
  XOR U4845 ( .A(DB[650]), .B(DB[643]), .Z(n1681) );
  AND U4846 ( .A(n1682), .B(n1683), .Z(n1680) );
  XOR U4847 ( .A(n1684), .B(n1685), .Z(n1683) );
  XOR U4848 ( .A(DB[643]), .B(DB[636]), .Z(n1685) );
  AND U4849 ( .A(n1686), .B(n1687), .Z(n1684) );
  XOR U4850 ( .A(n1688), .B(n1689), .Z(n1687) );
  XOR U4851 ( .A(DB[636]), .B(DB[629]), .Z(n1689) );
  AND U4852 ( .A(n1690), .B(n1691), .Z(n1688) );
  XOR U4853 ( .A(n1692), .B(n1693), .Z(n1691) );
  XOR U4854 ( .A(DB[629]), .B(DB[622]), .Z(n1693) );
  AND U4855 ( .A(n1694), .B(n1695), .Z(n1692) );
  XOR U4856 ( .A(n1696), .B(n1697), .Z(n1695) );
  XOR U4857 ( .A(DB[622]), .B(DB[615]), .Z(n1697) );
  AND U4858 ( .A(n1698), .B(n1699), .Z(n1696) );
  XOR U4859 ( .A(n1700), .B(n1701), .Z(n1699) );
  XOR U4860 ( .A(DB[615]), .B(DB[608]), .Z(n1701) );
  AND U4861 ( .A(n1702), .B(n1703), .Z(n1700) );
  XOR U4862 ( .A(n1704), .B(n1705), .Z(n1703) );
  XOR U4863 ( .A(DB[608]), .B(DB[601]), .Z(n1705) );
  AND U4864 ( .A(n1706), .B(n1707), .Z(n1704) );
  XOR U4865 ( .A(n1708), .B(n1709), .Z(n1707) );
  XOR U4866 ( .A(DB[601]), .B(DB[594]), .Z(n1709) );
  AND U4867 ( .A(n1710), .B(n1711), .Z(n1708) );
  XOR U4868 ( .A(n1712), .B(n1713), .Z(n1711) );
  XOR U4869 ( .A(DB[594]), .B(DB[587]), .Z(n1713) );
  AND U4870 ( .A(n1714), .B(n1715), .Z(n1712) );
  XOR U4871 ( .A(n1716), .B(n1717), .Z(n1715) );
  XOR U4872 ( .A(DB[587]), .B(DB[580]), .Z(n1717) );
  AND U4873 ( .A(n1718), .B(n1719), .Z(n1716) );
  XOR U4874 ( .A(n1720), .B(n1721), .Z(n1719) );
  XOR U4875 ( .A(DB[580]), .B(DB[573]), .Z(n1721) );
  AND U4876 ( .A(n1722), .B(n1723), .Z(n1720) );
  XOR U4877 ( .A(n1724), .B(n1725), .Z(n1723) );
  XOR U4878 ( .A(DB[573]), .B(DB[566]), .Z(n1725) );
  AND U4879 ( .A(n1726), .B(n1727), .Z(n1724) );
  XOR U4880 ( .A(n1728), .B(n1729), .Z(n1727) );
  XOR U4881 ( .A(DB[566]), .B(DB[559]), .Z(n1729) );
  AND U4882 ( .A(n1730), .B(n1731), .Z(n1728) );
  XOR U4883 ( .A(n1732), .B(n1733), .Z(n1731) );
  XOR U4884 ( .A(DB[559]), .B(DB[552]), .Z(n1733) );
  AND U4885 ( .A(n1734), .B(n1735), .Z(n1732) );
  XOR U4886 ( .A(n1736), .B(n1737), .Z(n1735) );
  XOR U4887 ( .A(DB[552]), .B(DB[545]), .Z(n1737) );
  AND U4888 ( .A(n1738), .B(n1739), .Z(n1736) );
  XOR U4889 ( .A(n1740), .B(n1741), .Z(n1739) );
  XOR U4890 ( .A(DB[545]), .B(DB[538]), .Z(n1741) );
  AND U4891 ( .A(n1742), .B(n1743), .Z(n1740) );
  XOR U4892 ( .A(n1744), .B(n1745), .Z(n1743) );
  XOR U4893 ( .A(DB[538]), .B(DB[531]), .Z(n1745) );
  AND U4894 ( .A(n1746), .B(n1747), .Z(n1744) );
  XOR U4895 ( .A(n1748), .B(n1749), .Z(n1747) );
  XOR U4896 ( .A(DB[531]), .B(DB[524]), .Z(n1749) );
  AND U4897 ( .A(n1750), .B(n1751), .Z(n1748) );
  XOR U4898 ( .A(n1752), .B(n1753), .Z(n1751) );
  XOR U4899 ( .A(DB[524]), .B(DB[517]), .Z(n1753) );
  AND U4900 ( .A(n1754), .B(n1755), .Z(n1752) );
  XOR U4901 ( .A(n1756), .B(n1757), .Z(n1755) );
  XOR U4902 ( .A(DB[517]), .B(DB[510]), .Z(n1757) );
  AND U4903 ( .A(n1758), .B(n1759), .Z(n1756) );
  XOR U4904 ( .A(n1760), .B(n1761), .Z(n1759) );
  XOR U4905 ( .A(DB[510]), .B(DB[503]), .Z(n1761) );
  AND U4906 ( .A(n1762), .B(n1763), .Z(n1760) );
  XOR U4907 ( .A(n1764), .B(n1765), .Z(n1763) );
  XOR U4908 ( .A(DB[503]), .B(DB[496]), .Z(n1765) );
  AND U4909 ( .A(n1766), .B(n1767), .Z(n1764) );
  XOR U4910 ( .A(n1768), .B(n1769), .Z(n1767) );
  XOR U4911 ( .A(DB[496]), .B(DB[489]), .Z(n1769) );
  AND U4912 ( .A(n1770), .B(n1771), .Z(n1768) );
  XOR U4913 ( .A(n1772), .B(n1773), .Z(n1771) );
  XOR U4914 ( .A(DB[489]), .B(DB[482]), .Z(n1773) );
  AND U4915 ( .A(n1774), .B(n1775), .Z(n1772) );
  XOR U4916 ( .A(n1776), .B(n1777), .Z(n1775) );
  XOR U4917 ( .A(DB[482]), .B(DB[475]), .Z(n1777) );
  AND U4918 ( .A(n1778), .B(n1779), .Z(n1776) );
  XOR U4919 ( .A(n1780), .B(n1781), .Z(n1779) );
  XOR U4920 ( .A(DB[475]), .B(DB[468]), .Z(n1781) );
  AND U4921 ( .A(n1782), .B(n1783), .Z(n1780) );
  XOR U4922 ( .A(n1784), .B(n1785), .Z(n1783) );
  XOR U4923 ( .A(DB[468]), .B(DB[461]), .Z(n1785) );
  AND U4924 ( .A(n1786), .B(n1787), .Z(n1784) );
  XOR U4925 ( .A(n1788), .B(n1789), .Z(n1787) );
  XOR U4926 ( .A(DB[461]), .B(DB[454]), .Z(n1789) );
  AND U4927 ( .A(n1790), .B(n1791), .Z(n1788) );
  XOR U4928 ( .A(n1792), .B(n1793), .Z(n1791) );
  XOR U4929 ( .A(DB[454]), .B(DB[447]), .Z(n1793) );
  AND U4930 ( .A(n1794), .B(n1795), .Z(n1792) );
  XOR U4931 ( .A(n1796), .B(n1797), .Z(n1795) );
  XOR U4932 ( .A(DB[447]), .B(DB[440]), .Z(n1797) );
  AND U4933 ( .A(n1798), .B(n1799), .Z(n1796) );
  XOR U4934 ( .A(n1800), .B(n1801), .Z(n1799) );
  XOR U4935 ( .A(DB[440]), .B(DB[433]), .Z(n1801) );
  AND U4936 ( .A(n1802), .B(n1803), .Z(n1800) );
  XOR U4937 ( .A(n1804), .B(n1805), .Z(n1803) );
  XOR U4938 ( .A(DB[433]), .B(DB[426]), .Z(n1805) );
  AND U4939 ( .A(n1806), .B(n1807), .Z(n1804) );
  XOR U4940 ( .A(n1808), .B(n1809), .Z(n1807) );
  XOR U4941 ( .A(DB[426]), .B(DB[419]), .Z(n1809) );
  AND U4942 ( .A(n1810), .B(n1811), .Z(n1808) );
  XOR U4943 ( .A(n1812), .B(n1813), .Z(n1811) );
  XOR U4944 ( .A(DB[419]), .B(DB[412]), .Z(n1813) );
  AND U4945 ( .A(n1814), .B(n1815), .Z(n1812) );
  XOR U4946 ( .A(n1816), .B(n1817), .Z(n1815) );
  XOR U4947 ( .A(DB[412]), .B(DB[405]), .Z(n1817) );
  AND U4948 ( .A(n1818), .B(n1819), .Z(n1816) );
  XOR U4949 ( .A(n1820), .B(n1821), .Z(n1819) );
  XOR U4950 ( .A(DB[405]), .B(DB[398]), .Z(n1821) );
  AND U4951 ( .A(n1822), .B(n1823), .Z(n1820) );
  XOR U4952 ( .A(n1824), .B(n1825), .Z(n1823) );
  XOR U4953 ( .A(DB[398]), .B(DB[391]), .Z(n1825) );
  AND U4954 ( .A(n1826), .B(n1827), .Z(n1824) );
  XOR U4955 ( .A(n1828), .B(n1829), .Z(n1827) );
  XOR U4956 ( .A(DB[391]), .B(DB[384]), .Z(n1829) );
  AND U4957 ( .A(n1830), .B(n1831), .Z(n1828) );
  XOR U4958 ( .A(n1832), .B(n1833), .Z(n1831) );
  XOR U4959 ( .A(DB[384]), .B(DB[377]), .Z(n1833) );
  AND U4960 ( .A(n1834), .B(n1835), .Z(n1832) );
  XOR U4961 ( .A(n1836), .B(n1837), .Z(n1835) );
  XOR U4962 ( .A(DB[377]), .B(DB[370]), .Z(n1837) );
  AND U4963 ( .A(n1838), .B(n1839), .Z(n1836) );
  XOR U4964 ( .A(n1840), .B(n1841), .Z(n1839) );
  XOR U4965 ( .A(DB[370]), .B(DB[363]), .Z(n1841) );
  AND U4966 ( .A(n1842), .B(n1843), .Z(n1840) );
  XOR U4967 ( .A(n1844), .B(n1845), .Z(n1843) );
  XOR U4968 ( .A(DB[363]), .B(DB[356]), .Z(n1845) );
  AND U4969 ( .A(n1846), .B(n1847), .Z(n1844) );
  XOR U4970 ( .A(n1848), .B(n1849), .Z(n1847) );
  XOR U4971 ( .A(DB[356]), .B(DB[349]), .Z(n1849) );
  AND U4972 ( .A(n1850), .B(n1851), .Z(n1848) );
  XOR U4973 ( .A(n1852), .B(n1853), .Z(n1851) );
  XOR U4974 ( .A(DB[349]), .B(DB[342]), .Z(n1853) );
  AND U4975 ( .A(n1854), .B(n1855), .Z(n1852) );
  XOR U4976 ( .A(n1856), .B(n1857), .Z(n1855) );
  XOR U4977 ( .A(DB[342]), .B(DB[335]), .Z(n1857) );
  AND U4978 ( .A(n1858), .B(n1859), .Z(n1856) );
  XOR U4979 ( .A(n1860), .B(n1861), .Z(n1859) );
  XOR U4980 ( .A(DB[335]), .B(DB[328]), .Z(n1861) );
  AND U4981 ( .A(n1862), .B(n1863), .Z(n1860) );
  XOR U4982 ( .A(n1864), .B(n1865), .Z(n1863) );
  XOR U4983 ( .A(DB[328]), .B(DB[321]), .Z(n1865) );
  AND U4984 ( .A(n1866), .B(n1867), .Z(n1864) );
  XOR U4985 ( .A(n1868), .B(n1869), .Z(n1867) );
  XOR U4986 ( .A(DB[321]), .B(DB[314]), .Z(n1869) );
  AND U4987 ( .A(n1870), .B(n1871), .Z(n1868) );
  XOR U4988 ( .A(n1872), .B(n1873), .Z(n1871) );
  XOR U4989 ( .A(DB[314]), .B(DB[307]), .Z(n1873) );
  AND U4990 ( .A(n1874), .B(n1875), .Z(n1872) );
  XOR U4991 ( .A(n1876), .B(n1877), .Z(n1875) );
  XOR U4992 ( .A(DB[307]), .B(DB[300]), .Z(n1877) );
  AND U4993 ( .A(n1878), .B(n1879), .Z(n1876) );
  XOR U4994 ( .A(n1880), .B(n1881), .Z(n1879) );
  XOR U4995 ( .A(DB[300]), .B(DB[293]), .Z(n1881) );
  AND U4996 ( .A(n1882), .B(n1883), .Z(n1880) );
  XOR U4997 ( .A(n1884), .B(n1885), .Z(n1883) );
  XOR U4998 ( .A(DB[293]), .B(DB[286]), .Z(n1885) );
  AND U4999 ( .A(n1886), .B(n1887), .Z(n1884) );
  XOR U5000 ( .A(n1888), .B(n1889), .Z(n1887) );
  XOR U5001 ( .A(DB[286]), .B(DB[279]), .Z(n1889) );
  AND U5002 ( .A(n1890), .B(n1891), .Z(n1888) );
  XOR U5003 ( .A(n1892), .B(n1893), .Z(n1891) );
  XOR U5004 ( .A(DB[279]), .B(DB[272]), .Z(n1893) );
  AND U5005 ( .A(n1894), .B(n1895), .Z(n1892) );
  XOR U5006 ( .A(n1896), .B(n1897), .Z(n1895) );
  XOR U5007 ( .A(DB[272]), .B(DB[265]), .Z(n1897) );
  AND U5008 ( .A(n1898), .B(n1899), .Z(n1896) );
  XOR U5009 ( .A(n1900), .B(n1901), .Z(n1899) );
  XOR U5010 ( .A(DB[265]), .B(DB[258]), .Z(n1901) );
  AND U5011 ( .A(n1902), .B(n1903), .Z(n1900) );
  XOR U5012 ( .A(n1904), .B(n1905), .Z(n1903) );
  XOR U5013 ( .A(DB[258]), .B(DB[251]), .Z(n1905) );
  AND U5014 ( .A(n1906), .B(n1907), .Z(n1904) );
  XOR U5015 ( .A(n1908), .B(n1909), .Z(n1907) );
  XOR U5016 ( .A(DB[251]), .B(DB[244]), .Z(n1909) );
  AND U5017 ( .A(n1910), .B(n1911), .Z(n1908) );
  XOR U5018 ( .A(n1912), .B(n1913), .Z(n1911) );
  XOR U5019 ( .A(DB[244]), .B(DB[237]), .Z(n1913) );
  AND U5020 ( .A(n1914), .B(n1915), .Z(n1912) );
  XOR U5021 ( .A(n1916), .B(n1917), .Z(n1915) );
  XOR U5022 ( .A(DB[237]), .B(DB[230]), .Z(n1917) );
  AND U5023 ( .A(n1918), .B(n1919), .Z(n1916) );
  XOR U5024 ( .A(n1920), .B(n1921), .Z(n1919) );
  XOR U5025 ( .A(DB[230]), .B(DB[223]), .Z(n1921) );
  AND U5026 ( .A(n1922), .B(n1923), .Z(n1920) );
  XOR U5027 ( .A(n1924), .B(n1925), .Z(n1923) );
  XOR U5028 ( .A(DB[223]), .B(DB[216]), .Z(n1925) );
  AND U5029 ( .A(n1926), .B(n1927), .Z(n1924) );
  XOR U5030 ( .A(n1928), .B(n1929), .Z(n1927) );
  XOR U5031 ( .A(DB[216]), .B(DB[209]), .Z(n1929) );
  AND U5032 ( .A(n1930), .B(n1931), .Z(n1928) );
  XOR U5033 ( .A(n1932), .B(n1933), .Z(n1931) );
  XOR U5034 ( .A(DB[209]), .B(DB[202]), .Z(n1933) );
  AND U5035 ( .A(n1934), .B(n1935), .Z(n1932) );
  XOR U5036 ( .A(n1936), .B(n1937), .Z(n1935) );
  XOR U5037 ( .A(DB[202]), .B(DB[195]), .Z(n1937) );
  AND U5038 ( .A(n1938), .B(n1939), .Z(n1936) );
  XOR U5039 ( .A(n1940), .B(n1941), .Z(n1939) );
  XOR U5040 ( .A(DB[195]), .B(DB[188]), .Z(n1941) );
  AND U5041 ( .A(n1942), .B(n1943), .Z(n1940) );
  XOR U5042 ( .A(n1944), .B(n1945), .Z(n1943) );
  XOR U5043 ( .A(DB[188]), .B(DB[181]), .Z(n1945) );
  AND U5044 ( .A(n1946), .B(n1947), .Z(n1944) );
  XOR U5045 ( .A(n1948), .B(n1949), .Z(n1947) );
  XOR U5046 ( .A(DB[181]), .B(DB[174]), .Z(n1949) );
  AND U5047 ( .A(n1950), .B(n1951), .Z(n1948) );
  XOR U5048 ( .A(n1952), .B(n1953), .Z(n1951) );
  XOR U5049 ( .A(DB[174]), .B(DB[167]), .Z(n1953) );
  AND U5050 ( .A(n1954), .B(n1955), .Z(n1952) );
  XOR U5051 ( .A(n1956), .B(n1957), .Z(n1955) );
  XOR U5052 ( .A(DB[167]), .B(DB[160]), .Z(n1957) );
  AND U5053 ( .A(n1958), .B(n1959), .Z(n1956) );
  XOR U5054 ( .A(n1960), .B(n1961), .Z(n1959) );
  XOR U5055 ( .A(DB[160]), .B(DB[153]), .Z(n1961) );
  AND U5056 ( .A(n1962), .B(n1963), .Z(n1960) );
  XOR U5057 ( .A(n1964), .B(n1965), .Z(n1963) );
  XOR U5058 ( .A(DB[153]), .B(DB[146]), .Z(n1965) );
  AND U5059 ( .A(n1966), .B(n1967), .Z(n1964) );
  XOR U5060 ( .A(n1968), .B(n1969), .Z(n1967) );
  XOR U5061 ( .A(DB[146]), .B(DB[139]), .Z(n1969) );
  AND U5062 ( .A(n1970), .B(n1971), .Z(n1968) );
  XOR U5063 ( .A(n1972), .B(n1973), .Z(n1971) );
  XOR U5064 ( .A(DB[139]), .B(DB[132]), .Z(n1973) );
  AND U5065 ( .A(n1974), .B(n1975), .Z(n1972) );
  XOR U5066 ( .A(n1976), .B(n1977), .Z(n1975) );
  XOR U5067 ( .A(DB[132]), .B(DB[125]), .Z(n1977) );
  AND U5068 ( .A(n1978), .B(n1979), .Z(n1976) );
  XOR U5069 ( .A(n1980), .B(n1981), .Z(n1979) );
  XOR U5070 ( .A(DB[125]), .B(DB[118]), .Z(n1981) );
  AND U5071 ( .A(n1982), .B(n1983), .Z(n1980) );
  XOR U5072 ( .A(n1984), .B(n1985), .Z(n1983) );
  XOR U5073 ( .A(DB[118]), .B(DB[111]), .Z(n1985) );
  AND U5074 ( .A(n1986), .B(n1987), .Z(n1984) );
  XOR U5075 ( .A(n1988), .B(n1989), .Z(n1987) );
  XOR U5076 ( .A(DB[111]), .B(DB[104]), .Z(n1989) );
  AND U5077 ( .A(n1990), .B(n1991), .Z(n1988) );
  XOR U5078 ( .A(n1992), .B(n1993), .Z(n1991) );
  XOR U5079 ( .A(DB[97]), .B(DB[104]), .Z(n1993) );
  AND U5080 ( .A(n1994), .B(n1995), .Z(n1992) );
  XOR U5081 ( .A(n1996), .B(n1997), .Z(n1995) );
  XOR U5082 ( .A(DB[97]), .B(DB[90]), .Z(n1997) );
  AND U5083 ( .A(n1998), .B(n1999), .Z(n1996) );
  XOR U5084 ( .A(n2000), .B(n2001), .Z(n1999) );
  XOR U5085 ( .A(DB[90]), .B(DB[83]), .Z(n2001) );
  AND U5086 ( .A(n2002), .B(n2003), .Z(n2000) );
  XOR U5087 ( .A(n2004), .B(n2005), .Z(n2003) );
  XOR U5088 ( .A(DB[83]), .B(DB[76]), .Z(n2005) );
  AND U5089 ( .A(n2006), .B(n2007), .Z(n2004) );
  XOR U5090 ( .A(n2008), .B(n2009), .Z(n2007) );
  XOR U5091 ( .A(DB[76]), .B(DB[69]), .Z(n2009) );
  AND U5092 ( .A(n2010), .B(n2011), .Z(n2008) );
  XOR U5093 ( .A(n2012), .B(n2013), .Z(n2011) );
  XOR U5094 ( .A(DB[69]), .B(DB[62]), .Z(n2013) );
  AND U5095 ( .A(n2014), .B(n2015), .Z(n2012) );
  XOR U5096 ( .A(n2016), .B(n2017), .Z(n2015) );
  XOR U5097 ( .A(DB[62]), .B(DB[55]), .Z(n2017) );
  AND U5098 ( .A(n2018), .B(n2019), .Z(n2016) );
  XOR U5099 ( .A(n2020), .B(n2021), .Z(n2019) );
  XOR U5100 ( .A(DB[55]), .B(DB[48]), .Z(n2021) );
  AND U5101 ( .A(n2022), .B(n2023), .Z(n2020) );
  XOR U5102 ( .A(n2024), .B(n2025), .Z(n2023) );
  XOR U5103 ( .A(DB[48]), .B(DB[41]), .Z(n2025) );
  AND U5104 ( .A(n2026), .B(n2027), .Z(n2024) );
  XOR U5105 ( .A(n2028), .B(n2029), .Z(n2027) );
  XOR U5106 ( .A(DB[41]), .B(DB[34]), .Z(n2029) );
  AND U5107 ( .A(n2030), .B(n2031), .Z(n2028) );
  XOR U5108 ( .A(n2032), .B(n2033), .Z(n2031) );
  XOR U5109 ( .A(DB[34]), .B(DB[27]), .Z(n2033) );
  AND U5110 ( .A(n2034), .B(n2035), .Z(n2032) );
  XOR U5111 ( .A(n2036), .B(n2037), .Z(n2035) );
  XOR U5112 ( .A(DB[27]), .B(DB[20]), .Z(n2037) );
  AND U5113 ( .A(n2038), .B(n2039), .Z(n2036) );
  XOR U5114 ( .A(n2040), .B(n2041), .Z(n2039) );
  XOR U5115 ( .A(DB[20]), .B(DB[13]), .Z(n2041) );
  AND U5116 ( .A(n2042), .B(n2043), .Z(n2040) );
  XOR U5117 ( .A(DB[6]), .B(DB[13]), .Z(n2043) );
  XOR U5118 ( .A(DB[3582]), .B(n2044), .Z(min_val_out[5]) );
  AND U5119 ( .A(n2), .B(n2045), .Z(n2044) );
  XOR U5120 ( .A(n2046), .B(n2047), .Z(n2045) );
  XOR U5121 ( .A(DB[3582]), .B(DB[3575]), .Z(n2047) );
  AND U5122 ( .A(n6), .B(n2048), .Z(n2046) );
  XOR U5123 ( .A(n2049), .B(n2050), .Z(n2048) );
  XOR U5124 ( .A(DB[3575]), .B(DB[3568]), .Z(n2050) );
  AND U5125 ( .A(n10), .B(n2051), .Z(n2049) );
  XOR U5126 ( .A(n2052), .B(n2053), .Z(n2051) );
  XOR U5127 ( .A(DB[3568]), .B(DB[3561]), .Z(n2053) );
  AND U5128 ( .A(n14), .B(n2054), .Z(n2052) );
  XOR U5129 ( .A(n2055), .B(n2056), .Z(n2054) );
  XOR U5130 ( .A(DB[3561]), .B(DB[3554]), .Z(n2056) );
  AND U5131 ( .A(n18), .B(n2057), .Z(n2055) );
  XOR U5132 ( .A(n2058), .B(n2059), .Z(n2057) );
  XOR U5133 ( .A(DB[3554]), .B(DB[3547]), .Z(n2059) );
  AND U5134 ( .A(n22), .B(n2060), .Z(n2058) );
  XOR U5135 ( .A(n2061), .B(n2062), .Z(n2060) );
  XOR U5136 ( .A(DB[3547]), .B(DB[3540]), .Z(n2062) );
  AND U5137 ( .A(n26), .B(n2063), .Z(n2061) );
  XOR U5138 ( .A(n2064), .B(n2065), .Z(n2063) );
  XOR U5139 ( .A(DB[3540]), .B(DB[3533]), .Z(n2065) );
  AND U5140 ( .A(n30), .B(n2066), .Z(n2064) );
  XOR U5141 ( .A(n2067), .B(n2068), .Z(n2066) );
  XOR U5142 ( .A(DB[3533]), .B(DB[3526]), .Z(n2068) );
  AND U5143 ( .A(n34), .B(n2069), .Z(n2067) );
  XOR U5144 ( .A(n2070), .B(n2071), .Z(n2069) );
  XOR U5145 ( .A(DB[3526]), .B(DB[3519]), .Z(n2071) );
  AND U5146 ( .A(n38), .B(n2072), .Z(n2070) );
  XOR U5147 ( .A(n2073), .B(n2074), .Z(n2072) );
  XOR U5148 ( .A(DB[3519]), .B(DB[3512]), .Z(n2074) );
  AND U5149 ( .A(n42), .B(n2075), .Z(n2073) );
  XOR U5150 ( .A(n2076), .B(n2077), .Z(n2075) );
  XOR U5151 ( .A(DB[3512]), .B(DB[3505]), .Z(n2077) );
  AND U5152 ( .A(n46), .B(n2078), .Z(n2076) );
  XOR U5153 ( .A(n2079), .B(n2080), .Z(n2078) );
  XOR U5154 ( .A(DB[3505]), .B(DB[3498]), .Z(n2080) );
  AND U5155 ( .A(n50), .B(n2081), .Z(n2079) );
  XOR U5156 ( .A(n2082), .B(n2083), .Z(n2081) );
  XOR U5157 ( .A(DB[3498]), .B(DB[3491]), .Z(n2083) );
  AND U5158 ( .A(n54), .B(n2084), .Z(n2082) );
  XOR U5159 ( .A(n2085), .B(n2086), .Z(n2084) );
  XOR U5160 ( .A(DB[3491]), .B(DB[3484]), .Z(n2086) );
  AND U5161 ( .A(n58), .B(n2087), .Z(n2085) );
  XOR U5162 ( .A(n2088), .B(n2089), .Z(n2087) );
  XOR U5163 ( .A(DB[3484]), .B(DB[3477]), .Z(n2089) );
  AND U5164 ( .A(n62), .B(n2090), .Z(n2088) );
  XOR U5165 ( .A(n2091), .B(n2092), .Z(n2090) );
  XOR U5166 ( .A(DB[3477]), .B(DB[3470]), .Z(n2092) );
  AND U5167 ( .A(n66), .B(n2093), .Z(n2091) );
  XOR U5168 ( .A(n2094), .B(n2095), .Z(n2093) );
  XOR U5169 ( .A(DB[3470]), .B(DB[3463]), .Z(n2095) );
  AND U5170 ( .A(n70), .B(n2096), .Z(n2094) );
  XOR U5171 ( .A(n2097), .B(n2098), .Z(n2096) );
  XOR U5172 ( .A(DB[3463]), .B(DB[3456]), .Z(n2098) );
  AND U5173 ( .A(n74), .B(n2099), .Z(n2097) );
  XOR U5174 ( .A(n2100), .B(n2101), .Z(n2099) );
  XOR U5175 ( .A(DB[3456]), .B(DB[3449]), .Z(n2101) );
  AND U5176 ( .A(n78), .B(n2102), .Z(n2100) );
  XOR U5177 ( .A(n2103), .B(n2104), .Z(n2102) );
  XOR U5178 ( .A(DB[3449]), .B(DB[3442]), .Z(n2104) );
  AND U5179 ( .A(n82), .B(n2105), .Z(n2103) );
  XOR U5180 ( .A(n2106), .B(n2107), .Z(n2105) );
  XOR U5181 ( .A(DB[3442]), .B(DB[3435]), .Z(n2107) );
  AND U5182 ( .A(n86), .B(n2108), .Z(n2106) );
  XOR U5183 ( .A(n2109), .B(n2110), .Z(n2108) );
  XOR U5184 ( .A(DB[3435]), .B(DB[3428]), .Z(n2110) );
  AND U5185 ( .A(n90), .B(n2111), .Z(n2109) );
  XOR U5186 ( .A(n2112), .B(n2113), .Z(n2111) );
  XOR U5187 ( .A(DB[3428]), .B(DB[3421]), .Z(n2113) );
  AND U5188 ( .A(n94), .B(n2114), .Z(n2112) );
  XOR U5189 ( .A(n2115), .B(n2116), .Z(n2114) );
  XOR U5190 ( .A(DB[3421]), .B(DB[3414]), .Z(n2116) );
  AND U5191 ( .A(n98), .B(n2117), .Z(n2115) );
  XOR U5192 ( .A(n2118), .B(n2119), .Z(n2117) );
  XOR U5193 ( .A(DB[3414]), .B(DB[3407]), .Z(n2119) );
  AND U5194 ( .A(n102), .B(n2120), .Z(n2118) );
  XOR U5195 ( .A(n2121), .B(n2122), .Z(n2120) );
  XOR U5196 ( .A(DB[3407]), .B(DB[3400]), .Z(n2122) );
  AND U5197 ( .A(n106), .B(n2123), .Z(n2121) );
  XOR U5198 ( .A(n2124), .B(n2125), .Z(n2123) );
  XOR U5199 ( .A(DB[3400]), .B(DB[3393]), .Z(n2125) );
  AND U5200 ( .A(n110), .B(n2126), .Z(n2124) );
  XOR U5201 ( .A(n2127), .B(n2128), .Z(n2126) );
  XOR U5202 ( .A(DB[3393]), .B(DB[3386]), .Z(n2128) );
  AND U5203 ( .A(n114), .B(n2129), .Z(n2127) );
  XOR U5204 ( .A(n2130), .B(n2131), .Z(n2129) );
  XOR U5205 ( .A(DB[3386]), .B(DB[3379]), .Z(n2131) );
  AND U5206 ( .A(n118), .B(n2132), .Z(n2130) );
  XOR U5207 ( .A(n2133), .B(n2134), .Z(n2132) );
  XOR U5208 ( .A(DB[3379]), .B(DB[3372]), .Z(n2134) );
  AND U5209 ( .A(n122), .B(n2135), .Z(n2133) );
  XOR U5210 ( .A(n2136), .B(n2137), .Z(n2135) );
  XOR U5211 ( .A(DB[3372]), .B(DB[3365]), .Z(n2137) );
  AND U5212 ( .A(n126), .B(n2138), .Z(n2136) );
  XOR U5213 ( .A(n2139), .B(n2140), .Z(n2138) );
  XOR U5214 ( .A(DB[3365]), .B(DB[3358]), .Z(n2140) );
  AND U5215 ( .A(n130), .B(n2141), .Z(n2139) );
  XOR U5216 ( .A(n2142), .B(n2143), .Z(n2141) );
  XOR U5217 ( .A(DB[3358]), .B(DB[3351]), .Z(n2143) );
  AND U5218 ( .A(n134), .B(n2144), .Z(n2142) );
  XOR U5219 ( .A(n2145), .B(n2146), .Z(n2144) );
  XOR U5220 ( .A(DB[3351]), .B(DB[3344]), .Z(n2146) );
  AND U5221 ( .A(n138), .B(n2147), .Z(n2145) );
  XOR U5222 ( .A(n2148), .B(n2149), .Z(n2147) );
  XOR U5223 ( .A(DB[3344]), .B(DB[3337]), .Z(n2149) );
  AND U5224 ( .A(n142), .B(n2150), .Z(n2148) );
  XOR U5225 ( .A(n2151), .B(n2152), .Z(n2150) );
  XOR U5226 ( .A(DB[3337]), .B(DB[3330]), .Z(n2152) );
  AND U5227 ( .A(n146), .B(n2153), .Z(n2151) );
  XOR U5228 ( .A(n2154), .B(n2155), .Z(n2153) );
  XOR U5229 ( .A(DB[3330]), .B(DB[3323]), .Z(n2155) );
  AND U5230 ( .A(n150), .B(n2156), .Z(n2154) );
  XOR U5231 ( .A(n2157), .B(n2158), .Z(n2156) );
  XOR U5232 ( .A(DB[3323]), .B(DB[3316]), .Z(n2158) );
  AND U5233 ( .A(n154), .B(n2159), .Z(n2157) );
  XOR U5234 ( .A(n2160), .B(n2161), .Z(n2159) );
  XOR U5235 ( .A(DB[3316]), .B(DB[3309]), .Z(n2161) );
  AND U5236 ( .A(n158), .B(n2162), .Z(n2160) );
  XOR U5237 ( .A(n2163), .B(n2164), .Z(n2162) );
  XOR U5238 ( .A(DB[3309]), .B(DB[3302]), .Z(n2164) );
  AND U5239 ( .A(n162), .B(n2165), .Z(n2163) );
  XOR U5240 ( .A(n2166), .B(n2167), .Z(n2165) );
  XOR U5241 ( .A(DB[3302]), .B(DB[3295]), .Z(n2167) );
  AND U5242 ( .A(n166), .B(n2168), .Z(n2166) );
  XOR U5243 ( .A(n2169), .B(n2170), .Z(n2168) );
  XOR U5244 ( .A(DB[3295]), .B(DB[3288]), .Z(n2170) );
  AND U5245 ( .A(n170), .B(n2171), .Z(n2169) );
  XOR U5246 ( .A(n2172), .B(n2173), .Z(n2171) );
  XOR U5247 ( .A(DB[3288]), .B(DB[3281]), .Z(n2173) );
  AND U5248 ( .A(n174), .B(n2174), .Z(n2172) );
  XOR U5249 ( .A(n2175), .B(n2176), .Z(n2174) );
  XOR U5250 ( .A(DB[3281]), .B(DB[3274]), .Z(n2176) );
  AND U5251 ( .A(n178), .B(n2177), .Z(n2175) );
  XOR U5252 ( .A(n2178), .B(n2179), .Z(n2177) );
  XOR U5253 ( .A(DB[3274]), .B(DB[3267]), .Z(n2179) );
  AND U5254 ( .A(n182), .B(n2180), .Z(n2178) );
  XOR U5255 ( .A(n2181), .B(n2182), .Z(n2180) );
  XOR U5256 ( .A(DB[3267]), .B(DB[3260]), .Z(n2182) );
  AND U5257 ( .A(n186), .B(n2183), .Z(n2181) );
  XOR U5258 ( .A(n2184), .B(n2185), .Z(n2183) );
  XOR U5259 ( .A(DB[3260]), .B(DB[3253]), .Z(n2185) );
  AND U5260 ( .A(n190), .B(n2186), .Z(n2184) );
  XOR U5261 ( .A(n2187), .B(n2188), .Z(n2186) );
  XOR U5262 ( .A(DB[3253]), .B(DB[3246]), .Z(n2188) );
  AND U5263 ( .A(n194), .B(n2189), .Z(n2187) );
  XOR U5264 ( .A(n2190), .B(n2191), .Z(n2189) );
  XOR U5265 ( .A(DB[3246]), .B(DB[3239]), .Z(n2191) );
  AND U5266 ( .A(n198), .B(n2192), .Z(n2190) );
  XOR U5267 ( .A(n2193), .B(n2194), .Z(n2192) );
  XOR U5268 ( .A(DB[3239]), .B(DB[3232]), .Z(n2194) );
  AND U5269 ( .A(n202), .B(n2195), .Z(n2193) );
  XOR U5270 ( .A(n2196), .B(n2197), .Z(n2195) );
  XOR U5271 ( .A(DB[3232]), .B(DB[3225]), .Z(n2197) );
  AND U5272 ( .A(n206), .B(n2198), .Z(n2196) );
  XOR U5273 ( .A(n2199), .B(n2200), .Z(n2198) );
  XOR U5274 ( .A(DB[3225]), .B(DB[3218]), .Z(n2200) );
  AND U5275 ( .A(n210), .B(n2201), .Z(n2199) );
  XOR U5276 ( .A(n2202), .B(n2203), .Z(n2201) );
  XOR U5277 ( .A(DB[3218]), .B(DB[3211]), .Z(n2203) );
  AND U5278 ( .A(n214), .B(n2204), .Z(n2202) );
  XOR U5279 ( .A(n2205), .B(n2206), .Z(n2204) );
  XOR U5280 ( .A(DB[3211]), .B(DB[3204]), .Z(n2206) );
  AND U5281 ( .A(n218), .B(n2207), .Z(n2205) );
  XOR U5282 ( .A(n2208), .B(n2209), .Z(n2207) );
  XOR U5283 ( .A(DB[3204]), .B(DB[3197]), .Z(n2209) );
  AND U5284 ( .A(n222), .B(n2210), .Z(n2208) );
  XOR U5285 ( .A(n2211), .B(n2212), .Z(n2210) );
  XOR U5286 ( .A(DB[3197]), .B(DB[3190]), .Z(n2212) );
  AND U5287 ( .A(n226), .B(n2213), .Z(n2211) );
  XOR U5288 ( .A(n2214), .B(n2215), .Z(n2213) );
  XOR U5289 ( .A(DB[3190]), .B(DB[3183]), .Z(n2215) );
  AND U5290 ( .A(n230), .B(n2216), .Z(n2214) );
  XOR U5291 ( .A(n2217), .B(n2218), .Z(n2216) );
  XOR U5292 ( .A(DB[3183]), .B(DB[3176]), .Z(n2218) );
  AND U5293 ( .A(n234), .B(n2219), .Z(n2217) );
  XOR U5294 ( .A(n2220), .B(n2221), .Z(n2219) );
  XOR U5295 ( .A(DB[3176]), .B(DB[3169]), .Z(n2221) );
  AND U5296 ( .A(n238), .B(n2222), .Z(n2220) );
  XOR U5297 ( .A(n2223), .B(n2224), .Z(n2222) );
  XOR U5298 ( .A(DB[3169]), .B(DB[3162]), .Z(n2224) );
  AND U5299 ( .A(n242), .B(n2225), .Z(n2223) );
  XOR U5300 ( .A(n2226), .B(n2227), .Z(n2225) );
  XOR U5301 ( .A(DB[3162]), .B(DB[3155]), .Z(n2227) );
  AND U5302 ( .A(n246), .B(n2228), .Z(n2226) );
  XOR U5303 ( .A(n2229), .B(n2230), .Z(n2228) );
  XOR U5304 ( .A(DB[3155]), .B(DB[3148]), .Z(n2230) );
  AND U5305 ( .A(n250), .B(n2231), .Z(n2229) );
  XOR U5306 ( .A(n2232), .B(n2233), .Z(n2231) );
  XOR U5307 ( .A(DB[3148]), .B(DB[3141]), .Z(n2233) );
  AND U5308 ( .A(n254), .B(n2234), .Z(n2232) );
  XOR U5309 ( .A(n2235), .B(n2236), .Z(n2234) );
  XOR U5310 ( .A(DB[3141]), .B(DB[3134]), .Z(n2236) );
  AND U5311 ( .A(n258), .B(n2237), .Z(n2235) );
  XOR U5312 ( .A(n2238), .B(n2239), .Z(n2237) );
  XOR U5313 ( .A(DB[3134]), .B(DB[3127]), .Z(n2239) );
  AND U5314 ( .A(n262), .B(n2240), .Z(n2238) );
  XOR U5315 ( .A(n2241), .B(n2242), .Z(n2240) );
  XOR U5316 ( .A(DB[3127]), .B(DB[3120]), .Z(n2242) );
  AND U5317 ( .A(n266), .B(n2243), .Z(n2241) );
  XOR U5318 ( .A(n2244), .B(n2245), .Z(n2243) );
  XOR U5319 ( .A(DB[3120]), .B(DB[3113]), .Z(n2245) );
  AND U5320 ( .A(n270), .B(n2246), .Z(n2244) );
  XOR U5321 ( .A(n2247), .B(n2248), .Z(n2246) );
  XOR U5322 ( .A(DB[3113]), .B(DB[3106]), .Z(n2248) );
  AND U5323 ( .A(n274), .B(n2249), .Z(n2247) );
  XOR U5324 ( .A(n2250), .B(n2251), .Z(n2249) );
  XOR U5325 ( .A(DB[3106]), .B(DB[3099]), .Z(n2251) );
  AND U5326 ( .A(n278), .B(n2252), .Z(n2250) );
  XOR U5327 ( .A(n2253), .B(n2254), .Z(n2252) );
  XOR U5328 ( .A(DB[3099]), .B(DB[3092]), .Z(n2254) );
  AND U5329 ( .A(n282), .B(n2255), .Z(n2253) );
  XOR U5330 ( .A(n2256), .B(n2257), .Z(n2255) );
  XOR U5331 ( .A(DB[3092]), .B(DB[3085]), .Z(n2257) );
  AND U5332 ( .A(n286), .B(n2258), .Z(n2256) );
  XOR U5333 ( .A(n2259), .B(n2260), .Z(n2258) );
  XOR U5334 ( .A(DB[3085]), .B(DB[3078]), .Z(n2260) );
  AND U5335 ( .A(n290), .B(n2261), .Z(n2259) );
  XOR U5336 ( .A(n2262), .B(n2263), .Z(n2261) );
  XOR U5337 ( .A(DB[3078]), .B(DB[3071]), .Z(n2263) );
  AND U5338 ( .A(n294), .B(n2264), .Z(n2262) );
  XOR U5339 ( .A(n2265), .B(n2266), .Z(n2264) );
  XOR U5340 ( .A(DB[3071]), .B(DB[3064]), .Z(n2266) );
  AND U5341 ( .A(n298), .B(n2267), .Z(n2265) );
  XOR U5342 ( .A(n2268), .B(n2269), .Z(n2267) );
  XOR U5343 ( .A(DB[3064]), .B(DB[3057]), .Z(n2269) );
  AND U5344 ( .A(n302), .B(n2270), .Z(n2268) );
  XOR U5345 ( .A(n2271), .B(n2272), .Z(n2270) );
  XOR U5346 ( .A(DB[3057]), .B(DB[3050]), .Z(n2272) );
  AND U5347 ( .A(n306), .B(n2273), .Z(n2271) );
  XOR U5348 ( .A(n2274), .B(n2275), .Z(n2273) );
  XOR U5349 ( .A(DB[3050]), .B(DB[3043]), .Z(n2275) );
  AND U5350 ( .A(n310), .B(n2276), .Z(n2274) );
  XOR U5351 ( .A(n2277), .B(n2278), .Z(n2276) );
  XOR U5352 ( .A(DB[3043]), .B(DB[3036]), .Z(n2278) );
  AND U5353 ( .A(n314), .B(n2279), .Z(n2277) );
  XOR U5354 ( .A(n2280), .B(n2281), .Z(n2279) );
  XOR U5355 ( .A(DB[3036]), .B(DB[3029]), .Z(n2281) );
  AND U5356 ( .A(n318), .B(n2282), .Z(n2280) );
  XOR U5357 ( .A(n2283), .B(n2284), .Z(n2282) );
  XOR U5358 ( .A(DB[3029]), .B(DB[3022]), .Z(n2284) );
  AND U5359 ( .A(n322), .B(n2285), .Z(n2283) );
  XOR U5360 ( .A(n2286), .B(n2287), .Z(n2285) );
  XOR U5361 ( .A(DB[3022]), .B(DB[3015]), .Z(n2287) );
  AND U5362 ( .A(n326), .B(n2288), .Z(n2286) );
  XOR U5363 ( .A(n2289), .B(n2290), .Z(n2288) );
  XOR U5364 ( .A(DB[3015]), .B(DB[3008]), .Z(n2290) );
  AND U5365 ( .A(n330), .B(n2291), .Z(n2289) );
  XOR U5366 ( .A(n2292), .B(n2293), .Z(n2291) );
  XOR U5367 ( .A(DB[3008]), .B(DB[3001]), .Z(n2293) );
  AND U5368 ( .A(n334), .B(n2294), .Z(n2292) );
  XOR U5369 ( .A(n2295), .B(n2296), .Z(n2294) );
  XOR U5370 ( .A(DB[3001]), .B(DB[2994]), .Z(n2296) );
  AND U5371 ( .A(n338), .B(n2297), .Z(n2295) );
  XOR U5372 ( .A(n2298), .B(n2299), .Z(n2297) );
  XOR U5373 ( .A(DB[2994]), .B(DB[2987]), .Z(n2299) );
  AND U5374 ( .A(n342), .B(n2300), .Z(n2298) );
  XOR U5375 ( .A(n2301), .B(n2302), .Z(n2300) );
  XOR U5376 ( .A(DB[2987]), .B(DB[2980]), .Z(n2302) );
  AND U5377 ( .A(n346), .B(n2303), .Z(n2301) );
  XOR U5378 ( .A(n2304), .B(n2305), .Z(n2303) );
  XOR U5379 ( .A(DB[2980]), .B(DB[2973]), .Z(n2305) );
  AND U5380 ( .A(n350), .B(n2306), .Z(n2304) );
  XOR U5381 ( .A(n2307), .B(n2308), .Z(n2306) );
  XOR U5382 ( .A(DB[2973]), .B(DB[2966]), .Z(n2308) );
  AND U5383 ( .A(n354), .B(n2309), .Z(n2307) );
  XOR U5384 ( .A(n2310), .B(n2311), .Z(n2309) );
  XOR U5385 ( .A(DB[2966]), .B(DB[2959]), .Z(n2311) );
  AND U5386 ( .A(n358), .B(n2312), .Z(n2310) );
  XOR U5387 ( .A(n2313), .B(n2314), .Z(n2312) );
  XOR U5388 ( .A(DB[2959]), .B(DB[2952]), .Z(n2314) );
  AND U5389 ( .A(n362), .B(n2315), .Z(n2313) );
  XOR U5390 ( .A(n2316), .B(n2317), .Z(n2315) );
  XOR U5391 ( .A(DB[2952]), .B(DB[2945]), .Z(n2317) );
  AND U5392 ( .A(n366), .B(n2318), .Z(n2316) );
  XOR U5393 ( .A(n2319), .B(n2320), .Z(n2318) );
  XOR U5394 ( .A(DB[2945]), .B(DB[2938]), .Z(n2320) );
  AND U5395 ( .A(n370), .B(n2321), .Z(n2319) );
  XOR U5396 ( .A(n2322), .B(n2323), .Z(n2321) );
  XOR U5397 ( .A(DB[2938]), .B(DB[2931]), .Z(n2323) );
  AND U5398 ( .A(n374), .B(n2324), .Z(n2322) );
  XOR U5399 ( .A(n2325), .B(n2326), .Z(n2324) );
  XOR U5400 ( .A(DB[2931]), .B(DB[2924]), .Z(n2326) );
  AND U5401 ( .A(n378), .B(n2327), .Z(n2325) );
  XOR U5402 ( .A(n2328), .B(n2329), .Z(n2327) );
  XOR U5403 ( .A(DB[2924]), .B(DB[2917]), .Z(n2329) );
  AND U5404 ( .A(n382), .B(n2330), .Z(n2328) );
  XOR U5405 ( .A(n2331), .B(n2332), .Z(n2330) );
  XOR U5406 ( .A(DB[2917]), .B(DB[2910]), .Z(n2332) );
  AND U5407 ( .A(n386), .B(n2333), .Z(n2331) );
  XOR U5408 ( .A(n2334), .B(n2335), .Z(n2333) );
  XOR U5409 ( .A(DB[2910]), .B(DB[2903]), .Z(n2335) );
  AND U5410 ( .A(n390), .B(n2336), .Z(n2334) );
  XOR U5411 ( .A(n2337), .B(n2338), .Z(n2336) );
  XOR U5412 ( .A(DB[2903]), .B(DB[2896]), .Z(n2338) );
  AND U5413 ( .A(n394), .B(n2339), .Z(n2337) );
  XOR U5414 ( .A(n2340), .B(n2341), .Z(n2339) );
  XOR U5415 ( .A(DB[2896]), .B(DB[2889]), .Z(n2341) );
  AND U5416 ( .A(n398), .B(n2342), .Z(n2340) );
  XOR U5417 ( .A(n2343), .B(n2344), .Z(n2342) );
  XOR U5418 ( .A(DB[2889]), .B(DB[2882]), .Z(n2344) );
  AND U5419 ( .A(n402), .B(n2345), .Z(n2343) );
  XOR U5420 ( .A(n2346), .B(n2347), .Z(n2345) );
  XOR U5421 ( .A(DB[2882]), .B(DB[2875]), .Z(n2347) );
  AND U5422 ( .A(n406), .B(n2348), .Z(n2346) );
  XOR U5423 ( .A(n2349), .B(n2350), .Z(n2348) );
  XOR U5424 ( .A(DB[2875]), .B(DB[2868]), .Z(n2350) );
  AND U5425 ( .A(n410), .B(n2351), .Z(n2349) );
  XOR U5426 ( .A(n2352), .B(n2353), .Z(n2351) );
  XOR U5427 ( .A(DB[2868]), .B(DB[2861]), .Z(n2353) );
  AND U5428 ( .A(n414), .B(n2354), .Z(n2352) );
  XOR U5429 ( .A(n2355), .B(n2356), .Z(n2354) );
  XOR U5430 ( .A(DB[2861]), .B(DB[2854]), .Z(n2356) );
  AND U5431 ( .A(n418), .B(n2357), .Z(n2355) );
  XOR U5432 ( .A(n2358), .B(n2359), .Z(n2357) );
  XOR U5433 ( .A(DB[2854]), .B(DB[2847]), .Z(n2359) );
  AND U5434 ( .A(n422), .B(n2360), .Z(n2358) );
  XOR U5435 ( .A(n2361), .B(n2362), .Z(n2360) );
  XOR U5436 ( .A(DB[2847]), .B(DB[2840]), .Z(n2362) );
  AND U5437 ( .A(n426), .B(n2363), .Z(n2361) );
  XOR U5438 ( .A(n2364), .B(n2365), .Z(n2363) );
  XOR U5439 ( .A(DB[2840]), .B(DB[2833]), .Z(n2365) );
  AND U5440 ( .A(n430), .B(n2366), .Z(n2364) );
  XOR U5441 ( .A(n2367), .B(n2368), .Z(n2366) );
  XOR U5442 ( .A(DB[2833]), .B(DB[2826]), .Z(n2368) );
  AND U5443 ( .A(n434), .B(n2369), .Z(n2367) );
  XOR U5444 ( .A(n2370), .B(n2371), .Z(n2369) );
  XOR U5445 ( .A(DB[2826]), .B(DB[2819]), .Z(n2371) );
  AND U5446 ( .A(n438), .B(n2372), .Z(n2370) );
  XOR U5447 ( .A(n2373), .B(n2374), .Z(n2372) );
  XOR U5448 ( .A(DB[2819]), .B(DB[2812]), .Z(n2374) );
  AND U5449 ( .A(n442), .B(n2375), .Z(n2373) );
  XOR U5450 ( .A(n2376), .B(n2377), .Z(n2375) );
  XOR U5451 ( .A(DB[2812]), .B(DB[2805]), .Z(n2377) );
  AND U5452 ( .A(n446), .B(n2378), .Z(n2376) );
  XOR U5453 ( .A(n2379), .B(n2380), .Z(n2378) );
  XOR U5454 ( .A(DB[2805]), .B(DB[2798]), .Z(n2380) );
  AND U5455 ( .A(n450), .B(n2381), .Z(n2379) );
  XOR U5456 ( .A(n2382), .B(n2383), .Z(n2381) );
  XOR U5457 ( .A(DB[2798]), .B(DB[2791]), .Z(n2383) );
  AND U5458 ( .A(n454), .B(n2384), .Z(n2382) );
  XOR U5459 ( .A(n2385), .B(n2386), .Z(n2384) );
  XOR U5460 ( .A(DB[2791]), .B(DB[2784]), .Z(n2386) );
  AND U5461 ( .A(n458), .B(n2387), .Z(n2385) );
  XOR U5462 ( .A(n2388), .B(n2389), .Z(n2387) );
  XOR U5463 ( .A(DB[2784]), .B(DB[2777]), .Z(n2389) );
  AND U5464 ( .A(n462), .B(n2390), .Z(n2388) );
  XOR U5465 ( .A(n2391), .B(n2392), .Z(n2390) );
  XOR U5466 ( .A(DB[2777]), .B(DB[2770]), .Z(n2392) );
  AND U5467 ( .A(n466), .B(n2393), .Z(n2391) );
  XOR U5468 ( .A(n2394), .B(n2395), .Z(n2393) );
  XOR U5469 ( .A(DB[2770]), .B(DB[2763]), .Z(n2395) );
  AND U5470 ( .A(n470), .B(n2396), .Z(n2394) );
  XOR U5471 ( .A(n2397), .B(n2398), .Z(n2396) );
  XOR U5472 ( .A(DB[2763]), .B(DB[2756]), .Z(n2398) );
  AND U5473 ( .A(n474), .B(n2399), .Z(n2397) );
  XOR U5474 ( .A(n2400), .B(n2401), .Z(n2399) );
  XOR U5475 ( .A(DB[2756]), .B(DB[2749]), .Z(n2401) );
  AND U5476 ( .A(n478), .B(n2402), .Z(n2400) );
  XOR U5477 ( .A(n2403), .B(n2404), .Z(n2402) );
  XOR U5478 ( .A(DB[2749]), .B(DB[2742]), .Z(n2404) );
  AND U5479 ( .A(n482), .B(n2405), .Z(n2403) );
  XOR U5480 ( .A(n2406), .B(n2407), .Z(n2405) );
  XOR U5481 ( .A(DB[2742]), .B(DB[2735]), .Z(n2407) );
  AND U5482 ( .A(n486), .B(n2408), .Z(n2406) );
  XOR U5483 ( .A(n2409), .B(n2410), .Z(n2408) );
  XOR U5484 ( .A(DB[2735]), .B(DB[2728]), .Z(n2410) );
  AND U5485 ( .A(n490), .B(n2411), .Z(n2409) );
  XOR U5486 ( .A(n2412), .B(n2413), .Z(n2411) );
  XOR U5487 ( .A(DB[2728]), .B(DB[2721]), .Z(n2413) );
  AND U5488 ( .A(n494), .B(n2414), .Z(n2412) );
  XOR U5489 ( .A(n2415), .B(n2416), .Z(n2414) );
  XOR U5490 ( .A(DB[2721]), .B(DB[2714]), .Z(n2416) );
  AND U5491 ( .A(n498), .B(n2417), .Z(n2415) );
  XOR U5492 ( .A(n2418), .B(n2419), .Z(n2417) );
  XOR U5493 ( .A(DB[2714]), .B(DB[2707]), .Z(n2419) );
  AND U5494 ( .A(n502), .B(n2420), .Z(n2418) );
  XOR U5495 ( .A(n2421), .B(n2422), .Z(n2420) );
  XOR U5496 ( .A(DB[2707]), .B(DB[2700]), .Z(n2422) );
  AND U5497 ( .A(n506), .B(n2423), .Z(n2421) );
  XOR U5498 ( .A(n2424), .B(n2425), .Z(n2423) );
  XOR U5499 ( .A(DB[2700]), .B(DB[2693]), .Z(n2425) );
  AND U5500 ( .A(n510), .B(n2426), .Z(n2424) );
  XOR U5501 ( .A(n2427), .B(n2428), .Z(n2426) );
  XOR U5502 ( .A(DB[2693]), .B(DB[2686]), .Z(n2428) );
  AND U5503 ( .A(n514), .B(n2429), .Z(n2427) );
  XOR U5504 ( .A(n2430), .B(n2431), .Z(n2429) );
  XOR U5505 ( .A(DB[2686]), .B(DB[2679]), .Z(n2431) );
  AND U5506 ( .A(n518), .B(n2432), .Z(n2430) );
  XOR U5507 ( .A(n2433), .B(n2434), .Z(n2432) );
  XOR U5508 ( .A(DB[2679]), .B(DB[2672]), .Z(n2434) );
  AND U5509 ( .A(n522), .B(n2435), .Z(n2433) );
  XOR U5510 ( .A(n2436), .B(n2437), .Z(n2435) );
  XOR U5511 ( .A(DB[2672]), .B(DB[2665]), .Z(n2437) );
  AND U5512 ( .A(n526), .B(n2438), .Z(n2436) );
  XOR U5513 ( .A(n2439), .B(n2440), .Z(n2438) );
  XOR U5514 ( .A(DB[2665]), .B(DB[2658]), .Z(n2440) );
  AND U5515 ( .A(n530), .B(n2441), .Z(n2439) );
  XOR U5516 ( .A(n2442), .B(n2443), .Z(n2441) );
  XOR U5517 ( .A(DB[2658]), .B(DB[2651]), .Z(n2443) );
  AND U5518 ( .A(n534), .B(n2444), .Z(n2442) );
  XOR U5519 ( .A(n2445), .B(n2446), .Z(n2444) );
  XOR U5520 ( .A(DB[2651]), .B(DB[2644]), .Z(n2446) );
  AND U5521 ( .A(n538), .B(n2447), .Z(n2445) );
  XOR U5522 ( .A(n2448), .B(n2449), .Z(n2447) );
  XOR U5523 ( .A(DB[2644]), .B(DB[2637]), .Z(n2449) );
  AND U5524 ( .A(n542), .B(n2450), .Z(n2448) );
  XOR U5525 ( .A(n2451), .B(n2452), .Z(n2450) );
  XOR U5526 ( .A(DB[2637]), .B(DB[2630]), .Z(n2452) );
  AND U5527 ( .A(n546), .B(n2453), .Z(n2451) );
  XOR U5528 ( .A(n2454), .B(n2455), .Z(n2453) );
  XOR U5529 ( .A(DB[2630]), .B(DB[2623]), .Z(n2455) );
  AND U5530 ( .A(n550), .B(n2456), .Z(n2454) );
  XOR U5531 ( .A(n2457), .B(n2458), .Z(n2456) );
  XOR U5532 ( .A(DB[2623]), .B(DB[2616]), .Z(n2458) );
  AND U5533 ( .A(n554), .B(n2459), .Z(n2457) );
  XOR U5534 ( .A(n2460), .B(n2461), .Z(n2459) );
  XOR U5535 ( .A(DB[2616]), .B(DB[2609]), .Z(n2461) );
  AND U5536 ( .A(n558), .B(n2462), .Z(n2460) );
  XOR U5537 ( .A(n2463), .B(n2464), .Z(n2462) );
  XOR U5538 ( .A(DB[2609]), .B(DB[2602]), .Z(n2464) );
  AND U5539 ( .A(n562), .B(n2465), .Z(n2463) );
  XOR U5540 ( .A(n2466), .B(n2467), .Z(n2465) );
  XOR U5541 ( .A(DB[2602]), .B(DB[2595]), .Z(n2467) );
  AND U5542 ( .A(n566), .B(n2468), .Z(n2466) );
  XOR U5543 ( .A(n2469), .B(n2470), .Z(n2468) );
  XOR U5544 ( .A(DB[2595]), .B(DB[2588]), .Z(n2470) );
  AND U5545 ( .A(n570), .B(n2471), .Z(n2469) );
  XOR U5546 ( .A(n2472), .B(n2473), .Z(n2471) );
  XOR U5547 ( .A(DB[2588]), .B(DB[2581]), .Z(n2473) );
  AND U5548 ( .A(n574), .B(n2474), .Z(n2472) );
  XOR U5549 ( .A(n2475), .B(n2476), .Z(n2474) );
  XOR U5550 ( .A(DB[2581]), .B(DB[2574]), .Z(n2476) );
  AND U5551 ( .A(n578), .B(n2477), .Z(n2475) );
  XOR U5552 ( .A(n2478), .B(n2479), .Z(n2477) );
  XOR U5553 ( .A(DB[2574]), .B(DB[2567]), .Z(n2479) );
  AND U5554 ( .A(n582), .B(n2480), .Z(n2478) );
  XOR U5555 ( .A(n2481), .B(n2482), .Z(n2480) );
  XOR U5556 ( .A(DB[2567]), .B(DB[2560]), .Z(n2482) );
  AND U5557 ( .A(n586), .B(n2483), .Z(n2481) );
  XOR U5558 ( .A(n2484), .B(n2485), .Z(n2483) );
  XOR U5559 ( .A(DB[2560]), .B(DB[2553]), .Z(n2485) );
  AND U5560 ( .A(n590), .B(n2486), .Z(n2484) );
  XOR U5561 ( .A(n2487), .B(n2488), .Z(n2486) );
  XOR U5562 ( .A(DB[2553]), .B(DB[2546]), .Z(n2488) );
  AND U5563 ( .A(n594), .B(n2489), .Z(n2487) );
  XOR U5564 ( .A(n2490), .B(n2491), .Z(n2489) );
  XOR U5565 ( .A(DB[2546]), .B(DB[2539]), .Z(n2491) );
  AND U5566 ( .A(n598), .B(n2492), .Z(n2490) );
  XOR U5567 ( .A(n2493), .B(n2494), .Z(n2492) );
  XOR U5568 ( .A(DB[2539]), .B(DB[2532]), .Z(n2494) );
  AND U5569 ( .A(n602), .B(n2495), .Z(n2493) );
  XOR U5570 ( .A(n2496), .B(n2497), .Z(n2495) );
  XOR U5571 ( .A(DB[2532]), .B(DB[2525]), .Z(n2497) );
  AND U5572 ( .A(n606), .B(n2498), .Z(n2496) );
  XOR U5573 ( .A(n2499), .B(n2500), .Z(n2498) );
  XOR U5574 ( .A(DB[2525]), .B(DB[2518]), .Z(n2500) );
  AND U5575 ( .A(n610), .B(n2501), .Z(n2499) );
  XOR U5576 ( .A(n2502), .B(n2503), .Z(n2501) );
  XOR U5577 ( .A(DB[2518]), .B(DB[2511]), .Z(n2503) );
  AND U5578 ( .A(n614), .B(n2504), .Z(n2502) );
  XOR U5579 ( .A(n2505), .B(n2506), .Z(n2504) );
  XOR U5580 ( .A(DB[2511]), .B(DB[2504]), .Z(n2506) );
  AND U5581 ( .A(n618), .B(n2507), .Z(n2505) );
  XOR U5582 ( .A(n2508), .B(n2509), .Z(n2507) );
  XOR U5583 ( .A(DB[2504]), .B(DB[2497]), .Z(n2509) );
  AND U5584 ( .A(n622), .B(n2510), .Z(n2508) );
  XOR U5585 ( .A(n2511), .B(n2512), .Z(n2510) );
  XOR U5586 ( .A(DB[2497]), .B(DB[2490]), .Z(n2512) );
  AND U5587 ( .A(n626), .B(n2513), .Z(n2511) );
  XOR U5588 ( .A(n2514), .B(n2515), .Z(n2513) );
  XOR U5589 ( .A(DB[2490]), .B(DB[2483]), .Z(n2515) );
  AND U5590 ( .A(n630), .B(n2516), .Z(n2514) );
  XOR U5591 ( .A(n2517), .B(n2518), .Z(n2516) );
  XOR U5592 ( .A(DB[2483]), .B(DB[2476]), .Z(n2518) );
  AND U5593 ( .A(n634), .B(n2519), .Z(n2517) );
  XOR U5594 ( .A(n2520), .B(n2521), .Z(n2519) );
  XOR U5595 ( .A(DB[2476]), .B(DB[2469]), .Z(n2521) );
  AND U5596 ( .A(n638), .B(n2522), .Z(n2520) );
  XOR U5597 ( .A(n2523), .B(n2524), .Z(n2522) );
  XOR U5598 ( .A(DB[2469]), .B(DB[2462]), .Z(n2524) );
  AND U5599 ( .A(n642), .B(n2525), .Z(n2523) );
  XOR U5600 ( .A(n2526), .B(n2527), .Z(n2525) );
  XOR U5601 ( .A(DB[2462]), .B(DB[2455]), .Z(n2527) );
  AND U5602 ( .A(n646), .B(n2528), .Z(n2526) );
  XOR U5603 ( .A(n2529), .B(n2530), .Z(n2528) );
  XOR U5604 ( .A(DB[2455]), .B(DB[2448]), .Z(n2530) );
  AND U5605 ( .A(n650), .B(n2531), .Z(n2529) );
  XOR U5606 ( .A(n2532), .B(n2533), .Z(n2531) );
  XOR U5607 ( .A(DB[2448]), .B(DB[2441]), .Z(n2533) );
  AND U5608 ( .A(n654), .B(n2534), .Z(n2532) );
  XOR U5609 ( .A(n2535), .B(n2536), .Z(n2534) );
  XOR U5610 ( .A(DB[2441]), .B(DB[2434]), .Z(n2536) );
  AND U5611 ( .A(n658), .B(n2537), .Z(n2535) );
  XOR U5612 ( .A(n2538), .B(n2539), .Z(n2537) );
  XOR U5613 ( .A(DB[2434]), .B(DB[2427]), .Z(n2539) );
  AND U5614 ( .A(n662), .B(n2540), .Z(n2538) );
  XOR U5615 ( .A(n2541), .B(n2542), .Z(n2540) );
  XOR U5616 ( .A(DB[2427]), .B(DB[2420]), .Z(n2542) );
  AND U5617 ( .A(n666), .B(n2543), .Z(n2541) );
  XOR U5618 ( .A(n2544), .B(n2545), .Z(n2543) );
  XOR U5619 ( .A(DB[2420]), .B(DB[2413]), .Z(n2545) );
  AND U5620 ( .A(n670), .B(n2546), .Z(n2544) );
  XOR U5621 ( .A(n2547), .B(n2548), .Z(n2546) );
  XOR U5622 ( .A(DB[2413]), .B(DB[2406]), .Z(n2548) );
  AND U5623 ( .A(n674), .B(n2549), .Z(n2547) );
  XOR U5624 ( .A(n2550), .B(n2551), .Z(n2549) );
  XOR U5625 ( .A(DB[2406]), .B(DB[2399]), .Z(n2551) );
  AND U5626 ( .A(n678), .B(n2552), .Z(n2550) );
  XOR U5627 ( .A(n2553), .B(n2554), .Z(n2552) );
  XOR U5628 ( .A(DB[2399]), .B(DB[2392]), .Z(n2554) );
  AND U5629 ( .A(n682), .B(n2555), .Z(n2553) );
  XOR U5630 ( .A(n2556), .B(n2557), .Z(n2555) );
  XOR U5631 ( .A(DB[2392]), .B(DB[2385]), .Z(n2557) );
  AND U5632 ( .A(n686), .B(n2558), .Z(n2556) );
  XOR U5633 ( .A(n2559), .B(n2560), .Z(n2558) );
  XOR U5634 ( .A(DB[2385]), .B(DB[2378]), .Z(n2560) );
  AND U5635 ( .A(n690), .B(n2561), .Z(n2559) );
  XOR U5636 ( .A(n2562), .B(n2563), .Z(n2561) );
  XOR U5637 ( .A(DB[2378]), .B(DB[2371]), .Z(n2563) );
  AND U5638 ( .A(n694), .B(n2564), .Z(n2562) );
  XOR U5639 ( .A(n2565), .B(n2566), .Z(n2564) );
  XOR U5640 ( .A(DB[2371]), .B(DB[2364]), .Z(n2566) );
  AND U5641 ( .A(n698), .B(n2567), .Z(n2565) );
  XOR U5642 ( .A(n2568), .B(n2569), .Z(n2567) );
  XOR U5643 ( .A(DB[2364]), .B(DB[2357]), .Z(n2569) );
  AND U5644 ( .A(n702), .B(n2570), .Z(n2568) );
  XOR U5645 ( .A(n2571), .B(n2572), .Z(n2570) );
  XOR U5646 ( .A(DB[2357]), .B(DB[2350]), .Z(n2572) );
  AND U5647 ( .A(n706), .B(n2573), .Z(n2571) );
  XOR U5648 ( .A(n2574), .B(n2575), .Z(n2573) );
  XOR U5649 ( .A(DB[2350]), .B(DB[2343]), .Z(n2575) );
  AND U5650 ( .A(n710), .B(n2576), .Z(n2574) );
  XOR U5651 ( .A(n2577), .B(n2578), .Z(n2576) );
  XOR U5652 ( .A(DB[2343]), .B(DB[2336]), .Z(n2578) );
  AND U5653 ( .A(n714), .B(n2579), .Z(n2577) );
  XOR U5654 ( .A(n2580), .B(n2581), .Z(n2579) );
  XOR U5655 ( .A(DB[2336]), .B(DB[2329]), .Z(n2581) );
  AND U5656 ( .A(n718), .B(n2582), .Z(n2580) );
  XOR U5657 ( .A(n2583), .B(n2584), .Z(n2582) );
  XOR U5658 ( .A(DB[2329]), .B(DB[2322]), .Z(n2584) );
  AND U5659 ( .A(n722), .B(n2585), .Z(n2583) );
  XOR U5660 ( .A(n2586), .B(n2587), .Z(n2585) );
  XOR U5661 ( .A(DB[2322]), .B(DB[2315]), .Z(n2587) );
  AND U5662 ( .A(n726), .B(n2588), .Z(n2586) );
  XOR U5663 ( .A(n2589), .B(n2590), .Z(n2588) );
  XOR U5664 ( .A(DB[2315]), .B(DB[2308]), .Z(n2590) );
  AND U5665 ( .A(n730), .B(n2591), .Z(n2589) );
  XOR U5666 ( .A(n2592), .B(n2593), .Z(n2591) );
  XOR U5667 ( .A(DB[2308]), .B(DB[2301]), .Z(n2593) );
  AND U5668 ( .A(n734), .B(n2594), .Z(n2592) );
  XOR U5669 ( .A(n2595), .B(n2596), .Z(n2594) );
  XOR U5670 ( .A(DB[2301]), .B(DB[2294]), .Z(n2596) );
  AND U5671 ( .A(n738), .B(n2597), .Z(n2595) );
  XOR U5672 ( .A(n2598), .B(n2599), .Z(n2597) );
  XOR U5673 ( .A(DB[2294]), .B(DB[2287]), .Z(n2599) );
  AND U5674 ( .A(n742), .B(n2600), .Z(n2598) );
  XOR U5675 ( .A(n2601), .B(n2602), .Z(n2600) );
  XOR U5676 ( .A(DB[2287]), .B(DB[2280]), .Z(n2602) );
  AND U5677 ( .A(n746), .B(n2603), .Z(n2601) );
  XOR U5678 ( .A(n2604), .B(n2605), .Z(n2603) );
  XOR U5679 ( .A(DB[2280]), .B(DB[2273]), .Z(n2605) );
  AND U5680 ( .A(n750), .B(n2606), .Z(n2604) );
  XOR U5681 ( .A(n2607), .B(n2608), .Z(n2606) );
  XOR U5682 ( .A(DB[2273]), .B(DB[2266]), .Z(n2608) );
  AND U5683 ( .A(n754), .B(n2609), .Z(n2607) );
  XOR U5684 ( .A(n2610), .B(n2611), .Z(n2609) );
  XOR U5685 ( .A(DB[2266]), .B(DB[2259]), .Z(n2611) );
  AND U5686 ( .A(n758), .B(n2612), .Z(n2610) );
  XOR U5687 ( .A(n2613), .B(n2614), .Z(n2612) );
  XOR U5688 ( .A(DB[2259]), .B(DB[2252]), .Z(n2614) );
  AND U5689 ( .A(n762), .B(n2615), .Z(n2613) );
  XOR U5690 ( .A(n2616), .B(n2617), .Z(n2615) );
  XOR U5691 ( .A(DB[2252]), .B(DB[2245]), .Z(n2617) );
  AND U5692 ( .A(n766), .B(n2618), .Z(n2616) );
  XOR U5693 ( .A(n2619), .B(n2620), .Z(n2618) );
  XOR U5694 ( .A(DB[2245]), .B(DB[2238]), .Z(n2620) );
  AND U5695 ( .A(n770), .B(n2621), .Z(n2619) );
  XOR U5696 ( .A(n2622), .B(n2623), .Z(n2621) );
  XOR U5697 ( .A(DB[2238]), .B(DB[2231]), .Z(n2623) );
  AND U5698 ( .A(n774), .B(n2624), .Z(n2622) );
  XOR U5699 ( .A(n2625), .B(n2626), .Z(n2624) );
  XOR U5700 ( .A(DB[2231]), .B(DB[2224]), .Z(n2626) );
  AND U5701 ( .A(n778), .B(n2627), .Z(n2625) );
  XOR U5702 ( .A(n2628), .B(n2629), .Z(n2627) );
  XOR U5703 ( .A(DB[2224]), .B(DB[2217]), .Z(n2629) );
  AND U5704 ( .A(n782), .B(n2630), .Z(n2628) );
  XOR U5705 ( .A(n2631), .B(n2632), .Z(n2630) );
  XOR U5706 ( .A(DB[2217]), .B(DB[2210]), .Z(n2632) );
  AND U5707 ( .A(n786), .B(n2633), .Z(n2631) );
  XOR U5708 ( .A(n2634), .B(n2635), .Z(n2633) );
  XOR U5709 ( .A(DB[2210]), .B(DB[2203]), .Z(n2635) );
  AND U5710 ( .A(n790), .B(n2636), .Z(n2634) );
  XOR U5711 ( .A(n2637), .B(n2638), .Z(n2636) );
  XOR U5712 ( .A(DB[2203]), .B(DB[2196]), .Z(n2638) );
  AND U5713 ( .A(n794), .B(n2639), .Z(n2637) );
  XOR U5714 ( .A(n2640), .B(n2641), .Z(n2639) );
  XOR U5715 ( .A(DB[2196]), .B(DB[2189]), .Z(n2641) );
  AND U5716 ( .A(n798), .B(n2642), .Z(n2640) );
  XOR U5717 ( .A(n2643), .B(n2644), .Z(n2642) );
  XOR U5718 ( .A(DB[2189]), .B(DB[2182]), .Z(n2644) );
  AND U5719 ( .A(n802), .B(n2645), .Z(n2643) );
  XOR U5720 ( .A(n2646), .B(n2647), .Z(n2645) );
  XOR U5721 ( .A(DB[2182]), .B(DB[2175]), .Z(n2647) );
  AND U5722 ( .A(n806), .B(n2648), .Z(n2646) );
  XOR U5723 ( .A(n2649), .B(n2650), .Z(n2648) );
  XOR U5724 ( .A(DB[2175]), .B(DB[2168]), .Z(n2650) );
  AND U5725 ( .A(n810), .B(n2651), .Z(n2649) );
  XOR U5726 ( .A(n2652), .B(n2653), .Z(n2651) );
  XOR U5727 ( .A(DB[2168]), .B(DB[2161]), .Z(n2653) );
  AND U5728 ( .A(n814), .B(n2654), .Z(n2652) );
  XOR U5729 ( .A(n2655), .B(n2656), .Z(n2654) );
  XOR U5730 ( .A(DB[2161]), .B(DB[2154]), .Z(n2656) );
  AND U5731 ( .A(n818), .B(n2657), .Z(n2655) );
  XOR U5732 ( .A(n2658), .B(n2659), .Z(n2657) );
  XOR U5733 ( .A(DB[2154]), .B(DB[2147]), .Z(n2659) );
  AND U5734 ( .A(n822), .B(n2660), .Z(n2658) );
  XOR U5735 ( .A(n2661), .B(n2662), .Z(n2660) );
  XOR U5736 ( .A(DB[2147]), .B(DB[2140]), .Z(n2662) );
  AND U5737 ( .A(n826), .B(n2663), .Z(n2661) );
  XOR U5738 ( .A(n2664), .B(n2665), .Z(n2663) );
  XOR U5739 ( .A(DB[2140]), .B(DB[2133]), .Z(n2665) );
  AND U5740 ( .A(n830), .B(n2666), .Z(n2664) );
  XOR U5741 ( .A(n2667), .B(n2668), .Z(n2666) );
  XOR U5742 ( .A(DB[2133]), .B(DB[2126]), .Z(n2668) );
  AND U5743 ( .A(n834), .B(n2669), .Z(n2667) );
  XOR U5744 ( .A(n2670), .B(n2671), .Z(n2669) );
  XOR U5745 ( .A(DB[2126]), .B(DB[2119]), .Z(n2671) );
  AND U5746 ( .A(n838), .B(n2672), .Z(n2670) );
  XOR U5747 ( .A(n2673), .B(n2674), .Z(n2672) );
  XOR U5748 ( .A(DB[2119]), .B(DB[2112]), .Z(n2674) );
  AND U5749 ( .A(n842), .B(n2675), .Z(n2673) );
  XOR U5750 ( .A(n2676), .B(n2677), .Z(n2675) );
  XOR U5751 ( .A(DB[2112]), .B(DB[2105]), .Z(n2677) );
  AND U5752 ( .A(n846), .B(n2678), .Z(n2676) );
  XOR U5753 ( .A(n2679), .B(n2680), .Z(n2678) );
  XOR U5754 ( .A(DB[2105]), .B(DB[2098]), .Z(n2680) );
  AND U5755 ( .A(n850), .B(n2681), .Z(n2679) );
  XOR U5756 ( .A(n2682), .B(n2683), .Z(n2681) );
  XOR U5757 ( .A(DB[2098]), .B(DB[2091]), .Z(n2683) );
  AND U5758 ( .A(n854), .B(n2684), .Z(n2682) );
  XOR U5759 ( .A(n2685), .B(n2686), .Z(n2684) );
  XOR U5760 ( .A(DB[2091]), .B(DB[2084]), .Z(n2686) );
  AND U5761 ( .A(n858), .B(n2687), .Z(n2685) );
  XOR U5762 ( .A(n2688), .B(n2689), .Z(n2687) );
  XOR U5763 ( .A(DB[2084]), .B(DB[2077]), .Z(n2689) );
  AND U5764 ( .A(n862), .B(n2690), .Z(n2688) );
  XOR U5765 ( .A(n2691), .B(n2692), .Z(n2690) );
  XOR U5766 ( .A(DB[2077]), .B(DB[2070]), .Z(n2692) );
  AND U5767 ( .A(n866), .B(n2693), .Z(n2691) );
  XOR U5768 ( .A(n2694), .B(n2695), .Z(n2693) );
  XOR U5769 ( .A(DB[2070]), .B(DB[2063]), .Z(n2695) );
  AND U5770 ( .A(n870), .B(n2696), .Z(n2694) );
  XOR U5771 ( .A(n2697), .B(n2698), .Z(n2696) );
  XOR U5772 ( .A(DB[2063]), .B(DB[2056]), .Z(n2698) );
  AND U5773 ( .A(n874), .B(n2699), .Z(n2697) );
  XOR U5774 ( .A(n2700), .B(n2701), .Z(n2699) );
  XOR U5775 ( .A(DB[2056]), .B(DB[2049]), .Z(n2701) );
  AND U5776 ( .A(n878), .B(n2702), .Z(n2700) );
  XOR U5777 ( .A(n2703), .B(n2704), .Z(n2702) );
  XOR U5778 ( .A(DB[2049]), .B(DB[2042]), .Z(n2704) );
  AND U5779 ( .A(n882), .B(n2705), .Z(n2703) );
  XOR U5780 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR U5781 ( .A(DB[2042]), .B(DB[2035]), .Z(n2707) );
  AND U5782 ( .A(n886), .B(n2708), .Z(n2706) );
  XOR U5783 ( .A(n2709), .B(n2710), .Z(n2708) );
  XOR U5784 ( .A(DB[2035]), .B(DB[2028]), .Z(n2710) );
  AND U5785 ( .A(n890), .B(n2711), .Z(n2709) );
  XOR U5786 ( .A(n2712), .B(n2713), .Z(n2711) );
  XOR U5787 ( .A(DB[2028]), .B(DB[2021]), .Z(n2713) );
  AND U5788 ( .A(n894), .B(n2714), .Z(n2712) );
  XOR U5789 ( .A(n2715), .B(n2716), .Z(n2714) );
  XOR U5790 ( .A(DB[2021]), .B(DB[2014]), .Z(n2716) );
  AND U5791 ( .A(n898), .B(n2717), .Z(n2715) );
  XOR U5792 ( .A(n2718), .B(n2719), .Z(n2717) );
  XOR U5793 ( .A(DB[2014]), .B(DB[2007]), .Z(n2719) );
  AND U5794 ( .A(n902), .B(n2720), .Z(n2718) );
  XOR U5795 ( .A(n2721), .B(n2722), .Z(n2720) );
  XOR U5796 ( .A(DB[2007]), .B(DB[2000]), .Z(n2722) );
  AND U5797 ( .A(n906), .B(n2723), .Z(n2721) );
  XOR U5798 ( .A(n2724), .B(n2725), .Z(n2723) );
  XOR U5799 ( .A(DB[2000]), .B(DB[1993]), .Z(n2725) );
  AND U5800 ( .A(n910), .B(n2726), .Z(n2724) );
  XOR U5801 ( .A(n2727), .B(n2728), .Z(n2726) );
  XOR U5802 ( .A(DB[1993]), .B(DB[1986]), .Z(n2728) );
  AND U5803 ( .A(n914), .B(n2729), .Z(n2727) );
  XOR U5804 ( .A(n2730), .B(n2731), .Z(n2729) );
  XOR U5805 ( .A(DB[1986]), .B(DB[1979]), .Z(n2731) );
  AND U5806 ( .A(n918), .B(n2732), .Z(n2730) );
  XOR U5807 ( .A(n2733), .B(n2734), .Z(n2732) );
  XOR U5808 ( .A(DB[1979]), .B(DB[1972]), .Z(n2734) );
  AND U5809 ( .A(n922), .B(n2735), .Z(n2733) );
  XOR U5810 ( .A(n2736), .B(n2737), .Z(n2735) );
  XOR U5811 ( .A(DB[1972]), .B(DB[1965]), .Z(n2737) );
  AND U5812 ( .A(n926), .B(n2738), .Z(n2736) );
  XOR U5813 ( .A(n2739), .B(n2740), .Z(n2738) );
  XOR U5814 ( .A(DB[1965]), .B(DB[1958]), .Z(n2740) );
  AND U5815 ( .A(n930), .B(n2741), .Z(n2739) );
  XOR U5816 ( .A(n2742), .B(n2743), .Z(n2741) );
  XOR U5817 ( .A(DB[1958]), .B(DB[1951]), .Z(n2743) );
  AND U5818 ( .A(n934), .B(n2744), .Z(n2742) );
  XOR U5819 ( .A(n2745), .B(n2746), .Z(n2744) );
  XOR U5820 ( .A(DB[1951]), .B(DB[1944]), .Z(n2746) );
  AND U5821 ( .A(n938), .B(n2747), .Z(n2745) );
  XOR U5822 ( .A(n2748), .B(n2749), .Z(n2747) );
  XOR U5823 ( .A(DB[1944]), .B(DB[1937]), .Z(n2749) );
  AND U5824 ( .A(n942), .B(n2750), .Z(n2748) );
  XOR U5825 ( .A(n2751), .B(n2752), .Z(n2750) );
  XOR U5826 ( .A(DB[1937]), .B(DB[1930]), .Z(n2752) );
  AND U5827 ( .A(n946), .B(n2753), .Z(n2751) );
  XOR U5828 ( .A(n2754), .B(n2755), .Z(n2753) );
  XOR U5829 ( .A(DB[1930]), .B(DB[1923]), .Z(n2755) );
  AND U5830 ( .A(n950), .B(n2756), .Z(n2754) );
  XOR U5831 ( .A(n2757), .B(n2758), .Z(n2756) );
  XOR U5832 ( .A(DB[1923]), .B(DB[1916]), .Z(n2758) );
  AND U5833 ( .A(n954), .B(n2759), .Z(n2757) );
  XOR U5834 ( .A(n2760), .B(n2761), .Z(n2759) );
  XOR U5835 ( .A(DB[1916]), .B(DB[1909]), .Z(n2761) );
  AND U5836 ( .A(n958), .B(n2762), .Z(n2760) );
  XOR U5837 ( .A(n2763), .B(n2764), .Z(n2762) );
  XOR U5838 ( .A(DB[1909]), .B(DB[1902]), .Z(n2764) );
  AND U5839 ( .A(n962), .B(n2765), .Z(n2763) );
  XOR U5840 ( .A(n2766), .B(n2767), .Z(n2765) );
  XOR U5841 ( .A(DB[1902]), .B(DB[1895]), .Z(n2767) );
  AND U5842 ( .A(n966), .B(n2768), .Z(n2766) );
  XOR U5843 ( .A(n2769), .B(n2770), .Z(n2768) );
  XOR U5844 ( .A(DB[1895]), .B(DB[1888]), .Z(n2770) );
  AND U5845 ( .A(n970), .B(n2771), .Z(n2769) );
  XOR U5846 ( .A(n2772), .B(n2773), .Z(n2771) );
  XOR U5847 ( .A(DB[1888]), .B(DB[1881]), .Z(n2773) );
  AND U5848 ( .A(n974), .B(n2774), .Z(n2772) );
  XOR U5849 ( .A(n2775), .B(n2776), .Z(n2774) );
  XOR U5850 ( .A(DB[1881]), .B(DB[1874]), .Z(n2776) );
  AND U5851 ( .A(n978), .B(n2777), .Z(n2775) );
  XOR U5852 ( .A(n2778), .B(n2779), .Z(n2777) );
  XOR U5853 ( .A(DB[1874]), .B(DB[1867]), .Z(n2779) );
  AND U5854 ( .A(n982), .B(n2780), .Z(n2778) );
  XOR U5855 ( .A(n2781), .B(n2782), .Z(n2780) );
  XOR U5856 ( .A(DB[1867]), .B(DB[1860]), .Z(n2782) );
  AND U5857 ( .A(n986), .B(n2783), .Z(n2781) );
  XOR U5858 ( .A(n2784), .B(n2785), .Z(n2783) );
  XOR U5859 ( .A(DB[1860]), .B(DB[1853]), .Z(n2785) );
  AND U5860 ( .A(n990), .B(n2786), .Z(n2784) );
  XOR U5861 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR U5862 ( .A(DB[1853]), .B(DB[1846]), .Z(n2788) );
  AND U5863 ( .A(n994), .B(n2789), .Z(n2787) );
  XOR U5864 ( .A(n2790), .B(n2791), .Z(n2789) );
  XOR U5865 ( .A(DB[1846]), .B(DB[1839]), .Z(n2791) );
  AND U5866 ( .A(n998), .B(n2792), .Z(n2790) );
  XOR U5867 ( .A(n2793), .B(n2794), .Z(n2792) );
  XOR U5868 ( .A(DB[1839]), .B(DB[1832]), .Z(n2794) );
  AND U5869 ( .A(n1002), .B(n2795), .Z(n2793) );
  XOR U5870 ( .A(n2796), .B(n2797), .Z(n2795) );
  XOR U5871 ( .A(DB[1832]), .B(DB[1825]), .Z(n2797) );
  AND U5872 ( .A(n1006), .B(n2798), .Z(n2796) );
  XOR U5873 ( .A(n2799), .B(n2800), .Z(n2798) );
  XOR U5874 ( .A(DB[1825]), .B(DB[1818]), .Z(n2800) );
  AND U5875 ( .A(n1010), .B(n2801), .Z(n2799) );
  XOR U5876 ( .A(n2802), .B(n2803), .Z(n2801) );
  XOR U5877 ( .A(DB[1818]), .B(DB[1811]), .Z(n2803) );
  AND U5878 ( .A(n1014), .B(n2804), .Z(n2802) );
  XOR U5879 ( .A(n2805), .B(n2806), .Z(n2804) );
  XOR U5880 ( .A(DB[1811]), .B(DB[1804]), .Z(n2806) );
  AND U5881 ( .A(n1018), .B(n2807), .Z(n2805) );
  XOR U5882 ( .A(n2808), .B(n2809), .Z(n2807) );
  XOR U5883 ( .A(DB[1804]), .B(DB[1797]), .Z(n2809) );
  AND U5884 ( .A(n1022), .B(n2810), .Z(n2808) );
  XOR U5885 ( .A(n2811), .B(n2812), .Z(n2810) );
  XOR U5886 ( .A(DB[1797]), .B(DB[1790]), .Z(n2812) );
  AND U5887 ( .A(n1026), .B(n2813), .Z(n2811) );
  XOR U5888 ( .A(n2814), .B(n2815), .Z(n2813) );
  XOR U5889 ( .A(DB[1790]), .B(DB[1783]), .Z(n2815) );
  AND U5890 ( .A(n1030), .B(n2816), .Z(n2814) );
  XOR U5891 ( .A(n2817), .B(n2818), .Z(n2816) );
  XOR U5892 ( .A(DB[1783]), .B(DB[1776]), .Z(n2818) );
  AND U5893 ( .A(n1034), .B(n2819), .Z(n2817) );
  XOR U5894 ( .A(n2820), .B(n2821), .Z(n2819) );
  XOR U5895 ( .A(DB[1776]), .B(DB[1769]), .Z(n2821) );
  AND U5896 ( .A(n1038), .B(n2822), .Z(n2820) );
  XOR U5897 ( .A(n2823), .B(n2824), .Z(n2822) );
  XOR U5898 ( .A(DB[1769]), .B(DB[1762]), .Z(n2824) );
  AND U5899 ( .A(n1042), .B(n2825), .Z(n2823) );
  XOR U5900 ( .A(n2826), .B(n2827), .Z(n2825) );
  XOR U5901 ( .A(DB[1762]), .B(DB[1755]), .Z(n2827) );
  AND U5902 ( .A(n1046), .B(n2828), .Z(n2826) );
  XOR U5903 ( .A(n2829), .B(n2830), .Z(n2828) );
  XOR U5904 ( .A(DB[1755]), .B(DB[1748]), .Z(n2830) );
  AND U5905 ( .A(n1050), .B(n2831), .Z(n2829) );
  XOR U5906 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U5907 ( .A(DB[1748]), .B(DB[1741]), .Z(n2833) );
  AND U5908 ( .A(n1054), .B(n2834), .Z(n2832) );
  XOR U5909 ( .A(n2835), .B(n2836), .Z(n2834) );
  XOR U5910 ( .A(DB[1741]), .B(DB[1734]), .Z(n2836) );
  AND U5911 ( .A(n1058), .B(n2837), .Z(n2835) );
  XOR U5912 ( .A(n2838), .B(n2839), .Z(n2837) );
  XOR U5913 ( .A(DB[1734]), .B(DB[1727]), .Z(n2839) );
  AND U5914 ( .A(n1062), .B(n2840), .Z(n2838) );
  XOR U5915 ( .A(n2841), .B(n2842), .Z(n2840) );
  XOR U5916 ( .A(DB[1727]), .B(DB[1720]), .Z(n2842) );
  AND U5917 ( .A(n1066), .B(n2843), .Z(n2841) );
  XOR U5918 ( .A(n2844), .B(n2845), .Z(n2843) );
  XOR U5919 ( .A(DB[1720]), .B(DB[1713]), .Z(n2845) );
  AND U5920 ( .A(n1070), .B(n2846), .Z(n2844) );
  XOR U5921 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR U5922 ( .A(DB[1713]), .B(DB[1706]), .Z(n2848) );
  AND U5923 ( .A(n1074), .B(n2849), .Z(n2847) );
  XOR U5924 ( .A(n2850), .B(n2851), .Z(n2849) );
  XOR U5925 ( .A(DB[1706]), .B(DB[1699]), .Z(n2851) );
  AND U5926 ( .A(n1078), .B(n2852), .Z(n2850) );
  XOR U5927 ( .A(n2853), .B(n2854), .Z(n2852) );
  XOR U5928 ( .A(DB[1699]), .B(DB[1692]), .Z(n2854) );
  AND U5929 ( .A(n1082), .B(n2855), .Z(n2853) );
  XOR U5930 ( .A(n2856), .B(n2857), .Z(n2855) );
  XOR U5931 ( .A(DB[1692]), .B(DB[1685]), .Z(n2857) );
  AND U5932 ( .A(n1086), .B(n2858), .Z(n2856) );
  XOR U5933 ( .A(n2859), .B(n2860), .Z(n2858) );
  XOR U5934 ( .A(DB[1685]), .B(DB[1678]), .Z(n2860) );
  AND U5935 ( .A(n1090), .B(n2861), .Z(n2859) );
  XOR U5936 ( .A(n2862), .B(n2863), .Z(n2861) );
  XOR U5937 ( .A(DB[1678]), .B(DB[1671]), .Z(n2863) );
  AND U5938 ( .A(n1094), .B(n2864), .Z(n2862) );
  XOR U5939 ( .A(n2865), .B(n2866), .Z(n2864) );
  XOR U5940 ( .A(DB[1671]), .B(DB[1664]), .Z(n2866) );
  AND U5941 ( .A(n1098), .B(n2867), .Z(n2865) );
  XOR U5942 ( .A(n2868), .B(n2869), .Z(n2867) );
  XOR U5943 ( .A(DB[1664]), .B(DB[1657]), .Z(n2869) );
  AND U5944 ( .A(n1102), .B(n2870), .Z(n2868) );
  XOR U5945 ( .A(n2871), .B(n2872), .Z(n2870) );
  XOR U5946 ( .A(DB[1657]), .B(DB[1650]), .Z(n2872) );
  AND U5947 ( .A(n1106), .B(n2873), .Z(n2871) );
  XOR U5948 ( .A(n2874), .B(n2875), .Z(n2873) );
  XOR U5949 ( .A(DB[1650]), .B(DB[1643]), .Z(n2875) );
  AND U5950 ( .A(n1110), .B(n2876), .Z(n2874) );
  XOR U5951 ( .A(n2877), .B(n2878), .Z(n2876) );
  XOR U5952 ( .A(DB[1643]), .B(DB[1636]), .Z(n2878) );
  AND U5953 ( .A(n1114), .B(n2879), .Z(n2877) );
  XOR U5954 ( .A(n2880), .B(n2881), .Z(n2879) );
  XOR U5955 ( .A(DB[1636]), .B(DB[1629]), .Z(n2881) );
  AND U5956 ( .A(n1118), .B(n2882), .Z(n2880) );
  XOR U5957 ( .A(n2883), .B(n2884), .Z(n2882) );
  XOR U5958 ( .A(DB[1629]), .B(DB[1622]), .Z(n2884) );
  AND U5959 ( .A(n1122), .B(n2885), .Z(n2883) );
  XOR U5960 ( .A(n2886), .B(n2887), .Z(n2885) );
  XOR U5961 ( .A(DB[1622]), .B(DB[1615]), .Z(n2887) );
  AND U5962 ( .A(n1126), .B(n2888), .Z(n2886) );
  XOR U5963 ( .A(n2889), .B(n2890), .Z(n2888) );
  XOR U5964 ( .A(DB[1615]), .B(DB[1608]), .Z(n2890) );
  AND U5965 ( .A(n1130), .B(n2891), .Z(n2889) );
  XOR U5966 ( .A(n2892), .B(n2893), .Z(n2891) );
  XOR U5967 ( .A(DB[1608]), .B(DB[1601]), .Z(n2893) );
  AND U5968 ( .A(n1134), .B(n2894), .Z(n2892) );
  XOR U5969 ( .A(n2895), .B(n2896), .Z(n2894) );
  XOR U5970 ( .A(DB[1601]), .B(DB[1594]), .Z(n2896) );
  AND U5971 ( .A(n1138), .B(n2897), .Z(n2895) );
  XOR U5972 ( .A(n2898), .B(n2899), .Z(n2897) );
  XOR U5973 ( .A(DB[1594]), .B(DB[1587]), .Z(n2899) );
  AND U5974 ( .A(n1142), .B(n2900), .Z(n2898) );
  XOR U5975 ( .A(n2901), .B(n2902), .Z(n2900) );
  XOR U5976 ( .A(DB[1587]), .B(DB[1580]), .Z(n2902) );
  AND U5977 ( .A(n1146), .B(n2903), .Z(n2901) );
  XOR U5978 ( .A(n2904), .B(n2905), .Z(n2903) );
  XOR U5979 ( .A(DB[1580]), .B(DB[1573]), .Z(n2905) );
  AND U5980 ( .A(n1150), .B(n2906), .Z(n2904) );
  XOR U5981 ( .A(n2907), .B(n2908), .Z(n2906) );
  XOR U5982 ( .A(DB[1573]), .B(DB[1566]), .Z(n2908) );
  AND U5983 ( .A(n1154), .B(n2909), .Z(n2907) );
  XOR U5984 ( .A(n2910), .B(n2911), .Z(n2909) );
  XOR U5985 ( .A(DB[1566]), .B(DB[1559]), .Z(n2911) );
  AND U5986 ( .A(n1158), .B(n2912), .Z(n2910) );
  XOR U5987 ( .A(n2913), .B(n2914), .Z(n2912) );
  XOR U5988 ( .A(DB[1559]), .B(DB[1552]), .Z(n2914) );
  AND U5989 ( .A(n1162), .B(n2915), .Z(n2913) );
  XOR U5990 ( .A(n2916), .B(n2917), .Z(n2915) );
  XOR U5991 ( .A(DB[1552]), .B(DB[1545]), .Z(n2917) );
  AND U5992 ( .A(n1166), .B(n2918), .Z(n2916) );
  XOR U5993 ( .A(n2919), .B(n2920), .Z(n2918) );
  XOR U5994 ( .A(DB[1545]), .B(DB[1538]), .Z(n2920) );
  AND U5995 ( .A(n1170), .B(n2921), .Z(n2919) );
  XOR U5996 ( .A(n2922), .B(n2923), .Z(n2921) );
  XOR U5997 ( .A(DB[1538]), .B(DB[1531]), .Z(n2923) );
  AND U5998 ( .A(n1174), .B(n2924), .Z(n2922) );
  XOR U5999 ( .A(n2925), .B(n2926), .Z(n2924) );
  XOR U6000 ( .A(DB[1531]), .B(DB[1524]), .Z(n2926) );
  AND U6001 ( .A(n1178), .B(n2927), .Z(n2925) );
  XOR U6002 ( .A(n2928), .B(n2929), .Z(n2927) );
  XOR U6003 ( .A(DB[1524]), .B(DB[1517]), .Z(n2929) );
  AND U6004 ( .A(n1182), .B(n2930), .Z(n2928) );
  XOR U6005 ( .A(n2931), .B(n2932), .Z(n2930) );
  XOR U6006 ( .A(DB[1517]), .B(DB[1510]), .Z(n2932) );
  AND U6007 ( .A(n1186), .B(n2933), .Z(n2931) );
  XOR U6008 ( .A(n2934), .B(n2935), .Z(n2933) );
  XOR U6009 ( .A(DB[1510]), .B(DB[1503]), .Z(n2935) );
  AND U6010 ( .A(n1190), .B(n2936), .Z(n2934) );
  XOR U6011 ( .A(n2937), .B(n2938), .Z(n2936) );
  XOR U6012 ( .A(DB[1503]), .B(DB[1496]), .Z(n2938) );
  AND U6013 ( .A(n1194), .B(n2939), .Z(n2937) );
  XOR U6014 ( .A(n2940), .B(n2941), .Z(n2939) );
  XOR U6015 ( .A(DB[1496]), .B(DB[1489]), .Z(n2941) );
  AND U6016 ( .A(n1198), .B(n2942), .Z(n2940) );
  XOR U6017 ( .A(n2943), .B(n2944), .Z(n2942) );
  XOR U6018 ( .A(DB[1489]), .B(DB[1482]), .Z(n2944) );
  AND U6019 ( .A(n1202), .B(n2945), .Z(n2943) );
  XOR U6020 ( .A(n2946), .B(n2947), .Z(n2945) );
  XOR U6021 ( .A(DB[1482]), .B(DB[1475]), .Z(n2947) );
  AND U6022 ( .A(n1206), .B(n2948), .Z(n2946) );
  XOR U6023 ( .A(n2949), .B(n2950), .Z(n2948) );
  XOR U6024 ( .A(DB[1475]), .B(DB[1468]), .Z(n2950) );
  AND U6025 ( .A(n1210), .B(n2951), .Z(n2949) );
  XOR U6026 ( .A(n2952), .B(n2953), .Z(n2951) );
  XOR U6027 ( .A(DB[1468]), .B(DB[1461]), .Z(n2953) );
  AND U6028 ( .A(n1214), .B(n2954), .Z(n2952) );
  XOR U6029 ( .A(n2955), .B(n2956), .Z(n2954) );
  XOR U6030 ( .A(DB[1461]), .B(DB[1454]), .Z(n2956) );
  AND U6031 ( .A(n1218), .B(n2957), .Z(n2955) );
  XOR U6032 ( .A(n2958), .B(n2959), .Z(n2957) );
  XOR U6033 ( .A(DB[1454]), .B(DB[1447]), .Z(n2959) );
  AND U6034 ( .A(n1222), .B(n2960), .Z(n2958) );
  XOR U6035 ( .A(n2961), .B(n2962), .Z(n2960) );
  XOR U6036 ( .A(DB[1447]), .B(DB[1440]), .Z(n2962) );
  AND U6037 ( .A(n1226), .B(n2963), .Z(n2961) );
  XOR U6038 ( .A(n2964), .B(n2965), .Z(n2963) );
  XOR U6039 ( .A(DB[1440]), .B(DB[1433]), .Z(n2965) );
  AND U6040 ( .A(n1230), .B(n2966), .Z(n2964) );
  XOR U6041 ( .A(n2967), .B(n2968), .Z(n2966) );
  XOR U6042 ( .A(DB[1433]), .B(DB[1426]), .Z(n2968) );
  AND U6043 ( .A(n1234), .B(n2969), .Z(n2967) );
  XOR U6044 ( .A(n2970), .B(n2971), .Z(n2969) );
  XOR U6045 ( .A(DB[1426]), .B(DB[1419]), .Z(n2971) );
  AND U6046 ( .A(n1238), .B(n2972), .Z(n2970) );
  XOR U6047 ( .A(n2973), .B(n2974), .Z(n2972) );
  XOR U6048 ( .A(DB[1419]), .B(DB[1412]), .Z(n2974) );
  AND U6049 ( .A(n1242), .B(n2975), .Z(n2973) );
  XOR U6050 ( .A(n2976), .B(n2977), .Z(n2975) );
  XOR U6051 ( .A(DB[1412]), .B(DB[1405]), .Z(n2977) );
  AND U6052 ( .A(n1246), .B(n2978), .Z(n2976) );
  XOR U6053 ( .A(n2979), .B(n2980), .Z(n2978) );
  XOR U6054 ( .A(DB[1405]), .B(DB[1398]), .Z(n2980) );
  AND U6055 ( .A(n1250), .B(n2981), .Z(n2979) );
  XOR U6056 ( .A(n2982), .B(n2983), .Z(n2981) );
  XOR U6057 ( .A(DB[1398]), .B(DB[1391]), .Z(n2983) );
  AND U6058 ( .A(n1254), .B(n2984), .Z(n2982) );
  XOR U6059 ( .A(n2985), .B(n2986), .Z(n2984) );
  XOR U6060 ( .A(DB[1391]), .B(DB[1384]), .Z(n2986) );
  AND U6061 ( .A(n1258), .B(n2987), .Z(n2985) );
  XOR U6062 ( .A(n2988), .B(n2989), .Z(n2987) );
  XOR U6063 ( .A(DB[1384]), .B(DB[1377]), .Z(n2989) );
  AND U6064 ( .A(n1262), .B(n2990), .Z(n2988) );
  XOR U6065 ( .A(n2991), .B(n2992), .Z(n2990) );
  XOR U6066 ( .A(DB[1377]), .B(DB[1370]), .Z(n2992) );
  AND U6067 ( .A(n1266), .B(n2993), .Z(n2991) );
  XOR U6068 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR U6069 ( .A(DB[1370]), .B(DB[1363]), .Z(n2995) );
  AND U6070 ( .A(n1270), .B(n2996), .Z(n2994) );
  XOR U6071 ( .A(n2997), .B(n2998), .Z(n2996) );
  XOR U6072 ( .A(DB[1363]), .B(DB[1356]), .Z(n2998) );
  AND U6073 ( .A(n1274), .B(n2999), .Z(n2997) );
  XOR U6074 ( .A(n3000), .B(n3001), .Z(n2999) );
  XOR U6075 ( .A(DB[1356]), .B(DB[1349]), .Z(n3001) );
  AND U6076 ( .A(n1278), .B(n3002), .Z(n3000) );
  XOR U6077 ( .A(n3003), .B(n3004), .Z(n3002) );
  XOR U6078 ( .A(DB[1349]), .B(DB[1342]), .Z(n3004) );
  AND U6079 ( .A(n1282), .B(n3005), .Z(n3003) );
  XOR U6080 ( .A(n3006), .B(n3007), .Z(n3005) );
  XOR U6081 ( .A(DB[1342]), .B(DB[1335]), .Z(n3007) );
  AND U6082 ( .A(n1286), .B(n3008), .Z(n3006) );
  XOR U6083 ( .A(n3009), .B(n3010), .Z(n3008) );
  XOR U6084 ( .A(DB[1335]), .B(DB[1328]), .Z(n3010) );
  AND U6085 ( .A(n1290), .B(n3011), .Z(n3009) );
  XOR U6086 ( .A(n3012), .B(n3013), .Z(n3011) );
  XOR U6087 ( .A(DB[1328]), .B(DB[1321]), .Z(n3013) );
  AND U6088 ( .A(n1294), .B(n3014), .Z(n3012) );
  XOR U6089 ( .A(n3015), .B(n3016), .Z(n3014) );
  XOR U6090 ( .A(DB[1321]), .B(DB[1314]), .Z(n3016) );
  AND U6091 ( .A(n1298), .B(n3017), .Z(n3015) );
  XOR U6092 ( .A(n3018), .B(n3019), .Z(n3017) );
  XOR U6093 ( .A(DB[1314]), .B(DB[1307]), .Z(n3019) );
  AND U6094 ( .A(n1302), .B(n3020), .Z(n3018) );
  XOR U6095 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR U6096 ( .A(DB[1307]), .B(DB[1300]), .Z(n3022) );
  AND U6097 ( .A(n1306), .B(n3023), .Z(n3021) );
  XOR U6098 ( .A(n3024), .B(n3025), .Z(n3023) );
  XOR U6099 ( .A(DB[1300]), .B(DB[1293]), .Z(n3025) );
  AND U6100 ( .A(n1310), .B(n3026), .Z(n3024) );
  XOR U6101 ( .A(n3027), .B(n3028), .Z(n3026) );
  XOR U6102 ( .A(DB[1293]), .B(DB[1286]), .Z(n3028) );
  AND U6103 ( .A(n1314), .B(n3029), .Z(n3027) );
  XOR U6104 ( .A(n3030), .B(n3031), .Z(n3029) );
  XOR U6105 ( .A(DB[1286]), .B(DB[1279]), .Z(n3031) );
  AND U6106 ( .A(n1318), .B(n3032), .Z(n3030) );
  XOR U6107 ( .A(n3033), .B(n3034), .Z(n3032) );
  XOR U6108 ( .A(DB[1279]), .B(DB[1272]), .Z(n3034) );
  AND U6109 ( .A(n1322), .B(n3035), .Z(n3033) );
  XOR U6110 ( .A(n3036), .B(n3037), .Z(n3035) );
  XOR U6111 ( .A(DB[1272]), .B(DB[1265]), .Z(n3037) );
  AND U6112 ( .A(n1326), .B(n3038), .Z(n3036) );
  XOR U6113 ( .A(n3039), .B(n3040), .Z(n3038) );
  XOR U6114 ( .A(DB[1265]), .B(DB[1258]), .Z(n3040) );
  AND U6115 ( .A(n1330), .B(n3041), .Z(n3039) );
  XOR U6116 ( .A(n3042), .B(n3043), .Z(n3041) );
  XOR U6117 ( .A(DB[1258]), .B(DB[1251]), .Z(n3043) );
  AND U6118 ( .A(n1334), .B(n3044), .Z(n3042) );
  XOR U6119 ( .A(n3045), .B(n3046), .Z(n3044) );
  XOR U6120 ( .A(DB[1251]), .B(DB[1244]), .Z(n3046) );
  AND U6121 ( .A(n1338), .B(n3047), .Z(n3045) );
  XOR U6122 ( .A(n3048), .B(n3049), .Z(n3047) );
  XOR U6123 ( .A(DB[1244]), .B(DB[1237]), .Z(n3049) );
  AND U6124 ( .A(n1342), .B(n3050), .Z(n3048) );
  XOR U6125 ( .A(n3051), .B(n3052), .Z(n3050) );
  XOR U6126 ( .A(DB[1237]), .B(DB[1230]), .Z(n3052) );
  AND U6127 ( .A(n1346), .B(n3053), .Z(n3051) );
  XOR U6128 ( .A(n3054), .B(n3055), .Z(n3053) );
  XOR U6129 ( .A(DB[1230]), .B(DB[1223]), .Z(n3055) );
  AND U6130 ( .A(n1350), .B(n3056), .Z(n3054) );
  XOR U6131 ( .A(n3057), .B(n3058), .Z(n3056) );
  XOR U6132 ( .A(DB[1223]), .B(DB[1216]), .Z(n3058) );
  AND U6133 ( .A(n1354), .B(n3059), .Z(n3057) );
  XOR U6134 ( .A(n3060), .B(n3061), .Z(n3059) );
  XOR U6135 ( .A(DB[1216]), .B(DB[1209]), .Z(n3061) );
  AND U6136 ( .A(n1358), .B(n3062), .Z(n3060) );
  XOR U6137 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR U6138 ( .A(DB[1209]), .B(DB[1202]), .Z(n3064) );
  AND U6139 ( .A(n1362), .B(n3065), .Z(n3063) );
  XOR U6140 ( .A(n3066), .B(n3067), .Z(n3065) );
  XOR U6141 ( .A(DB[1202]), .B(DB[1195]), .Z(n3067) );
  AND U6142 ( .A(n1366), .B(n3068), .Z(n3066) );
  XOR U6143 ( .A(n3069), .B(n3070), .Z(n3068) );
  XOR U6144 ( .A(DB[1195]), .B(DB[1188]), .Z(n3070) );
  AND U6145 ( .A(n1370), .B(n3071), .Z(n3069) );
  XOR U6146 ( .A(n3072), .B(n3073), .Z(n3071) );
  XOR U6147 ( .A(DB[1188]), .B(DB[1181]), .Z(n3073) );
  AND U6148 ( .A(n1374), .B(n3074), .Z(n3072) );
  XOR U6149 ( .A(n3075), .B(n3076), .Z(n3074) );
  XOR U6150 ( .A(DB[1181]), .B(DB[1174]), .Z(n3076) );
  AND U6151 ( .A(n1378), .B(n3077), .Z(n3075) );
  XOR U6152 ( .A(n3078), .B(n3079), .Z(n3077) );
  XOR U6153 ( .A(DB[1174]), .B(DB[1167]), .Z(n3079) );
  AND U6154 ( .A(n1382), .B(n3080), .Z(n3078) );
  XOR U6155 ( .A(n3081), .B(n3082), .Z(n3080) );
  XOR U6156 ( .A(DB[1167]), .B(DB[1160]), .Z(n3082) );
  AND U6157 ( .A(n1386), .B(n3083), .Z(n3081) );
  XOR U6158 ( .A(n3084), .B(n3085), .Z(n3083) );
  XOR U6159 ( .A(DB[1160]), .B(DB[1153]), .Z(n3085) );
  AND U6160 ( .A(n1390), .B(n3086), .Z(n3084) );
  XOR U6161 ( .A(n3087), .B(n3088), .Z(n3086) );
  XOR U6162 ( .A(DB[1153]), .B(DB[1146]), .Z(n3088) );
  AND U6163 ( .A(n1394), .B(n3089), .Z(n3087) );
  XOR U6164 ( .A(n3090), .B(n3091), .Z(n3089) );
  XOR U6165 ( .A(DB[1146]), .B(DB[1139]), .Z(n3091) );
  AND U6166 ( .A(n1398), .B(n3092), .Z(n3090) );
  XOR U6167 ( .A(n3093), .B(n3094), .Z(n3092) );
  XOR U6168 ( .A(DB[1139]), .B(DB[1132]), .Z(n3094) );
  AND U6169 ( .A(n1402), .B(n3095), .Z(n3093) );
  XOR U6170 ( .A(n3096), .B(n3097), .Z(n3095) );
  XOR U6171 ( .A(DB[1132]), .B(DB[1125]), .Z(n3097) );
  AND U6172 ( .A(n1406), .B(n3098), .Z(n3096) );
  XOR U6173 ( .A(n3099), .B(n3100), .Z(n3098) );
  XOR U6174 ( .A(DB[1125]), .B(DB[1118]), .Z(n3100) );
  AND U6175 ( .A(n1410), .B(n3101), .Z(n3099) );
  XOR U6176 ( .A(n3102), .B(n3103), .Z(n3101) );
  XOR U6177 ( .A(DB[1118]), .B(DB[1111]), .Z(n3103) );
  AND U6178 ( .A(n1414), .B(n3104), .Z(n3102) );
  XOR U6179 ( .A(n3105), .B(n3106), .Z(n3104) );
  XOR U6180 ( .A(DB[1111]), .B(DB[1104]), .Z(n3106) );
  AND U6181 ( .A(n1418), .B(n3107), .Z(n3105) );
  XOR U6182 ( .A(n3108), .B(n3109), .Z(n3107) );
  XOR U6183 ( .A(DB[1104]), .B(DB[1097]), .Z(n3109) );
  AND U6184 ( .A(n1422), .B(n3110), .Z(n3108) );
  XOR U6185 ( .A(n3111), .B(n3112), .Z(n3110) );
  XOR U6186 ( .A(DB[1097]), .B(DB[1090]), .Z(n3112) );
  AND U6187 ( .A(n1426), .B(n3113), .Z(n3111) );
  XOR U6188 ( .A(n3114), .B(n3115), .Z(n3113) );
  XOR U6189 ( .A(DB[1090]), .B(DB[1083]), .Z(n3115) );
  AND U6190 ( .A(n1430), .B(n3116), .Z(n3114) );
  XOR U6191 ( .A(n3117), .B(n3118), .Z(n3116) );
  XOR U6192 ( .A(DB[1083]), .B(DB[1076]), .Z(n3118) );
  AND U6193 ( .A(n1434), .B(n3119), .Z(n3117) );
  XOR U6194 ( .A(n3120), .B(n3121), .Z(n3119) );
  XOR U6195 ( .A(DB[1076]), .B(DB[1069]), .Z(n3121) );
  AND U6196 ( .A(n1438), .B(n3122), .Z(n3120) );
  XOR U6197 ( .A(n3123), .B(n3124), .Z(n3122) );
  XOR U6198 ( .A(DB[1069]), .B(DB[1062]), .Z(n3124) );
  AND U6199 ( .A(n1442), .B(n3125), .Z(n3123) );
  XOR U6200 ( .A(n3126), .B(n3127), .Z(n3125) );
  XOR U6201 ( .A(DB[1062]), .B(DB[1055]), .Z(n3127) );
  AND U6202 ( .A(n1446), .B(n3128), .Z(n3126) );
  XOR U6203 ( .A(n3129), .B(n3130), .Z(n3128) );
  XOR U6204 ( .A(DB[1055]), .B(DB[1048]), .Z(n3130) );
  AND U6205 ( .A(n1450), .B(n3131), .Z(n3129) );
  XOR U6206 ( .A(n3132), .B(n3133), .Z(n3131) );
  XOR U6207 ( .A(DB[1048]), .B(DB[1041]), .Z(n3133) );
  AND U6208 ( .A(n1454), .B(n3134), .Z(n3132) );
  XOR U6209 ( .A(n3135), .B(n3136), .Z(n3134) );
  XOR U6210 ( .A(DB[1041]), .B(DB[1034]), .Z(n3136) );
  AND U6211 ( .A(n1458), .B(n3137), .Z(n3135) );
  XOR U6212 ( .A(n3138), .B(n3139), .Z(n3137) );
  XOR U6213 ( .A(DB[1034]), .B(DB[1027]), .Z(n3139) );
  AND U6214 ( .A(n1462), .B(n3140), .Z(n3138) );
  XOR U6215 ( .A(n3141), .B(n3142), .Z(n3140) );
  XOR U6216 ( .A(DB[1027]), .B(DB[1020]), .Z(n3142) );
  AND U6217 ( .A(n1466), .B(n3143), .Z(n3141) );
  XOR U6218 ( .A(n3144), .B(n3145), .Z(n3143) );
  XOR U6219 ( .A(DB[1020]), .B(DB[1013]), .Z(n3145) );
  AND U6220 ( .A(n1470), .B(n3146), .Z(n3144) );
  XOR U6221 ( .A(n3147), .B(n3148), .Z(n3146) );
  XOR U6222 ( .A(DB[1013]), .B(DB[1006]), .Z(n3148) );
  AND U6223 ( .A(n1474), .B(n3149), .Z(n3147) );
  XOR U6224 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U6225 ( .A(DB[999]), .B(DB[1006]), .Z(n3151) );
  AND U6226 ( .A(n1478), .B(n3152), .Z(n3150) );
  XOR U6227 ( .A(n3153), .B(n3154), .Z(n3152) );
  XOR U6228 ( .A(DB[999]), .B(DB[992]), .Z(n3154) );
  AND U6229 ( .A(n1482), .B(n3155), .Z(n3153) );
  XOR U6230 ( .A(n3156), .B(n3157), .Z(n3155) );
  XOR U6231 ( .A(DB[992]), .B(DB[985]), .Z(n3157) );
  AND U6232 ( .A(n1486), .B(n3158), .Z(n3156) );
  XOR U6233 ( .A(n3159), .B(n3160), .Z(n3158) );
  XOR U6234 ( .A(DB[985]), .B(DB[978]), .Z(n3160) );
  AND U6235 ( .A(n1490), .B(n3161), .Z(n3159) );
  XOR U6236 ( .A(n3162), .B(n3163), .Z(n3161) );
  XOR U6237 ( .A(DB[978]), .B(DB[971]), .Z(n3163) );
  AND U6238 ( .A(n1494), .B(n3164), .Z(n3162) );
  XOR U6239 ( .A(n3165), .B(n3166), .Z(n3164) );
  XOR U6240 ( .A(DB[971]), .B(DB[964]), .Z(n3166) );
  AND U6241 ( .A(n1498), .B(n3167), .Z(n3165) );
  XOR U6242 ( .A(n3168), .B(n3169), .Z(n3167) );
  XOR U6243 ( .A(DB[964]), .B(DB[957]), .Z(n3169) );
  AND U6244 ( .A(n1502), .B(n3170), .Z(n3168) );
  XOR U6245 ( .A(n3171), .B(n3172), .Z(n3170) );
  XOR U6246 ( .A(DB[957]), .B(DB[950]), .Z(n3172) );
  AND U6247 ( .A(n1506), .B(n3173), .Z(n3171) );
  XOR U6248 ( .A(n3174), .B(n3175), .Z(n3173) );
  XOR U6249 ( .A(DB[950]), .B(DB[943]), .Z(n3175) );
  AND U6250 ( .A(n1510), .B(n3176), .Z(n3174) );
  XOR U6251 ( .A(n3177), .B(n3178), .Z(n3176) );
  XOR U6252 ( .A(DB[943]), .B(DB[936]), .Z(n3178) );
  AND U6253 ( .A(n1514), .B(n3179), .Z(n3177) );
  XOR U6254 ( .A(n3180), .B(n3181), .Z(n3179) );
  XOR U6255 ( .A(DB[936]), .B(DB[929]), .Z(n3181) );
  AND U6256 ( .A(n1518), .B(n3182), .Z(n3180) );
  XOR U6257 ( .A(n3183), .B(n3184), .Z(n3182) );
  XOR U6258 ( .A(DB[929]), .B(DB[922]), .Z(n3184) );
  AND U6259 ( .A(n1522), .B(n3185), .Z(n3183) );
  XOR U6260 ( .A(n3186), .B(n3187), .Z(n3185) );
  XOR U6261 ( .A(DB[922]), .B(DB[915]), .Z(n3187) );
  AND U6262 ( .A(n1526), .B(n3188), .Z(n3186) );
  XOR U6263 ( .A(n3189), .B(n3190), .Z(n3188) );
  XOR U6264 ( .A(DB[915]), .B(DB[908]), .Z(n3190) );
  AND U6265 ( .A(n1530), .B(n3191), .Z(n3189) );
  XOR U6266 ( .A(n3192), .B(n3193), .Z(n3191) );
  XOR U6267 ( .A(DB[908]), .B(DB[901]), .Z(n3193) );
  AND U6268 ( .A(n1534), .B(n3194), .Z(n3192) );
  XOR U6269 ( .A(n3195), .B(n3196), .Z(n3194) );
  XOR U6270 ( .A(DB[901]), .B(DB[894]), .Z(n3196) );
  AND U6271 ( .A(n1538), .B(n3197), .Z(n3195) );
  XOR U6272 ( .A(n3198), .B(n3199), .Z(n3197) );
  XOR U6273 ( .A(DB[894]), .B(DB[887]), .Z(n3199) );
  AND U6274 ( .A(n1542), .B(n3200), .Z(n3198) );
  XOR U6275 ( .A(n3201), .B(n3202), .Z(n3200) );
  XOR U6276 ( .A(DB[887]), .B(DB[880]), .Z(n3202) );
  AND U6277 ( .A(n1546), .B(n3203), .Z(n3201) );
  XOR U6278 ( .A(n3204), .B(n3205), .Z(n3203) );
  XOR U6279 ( .A(DB[880]), .B(DB[873]), .Z(n3205) );
  AND U6280 ( .A(n1550), .B(n3206), .Z(n3204) );
  XOR U6281 ( .A(n3207), .B(n3208), .Z(n3206) );
  XOR U6282 ( .A(DB[873]), .B(DB[866]), .Z(n3208) );
  AND U6283 ( .A(n1554), .B(n3209), .Z(n3207) );
  XOR U6284 ( .A(n3210), .B(n3211), .Z(n3209) );
  XOR U6285 ( .A(DB[866]), .B(DB[859]), .Z(n3211) );
  AND U6286 ( .A(n1558), .B(n3212), .Z(n3210) );
  XOR U6287 ( .A(n3213), .B(n3214), .Z(n3212) );
  XOR U6288 ( .A(DB[859]), .B(DB[852]), .Z(n3214) );
  AND U6289 ( .A(n1562), .B(n3215), .Z(n3213) );
  XOR U6290 ( .A(n3216), .B(n3217), .Z(n3215) );
  XOR U6291 ( .A(DB[852]), .B(DB[845]), .Z(n3217) );
  AND U6292 ( .A(n1566), .B(n3218), .Z(n3216) );
  XOR U6293 ( .A(n3219), .B(n3220), .Z(n3218) );
  XOR U6294 ( .A(DB[845]), .B(DB[838]), .Z(n3220) );
  AND U6295 ( .A(n1570), .B(n3221), .Z(n3219) );
  XOR U6296 ( .A(n3222), .B(n3223), .Z(n3221) );
  XOR U6297 ( .A(DB[838]), .B(DB[831]), .Z(n3223) );
  AND U6298 ( .A(n1574), .B(n3224), .Z(n3222) );
  XOR U6299 ( .A(n3225), .B(n3226), .Z(n3224) );
  XOR U6300 ( .A(DB[831]), .B(DB[824]), .Z(n3226) );
  AND U6301 ( .A(n1578), .B(n3227), .Z(n3225) );
  XOR U6302 ( .A(n3228), .B(n3229), .Z(n3227) );
  XOR U6303 ( .A(DB[824]), .B(DB[817]), .Z(n3229) );
  AND U6304 ( .A(n1582), .B(n3230), .Z(n3228) );
  XOR U6305 ( .A(n3231), .B(n3232), .Z(n3230) );
  XOR U6306 ( .A(DB[817]), .B(DB[810]), .Z(n3232) );
  AND U6307 ( .A(n1586), .B(n3233), .Z(n3231) );
  XOR U6308 ( .A(n3234), .B(n3235), .Z(n3233) );
  XOR U6309 ( .A(DB[810]), .B(DB[803]), .Z(n3235) );
  AND U6310 ( .A(n1590), .B(n3236), .Z(n3234) );
  XOR U6311 ( .A(n3237), .B(n3238), .Z(n3236) );
  XOR U6312 ( .A(DB[803]), .B(DB[796]), .Z(n3238) );
  AND U6313 ( .A(n1594), .B(n3239), .Z(n3237) );
  XOR U6314 ( .A(n3240), .B(n3241), .Z(n3239) );
  XOR U6315 ( .A(DB[796]), .B(DB[789]), .Z(n3241) );
  AND U6316 ( .A(n1598), .B(n3242), .Z(n3240) );
  XOR U6317 ( .A(n3243), .B(n3244), .Z(n3242) );
  XOR U6318 ( .A(DB[789]), .B(DB[782]), .Z(n3244) );
  AND U6319 ( .A(n1602), .B(n3245), .Z(n3243) );
  XOR U6320 ( .A(n3246), .B(n3247), .Z(n3245) );
  XOR U6321 ( .A(DB[782]), .B(DB[775]), .Z(n3247) );
  AND U6322 ( .A(n1606), .B(n3248), .Z(n3246) );
  XOR U6323 ( .A(n3249), .B(n3250), .Z(n3248) );
  XOR U6324 ( .A(DB[775]), .B(DB[768]), .Z(n3250) );
  AND U6325 ( .A(n1610), .B(n3251), .Z(n3249) );
  XOR U6326 ( .A(n3252), .B(n3253), .Z(n3251) );
  XOR U6327 ( .A(DB[768]), .B(DB[761]), .Z(n3253) );
  AND U6328 ( .A(n1614), .B(n3254), .Z(n3252) );
  XOR U6329 ( .A(n3255), .B(n3256), .Z(n3254) );
  XOR U6330 ( .A(DB[761]), .B(DB[754]), .Z(n3256) );
  AND U6331 ( .A(n1618), .B(n3257), .Z(n3255) );
  XOR U6332 ( .A(n3258), .B(n3259), .Z(n3257) );
  XOR U6333 ( .A(DB[754]), .B(DB[747]), .Z(n3259) );
  AND U6334 ( .A(n1622), .B(n3260), .Z(n3258) );
  XOR U6335 ( .A(n3261), .B(n3262), .Z(n3260) );
  XOR U6336 ( .A(DB[747]), .B(DB[740]), .Z(n3262) );
  AND U6337 ( .A(n1626), .B(n3263), .Z(n3261) );
  XOR U6338 ( .A(n3264), .B(n3265), .Z(n3263) );
  XOR U6339 ( .A(DB[740]), .B(DB[733]), .Z(n3265) );
  AND U6340 ( .A(n1630), .B(n3266), .Z(n3264) );
  XOR U6341 ( .A(n3267), .B(n3268), .Z(n3266) );
  XOR U6342 ( .A(DB[733]), .B(DB[726]), .Z(n3268) );
  AND U6343 ( .A(n1634), .B(n3269), .Z(n3267) );
  XOR U6344 ( .A(n3270), .B(n3271), .Z(n3269) );
  XOR U6345 ( .A(DB[726]), .B(DB[719]), .Z(n3271) );
  AND U6346 ( .A(n1638), .B(n3272), .Z(n3270) );
  XOR U6347 ( .A(n3273), .B(n3274), .Z(n3272) );
  XOR U6348 ( .A(DB[719]), .B(DB[712]), .Z(n3274) );
  AND U6349 ( .A(n1642), .B(n3275), .Z(n3273) );
  XOR U6350 ( .A(n3276), .B(n3277), .Z(n3275) );
  XOR U6351 ( .A(DB[712]), .B(DB[705]), .Z(n3277) );
  AND U6352 ( .A(n1646), .B(n3278), .Z(n3276) );
  XOR U6353 ( .A(n3279), .B(n3280), .Z(n3278) );
  XOR U6354 ( .A(DB[705]), .B(DB[698]), .Z(n3280) );
  AND U6355 ( .A(n1650), .B(n3281), .Z(n3279) );
  XOR U6356 ( .A(n3282), .B(n3283), .Z(n3281) );
  XOR U6357 ( .A(DB[698]), .B(DB[691]), .Z(n3283) );
  AND U6358 ( .A(n1654), .B(n3284), .Z(n3282) );
  XOR U6359 ( .A(n3285), .B(n3286), .Z(n3284) );
  XOR U6360 ( .A(DB[691]), .B(DB[684]), .Z(n3286) );
  AND U6361 ( .A(n1658), .B(n3287), .Z(n3285) );
  XOR U6362 ( .A(n3288), .B(n3289), .Z(n3287) );
  XOR U6363 ( .A(DB[684]), .B(DB[677]), .Z(n3289) );
  AND U6364 ( .A(n1662), .B(n3290), .Z(n3288) );
  XOR U6365 ( .A(n3291), .B(n3292), .Z(n3290) );
  XOR U6366 ( .A(DB[677]), .B(DB[670]), .Z(n3292) );
  AND U6367 ( .A(n1666), .B(n3293), .Z(n3291) );
  XOR U6368 ( .A(n3294), .B(n3295), .Z(n3293) );
  XOR U6369 ( .A(DB[670]), .B(DB[663]), .Z(n3295) );
  AND U6370 ( .A(n1670), .B(n3296), .Z(n3294) );
  XOR U6371 ( .A(n3297), .B(n3298), .Z(n3296) );
  XOR U6372 ( .A(DB[663]), .B(DB[656]), .Z(n3298) );
  AND U6373 ( .A(n1674), .B(n3299), .Z(n3297) );
  XOR U6374 ( .A(n3300), .B(n3301), .Z(n3299) );
  XOR U6375 ( .A(DB[656]), .B(DB[649]), .Z(n3301) );
  AND U6376 ( .A(n1678), .B(n3302), .Z(n3300) );
  XOR U6377 ( .A(n3303), .B(n3304), .Z(n3302) );
  XOR U6378 ( .A(DB[649]), .B(DB[642]), .Z(n3304) );
  AND U6379 ( .A(n1682), .B(n3305), .Z(n3303) );
  XOR U6380 ( .A(n3306), .B(n3307), .Z(n3305) );
  XOR U6381 ( .A(DB[642]), .B(DB[635]), .Z(n3307) );
  AND U6382 ( .A(n1686), .B(n3308), .Z(n3306) );
  XOR U6383 ( .A(n3309), .B(n3310), .Z(n3308) );
  XOR U6384 ( .A(DB[635]), .B(DB[628]), .Z(n3310) );
  AND U6385 ( .A(n1690), .B(n3311), .Z(n3309) );
  XOR U6386 ( .A(n3312), .B(n3313), .Z(n3311) );
  XOR U6387 ( .A(DB[628]), .B(DB[621]), .Z(n3313) );
  AND U6388 ( .A(n1694), .B(n3314), .Z(n3312) );
  XOR U6389 ( .A(n3315), .B(n3316), .Z(n3314) );
  XOR U6390 ( .A(DB[621]), .B(DB[614]), .Z(n3316) );
  AND U6391 ( .A(n1698), .B(n3317), .Z(n3315) );
  XOR U6392 ( .A(n3318), .B(n3319), .Z(n3317) );
  XOR U6393 ( .A(DB[614]), .B(DB[607]), .Z(n3319) );
  AND U6394 ( .A(n1702), .B(n3320), .Z(n3318) );
  XOR U6395 ( .A(n3321), .B(n3322), .Z(n3320) );
  XOR U6396 ( .A(DB[607]), .B(DB[600]), .Z(n3322) );
  AND U6397 ( .A(n1706), .B(n3323), .Z(n3321) );
  XOR U6398 ( .A(n3324), .B(n3325), .Z(n3323) );
  XOR U6399 ( .A(DB[600]), .B(DB[593]), .Z(n3325) );
  AND U6400 ( .A(n1710), .B(n3326), .Z(n3324) );
  XOR U6401 ( .A(n3327), .B(n3328), .Z(n3326) );
  XOR U6402 ( .A(DB[593]), .B(DB[586]), .Z(n3328) );
  AND U6403 ( .A(n1714), .B(n3329), .Z(n3327) );
  XOR U6404 ( .A(n3330), .B(n3331), .Z(n3329) );
  XOR U6405 ( .A(DB[586]), .B(DB[579]), .Z(n3331) );
  AND U6406 ( .A(n1718), .B(n3332), .Z(n3330) );
  XOR U6407 ( .A(n3333), .B(n3334), .Z(n3332) );
  XOR U6408 ( .A(DB[579]), .B(DB[572]), .Z(n3334) );
  AND U6409 ( .A(n1722), .B(n3335), .Z(n3333) );
  XOR U6410 ( .A(n3336), .B(n3337), .Z(n3335) );
  XOR U6411 ( .A(DB[572]), .B(DB[565]), .Z(n3337) );
  AND U6412 ( .A(n1726), .B(n3338), .Z(n3336) );
  XOR U6413 ( .A(n3339), .B(n3340), .Z(n3338) );
  XOR U6414 ( .A(DB[565]), .B(DB[558]), .Z(n3340) );
  AND U6415 ( .A(n1730), .B(n3341), .Z(n3339) );
  XOR U6416 ( .A(n3342), .B(n3343), .Z(n3341) );
  XOR U6417 ( .A(DB[558]), .B(DB[551]), .Z(n3343) );
  AND U6418 ( .A(n1734), .B(n3344), .Z(n3342) );
  XOR U6419 ( .A(n3345), .B(n3346), .Z(n3344) );
  XOR U6420 ( .A(DB[551]), .B(DB[544]), .Z(n3346) );
  AND U6421 ( .A(n1738), .B(n3347), .Z(n3345) );
  XOR U6422 ( .A(n3348), .B(n3349), .Z(n3347) );
  XOR U6423 ( .A(DB[544]), .B(DB[537]), .Z(n3349) );
  AND U6424 ( .A(n1742), .B(n3350), .Z(n3348) );
  XOR U6425 ( .A(n3351), .B(n3352), .Z(n3350) );
  XOR U6426 ( .A(DB[537]), .B(DB[530]), .Z(n3352) );
  AND U6427 ( .A(n1746), .B(n3353), .Z(n3351) );
  XOR U6428 ( .A(n3354), .B(n3355), .Z(n3353) );
  XOR U6429 ( .A(DB[530]), .B(DB[523]), .Z(n3355) );
  AND U6430 ( .A(n1750), .B(n3356), .Z(n3354) );
  XOR U6431 ( .A(n3357), .B(n3358), .Z(n3356) );
  XOR U6432 ( .A(DB[523]), .B(DB[516]), .Z(n3358) );
  AND U6433 ( .A(n1754), .B(n3359), .Z(n3357) );
  XOR U6434 ( .A(n3360), .B(n3361), .Z(n3359) );
  XOR U6435 ( .A(DB[516]), .B(DB[509]), .Z(n3361) );
  AND U6436 ( .A(n1758), .B(n3362), .Z(n3360) );
  XOR U6437 ( .A(n3363), .B(n3364), .Z(n3362) );
  XOR U6438 ( .A(DB[509]), .B(DB[502]), .Z(n3364) );
  AND U6439 ( .A(n1762), .B(n3365), .Z(n3363) );
  XOR U6440 ( .A(n3366), .B(n3367), .Z(n3365) );
  XOR U6441 ( .A(DB[502]), .B(DB[495]), .Z(n3367) );
  AND U6442 ( .A(n1766), .B(n3368), .Z(n3366) );
  XOR U6443 ( .A(n3369), .B(n3370), .Z(n3368) );
  XOR U6444 ( .A(DB[495]), .B(DB[488]), .Z(n3370) );
  AND U6445 ( .A(n1770), .B(n3371), .Z(n3369) );
  XOR U6446 ( .A(n3372), .B(n3373), .Z(n3371) );
  XOR U6447 ( .A(DB[488]), .B(DB[481]), .Z(n3373) );
  AND U6448 ( .A(n1774), .B(n3374), .Z(n3372) );
  XOR U6449 ( .A(n3375), .B(n3376), .Z(n3374) );
  XOR U6450 ( .A(DB[481]), .B(DB[474]), .Z(n3376) );
  AND U6451 ( .A(n1778), .B(n3377), .Z(n3375) );
  XOR U6452 ( .A(n3378), .B(n3379), .Z(n3377) );
  XOR U6453 ( .A(DB[474]), .B(DB[467]), .Z(n3379) );
  AND U6454 ( .A(n1782), .B(n3380), .Z(n3378) );
  XOR U6455 ( .A(n3381), .B(n3382), .Z(n3380) );
  XOR U6456 ( .A(DB[467]), .B(DB[460]), .Z(n3382) );
  AND U6457 ( .A(n1786), .B(n3383), .Z(n3381) );
  XOR U6458 ( .A(n3384), .B(n3385), .Z(n3383) );
  XOR U6459 ( .A(DB[460]), .B(DB[453]), .Z(n3385) );
  AND U6460 ( .A(n1790), .B(n3386), .Z(n3384) );
  XOR U6461 ( .A(n3387), .B(n3388), .Z(n3386) );
  XOR U6462 ( .A(DB[453]), .B(DB[446]), .Z(n3388) );
  AND U6463 ( .A(n1794), .B(n3389), .Z(n3387) );
  XOR U6464 ( .A(n3390), .B(n3391), .Z(n3389) );
  XOR U6465 ( .A(DB[446]), .B(DB[439]), .Z(n3391) );
  AND U6466 ( .A(n1798), .B(n3392), .Z(n3390) );
  XOR U6467 ( .A(n3393), .B(n3394), .Z(n3392) );
  XOR U6468 ( .A(DB[439]), .B(DB[432]), .Z(n3394) );
  AND U6469 ( .A(n1802), .B(n3395), .Z(n3393) );
  XOR U6470 ( .A(n3396), .B(n3397), .Z(n3395) );
  XOR U6471 ( .A(DB[432]), .B(DB[425]), .Z(n3397) );
  AND U6472 ( .A(n1806), .B(n3398), .Z(n3396) );
  XOR U6473 ( .A(n3399), .B(n3400), .Z(n3398) );
  XOR U6474 ( .A(DB[425]), .B(DB[418]), .Z(n3400) );
  AND U6475 ( .A(n1810), .B(n3401), .Z(n3399) );
  XOR U6476 ( .A(n3402), .B(n3403), .Z(n3401) );
  XOR U6477 ( .A(DB[418]), .B(DB[411]), .Z(n3403) );
  AND U6478 ( .A(n1814), .B(n3404), .Z(n3402) );
  XOR U6479 ( .A(n3405), .B(n3406), .Z(n3404) );
  XOR U6480 ( .A(DB[411]), .B(DB[404]), .Z(n3406) );
  AND U6481 ( .A(n1818), .B(n3407), .Z(n3405) );
  XOR U6482 ( .A(n3408), .B(n3409), .Z(n3407) );
  XOR U6483 ( .A(DB[404]), .B(DB[397]), .Z(n3409) );
  AND U6484 ( .A(n1822), .B(n3410), .Z(n3408) );
  XOR U6485 ( .A(n3411), .B(n3412), .Z(n3410) );
  XOR U6486 ( .A(DB[397]), .B(DB[390]), .Z(n3412) );
  AND U6487 ( .A(n1826), .B(n3413), .Z(n3411) );
  XOR U6488 ( .A(n3414), .B(n3415), .Z(n3413) );
  XOR U6489 ( .A(DB[390]), .B(DB[383]), .Z(n3415) );
  AND U6490 ( .A(n1830), .B(n3416), .Z(n3414) );
  XOR U6491 ( .A(n3417), .B(n3418), .Z(n3416) );
  XOR U6492 ( .A(DB[383]), .B(DB[376]), .Z(n3418) );
  AND U6493 ( .A(n1834), .B(n3419), .Z(n3417) );
  XOR U6494 ( .A(n3420), .B(n3421), .Z(n3419) );
  XOR U6495 ( .A(DB[376]), .B(DB[369]), .Z(n3421) );
  AND U6496 ( .A(n1838), .B(n3422), .Z(n3420) );
  XOR U6497 ( .A(n3423), .B(n3424), .Z(n3422) );
  XOR U6498 ( .A(DB[369]), .B(DB[362]), .Z(n3424) );
  AND U6499 ( .A(n1842), .B(n3425), .Z(n3423) );
  XOR U6500 ( .A(n3426), .B(n3427), .Z(n3425) );
  XOR U6501 ( .A(DB[362]), .B(DB[355]), .Z(n3427) );
  AND U6502 ( .A(n1846), .B(n3428), .Z(n3426) );
  XOR U6503 ( .A(n3429), .B(n3430), .Z(n3428) );
  XOR U6504 ( .A(DB[355]), .B(DB[348]), .Z(n3430) );
  AND U6505 ( .A(n1850), .B(n3431), .Z(n3429) );
  XOR U6506 ( .A(n3432), .B(n3433), .Z(n3431) );
  XOR U6507 ( .A(DB[348]), .B(DB[341]), .Z(n3433) );
  AND U6508 ( .A(n1854), .B(n3434), .Z(n3432) );
  XOR U6509 ( .A(n3435), .B(n3436), .Z(n3434) );
  XOR U6510 ( .A(DB[341]), .B(DB[334]), .Z(n3436) );
  AND U6511 ( .A(n1858), .B(n3437), .Z(n3435) );
  XOR U6512 ( .A(n3438), .B(n3439), .Z(n3437) );
  XOR U6513 ( .A(DB[334]), .B(DB[327]), .Z(n3439) );
  AND U6514 ( .A(n1862), .B(n3440), .Z(n3438) );
  XOR U6515 ( .A(n3441), .B(n3442), .Z(n3440) );
  XOR U6516 ( .A(DB[327]), .B(DB[320]), .Z(n3442) );
  AND U6517 ( .A(n1866), .B(n3443), .Z(n3441) );
  XOR U6518 ( .A(n3444), .B(n3445), .Z(n3443) );
  XOR U6519 ( .A(DB[320]), .B(DB[313]), .Z(n3445) );
  AND U6520 ( .A(n1870), .B(n3446), .Z(n3444) );
  XOR U6521 ( .A(n3447), .B(n3448), .Z(n3446) );
  XOR U6522 ( .A(DB[313]), .B(DB[306]), .Z(n3448) );
  AND U6523 ( .A(n1874), .B(n3449), .Z(n3447) );
  XOR U6524 ( .A(n3450), .B(n3451), .Z(n3449) );
  XOR U6525 ( .A(DB[306]), .B(DB[299]), .Z(n3451) );
  AND U6526 ( .A(n1878), .B(n3452), .Z(n3450) );
  XOR U6527 ( .A(n3453), .B(n3454), .Z(n3452) );
  XOR U6528 ( .A(DB[299]), .B(DB[292]), .Z(n3454) );
  AND U6529 ( .A(n1882), .B(n3455), .Z(n3453) );
  XOR U6530 ( .A(n3456), .B(n3457), .Z(n3455) );
  XOR U6531 ( .A(DB[292]), .B(DB[285]), .Z(n3457) );
  AND U6532 ( .A(n1886), .B(n3458), .Z(n3456) );
  XOR U6533 ( .A(n3459), .B(n3460), .Z(n3458) );
  XOR U6534 ( .A(DB[285]), .B(DB[278]), .Z(n3460) );
  AND U6535 ( .A(n1890), .B(n3461), .Z(n3459) );
  XOR U6536 ( .A(n3462), .B(n3463), .Z(n3461) );
  XOR U6537 ( .A(DB[278]), .B(DB[271]), .Z(n3463) );
  AND U6538 ( .A(n1894), .B(n3464), .Z(n3462) );
  XOR U6539 ( .A(n3465), .B(n3466), .Z(n3464) );
  XOR U6540 ( .A(DB[271]), .B(DB[264]), .Z(n3466) );
  AND U6541 ( .A(n1898), .B(n3467), .Z(n3465) );
  XOR U6542 ( .A(n3468), .B(n3469), .Z(n3467) );
  XOR U6543 ( .A(DB[264]), .B(DB[257]), .Z(n3469) );
  AND U6544 ( .A(n1902), .B(n3470), .Z(n3468) );
  XOR U6545 ( .A(n3471), .B(n3472), .Z(n3470) );
  XOR U6546 ( .A(DB[257]), .B(DB[250]), .Z(n3472) );
  AND U6547 ( .A(n1906), .B(n3473), .Z(n3471) );
  XOR U6548 ( .A(n3474), .B(n3475), .Z(n3473) );
  XOR U6549 ( .A(DB[250]), .B(DB[243]), .Z(n3475) );
  AND U6550 ( .A(n1910), .B(n3476), .Z(n3474) );
  XOR U6551 ( .A(n3477), .B(n3478), .Z(n3476) );
  XOR U6552 ( .A(DB[243]), .B(DB[236]), .Z(n3478) );
  AND U6553 ( .A(n1914), .B(n3479), .Z(n3477) );
  XOR U6554 ( .A(n3480), .B(n3481), .Z(n3479) );
  XOR U6555 ( .A(DB[236]), .B(DB[229]), .Z(n3481) );
  AND U6556 ( .A(n1918), .B(n3482), .Z(n3480) );
  XOR U6557 ( .A(n3483), .B(n3484), .Z(n3482) );
  XOR U6558 ( .A(DB[229]), .B(DB[222]), .Z(n3484) );
  AND U6559 ( .A(n1922), .B(n3485), .Z(n3483) );
  XOR U6560 ( .A(n3486), .B(n3487), .Z(n3485) );
  XOR U6561 ( .A(DB[222]), .B(DB[215]), .Z(n3487) );
  AND U6562 ( .A(n1926), .B(n3488), .Z(n3486) );
  XOR U6563 ( .A(n3489), .B(n3490), .Z(n3488) );
  XOR U6564 ( .A(DB[215]), .B(DB[208]), .Z(n3490) );
  AND U6565 ( .A(n1930), .B(n3491), .Z(n3489) );
  XOR U6566 ( .A(n3492), .B(n3493), .Z(n3491) );
  XOR U6567 ( .A(DB[208]), .B(DB[201]), .Z(n3493) );
  AND U6568 ( .A(n1934), .B(n3494), .Z(n3492) );
  XOR U6569 ( .A(n3495), .B(n3496), .Z(n3494) );
  XOR U6570 ( .A(DB[201]), .B(DB[194]), .Z(n3496) );
  AND U6571 ( .A(n1938), .B(n3497), .Z(n3495) );
  XOR U6572 ( .A(n3498), .B(n3499), .Z(n3497) );
  XOR U6573 ( .A(DB[194]), .B(DB[187]), .Z(n3499) );
  AND U6574 ( .A(n1942), .B(n3500), .Z(n3498) );
  XOR U6575 ( .A(n3501), .B(n3502), .Z(n3500) );
  XOR U6576 ( .A(DB[187]), .B(DB[180]), .Z(n3502) );
  AND U6577 ( .A(n1946), .B(n3503), .Z(n3501) );
  XOR U6578 ( .A(n3504), .B(n3505), .Z(n3503) );
  XOR U6579 ( .A(DB[180]), .B(DB[173]), .Z(n3505) );
  AND U6580 ( .A(n1950), .B(n3506), .Z(n3504) );
  XOR U6581 ( .A(n3507), .B(n3508), .Z(n3506) );
  XOR U6582 ( .A(DB[173]), .B(DB[166]), .Z(n3508) );
  AND U6583 ( .A(n1954), .B(n3509), .Z(n3507) );
  XOR U6584 ( .A(n3510), .B(n3511), .Z(n3509) );
  XOR U6585 ( .A(DB[166]), .B(DB[159]), .Z(n3511) );
  AND U6586 ( .A(n1958), .B(n3512), .Z(n3510) );
  XOR U6587 ( .A(n3513), .B(n3514), .Z(n3512) );
  XOR U6588 ( .A(DB[159]), .B(DB[152]), .Z(n3514) );
  AND U6589 ( .A(n1962), .B(n3515), .Z(n3513) );
  XOR U6590 ( .A(n3516), .B(n3517), .Z(n3515) );
  XOR U6591 ( .A(DB[152]), .B(DB[145]), .Z(n3517) );
  AND U6592 ( .A(n1966), .B(n3518), .Z(n3516) );
  XOR U6593 ( .A(n3519), .B(n3520), .Z(n3518) );
  XOR U6594 ( .A(DB[145]), .B(DB[138]), .Z(n3520) );
  AND U6595 ( .A(n1970), .B(n3521), .Z(n3519) );
  XOR U6596 ( .A(n3522), .B(n3523), .Z(n3521) );
  XOR U6597 ( .A(DB[138]), .B(DB[131]), .Z(n3523) );
  AND U6598 ( .A(n1974), .B(n3524), .Z(n3522) );
  XOR U6599 ( .A(n3525), .B(n3526), .Z(n3524) );
  XOR U6600 ( .A(DB[131]), .B(DB[124]), .Z(n3526) );
  AND U6601 ( .A(n1978), .B(n3527), .Z(n3525) );
  XOR U6602 ( .A(n3528), .B(n3529), .Z(n3527) );
  XOR U6603 ( .A(DB[124]), .B(DB[117]), .Z(n3529) );
  AND U6604 ( .A(n1982), .B(n3530), .Z(n3528) );
  XOR U6605 ( .A(n3531), .B(n3532), .Z(n3530) );
  XOR U6606 ( .A(DB[117]), .B(DB[110]), .Z(n3532) );
  AND U6607 ( .A(n1986), .B(n3533), .Z(n3531) );
  XOR U6608 ( .A(n3534), .B(n3535), .Z(n3533) );
  XOR U6609 ( .A(DB[110]), .B(DB[103]), .Z(n3535) );
  AND U6610 ( .A(n1990), .B(n3536), .Z(n3534) );
  XOR U6611 ( .A(n3537), .B(n3538), .Z(n3536) );
  XOR U6612 ( .A(DB[96]), .B(DB[103]), .Z(n3538) );
  AND U6613 ( .A(n1994), .B(n3539), .Z(n3537) );
  XOR U6614 ( .A(n3540), .B(n3541), .Z(n3539) );
  XOR U6615 ( .A(DB[96]), .B(DB[89]), .Z(n3541) );
  AND U6616 ( .A(n1998), .B(n3542), .Z(n3540) );
  XOR U6617 ( .A(n3543), .B(n3544), .Z(n3542) );
  XOR U6618 ( .A(DB[89]), .B(DB[82]), .Z(n3544) );
  AND U6619 ( .A(n2002), .B(n3545), .Z(n3543) );
  XOR U6620 ( .A(n3546), .B(n3547), .Z(n3545) );
  XOR U6621 ( .A(DB[82]), .B(DB[75]), .Z(n3547) );
  AND U6622 ( .A(n2006), .B(n3548), .Z(n3546) );
  XOR U6623 ( .A(n3549), .B(n3550), .Z(n3548) );
  XOR U6624 ( .A(DB[75]), .B(DB[68]), .Z(n3550) );
  AND U6625 ( .A(n2010), .B(n3551), .Z(n3549) );
  XOR U6626 ( .A(n3552), .B(n3553), .Z(n3551) );
  XOR U6627 ( .A(DB[68]), .B(DB[61]), .Z(n3553) );
  AND U6628 ( .A(n2014), .B(n3554), .Z(n3552) );
  XOR U6629 ( .A(n3555), .B(n3556), .Z(n3554) );
  XOR U6630 ( .A(DB[61]), .B(DB[54]), .Z(n3556) );
  AND U6631 ( .A(n2018), .B(n3557), .Z(n3555) );
  XOR U6632 ( .A(n3558), .B(n3559), .Z(n3557) );
  XOR U6633 ( .A(DB[54]), .B(DB[47]), .Z(n3559) );
  AND U6634 ( .A(n2022), .B(n3560), .Z(n3558) );
  XOR U6635 ( .A(n3561), .B(n3562), .Z(n3560) );
  XOR U6636 ( .A(DB[47]), .B(DB[40]), .Z(n3562) );
  AND U6637 ( .A(n2026), .B(n3563), .Z(n3561) );
  XOR U6638 ( .A(n3564), .B(n3565), .Z(n3563) );
  XOR U6639 ( .A(DB[40]), .B(DB[33]), .Z(n3565) );
  AND U6640 ( .A(n2030), .B(n3566), .Z(n3564) );
  XOR U6641 ( .A(n3567), .B(n3568), .Z(n3566) );
  XOR U6642 ( .A(DB[33]), .B(DB[26]), .Z(n3568) );
  AND U6643 ( .A(n2034), .B(n3569), .Z(n3567) );
  XOR U6644 ( .A(n3570), .B(n3571), .Z(n3569) );
  XOR U6645 ( .A(DB[26]), .B(DB[19]), .Z(n3571) );
  AND U6646 ( .A(n2038), .B(n3572), .Z(n3570) );
  XOR U6647 ( .A(n3573), .B(n3574), .Z(n3572) );
  XOR U6648 ( .A(DB[19]), .B(DB[12]), .Z(n3574) );
  AND U6649 ( .A(n2042), .B(n3575), .Z(n3573) );
  XOR U6650 ( .A(DB[5]), .B(DB[12]), .Z(n3575) );
  XOR U6651 ( .A(DB[3581]), .B(n3576), .Z(min_val_out[4]) );
  AND U6652 ( .A(n2), .B(n3577), .Z(n3576) );
  XOR U6653 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR U6654 ( .A(DB[3581]), .B(DB[3574]), .Z(n3579) );
  AND U6655 ( .A(n6), .B(n3580), .Z(n3578) );
  XOR U6656 ( .A(n3581), .B(n3582), .Z(n3580) );
  XOR U6657 ( .A(DB[3574]), .B(DB[3567]), .Z(n3582) );
  AND U6658 ( .A(n10), .B(n3583), .Z(n3581) );
  XOR U6659 ( .A(n3584), .B(n3585), .Z(n3583) );
  XOR U6660 ( .A(DB[3567]), .B(DB[3560]), .Z(n3585) );
  AND U6661 ( .A(n14), .B(n3586), .Z(n3584) );
  XOR U6662 ( .A(n3587), .B(n3588), .Z(n3586) );
  XOR U6663 ( .A(DB[3560]), .B(DB[3553]), .Z(n3588) );
  AND U6664 ( .A(n18), .B(n3589), .Z(n3587) );
  XOR U6665 ( .A(n3590), .B(n3591), .Z(n3589) );
  XOR U6666 ( .A(DB[3553]), .B(DB[3546]), .Z(n3591) );
  AND U6667 ( .A(n22), .B(n3592), .Z(n3590) );
  XOR U6668 ( .A(n3593), .B(n3594), .Z(n3592) );
  XOR U6669 ( .A(DB[3546]), .B(DB[3539]), .Z(n3594) );
  AND U6670 ( .A(n26), .B(n3595), .Z(n3593) );
  XOR U6671 ( .A(n3596), .B(n3597), .Z(n3595) );
  XOR U6672 ( .A(DB[3539]), .B(DB[3532]), .Z(n3597) );
  AND U6673 ( .A(n30), .B(n3598), .Z(n3596) );
  XOR U6674 ( .A(n3599), .B(n3600), .Z(n3598) );
  XOR U6675 ( .A(DB[3532]), .B(DB[3525]), .Z(n3600) );
  AND U6676 ( .A(n34), .B(n3601), .Z(n3599) );
  XOR U6677 ( .A(n3602), .B(n3603), .Z(n3601) );
  XOR U6678 ( .A(DB[3525]), .B(DB[3518]), .Z(n3603) );
  AND U6679 ( .A(n38), .B(n3604), .Z(n3602) );
  XOR U6680 ( .A(n3605), .B(n3606), .Z(n3604) );
  XOR U6681 ( .A(DB[3518]), .B(DB[3511]), .Z(n3606) );
  AND U6682 ( .A(n42), .B(n3607), .Z(n3605) );
  XOR U6683 ( .A(n3608), .B(n3609), .Z(n3607) );
  XOR U6684 ( .A(DB[3511]), .B(DB[3504]), .Z(n3609) );
  AND U6685 ( .A(n46), .B(n3610), .Z(n3608) );
  XOR U6686 ( .A(n3611), .B(n3612), .Z(n3610) );
  XOR U6687 ( .A(DB[3504]), .B(DB[3497]), .Z(n3612) );
  AND U6688 ( .A(n50), .B(n3613), .Z(n3611) );
  XOR U6689 ( .A(n3614), .B(n3615), .Z(n3613) );
  XOR U6690 ( .A(DB[3497]), .B(DB[3490]), .Z(n3615) );
  AND U6691 ( .A(n54), .B(n3616), .Z(n3614) );
  XOR U6692 ( .A(n3617), .B(n3618), .Z(n3616) );
  XOR U6693 ( .A(DB[3490]), .B(DB[3483]), .Z(n3618) );
  AND U6694 ( .A(n58), .B(n3619), .Z(n3617) );
  XOR U6695 ( .A(n3620), .B(n3621), .Z(n3619) );
  XOR U6696 ( .A(DB[3483]), .B(DB[3476]), .Z(n3621) );
  AND U6697 ( .A(n62), .B(n3622), .Z(n3620) );
  XOR U6698 ( .A(n3623), .B(n3624), .Z(n3622) );
  XOR U6699 ( .A(DB[3476]), .B(DB[3469]), .Z(n3624) );
  AND U6700 ( .A(n66), .B(n3625), .Z(n3623) );
  XOR U6701 ( .A(n3626), .B(n3627), .Z(n3625) );
  XOR U6702 ( .A(DB[3469]), .B(DB[3462]), .Z(n3627) );
  AND U6703 ( .A(n70), .B(n3628), .Z(n3626) );
  XOR U6704 ( .A(n3629), .B(n3630), .Z(n3628) );
  XOR U6705 ( .A(DB[3462]), .B(DB[3455]), .Z(n3630) );
  AND U6706 ( .A(n74), .B(n3631), .Z(n3629) );
  XOR U6707 ( .A(n3632), .B(n3633), .Z(n3631) );
  XOR U6708 ( .A(DB[3455]), .B(DB[3448]), .Z(n3633) );
  AND U6709 ( .A(n78), .B(n3634), .Z(n3632) );
  XOR U6710 ( .A(n3635), .B(n3636), .Z(n3634) );
  XOR U6711 ( .A(DB[3448]), .B(DB[3441]), .Z(n3636) );
  AND U6712 ( .A(n82), .B(n3637), .Z(n3635) );
  XOR U6713 ( .A(n3638), .B(n3639), .Z(n3637) );
  XOR U6714 ( .A(DB[3441]), .B(DB[3434]), .Z(n3639) );
  AND U6715 ( .A(n86), .B(n3640), .Z(n3638) );
  XOR U6716 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U6717 ( .A(DB[3434]), .B(DB[3427]), .Z(n3642) );
  AND U6718 ( .A(n90), .B(n3643), .Z(n3641) );
  XOR U6719 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U6720 ( .A(DB[3427]), .B(DB[3420]), .Z(n3645) );
  AND U6721 ( .A(n94), .B(n3646), .Z(n3644) );
  XOR U6722 ( .A(n3647), .B(n3648), .Z(n3646) );
  XOR U6723 ( .A(DB[3420]), .B(DB[3413]), .Z(n3648) );
  AND U6724 ( .A(n98), .B(n3649), .Z(n3647) );
  XOR U6725 ( .A(n3650), .B(n3651), .Z(n3649) );
  XOR U6726 ( .A(DB[3413]), .B(DB[3406]), .Z(n3651) );
  AND U6727 ( .A(n102), .B(n3652), .Z(n3650) );
  XOR U6728 ( .A(n3653), .B(n3654), .Z(n3652) );
  XOR U6729 ( .A(DB[3406]), .B(DB[3399]), .Z(n3654) );
  AND U6730 ( .A(n106), .B(n3655), .Z(n3653) );
  XOR U6731 ( .A(n3656), .B(n3657), .Z(n3655) );
  XOR U6732 ( .A(DB[3399]), .B(DB[3392]), .Z(n3657) );
  AND U6733 ( .A(n110), .B(n3658), .Z(n3656) );
  XOR U6734 ( .A(n3659), .B(n3660), .Z(n3658) );
  XOR U6735 ( .A(DB[3392]), .B(DB[3385]), .Z(n3660) );
  AND U6736 ( .A(n114), .B(n3661), .Z(n3659) );
  XOR U6737 ( .A(n3662), .B(n3663), .Z(n3661) );
  XOR U6738 ( .A(DB[3385]), .B(DB[3378]), .Z(n3663) );
  AND U6739 ( .A(n118), .B(n3664), .Z(n3662) );
  XOR U6740 ( .A(n3665), .B(n3666), .Z(n3664) );
  XOR U6741 ( .A(DB[3378]), .B(DB[3371]), .Z(n3666) );
  AND U6742 ( .A(n122), .B(n3667), .Z(n3665) );
  XOR U6743 ( .A(n3668), .B(n3669), .Z(n3667) );
  XOR U6744 ( .A(DB[3371]), .B(DB[3364]), .Z(n3669) );
  AND U6745 ( .A(n126), .B(n3670), .Z(n3668) );
  XOR U6746 ( .A(n3671), .B(n3672), .Z(n3670) );
  XOR U6747 ( .A(DB[3364]), .B(DB[3357]), .Z(n3672) );
  AND U6748 ( .A(n130), .B(n3673), .Z(n3671) );
  XOR U6749 ( .A(n3674), .B(n3675), .Z(n3673) );
  XOR U6750 ( .A(DB[3357]), .B(DB[3350]), .Z(n3675) );
  AND U6751 ( .A(n134), .B(n3676), .Z(n3674) );
  XOR U6752 ( .A(n3677), .B(n3678), .Z(n3676) );
  XOR U6753 ( .A(DB[3350]), .B(DB[3343]), .Z(n3678) );
  AND U6754 ( .A(n138), .B(n3679), .Z(n3677) );
  XOR U6755 ( .A(n3680), .B(n3681), .Z(n3679) );
  XOR U6756 ( .A(DB[3343]), .B(DB[3336]), .Z(n3681) );
  AND U6757 ( .A(n142), .B(n3682), .Z(n3680) );
  XOR U6758 ( .A(n3683), .B(n3684), .Z(n3682) );
  XOR U6759 ( .A(DB[3336]), .B(DB[3329]), .Z(n3684) );
  AND U6760 ( .A(n146), .B(n3685), .Z(n3683) );
  XOR U6761 ( .A(n3686), .B(n3687), .Z(n3685) );
  XOR U6762 ( .A(DB[3329]), .B(DB[3322]), .Z(n3687) );
  AND U6763 ( .A(n150), .B(n3688), .Z(n3686) );
  XOR U6764 ( .A(n3689), .B(n3690), .Z(n3688) );
  XOR U6765 ( .A(DB[3322]), .B(DB[3315]), .Z(n3690) );
  AND U6766 ( .A(n154), .B(n3691), .Z(n3689) );
  XOR U6767 ( .A(n3692), .B(n3693), .Z(n3691) );
  XOR U6768 ( .A(DB[3315]), .B(DB[3308]), .Z(n3693) );
  AND U6769 ( .A(n158), .B(n3694), .Z(n3692) );
  XOR U6770 ( .A(n3695), .B(n3696), .Z(n3694) );
  XOR U6771 ( .A(DB[3308]), .B(DB[3301]), .Z(n3696) );
  AND U6772 ( .A(n162), .B(n3697), .Z(n3695) );
  XOR U6773 ( .A(n3698), .B(n3699), .Z(n3697) );
  XOR U6774 ( .A(DB[3301]), .B(DB[3294]), .Z(n3699) );
  AND U6775 ( .A(n166), .B(n3700), .Z(n3698) );
  XOR U6776 ( .A(n3701), .B(n3702), .Z(n3700) );
  XOR U6777 ( .A(DB[3294]), .B(DB[3287]), .Z(n3702) );
  AND U6778 ( .A(n170), .B(n3703), .Z(n3701) );
  XOR U6779 ( .A(n3704), .B(n3705), .Z(n3703) );
  XOR U6780 ( .A(DB[3287]), .B(DB[3280]), .Z(n3705) );
  AND U6781 ( .A(n174), .B(n3706), .Z(n3704) );
  XOR U6782 ( .A(n3707), .B(n3708), .Z(n3706) );
  XOR U6783 ( .A(DB[3280]), .B(DB[3273]), .Z(n3708) );
  AND U6784 ( .A(n178), .B(n3709), .Z(n3707) );
  XOR U6785 ( .A(n3710), .B(n3711), .Z(n3709) );
  XOR U6786 ( .A(DB[3273]), .B(DB[3266]), .Z(n3711) );
  AND U6787 ( .A(n182), .B(n3712), .Z(n3710) );
  XOR U6788 ( .A(n3713), .B(n3714), .Z(n3712) );
  XOR U6789 ( .A(DB[3266]), .B(DB[3259]), .Z(n3714) );
  AND U6790 ( .A(n186), .B(n3715), .Z(n3713) );
  XOR U6791 ( .A(n3716), .B(n3717), .Z(n3715) );
  XOR U6792 ( .A(DB[3259]), .B(DB[3252]), .Z(n3717) );
  AND U6793 ( .A(n190), .B(n3718), .Z(n3716) );
  XOR U6794 ( .A(n3719), .B(n3720), .Z(n3718) );
  XOR U6795 ( .A(DB[3252]), .B(DB[3245]), .Z(n3720) );
  AND U6796 ( .A(n194), .B(n3721), .Z(n3719) );
  XOR U6797 ( .A(n3722), .B(n3723), .Z(n3721) );
  XOR U6798 ( .A(DB[3245]), .B(DB[3238]), .Z(n3723) );
  AND U6799 ( .A(n198), .B(n3724), .Z(n3722) );
  XOR U6800 ( .A(n3725), .B(n3726), .Z(n3724) );
  XOR U6801 ( .A(DB[3238]), .B(DB[3231]), .Z(n3726) );
  AND U6802 ( .A(n202), .B(n3727), .Z(n3725) );
  XOR U6803 ( .A(n3728), .B(n3729), .Z(n3727) );
  XOR U6804 ( .A(DB[3231]), .B(DB[3224]), .Z(n3729) );
  AND U6805 ( .A(n206), .B(n3730), .Z(n3728) );
  XOR U6806 ( .A(n3731), .B(n3732), .Z(n3730) );
  XOR U6807 ( .A(DB[3224]), .B(DB[3217]), .Z(n3732) );
  AND U6808 ( .A(n210), .B(n3733), .Z(n3731) );
  XOR U6809 ( .A(n3734), .B(n3735), .Z(n3733) );
  XOR U6810 ( .A(DB[3217]), .B(DB[3210]), .Z(n3735) );
  AND U6811 ( .A(n214), .B(n3736), .Z(n3734) );
  XOR U6812 ( .A(n3737), .B(n3738), .Z(n3736) );
  XOR U6813 ( .A(DB[3210]), .B(DB[3203]), .Z(n3738) );
  AND U6814 ( .A(n218), .B(n3739), .Z(n3737) );
  XOR U6815 ( .A(n3740), .B(n3741), .Z(n3739) );
  XOR U6816 ( .A(DB[3203]), .B(DB[3196]), .Z(n3741) );
  AND U6817 ( .A(n222), .B(n3742), .Z(n3740) );
  XOR U6818 ( .A(n3743), .B(n3744), .Z(n3742) );
  XOR U6819 ( .A(DB[3196]), .B(DB[3189]), .Z(n3744) );
  AND U6820 ( .A(n226), .B(n3745), .Z(n3743) );
  XOR U6821 ( .A(n3746), .B(n3747), .Z(n3745) );
  XOR U6822 ( .A(DB[3189]), .B(DB[3182]), .Z(n3747) );
  AND U6823 ( .A(n230), .B(n3748), .Z(n3746) );
  XOR U6824 ( .A(n3749), .B(n3750), .Z(n3748) );
  XOR U6825 ( .A(DB[3182]), .B(DB[3175]), .Z(n3750) );
  AND U6826 ( .A(n234), .B(n3751), .Z(n3749) );
  XOR U6827 ( .A(n3752), .B(n3753), .Z(n3751) );
  XOR U6828 ( .A(DB[3175]), .B(DB[3168]), .Z(n3753) );
  AND U6829 ( .A(n238), .B(n3754), .Z(n3752) );
  XOR U6830 ( .A(n3755), .B(n3756), .Z(n3754) );
  XOR U6831 ( .A(DB[3168]), .B(DB[3161]), .Z(n3756) );
  AND U6832 ( .A(n242), .B(n3757), .Z(n3755) );
  XOR U6833 ( .A(n3758), .B(n3759), .Z(n3757) );
  XOR U6834 ( .A(DB[3161]), .B(DB[3154]), .Z(n3759) );
  AND U6835 ( .A(n246), .B(n3760), .Z(n3758) );
  XOR U6836 ( .A(n3761), .B(n3762), .Z(n3760) );
  XOR U6837 ( .A(DB[3154]), .B(DB[3147]), .Z(n3762) );
  AND U6838 ( .A(n250), .B(n3763), .Z(n3761) );
  XOR U6839 ( .A(n3764), .B(n3765), .Z(n3763) );
  XOR U6840 ( .A(DB[3147]), .B(DB[3140]), .Z(n3765) );
  AND U6841 ( .A(n254), .B(n3766), .Z(n3764) );
  XOR U6842 ( .A(n3767), .B(n3768), .Z(n3766) );
  XOR U6843 ( .A(DB[3140]), .B(DB[3133]), .Z(n3768) );
  AND U6844 ( .A(n258), .B(n3769), .Z(n3767) );
  XOR U6845 ( .A(n3770), .B(n3771), .Z(n3769) );
  XOR U6846 ( .A(DB[3133]), .B(DB[3126]), .Z(n3771) );
  AND U6847 ( .A(n262), .B(n3772), .Z(n3770) );
  XOR U6848 ( .A(n3773), .B(n3774), .Z(n3772) );
  XOR U6849 ( .A(DB[3126]), .B(DB[3119]), .Z(n3774) );
  AND U6850 ( .A(n266), .B(n3775), .Z(n3773) );
  XOR U6851 ( .A(n3776), .B(n3777), .Z(n3775) );
  XOR U6852 ( .A(DB[3119]), .B(DB[3112]), .Z(n3777) );
  AND U6853 ( .A(n270), .B(n3778), .Z(n3776) );
  XOR U6854 ( .A(n3779), .B(n3780), .Z(n3778) );
  XOR U6855 ( .A(DB[3112]), .B(DB[3105]), .Z(n3780) );
  AND U6856 ( .A(n274), .B(n3781), .Z(n3779) );
  XOR U6857 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U6858 ( .A(DB[3105]), .B(DB[3098]), .Z(n3783) );
  AND U6859 ( .A(n278), .B(n3784), .Z(n3782) );
  XOR U6860 ( .A(n3785), .B(n3786), .Z(n3784) );
  XOR U6861 ( .A(DB[3098]), .B(DB[3091]), .Z(n3786) );
  AND U6862 ( .A(n282), .B(n3787), .Z(n3785) );
  XOR U6863 ( .A(n3788), .B(n3789), .Z(n3787) );
  XOR U6864 ( .A(DB[3091]), .B(DB[3084]), .Z(n3789) );
  AND U6865 ( .A(n286), .B(n3790), .Z(n3788) );
  XOR U6866 ( .A(n3791), .B(n3792), .Z(n3790) );
  XOR U6867 ( .A(DB[3084]), .B(DB[3077]), .Z(n3792) );
  AND U6868 ( .A(n290), .B(n3793), .Z(n3791) );
  XOR U6869 ( .A(n3794), .B(n3795), .Z(n3793) );
  XOR U6870 ( .A(DB[3077]), .B(DB[3070]), .Z(n3795) );
  AND U6871 ( .A(n294), .B(n3796), .Z(n3794) );
  XOR U6872 ( .A(n3797), .B(n3798), .Z(n3796) );
  XOR U6873 ( .A(DB[3070]), .B(DB[3063]), .Z(n3798) );
  AND U6874 ( .A(n298), .B(n3799), .Z(n3797) );
  XOR U6875 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U6876 ( .A(DB[3063]), .B(DB[3056]), .Z(n3801) );
  AND U6877 ( .A(n302), .B(n3802), .Z(n3800) );
  XOR U6878 ( .A(n3803), .B(n3804), .Z(n3802) );
  XOR U6879 ( .A(DB[3056]), .B(DB[3049]), .Z(n3804) );
  AND U6880 ( .A(n306), .B(n3805), .Z(n3803) );
  XOR U6881 ( .A(n3806), .B(n3807), .Z(n3805) );
  XOR U6882 ( .A(DB[3049]), .B(DB[3042]), .Z(n3807) );
  AND U6883 ( .A(n310), .B(n3808), .Z(n3806) );
  XOR U6884 ( .A(n3809), .B(n3810), .Z(n3808) );
  XOR U6885 ( .A(DB[3042]), .B(DB[3035]), .Z(n3810) );
  AND U6886 ( .A(n314), .B(n3811), .Z(n3809) );
  XOR U6887 ( .A(n3812), .B(n3813), .Z(n3811) );
  XOR U6888 ( .A(DB[3035]), .B(DB[3028]), .Z(n3813) );
  AND U6889 ( .A(n318), .B(n3814), .Z(n3812) );
  XOR U6890 ( .A(n3815), .B(n3816), .Z(n3814) );
  XOR U6891 ( .A(DB[3028]), .B(DB[3021]), .Z(n3816) );
  AND U6892 ( .A(n322), .B(n3817), .Z(n3815) );
  XOR U6893 ( .A(n3818), .B(n3819), .Z(n3817) );
  XOR U6894 ( .A(DB[3021]), .B(DB[3014]), .Z(n3819) );
  AND U6895 ( .A(n326), .B(n3820), .Z(n3818) );
  XOR U6896 ( .A(n3821), .B(n3822), .Z(n3820) );
  XOR U6897 ( .A(DB[3014]), .B(DB[3007]), .Z(n3822) );
  AND U6898 ( .A(n330), .B(n3823), .Z(n3821) );
  XOR U6899 ( .A(n3824), .B(n3825), .Z(n3823) );
  XOR U6900 ( .A(DB[3007]), .B(DB[3000]), .Z(n3825) );
  AND U6901 ( .A(n334), .B(n3826), .Z(n3824) );
  XOR U6902 ( .A(n3827), .B(n3828), .Z(n3826) );
  XOR U6903 ( .A(DB[3000]), .B(DB[2993]), .Z(n3828) );
  AND U6904 ( .A(n338), .B(n3829), .Z(n3827) );
  XOR U6905 ( .A(n3830), .B(n3831), .Z(n3829) );
  XOR U6906 ( .A(DB[2993]), .B(DB[2986]), .Z(n3831) );
  AND U6907 ( .A(n342), .B(n3832), .Z(n3830) );
  XOR U6908 ( .A(n3833), .B(n3834), .Z(n3832) );
  XOR U6909 ( .A(DB[2986]), .B(DB[2979]), .Z(n3834) );
  AND U6910 ( .A(n346), .B(n3835), .Z(n3833) );
  XOR U6911 ( .A(n3836), .B(n3837), .Z(n3835) );
  XOR U6912 ( .A(DB[2979]), .B(DB[2972]), .Z(n3837) );
  AND U6913 ( .A(n350), .B(n3838), .Z(n3836) );
  XOR U6914 ( .A(n3839), .B(n3840), .Z(n3838) );
  XOR U6915 ( .A(DB[2972]), .B(DB[2965]), .Z(n3840) );
  AND U6916 ( .A(n354), .B(n3841), .Z(n3839) );
  XOR U6917 ( .A(n3842), .B(n3843), .Z(n3841) );
  XOR U6918 ( .A(DB[2965]), .B(DB[2958]), .Z(n3843) );
  AND U6919 ( .A(n358), .B(n3844), .Z(n3842) );
  XOR U6920 ( .A(n3845), .B(n3846), .Z(n3844) );
  XOR U6921 ( .A(DB[2958]), .B(DB[2951]), .Z(n3846) );
  AND U6922 ( .A(n362), .B(n3847), .Z(n3845) );
  XOR U6923 ( .A(n3848), .B(n3849), .Z(n3847) );
  XOR U6924 ( .A(DB[2951]), .B(DB[2944]), .Z(n3849) );
  AND U6925 ( .A(n366), .B(n3850), .Z(n3848) );
  XOR U6926 ( .A(n3851), .B(n3852), .Z(n3850) );
  XOR U6927 ( .A(DB[2944]), .B(DB[2937]), .Z(n3852) );
  AND U6928 ( .A(n370), .B(n3853), .Z(n3851) );
  XOR U6929 ( .A(n3854), .B(n3855), .Z(n3853) );
  XOR U6930 ( .A(DB[2937]), .B(DB[2930]), .Z(n3855) );
  AND U6931 ( .A(n374), .B(n3856), .Z(n3854) );
  XOR U6932 ( .A(n3857), .B(n3858), .Z(n3856) );
  XOR U6933 ( .A(DB[2930]), .B(DB[2923]), .Z(n3858) );
  AND U6934 ( .A(n378), .B(n3859), .Z(n3857) );
  XOR U6935 ( .A(n3860), .B(n3861), .Z(n3859) );
  XOR U6936 ( .A(DB[2923]), .B(DB[2916]), .Z(n3861) );
  AND U6937 ( .A(n382), .B(n3862), .Z(n3860) );
  XOR U6938 ( .A(n3863), .B(n3864), .Z(n3862) );
  XOR U6939 ( .A(DB[2916]), .B(DB[2909]), .Z(n3864) );
  AND U6940 ( .A(n386), .B(n3865), .Z(n3863) );
  XOR U6941 ( .A(n3866), .B(n3867), .Z(n3865) );
  XOR U6942 ( .A(DB[2909]), .B(DB[2902]), .Z(n3867) );
  AND U6943 ( .A(n390), .B(n3868), .Z(n3866) );
  XOR U6944 ( .A(n3869), .B(n3870), .Z(n3868) );
  XOR U6945 ( .A(DB[2902]), .B(DB[2895]), .Z(n3870) );
  AND U6946 ( .A(n394), .B(n3871), .Z(n3869) );
  XOR U6947 ( .A(n3872), .B(n3873), .Z(n3871) );
  XOR U6948 ( .A(DB[2895]), .B(DB[2888]), .Z(n3873) );
  AND U6949 ( .A(n398), .B(n3874), .Z(n3872) );
  XOR U6950 ( .A(n3875), .B(n3876), .Z(n3874) );
  XOR U6951 ( .A(DB[2888]), .B(DB[2881]), .Z(n3876) );
  AND U6952 ( .A(n402), .B(n3877), .Z(n3875) );
  XOR U6953 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR U6954 ( .A(DB[2881]), .B(DB[2874]), .Z(n3879) );
  AND U6955 ( .A(n406), .B(n3880), .Z(n3878) );
  XOR U6956 ( .A(n3881), .B(n3882), .Z(n3880) );
  XOR U6957 ( .A(DB[2874]), .B(DB[2867]), .Z(n3882) );
  AND U6958 ( .A(n410), .B(n3883), .Z(n3881) );
  XOR U6959 ( .A(n3884), .B(n3885), .Z(n3883) );
  XOR U6960 ( .A(DB[2867]), .B(DB[2860]), .Z(n3885) );
  AND U6961 ( .A(n414), .B(n3886), .Z(n3884) );
  XOR U6962 ( .A(n3887), .B(n3888), .Z(n3886) );
  XOR U6963 ( .A(DB[2860]), .B(DB[2853]), .Z(n3888) );
  AND U6964 ( .A(n418), .B(n3889), .Z(n3887) );
  XOR U6965 ( .A(n3890), .B(n3891), .Z(n3889) );
  XOR U6966 ( .A(DB[2853]), .B(DB[2846]), .Z(n3891) );
  AND U6967 ( .A(n422), .B(n3892), .Z(n3890) );
  XOR U6968 ( .A(n3893), .B(n3894), .Z(n3892) );
  XOR U6969 ( .A(DB[2846]), .B(DB[2839]), .Z(n3894) );
  AND U6970 ( .A(n426), .B(n3895), .Z(n3893) );
  XOR U6971 ( .A(n3896), .B(n3897), .Z(n3895) );
  XOR U6972 ( .A(DB[2839]), .B(DB[2832]), .Z(n3897) );
  AND U6973 ( .A(n430), .B(n3898), .Z(n3896) );
  XOR U6974 ( .A(n3899), .B(n3900), .Z(n3898) );
  XOR U6975 ( .A(DB[2832]), .B(DB[2825]), .Z(n3900) );
  AND U6976 ( .A(n434), .B(n3901), .Z(n3899) );
  XOR U6977 ( .A(n3902), .B(n3903), .Z(n3901) );
  XOR U6978 ( .A(DB[2825]), .B(DB[2818]), .Z(n3903) );
  AND U6979 ( .A(n438), .B(n3904), .Z(n3902) );
  XOR U6980 ( .A(n3905), .B(n3906), .Z(n3904) );
  XOR U6981 ( .A(DB[2818]), .B(DB[2811]), .Z(n3906) );
  AND U6982 ( .A(n442), .B(n3907), .Z(n3905) );
  XOR U6983 ( .A(n3908), .B(n3909), .Z(n3907) );
  XOR U6984 ( .A(DB[2811]), .B(DB[2804]), .Z(n3909) );
  AND U6985 ( .A(n446), .B(n3910), .Z(n3908) );
  XOR U6986 ( .A(n3911), .B(n3912), .Z(n3910) );
  XOR U6987 ( .A(DB[2804]), .B(DB[2797]), .Z(n3912) );
  AND U6988 ( .A(n450), .B(n3913), .Z(n3911) );
  XOR U6989 ( .A(n3914), .B(n3915), .Z(n3913) );
  XOR U6990 ( .A(DB[2797]), .B(DB[2790]), .Z(n3915) );
  AND U6991 ( .A(n454), .B(n3916), .Z(n3914) );
  XOR U6992 ( .A(n3917), .B(n3918), .Z(n3916) );
  XOR U6993 ( .A(DB[2790]), .B(DB[2783]), .Z(n3918) );
  AND U6994 ( .A(n458), .B(n3919), .Z(n3917) );
  XOR U6995 ( .A(n3920), .B(n3921), .Z(n3919) );
  XOR U6996 ( .A(DB[2783]), .B(DB[2776]), .Z(n3921) );
  AND U6997 ( .A(n462), .B(n3922), .Z(n3920) );
  XOR U6998 ( .A(n3923), .B(n3924), .Z(n3922) );
  XOR U6999 ( .A(DB[2776]), .B(DB[2769]), .Z(n3924) );
  AND U7000 ( .A(n466), .B(n3925), .Z(n3923) );
  XOR U7001 ( .A(n3926), .B(n3927), .Z(n3925) );
  XOR U7002 ( .A(DB[2769]), .B(DB[2762]), .Z(n3927) );
  AND U7003 ( .A(n470), .B(n3928), .Z(n3926) );
  XOR U7004 ( .A(n3929), .B(n3930), .Z(n3928) );
  XOR U7005 ( .A(DB[2762]), .B(DB[2755]), .Z(n3930) );
  AND U7006 ( .A(n474), .B(n3931), .Z(n3929) );
  XOR U7007 ( .A(n3932), .B(n3933), .Z(n3931) );
  XOR U7008 ( .A(DB[2755]), .B(DB[2748]), .Z(n3933) );
  AND U7009 ( .A(n478), .B(n3934), .Z(n3932) );
  XOR U7010 ( .A(n3935), .B(n3936), .Z(n3934) );
  XOR U7011 ( .A(DB[2748]), .B(DB[2741]), .Z(n3936) );
  AND U7012 ( .A(n482), .B(n3937), .Z(n3935) );
  XOR U7013 ( .A(n3938), .B(n3939), .Z(n3937) );
  XOR U7014 ( .A(DB[2741]), .B(DB[2734]), .Z(n3939) );
  AND U7015 ( .A(n486), .B(n3940), .Z(n3938) );
  XOR U7016 ( .A(n3941), .B(n3942), .Z(n3940) );
  XOR U7017 ( .A(DB[2734]), .B(DB[2727]), .Z(n3942) );
  AND U7018 ( .A(n490), .B(n3943), .Z(n3941) );
  XOR U7019 ( .A(n3944), .B(n3945), .Z(n3943) );
  XOR U7020 ( .A(DB[2727]), .B(DB[2720]), .Z(n3945) );
  AND U7021 ( .A(n494), .B(n3946), .Z(n3944) );
  XOR U7022 ( .A(n3947), .B(n3948), .Z(n3946) );
  XOR U7023 ( .A(DB[2720]), .B(DB[2713]), .Z(n3948) );
  AND U7024 ( .A(n498), .B(n3949), .Z(n3947) );
  XOR U7025 ( .A(n3950), .B(n3951), .Z(n3949) );
  XOR U7026 ( .A(DB[2713]), .B(DB[2706]), .Z(n3951) );
  AND U7027 ( .A(n502), .B(n3952), .Z(n3950) );
  XOR U7028 ( .A(n3953), .B(n3954), .Z(n3952) );
  XOR U7029 ( .A(DB[2706]), .B(DB[2699]), .Z(n3954) );
  AND U7030 ( .A(n506), .B(n3955), .Z(n3953) );
  XOR U7031 ( .A(n3956), .B(n3957), .Z(n3955) );
  XOR U7032 ( .A(DB[2699]), .B(DB[2692]), .Z(n3957) );
  AND U7033 ( .A(n510), .B(n3958), .Z(n3956) );
  XOR U7034 ( .A(n3959), .B(n3960), .Z(n3958) );
  XOR U7035 ( .A(DB[2692]), .B(DB[2685]), .Z(n3960) );
  AND U7036 ( .A(n514), .B(n3961), .Z(n3959) );
  XOR U7037 ( .A(n3962), .B(n3963), .Z(n3961) );
  XOR U7038 ( .A(DB[2685]), .B(DB[2678]), .Z(n3963) );
  AND U7039 ( .A(n518), .B(n3964), .Z(n3962) );
  XOR U7040 ( .A(n3965), .B(n3966), .Z(n3964) );
  XOR U7041 ( .A(DB[2678]), .B(DB[2671]), .Z(n3966) );
  AND U7042 ( .A(n522), .B(n3967), .Z(n3965) );
  XOR U7043 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR U7044 ( .A(DB[2671]), .B(DB[2664]), .Z(n3969) );
  AND U7045 ( .A(n526), .B(n3970), .Z(n3968) );
  XOR U7046 ( .A(n3971), .B(n3972), .Z(n3970) );
  XOR U7047 ( .A(DB[2664]), .B(DB[2657]), .Z(n3972) );
  AND U7048 ( .A(n530), .B(n3973), .Z(n3971) );
  XOR U7049 ( .A(n3974), .B(n3975), .Z(n3973) );
  XOR U7050 ( .A(DB[2657]), .B(DB[2650]), .Z(n3975) );
  AND U7051 ( .A(n534), .B(n3976), .Z(n3974) );
  XOR U7052 ( .A(n3977), .B(n3978), .Z(n3976) );
  XOR U7053 ( .A(DB[2650]), .B(DB[2643]), .Z(n3978) );
  AND U7054 ( .A(n538), .B(n3979), .Z(n3977) );
  XOR U7055 ( .A(n3980), .B(n3981), .Z(n3979) );
  XOR U7056 ( .A(DB[2643]), .B(DB[2636]), .Z(n3981) );
  AND U7057 ( .A(n542), .B(n3982), .Z(n3980) );
  XOR U7058 ( .A(n3983), .B(n3984), .Z(n3982) );
  XOR U7059 ( .A(DB[2636]), .B(DB[2629]), .Z(n3984) );
  AND U7060 ( .A(n546), .B(n3985), .Z(n3983) );
  XOR U7061 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U7062 ( .A(DB[2629]), .B(DB[2622]), .Z(n3987) );
  AND U7063 ( .A(n550), .B(n3988), .Z(n3986) );
  XOR U7064 ( .A(n3989), .B(n3990), .Z(n3988) );
  XOR U7065 ( .A(DB[2622]), .B(DB[2615]), .Z(n3990) );
  AND U7066 ( .A(n554), .B(n3991), .Z(n3989) );
  XOR U7067 ( .A(n3992), .B(n3993), .Z(n3991) );
  XOR U7068 ( .A(DB[2615]), .B(DB[2608]), .Z(n3993) );
  AND U7069 ( .A(n558), .B(n3994), .Z(n3992) );
  XOR U7070 ( .A(n3995), .B(n3996), .Z(n3994) );
  XOR U7071 ( .A(DB[2608]), .B(DB[2601]), .Z(n3996) );
  AND U7072 ( .A(n562), .B(n3997), .Z(n3995) );
  XOR U7073 ( .A(n3998), .B(n3999), .Z(n3997) );
  XOR U7074 ( .A(DB[2601]), .B(DB[2594]), .Z(n3999) );
  AND U7075 ( .A(n566), .B(n4000), .Z(n3998) );
  XOR U7076 ( .A(n4001), .B(n4002), .Z(n4000) );
  XOR U7077 ( .A(DB[2594]), .B(DB[2587]), .Z(n4002) );
  AND U7078 ( .A(n570), .B(n4003), .Z(n4001) );
  XOR U7079 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U7080 ( .A(DB[2587]), .B(DB[2580]), .Z(n4005) );
  AND U7081 ( .A(n574), .B(n4006), .Z(n4004) );
  XOR U7082 ( .A(n4007), .B(n4008), .Z(n4006) );
  XOR U7083 ( .A(DB[2580]), .B(DB[2573]), .Z(n4008) );
  AND U7084 ( .A(n578), .B(n4009), .Z(n4007) );
  XOR U7085 ( .A(n4010), .B(n4011), .Z(n4009) );
  XOR U7086 ( .A(DB[2573]), .B(DB[2566]), .Z(n4011) );
  AND U7087 ( .A(n582), .B(n4012), .Z(n4010) );
  XOR U7088 ( .A(n4013), .B(n4014), .Z(n4012) );
  XOR U7089 ( .A(DB[2566]), .B(DB[2559]), .Z(n4014) );
  AND U7090 ( .A(n586), .B(n4015), .Z(n4013) );
  XOR U7091 ( .A(n4016), .B(n4017), .Z(n4015) );
  XOR U7092 ( .A(DB[2559]), .B(DB[2552]), .Z(n4017) );
  AND U7093 ( .A(n590), .B(n4018), .Z(n4016) );
  XOR U7094 ( .A(n4019), .B(n4020), .Z(n4018) );
  XOR U7095 ( .A(DB[2552]), .B(DB[2545]), .Z(n4020) );
  AND U7096 ( .A(n594), .B(n4021), .Z(n4019) );
  XOR U7097 ( .A(n4022), .B(n4023), .Z(n4021) );
  XOR U7098 ( .A(DB[2545]), .B(DB[2538]), .Z(n4023) );
  AND U7099 ( .A(n598), .B(n4024), .Z(n4022) );
  XOR U7100 ( .A(n4025), .B(n4026), .Z(n4024) );
  XOR U7101 ( .A(DB[2538]), .B(DB[2531]), .Z(n4026) );
  AND U7102 ( .A(n602), .B(n4027), .Z(n4025) );
  XOR U7103 ( .A(n4028), .B(n4029), .Z(n4027) );
  XOR U7104 ( .A(DB[2531]), .B(DB[2524]), .Z(n4029) );
  AND U7105 ( .A(n606), .B(n4030), .Z(n4028) );
  XOR U7106 ( .A(n4031), .B(n4032), .Z(n4030) );
  XOR U7107 ( .A(DB[2524]), .B(DB[2517]), .Z(n4032) );
  AND U7108 ( .A(n610), .B(n4033), .Z(n4031) );
  XOR U7109 ( .A(n4034), .B(n4035), .Z(n4033) );
  XOR U7110 ( .A(DB[2517]), .B(DB[2510]), .Z(n4035) );
  AND U7111 ( .A(n614), .B(n4036), .Z(n4034) );
  XOR U7112 ( .A(n4037), .B(n4038), .Z(n4036) );
  XOR U7113 ( .A(DB[2510]), .B(DB[2503]), .Z(n4038) );
  AND U7114 ( .A(n618), .B(n4039), .Z(n4037) );
  XOR U7115 ( .A(n4040), .B(n4041), .Z(n4039) );
  XOR U7116 ( .A(DB[2503]), .B(DB[2496]), .Z(n4041) );
  AND U7117 ( .A(n622), .B(n4042), .Z(n4040) );
  XOR U7118 ( .A(n4043), .B(n4044), .Z(n4042) );
  XOR U7119 ( .A(DB[2496]), .B(DB[2489]), .Z(n4044) );
  AND U7120 ( .A(n626), .B(n4045), .Z(n4043) );
  XOR U7121 ( .A(n4046), .B(n4047), .Z(n4045) );
  XOR U7122 ( .A(DB[2489]), .B(DB[2482]), .Z(n4047) );
  AND U7123 ( .A(n630), .B(n4048), .Z(n4046) );
  XOR U7124 ( .A(n4049), .B(n4050), .Z(n4048) );
  XOR U7125 ( .A(DB[2482]), .B(DB[2475]), .Z(n4050) );
  AND U7126 ( .A(n634), .B(n4051), .Z(n4049) );
  XOR U7127 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U7128 ( .A(DB[2475]), .B(DB[2468]), .Z(n4053) );
  AND U7129 ( .A(n638), .B(n4054), .Z(n4052) );
  XOR U7130 ( .A(n4055), .B(n4056), .Z(n4054) );
  XOR U7131 ( .A(DB[2468]), .B(DB[2461]), .Z(n4056) );
  AND U7132 ( .A(n642), .B(n4057), .Z(n4055) );
  XOR U7133 ( .A(n4058), .B(n4059), .Z(n4057) );
  XOR U7134 ( .A(DB[2461]), .B(DB[2454]), .Z(n4059) );
  AND U7135 ( .A(n646), .B(n4060), .Z(n4058) );
  XOR U7136 ( .A(n4061), .B(n4062), .Z(n4060) );
  XOR U7137 ( .A(DB[2454]), .B(DB[2447]), .Z(n4062) );
  AND U7138 ( .A(n650), .B(n4063), .Z(n4061) );
  XOR U7139 ( .A(n4064), .B(n4065), .Z(n4063) );
  XOR U7140 ( .A(DB[2447]), .B(DB[2440]), .Z(n4065) );
  AND U7141 ( .A(n654), .B(n4066), .Z(n4064) );
  XOR U7142 ( .A(n4067), .B(n4068), .Z(n4066) );
  XOR U7143 ( .A(DB[2440]), .B(DB[2433]), .Z(n4068) );
  AND U7144 ( .A(n658), .B(n4069), .Z(n4067) );
  XOR U7145 ( .A(n4070), .B(n4071), .Z(n4069) );
  XOR U7146 ( .A(DB[2433]), .B(DB[2426]), .Z(n4071) );
  AND U7147 ( .A(n662), .B(n4072), .Z(n4070) );
  XOR U7148 ( .A(n4073), .B(n4074), .Z(n4072) );
  XOR U7149 ( .A(DB[2426]), .B(DB[2419]), .Z(n4074) );
  AND U7150 ( .A(n666), .B(n4075), .Z(n4073) );
  XOR U7151 ( .A(n4076), .B(n4077), .Z(n4075) );
  XOR U7152 ( .A(DB[2419]), .B(DB[2412]), .Z(n4077) );
  AND U7153 ( .A(n670), .B(n4078), .Z(n4076) );
  XOR U7154 ( .A(n4079), .B(n4080), .Z(n4078) );
  XOR U7155 ( .A(DB[2412]), .B(DB[2405]), .Z(n4080) );
  AND U7156 ( .A(n674), .B(n4081), .Z(n4079) );
  XOR U7157 ( .A(n4082), .B(n4083), .Z(n4081) );
  XOR U7158 ( .A(DB[2405]), .B(DB[2398]), .Z(n4083) );
  AND U7159 ( .A(n678), .B(n4084), .Z(n4082) );
  XOR U7160 ( .A(n4085), .B(n4086), .Z(n4084) );
  XOR U7161 ( .A(DB[2398]), .B(DB[2391]), .Z(n4086) );
  AND U7162 ( .A(n682), .B(n4087), .Z(n4085) );
  XOR U7163 ( .A(n4088), .B(n4089), .Z(n4087) );
  XOR U7164 ( .A(DB[2391]), .B(DB[2384]), .Z(n4089) );
  AND U7165 ( .A(n686), .B(n4090), .Z(n4088) );
  XOR U7166 ( .A(n4091), .B(n4092), .Z(n4090) );
  XOR U7167 ( .A(DB[2384]), .B(DB[2377]), .Z(n4092) );
  AND U7168 ( .A(n690), .B(n4093), .Z(n4091) );
  XOR U7169 ( .A(n4094), .B(n4095), .Z(n4093) );
  XOR U7170 ( .A(DB[2377]), .B(DB[2370]), .Z(n4095) );
  AND U7171 ( .A(n694), .B(n4096), .Z(n4094) );
  XOR U7172 ( .A(n4097), .B(n4098), .Z(n4096) );
  XOR U7173 ( .A(DB[2370]), .B(DB[2363]), .Z(n4098) );
  AND U7174 ( .A(n698), .B(n4099), .Z(n4097) );
  XOR U7175 ( .A(n4100), .B(n4101), .Z(n4099) );
  XOR U7176 ( .A(DB[2363]), .B(DB[2356]), .Z(n4101) );
  AND U7177 ( .A(n702), .B(n4102), .Z(n4100) );
  XOR U7178 ( .A(n4103), .B(n4104), .Z(n4102) );
  XOR U7179 ( .A(DB[2356]), .B(DB[2349]), .Z(n4104) );
  AND U7180 ( .A(n706), .B(n4105), .Z(n4103) );
  XOR U7181 ( .A(n4106), .B(n4107), .Z(n4105) );
  XOR U7182 ( .A(DB[2349]), .B(DB[2342]), .Z(n4107) );
  AND U7183 ( .A(n710), .B(n4108), .Z(n4106) );
  XOR U7184 ( .A(n4109), .B(n4110), .Z(n4108) );
  XOR U7185 ( .A(DB[2342]), .B(DB[2335]), .Z(n4110) );
  AND U7186 ( .A(n714), .B(n4111), .Z(n4109) );
  XOR U7187 ( .A(n4112), .B(n4113), .Z(n4111) );
  XOR U7188 ( .A(DB[2335]), .B(DB[2328]), .Z(n4113) );
  AND U7189 ( .A(n718), .B(n4114), .Z(n4112) );
  XOR U7190 ( .A(n4115), .B(n4116), .Z(n4114) );
  XOR U7191 ( .A(DB[2328]), .B(DB[2321]), .Z(n4116) );
  AND U7192 ( .A(n722), .B(n4117), .Z(n4115) );
  XOR U7193 ( .A(n4118), .B(n4119), .Z(n4117) );
  XOR U7194 ( .A(DB[2321]), .B(DB[2314]), .Z(n4119) );
  AND U7195 ( .A(n726), .B(n4120), .Z(n4118) );
  XOR U7196 ( .A(n4121), .B(n4122), .Z(n4120) );
  XOR U7197 ( .A(DB[2314]), .B(DB[2307]), .Z(n4122) );
  AND U7198 ( .A(n730), .B(n4123), .Z(n4121) );
  XOR U7199 ( .A(n4124), .B(n4125), .Z(n4123) );
  XOR U7200 ( .A(DB[2307]), .B(DB[2300]), .Z(n4125) );
  AND U7201 ( .A(n734), .B(n4126), .Z(n4124) );
  XOR U7202 ( .A(n4127), .B(n4128), .Z(n4126) );
  XOR U7203 ( .A(DB[2300]), .B(DB[2293]), .Z(n4128) );
  AND U7204 ( .A(n738), .B(n4129), .Z(n4127) );
  XOR U7205 ( .A(n4130), .B(n4131), .Z(n4129) );
  XOR U7206 ( .A(DB[2293]), .B(DB[2286]), .Z(n4131) );
  AND U7207 ( .A(n742), .B(n4132), .Z(n4130) );
  XOR U7208 ( .A(n4133), .B(n4134), .Z(n4132) );
  XOR U7209 ( .A(DB[2286]), .B(DB[2279]), .Z(n4134) );
  AND U7210 ( .A(n746), .B(n4135), .Z(n4133) );
  XOR U7211 ( .A(n4136), .B(n4137), .Z(n4135) );
  XOR U7212 ( .A(DB[2279]), .B(DB[2272]), .Z(n4137) );
  AND U7213 ( .A(n750), .B(n4138), .Z(n4136) );
  XOR U7214 ( .A(n4139), .B(n4140), .Z(n4138) );
  XOR U7215 ( .A(DB[2272]), .B(DB[2265]), .Z(n4140) );
  AND U7216 ( .A(n754), .B(n4141), .Z(n4139) );
  XOR U7217 ( .A(n4142), .B(n4143), .Z(n4141) );
  XOR U7218 ( .A(DB[2265]), .B(DB[2258]), .Z(n4143) );
  AND U7219 ( .A(n758), .B(n4144), .Z(n4142) );
  XOR U7220 ( .A(n4145), .B(n4146), .Z(n4144) );
  XOR U7221 ( .A(DB[2258]), .B(DB[2251]), .Z(n4146) );
  AND U7222 ( .A(n762), .B(n4147), .Z(n4145) );
  XOR U7223 ( .A(n4148), .B(n4149), .Z(n4147) );
  XOR U7224 ( .A(DB[2251]), .B(DB[2244]), .Z(n4149) );
  AND U7225 ( .A(n766), .B(n4150), .Z(n4148) );
  XOR U7226 ( .A(n4151), .B(n4152), .Z(n4150) );
  XOR U7227 ( .A(DB[2244]), .B(DB[2237]), .Z(n4152) );
  AND U7228 ( .A(n770), .B(n4153), .Z(n4151) );
  XOR U7229 ( .A(n4154), .B(n4155), .Z(n4153) );
  XOR U7230 ( .A(DB[2237]), .B(DB[2230]), .Z(n4155) );
  AND U7231 ( .A(n774), .B(n4156), .Z(n4154) );
  XOR U7232 ( .A(n4157), .B(n4158), .Z(n4156) );
  XOR U7233 ( .A(DB[2230]), .B(DB[2223]), .Z(n4158) );
  AND U7234 ( .A(n778), .B(n4159), .Z(n4157) );
  XOR U7235 ( .A(n4160), .B(n4161), .Z(n4159) );
  XOR U7236 ( .A(DB[2223]), .B(DB[2216]), .Z(n4161) );
  AND U7237 ( .A(n782), .B(n4162), .Z(n4160) );
  XOR U7238 ( .A(n4163), .B(n4164), .Z(n4162) );
  XOR U7239 ( .A(DB[2216]), .B(DB[2209]), .Z(n4164) );
  AND U7240 ( .A(n786), .B(n4165), .Z(n4163) );
  XOR U7241 ( .A(n4166), .B(n4167), .Z(n4165) );
  XOR U7242 ( .A(DB[2209]), .B(DB[2202]), .Z(n4167) );
  AND U7243 ( .A(n790), .B(n4168), .Z(n4166) );
  XOR U7244 ( .A(n4169), .B(n4170), .Z(n4168) );
  XOR U7245 ( .A(DB[2202]), .B(DB[2195]), .Z(n4170) );
  AND U7246 ( .A(n794), .B(n4171), .Z(n4169) );
  XOR U7247 ( .A(n4172), .B(n4173), .Z(n4171) );
  XOR U7248 ( .A(DB[2195]), .B(DB[2188]), .Z(n4173) );
  AND U7249 ( .A(n798), .B(n4174), .Z(n4172) );
  XOR U7250 ( .A(n4175), .B(n4176), .Z(n4174) );
  XOR U7251 ( .A(DB[2188]), .B(DB[2181]), .Z(n4176) );
  AND U7252 ( .A(n802), .B(n4177), .Z(n4175) );
  XOR U7253 ( .A(n4178), .B(n4179), .Z(n4177) );
  XOR U7254 ( .A(DB[2181]), .B(DB[2174]), .Z(n4179) );
  AND U7255 ( .A(n806), .B(n4180), .Z(n4178) );
  XOR U7256 ( .A(n4181), .B(n4182), .Z(n4180) );
  XOR U7257 ( .A(DB[2174]), .B(DB[2167]), .Z(n4182) );
  AND U7258 ( .A(n810), .B(n4183), .Z(n4181) );
  XOR U7259 ( .A(n4184), .B(n4185), .Z(n4183) );
  XOR U7260 ( .A(DB[2167]), .B(DB[2160]), .Z(n4185) );
  AND U7261 ( .A(n814), .B(n4186), .Z(n4184) );
  XOR U7262 ( .A(n4187), .B(n4188), .Z(n4186) );
  XOR U7263 ( .A(DB[2160]), .B(DB[2153]), .Z(n4188) );
  AND U7264 ( .A(n818), .B(n4189), .Z(n4187) );
  XOR U7265 ( .A(n4190), .B(n4191), .Z(n4189) );
  XOR U7266 ( .A(DB[2153]), .B(DB[2146]), .Z(n4191) );
  AND U7267 ( .A(n822), .B(n4192), .Z(n4190) );
  XOR U7268 ( .A(n4193), .B(n4194), .Z(n4192) );
  XOR U7269 ( .A(DB[2146]), .B(DB[2139]), .Z(n4194) );
  AND U7270 ( .A(n826), .B(n4195), .Z(n4193) );
  XOR U7271 ( .A(n4196), .B(n4197), .Z(n4195) );
  XOR U7272 ( .A(DB[2139]), .B(DB[2132]), .Z(n4197) );
  AND U7273 ( .A(n830), .B(n4198), .Z(n4196) );
  XOR U7274 ( .A(n4199), .B(n4200), .Z(n4198) );
  XOR U7275 ( .A(DB[2132]), .B(DB[2125]), .Z(n4200) );
  AND U7276 ( .A(n834), .B(n4201), .Z(n4199) );
  XOR U7277 ( .A(n4202), .B(n4203), .Z(n4201) );
  XOR U7278 ( .A(DB[2125]), .B(DB[2118]), .Z(n4203) );
  AND U7279 ( .A(n838), .B(n4204), .Z(n4202) );
  XOR U7280 ( .A(n4205), .B(n4206), .Z(n4204) );
  XOR U7281 ( .A(DB[2118]), .B(DB[2111]), .Z(n4206) );
  AND U7282 ( .A(n842), .B(n4207), .Z(n4205) );
  XOR U7283 ( .A(n4208), .B(n4209), .Z(n4207) );
  XOR U7284 ( .A(DB[2111]), .B(DB[2104]), .Z(n4209) );
  AND U7285 ( .A(n846), .B(n4210), .Z(n4208) );
  XOR U7286 ( .A(n4211), .B(n4212), .Z(n4210) );
  XOR U7287 ( .A(DB[2104]), .B(DB[2097]), .Z(n4212) );
  AND U7288 ( .A(n850), .B(n4213), .Z(n4211) );
  XOR U7289 ( .A(n4214), .B(n4215), .Z(n4213) );
  XOR U7290 ( .A(DB[2097]), .B(DB[2090]), .Z(n4215) );
  AND U7291 ( .A(n854), .B(n4216), .Z(n4214) );
  XOR U7292 ( .A(n4217), .B(n4218), .Z(n4216) );
  XOR U7293 ( .A(DB[2090]), .B(DB[2083]), .Z(n4218) );
  AND U7294 ( .A(n858), .B(n4219), .Z(n4217) );
  XOR U7295 ( .A(n4220), .B(n4221), .Z(n4219) );
  XOR U7296 ( .A(DB[2083]), .B(DB[2076]), .Z(n4221) );
  AND U7297 ( .A(n862), .B(n4222), .Z(n4220) );
  XOR U7298 ( .A(n4223), .B(n4224), .Z(n4222) );
  XOR U7299 ( .A(DB[2076]), .B(DB[2069]), .Z(n4224) );
  AND U7300 ( .A(n866), .B(n4225), .Z(n4223) );
  XOR U7301 ( .A(n4226), .B(n4227), .Z(n4225) );
  XOR U7302 ( .A(DB[2069]), .B(DB[2062]), .Z(n4227) );
  AND U7303 ( .A(n870), .B(n4228), .Z(n4226) );
  XOR U7304 ( .A(n4229), .B(n4230), .Z(n4228) );
  XOR U7305 ( .A(DB[2062]), .B(DB[2055]), .Z(n4230) );
  AND U7306 ( .A(n874), .B(n4231), .Z(n4229) );
  XOR U7307 ( .A(n4232), .B(n4233), .Z(n4231) );
  XOR U7308 ( .A(DB[2055]), .B(DB[2048]), .Z(n4233) );
  AND U7309 ( .A(n878), .B(n4234), .Z(n4232) );
  XOR U7310 ( .A(n4235), .B(n4236), .Z(n4234) );
  XOR U7311 ( .A(DB[2048]), .B(DB[2041]), .Z(n4236) );
  AND U7312 ( .A(n882), .B(n4237), .Z(n4235) );
  XOR U7313 ( .A(n4238), .B(n4239), .Z(n4237) );
  XOR U7314 ( .A(DB[2041]), .B(DB[2034]), .Z(n4239) );
  AND U7315 ( .A(n886), .B(n4240), .Z(n4238) );
  XOR U7316 ( .A(n4241), .B(n4242), .Z(n4240) );
  XOR U7317 ( .A(DB[2034]), .B(DB[2027]), .Z(n4242) );
  AND U7318 ( .A(n890), .B(n4243), .Z(n4241) );
  XOR U7319 ( .A(n4244), .B(n4245), .Z(n4243) );
  XOR U7320 ( .A(DB[2027]), .B(DB[2020]), .Z(n4245) );
  AND U7321 ( .A(n894), .B(n4246), .Z(n4244) );
  XOR U7322 ( .A(n4247), .B(n4248), .Z(n4246) );
  XOR U7323 ( .A(DB[2020]), .B(DB[2013]), .Z(n4248) );
  AND U7324 ( .A(n898), .B(n4249), .Z(n4247) );
  XOR U7325 ( .A(n4250), .B(n4251), .Z(n4249) );
  XOR U7326 ( .A(DB[2013]), .B(DB[2006]), .Z(n4251) );
  AND U7327 ( .A(n902), .B(n4252), .Z(n4250) );
  XOR U7328 ( .A(n4253), .B(n4254), .Z(n4252) );
  XOR U7329 ( .A(DB[2006]), .B(DB[1999]), .Z(n4254) );
  AND U7330 ( .A(n906), .B(n4255), .Z(n4253) );
  XOR U7331 ( .A(n4256), .B(n4257), .Z(n4255) );
  XOR U7332 ( .A(DB[1999]), .B(DB[1992]), .Z(n4257) );
  AND U7333 ( .A(n910), .B(n4258), .Z(n4256) );
  XOR U7334 ( .A(n4259), .B(n4260), .Z(n4258) );
  XOR U7335 ( .A(DB[1992]), .B(DB[1985]), .Z(n4260) );
  AND U7336 ( .A(n914), .B(n4261), .Z(n4259) );
  XOR U7337 ( .A(n4262), .B(n4263), .Z(n4261) );
  XOR U7338 ( .A(DB[1985]), .B(DB[1978]), .Z(n4263) );
  AND U7339 ( .A(n918), .B(n4264), .Z(n4262) );
  XOR U7340 ( .A(n4265), .B(n4266), .Z(n4264) );
  XOR U7341 ( .A(DB[1978]), .B(DB[1971]), .Z(n4266) );
  AND U7342 ( .A(n922), .B(n4267), .Z(n4265) );
  XOR U7343 ( .A(n4268), .B(n4269), .Z(n4267) );
  XOR U7344 ( .A(DB[1971]), .B(DB[1964]), .Z(n4269) );
  AND U7345 ( .A(n926), .B(n4270), .Z(n4268) );
  XOR U7346 ( .A(n4271), .B(n4272), .Z(n4270) );
  XOR U7347 ( .A(DB[1964]), .B(DB[1957]), .Z(n4272) );
  AND U7348 ( .A(n930), .B(n4273), .Z(n4271) );
  XOR U7349 ( .A(n4274), .B(n4275), .Z(n4273) );
  XOR U7350 ( .A(DB[1957]), .B(DB[1950]), .Z(n4275) );
  AND U7351 ( .A(n934), .B(n4276), .Z(n4274) );
  XOR U7352 ( .A(n4277), .B(n4278), .Z(n4276) );
  XOR U7353 ( .A(DB[1950]), .B(DB[1943]), .Z(n4278) );
  AND U7354 ( .A(n938), .B(n4279), .Z(n4277) );
  XOR U7355 ( .A(n4280), .B(n4281), .Z(n4279) );
  XOR U7356 ( .A(DB[1943]), .B(DB[1936]), .Z(n4281) );
  AND U7357 ( .A(n942), .B(n4282), .Z(n4280) );
  XOR U7358 ( .A(n4283), .B(n4284), .Z(n4282) );
  XOR U7359 ( .A(DB[1936]), .B(DB[1929]), .Z(n4284) );
  AND U7360 ( .A(n946), .B(n4285), .Z(n4283) );
  XOR U7361 ( .A(n4286), .B(n4287), .Z(n4285) );
  XOR U7362 ( .A(DB[1929]), .B(DB[1922]), .Z(n4287) );
  AND U7363 ( .A(n950), .B(n4288), .Z(n4286) );
  XOR U7364 ( .A(n4289), .B(n4290), .Z(n4288) );
  XOR U7365 ( .A(DB[1922]), .B(DB[1915]), .Z(n4290) );
  AND U7366 ( .A(n954), .B(n4291), .Z(n4289) );
  XOR U7367 ( .A(n4292), .B(n4293), .Z(n4291) );
  XOR U7368 ( .A(DB[1915]), .B(DB[1908]), .Z(n4293) );
  AND U7369 ( .A(n958), .B(n4294), .Z(n4292) );
  XOR U7370 ( .A(n4295), .B(n4296), .Z(n4294) );
  XOR U7371 ( .A(DB[1908]), .B(DB[1901]), .Z(n4296) );
  AND U7372 ( .A(n962), .B(n4297), .Z(n4295) );
  XOR U7373 ( .A(n4298), .B(n4299), .Z(n4297) );
  XOR U7374 ( .A(DB[1901]), .B(DB[1894]), .Z(n4299) );
  AND U7375 ( .A(n966), .B(n4300), .Z(n4298) );
  XOR U7376 ( .A(n4301), .B(n4302), .Z(n4300) );
  XOR U7377 ( .A(DB[1894]), .B(DB[1887]), .Z(n4302) );
  AND U7378 ( .A(n970), .B(n4303), .Z(n4301) );
  XOR U7379 ( .A(n4304), .B(n4305), .Z(n4303) );
  XOR U7380 ( .A(DB[1887]), .B(DB[1880]), .Z(n4305) );
  AND U7381 ( .A(n974), .B(n4306), .Z(n4304) );
  XOR U7382 ( .A(n4307), .B(n4308), .Z(n4306) );
  XOR U7383 ( .A(DB[1880]), .B(DB[1873]), .Z(n4308) );
  AND U7384 ( .A(n978), .B(n4309), .Z(n4307) );
  XOR U7385 ( .A(n4310), .B(n4311), .Z(n4309) );
  XOR U7386 ( .A(DB[1873]), .B(DB[1866]), .Z(n4311) );
  AND U7387 ( .A(n982), .B(n4312), .Z(n4310) );
  XOR U7388 ( .A(n4313), .B(n4314), .Z(n4312) );
  XOR U7389 ( .A(DB[1866]), .B(DB[1859]), .Z(n4314) );
  AND U7390 ( .A(n986), .B(n4315), .Z(n4313) );
  XOR U7391 ( .A(n4316), .B(n4317), .Z(n4315) );
  XOR U7392 ( .A(DB[1859]), .B(DB[1852]), .Z(n4317) );
  AND U7393 ( .A(n990), .B(n4318), .Z(n4316) );
  XOR U7394 ( .A(n4319), .B(n4320), .Z(n4318) );
  XOR U7395 ( .A(DB[1852]), .B(DB[1845]), .Z(n4320) );
  AND U7396 ( .A(n994), .B(n4321), .Z(n4319) );
  XOR U7397 ( .A(n4322), .B(n4323), .Z(n4321) );
  XOR U7398 ( .A(DB[1845]), .B(DB[1838]), .Z(n4323) );
  AND U7399 ( .A(n998), .B(n4324), .Z(n4322) );
  XOR U7400 ( .A(n4325), .B(n4326), .Z(n4324) );
  XOR U7401 ( .A(DB[1838]), .B(DB[1831]), .Z(n4326) );
  AND U7402 ( .A(n1002), .B(n4327), .Z(n4325) );
  XOR U7403 ( .A(n4328), .B(n4329), .Z(n4327) );
  XOR U7404 ( .A(DB[1831]), .B(DB[1824]), .Z(n4329) );
  AND U7405 ( .A(n1006), .B(n4330), .Z(n4328) );
  XOR U7406 ( .A(n4331), .B(n4332), .Z(n4330) );
  XOR U7407 ( .A(DB[1824]), .B(DB[1817]), .Z(n4332) );
  AND U7408 ( .A(n1010), .B(n4333), .Z(n4331) );
  XOR U7409 ( .A(n4334), .B(n4335), .Z(n4333) );
  XOR U7410 ( .A(DB[1817]), .B(DB[1810]), .Z(n4335) );
  AND U7411 ( .A(n1014), .B(n4336), .Z(n4334) );
  XOR U7412 ( .A(n4337), .B(n4338), .Z(n4336) );
  XOR U7413 ( .A(DB[1810]), .B(DB[1803]), .Z(n4338) );
  AND U7414 ( .A(n1018), .B(n4339), .Z(n4337) );
  XOR U7415 ( .A(n4340), .B(n4341), .Z(n4339) );
  XOR U7416 ( .A(DB[1803]), .B(DB[1796]), .Z(n4341) );
  AND U7417 ( .A(n1022), .B(n4342), .Z(n4340) );
  XOR U7418 ( .A(n4343), .B(n4344), .Z(n4342) );
  XOR U7419 ( .A(DB[1796]), .B(DB[1789]), .Z(n4344) );
  AND U7420 ( .A(n1026), .B(n4345), .Z(n4343) );
  XOR U7421 ( .A(n4346), .B(n4347), .Z(n4345) );
  XOR U7422 ( .A(DB[1789]), .B(DB[1782]), .Z(n4347) );
  AND U7423 ( .A(n1030), .B(n4348), .Z(n4346) );
  XOR U7424 ( .A(n4349), .B(n4350), .Z(n4348) );
  XOR U7425 ( .A(DB[1782]), .B(DB[1775]), .Z(n4350) );
  AND U7426 ( .A(n1034), .B(n4351), .Z(n4349) );
  XOR U7427 ( .A(n4352), .B(n4353), .Z(n4351) );
  XOR U7428 ( .A(DB[1775]), .B(DB[1768]), .Z(n4353) );
  AND U7429 ( .A(n1038), .B(n4354), .Z(n4352) );
  XOR U7430 ( .A(n4355), .B(n4356), .Z(n4354) );
  XOR U7431 ( .A(DB[1768]), .B(DB[1761]), .Z(n4356) );
  AND U7432 ( .A(n1042), .B(n4357), .Z(n4355) );
  XOR U7433 ( .A(n4358), .B(n4359), .Z(n4357) );
  XOR U7434 ( .A(DB[1761]), .B(DB[1754]), .Z(n4359) );
  AND U7435 ( .A(n1046), .B(n4360), .Z(n4358) );
  XOR U7436 ( .A(n4361), .B(n4362), .Z(n4360) );
  XOR U7437 ( .A(DB[1754]), .B(DB[1747]), .Z(n4362) );
  AND U7438 ( .A(n1050), .B(n4363), .Z(n4361) );
  XOR U7439 ( .A(n4364), .B(n4365), .Z(n4363) );
  XOR U7440 ( .A(DB[1747]), .B(DB[1740]), .Z(n4365) );
  AND U7441 ( .A(n1054), .B(n4366), .Z(n4364) );
  XOR U7442 ( .A(n4367), .B(n4368), .Z(n4366) );
  XOR U7443 ( .A(DB[1740]), .B(DB[1733]), .Z(n4368) );
  AND U7444 ( .A(n1058), .B(n4369), .Z(n4367) );
  XOR U7445 ( .A(n4370), .B(n4371), .Z(n4369) );
  XOR U7446 ( .A(DB[1733]), .B(DB[1726]), .Z(n4371) );
  AND U7447 ( .A(n1062), .B(n4372), .Z(n4370) );
  XOR U7448 ( .A(n4373), .B(n4374), .Z(n4372) );
  XOR U7449 ( .A(DB[1726]), .B(DB[1719]), .Z(n4374) );
  AND U7450 ( .A(n1066), .B(n4375), .Z(n4373) );
  XOR U7451 ( .A(n4376), .B(n4377), .Z(n4375) );
  XOR U7452 ( .A(DB[1719]), .B(DB[1712]), .Z(n4377) );
  AND U7453 ( .A(n1070), .B(n4378), .Z(n4376) );
  XOR U7454 ( .A(n4379), .B(n4380), .Z(n4378) );
  XOR U7455 ( .A(DB[1712]), .B(DB[1705]), .Z(n4380) );
  AND U7456 ( .A(n1074), .B(n4381), .Z(n4379) );
  XOR U7457 ( .A(n4382), .B(n4383), .Z(n4381) );
  XOR U7458 ( .A(DB[1705]), .B(DB[1698]), .Z(n4383) );
  AND U7459 ( .A(n1078), .B(n4384), .Z(n4382) );
  XOR U7460 ( .A(n4385), .B(n4386), .Z(n4384) );
  XOR U7461 ( .A(DB[1698]), .B(DB[1691]), .Z(n4386) );
  AND U7462 ( .A(n1082), .B(n4387), .Z(n4385) );
  XOR U7463 ( .A(n4388), .B(n4389), .Z(n4387) );
  XOR U7464 ( .A(DB[1691]), .B(DB[1684]), .Z(n4389) );
  AND U7465 ( .A(n1086), .B(n4390), .Z(n4388) );
  XOR U7466 ( .A(n4391), .B(n4392), .Z(n4390) );
  XOR U7467 ( .A(DB[1684]), .B(DB[1677]), .Z(n4392) );
  AND U7468 ( .A(n1090), .B(n4393), .Z(n4391) );
  XOR U7469 ( .A(n4394), .B(n4395), .Z(n4393) );
  XOR U7470 ( .A(DB[1677]), .B(DB[1670]), .Z(n4395) );
  AND U7471 ( .A(n1094), .B(n4396), .Z(n4394) );
  XOR U7472 ( .A(n4397), .B(n4398), .Z(n4396) );
  XOR U7473 ( .A(DB[1670]), .B(DB[1663]), .Z(n4398) );
  AND U7474 ( .A(n1098), .B(n4399), .Z(n4397) );
  XOR U7475 ( .A(n4400), .B(n4401), .Z(n4399) );
  XOR U7476 ( .A(DB[1663]), .B(DB[1656]), .Z(n4401) );
  AND U7477 ( .A(n1102), .B(n4402), .Z(n4400) );
  XOR U7478 ( .A(n4403), .B(n4404), .Z(n4402) );
  XOR U7479 ( .A(DB[1656]), .B(DB[1649]), .Z(n4404) );
  AND U7480 ( .A(n1106), .B(n4405), .Z(n4403) );
  XOR U7481 ( .A(n4406), .B(n4407), .Z(n4405) );
  XOR U7482 ( .A(DB[1649]), .B(DB[1642]), .Z(n4407) );
  AND U7483 ( .A(n1110), .B(n4408), .Z(n4406) );
  XOR U7484 ( .A(n4409), .B(n4410), .Z(n4408) );
  XOR U7485 ( .A(DB[1642]), .B(DB[1635]), .Z(n4410) );
  AND U7486 ( .A(n1114), .B(n4411), .Z(n4409) );
  XOR U7487 ( .A(n4412), .B(n4413), .Z(n4411) );
  XOR U7488 ( .A(DB[1635]), .B(DB[1628]), .Z(n4413) );
  AND U7489 ( .A(n1118), .B(n4414), .Z(n4412) );
  XOR U7490 ( .A(n4415), .B(n4416), .Z(n4414) );
  XOR U7491 ( .A(DB[1628]), .B(DB[1621]), .Z(n4416) );
  AND U7492 ( .A(n1122), .B(n4417), .Z(n4415) );
  XOR U7493 ( .A(n4418), .B(n4419), .Z(n4417) );
  XOR U7494 ( .A(DB[1621]), .B(DB[1614]), .Z(n4419) );
  AND U7495 ( .A(n1126), .B(n4420), .Z(n4418) );
  XOR U7496 ( .A(n4421), .B(n4422), .Z(n4420) );
  XOR U7497 ( .A(DB[1614]), .B(DB[1607]), .Z(n4422) );
  AND U7498 ( .A(n1130), .B(n4423), .Z(n4421) );
  XOR U7499 ( .A(n4424), .B(n4425), .Z(n4423) );
  XOR U7500 ( .A(DB[1607]), .B(DB[1600]), .Z(n4425) );
  AND U7501 ( .A(n1134), .B(n4426), .Z(n4424) );
  XOR U7502 ( .A(n4427), .B(n4428), .Z(n4426) );
  XOR U7503 ( .A(DB[1600]), .B(DB[1593]), .Z(n4428) );
  AND U7504 ( .A(n1138), .B(n4429), .Z(n4427) );
  XOR U7505 ( .A(n4430), .B(n4431), .Z(n4429) );
  XOR U7506 ( .A(DB[1593]), .B(DB[1586]), .Z(n4431) );
  AND U7507 ( .A(n1142), .B(n4432), .Z(n4430) );
  XOR U7508 ( .A(n4433), .B(n4434), .Z(n4432) );
  XOR U7509 ( .A(DB[1586]), .B(DB[1579]), .Z(n4434) );
  AND U7510 ( .A(n1146), .B(n4435), .Z(n4433) );
  XOR U7511 ( .A(n4436), .B(n4437), .Z(n4435) );
  XOR U7512 ( .A(DB[1579]), .B(DB[1572]), .Z(n4437) );
  AND U7513 ( .A(n1150), .B(n4438), .Z(n4436) );
  XOR U7514 ( .A(n4439), .B(n4440), .Z(n4438) );
  XOR U7515 ( .A(DB[1572]), .B(DB[1565]), .Z(n4440) );
  AND U7516 ( .A(n1154), .B(n4441), .Z(n4439) );
  XOR U7517 ( .A(n4442), .B(n4443), .Z(n4441) );
  XOR U7518 ( .A(DB[1565]), .B(DB[1558]), .Z(n4443) );
  AND U7519 ( .A(n1158), .B(n4444), .Z(n4442) );
  XOR U7520 ( .A(n4445), .B(n4446), .Z(n4444) );
  XOR U7521 ( .A(DB[1558]), .B(DB[1551]), .Z(n4446) );
  AND U7522 ( .A(n1162), .B(n4447), .Z(n4445) );
  XOR U7523 ( .A(n4448), .B(n4449), .Z(n4447) );
  XOR U7524 ( .A(DB[1551]), .B(DB[1544]), .Z(n4449) );
  AND U7525 ( .A(n1166), .B(n4450), .Z(n4448) );
  XOR U7526 ( .A(n4451), .B(n4452), .Z(n4450) );
  XOR U7527 ( .A(DB[1544]), .B(DB[1537]), .Z(n4452) );
  AND U7528 ( .A(n1170), .B(n4453), .Z(n4451) );
  XOR U7529 ( .A(n4454), .B(n4455), .Z(n4453) );
  XOR U7530 ( .A(DB[1537]), .B(DB[1530]), .Z(n4455) );
  AND U7531 ( .A(n1174), .B(n4456), .Z(n4454) );
  XOR U7532 ( .A(n4457), .B(n4458), .Z(n4456) );
  XOR U7533 ( .A(DB[1530]), .B(DB[1523]), .Z(n4458) );
  AND U7534 ( .A(n1178), .B(n4459), .Z(n4457) );
  XOR U7535 ( .A(n4460), .B(n4461), .Z(n4459) );
  XOR U7536 ( .A(DB[1523]), .B(DB[1516]), .Z(n4461) );
  AND U7537 ( .A(n1182), .B(n4462), .Z(n4460) );
  XOR U7538 ( .A(n4463), .B(n4464), .Z(n4462) );
  XOR U7539 ( .A(DB[1516]), .B(DB[1509]), .Z(n4464) );
  AND U7540 ( .A(n1186), .B(n4465), .Z(n4463) );
  XOR U7541 ( .A(n4466), .B(n4467), .Z(n4465) );
  XOR U7542 ( .A(DB[1509]), .B(DB[1502]), .Z(n4467) );
  AND U7543 ( .A(n1190), .B(n4468), .Z(n4466) );
  XOR U7544 ( .A(n4469), .B(n4470), .Z(n4468) );
  XOR U7545 ( .A(DB[1502]), .B(DB[1495]), .Z(n4470) );
  AND U7546 ( .A(n1194), .B(n4471), .Z(n4469) );
  XOR U7547 ( .A(n4472), .B(n4473), .Z(n4471) );
  XOR U7548 ( .A(DB[1495]), .B(DB[1488]), .Z(n4473) );
  AND U7549 ( .A(n1198), .B(n4474), .Z(n4472) );
  XOR U7550 ( .A(n4475), .B(n4476), .Z(n4474) );
  XOR U7551 ( .A(DB[1488]), .B(DB[1481]), .Z(n4476) );
  AND U7552 ( .A(n1202), .B(n4477), .Z(n4475) );
  XOR U7553 ( .A(n4478), .B(n4479), .Z(n4477) );
  XOR U7554 ( .A(DB[1481]), .B(DB[1474]), .Z(n4479) );
  AND U7555 ( .A(n1206), .B(n4480), .Z(n4478) );
  XOR U7556 ( .A(n4481), .B(n4482), .Z(n4480) );
  XOR U7557 ( .A(DB[1474]), .B(DB[1467]), .Z(n4482) );
  AND U7558 ( .A(n1210), .B(n4483), .Z(n4481) );
  XOR U7559 ( .A(n4484), .B(n4485), .Z(n4483) );
  XOR U7560 ( .A(DB[1467]), .B(DB[1460]), .Z(n4485) );
  AND U7561 ( .A(n1214), .B(n4486), .Z(n4484) );
  XOR U7562 ( .A(n4487), .B(n4488), .Z(n4486) );
  XOR U7563 ( .A(DB[1460]), .B(DB[1453]), .Z(n4488) );
  AND U7564 ( .A(n1218), .B(n4489), .Z(n4487) );
  XOR U7565 ( .A(n4490), .B(n4491), .Z(n4489) );
  XOR U7566 ( .A(DB[1453]), .B(DB[1446]), .Z(n4491) );
  AND U7567 ( .A(n1222), .B(n4492), .Z(n4490) );
  XOR U7568 ( .A(n4493), .B(n4494), .Z(n4492) );
  XOR U7569 ( .A(DB[1446]), .B(DB[1439]), .Z(n4494) );
  AND U7570 ( .A(n1226), .B(n4495), .Z(n4493) );
  XOR U7571 ( .A(n4496), .B(n4497), .Z(n4495) );
  XOR U7572 ( .A(DB[1439]), .B(DB[1432]), .Z(n4497) );
  AND U7573 ( .A(n1230), .B(n4498), .Z(n4496) );
  XOR U7574 ( .A(n4499), .B(n4500), .Z(n4498) );
  XOR U7575 ( .A(DB[1432]), .B(DB[1425]), .Z(n4500) );
  AND U7576 ( .A(n1234), .B(n4501), .Z(n4499) );
  XOR U7577 ( .A(n4502), .B(n4503), .Z(n4501) );
  XOR U7578 ( .A(DB[1425]), .B(DB[1418]), .Z(n4503) );
  AND U7579 ( .A(n1238), .B(n4504), .Z(n4502) );
  XOR U7580 ( .A(n4505), .B(n4506), .Z(n4504) );
  XOR U7581 ( .A(DB[1418]), .B(DB[1411]), .Z(n4506) );
  AND U7582 ( .A(n1242), .B(n4507), .Z(n4505) );
  XOR U7583 ( .A(n4508), .B(n4509), .Z(n4507) );
  XOR U7584 ( .A(DB[1411]), .B(DB[1404]), .Z(n4509) );
  AND U7585 ( .A(n1246), .B(n4510), .Z(n4508) );
  XOR U7586 ( .A(n4511), .B(n4512), .Z(n4510) );
  XOR U7587 ( .A(DB[1404]), .B(DB[1397]), .Z(n4512) );
  AND U7588 ( .A(n1250), .B(n4513), .Z(n4511) );
  XOR U7589 ( .A(n4514), .B(n4515), .Z(n4513) );
  XOR U7590 ( .A(DB[1397]), .B(DB[1390]), .Z(n4515) );
  AND U7591 ( .A(n1254), .B(n4516), .Z(n4514) );
  XOR U7592 ( .A(n4517), .B(n4518), .Z(n4516) );
  XOR U7593 ( .A(DB[1390]), .B(DB[1383]), .Z(n4518) );
  AND U7594 ( .A(n1258), .B(n4519), .Z(n4517) );
  XOR U7595 ( .A(n4520), .B(n4521), .Z(n4519) );
  XOR U7596 ( .A(DB[1383]), .B(DB[1376]), .Z(n4521) );
  AND U7597 ( .A(n1262), .B(n4522), .Z(n4520) );
  XOR U7598 ( .A(n4523), .B(n4524), .Z(n4522) );
  XOR U7599 ( .A(DB[1376]), .B(DB[1369]), .Z(n4524) );
  AND U7600 ( .A(n1266), .B(n4525), .Z(n4523) );
  XOR U7601 ( .A(n4526), .B(n4527), .Z(n4525) );
  XOR U7602 ( .A(DB[1369]), .B(DB[1362]), .Z(n4527) );
  AND U7603 ( .A(n1270), .B(n4528), .Z(n4526) );
  XOR U7604 ( .A(n4529), .B(n4530), .Z(n4528) );
  XOR U7605 ( .A(DB[1362]), .B(DB[1355]), .Z(n4530) );
  AND U7606 ( .A(n1274), .B(n4531), .Z(n4529) );
  XOR U7607 ( .A(n4532), .B(n4533), .Z(n4531) );
  XOR U7608 ( .A(DB[1355]), .B(DB[1348]), .Z(n4533) );
  AND U7609 ( .A(n1278), .B(n4534), .Z(n4532) );
  XOR U7610 ( .A(n4535), .B(n4536), .Z(n4534) );
  XOR U7611 ( .A(DB[1348]), .B(DB[1341]), .Z(n4536) );
  AND U7612 ( .A(n1282), .B(n4537), .Z(n4535) );
  XOR U7613 ( .A(n4538), .B(n4539), .Z(n4537) );
  XOR U7614 ( .A(DB[1341]), .B(DB[1334]), .Z(n4539) );
  AND U7615 ( .A(n1286), .B(n4540), .Z(n4538) );
  XOR U7616 ( .A(n4541), .B(n4542), .Z(n4540) );
  XOR U7617 ( .A(DB[1334]), .B(DB[1327]), .Z(n4542) );
  AND U7618 ( .A(n1290), .B(n4543), .Z(n4541) );
  XOR U7619 ( .A(n4544), .B(n4545), .Z(n4543) );
  XOR U7620 ( .A(DB[1327]), .B(DB[1320]), .Z(n4545) );
  AND U7621 ( .A(n1294), .B(n4546), .Z(n4544) );
  XOR U7622 ( .A(n4547), .B(n4548), .Z(n4546) );
  XOR U7623 ( .A(DB[1320]), .B(DB[1313]), .Z(n4548) );
  AND U7624 ( .A(n1298), .B(n4549), .Z(n4547) );
  XOR U7625 ( .A(n4550), .B(n4551), .Z(n4549) );
  XOR U7626 ( .A(DB[1313]), .B(DB[1306]), .Z(n4551) );
  AND U7627 ( .A(n1302), .B(n4552), .Z(n4550) );
  XOR U7628 ( .A(n4553), .B(n4554), .Z(n4552) );
  XOR U7629 ( .A(DB[1306]), .B(DB[1299]), .Z(n4554) );
  AND U7630 ( .A(n1306), .B(n4555), .Z(n4553) );
  XOR U7631 ( .A(n4556), .B(n4557), .Z(n4555) );
  XOR U7632 ( .A(DB[1299]), .B(DB[1292]), .Z(n4557) );
  AND U7633 ( .A(n1310), .B(n4558), .Z(n4556) );
  XOR U7634 ( .A(n4559), .B(n4560), .Z(n4558) );
  XOR U7635 ( .A(DB[1292]), .B(DB[1285]), .Z(n4560) );
  AND U7636 ( .A(n1314), .B(n4561), .Z(n4559) );
  XOR U7637 ( .A(n4562), .B(n4563), .Z(n4561) );
  XOR U7638 ( .A(DB[1285]), .B(DB[1278]), .Z(n4563) );
  AND U7639 ( .A(n1318), .B(n4564), .Z(n4562) );
  XOR U7640 ( .A(n4565), .B(n4566), .Z(n4564) );
  XOR U7641 ( .A(DB[1278]), .B(DB[1271]), .Z(n4566) );
  AND U7642 ( .A(n1322), .B(n4567), .Z(n4565) );
  XOR U7643 ( .A(n4568), .B(n4569), .Z(n4567) );
  XOR U7644 ( .A(DB[1271]), .B(DB[1264]), .Z(n4569) );
  AND U7645 ( .A(n1326), .B(n4570), .Z(n4568) );
  XOR U7646 ( .A(n4571), .B(n4572), .Z(n4570) );
  XOR U7647 ( .A(DB[1264]), .B(DB[1257]), .Z(n4572) );
  AND U7648 ( .A(n1330), .B(n4573), .Z(n4571) );
  XOR U7649 ( .A(n4574), .B(n4575), .Z(n4573) );
  XOR U7650 ( .A(DB[1257]), .B(DB[1250]), .Z(n4575) );
  AND U7651 ( .A(n1334), .B(n4576), .Z(n4574) );
  XOR U7652 ( .A(n4577), .B(n4578), .Z(n4576) );
  XOR U7653 ( .A(DB[1250]), .B(DB[1243]), .Z(n4578) );
  AND U7654 ( .A(n1338), .B(n4579), .Z(n4577) );
  XOR U7655 ( .A(n4580), .B(n4581), .Z(n4579) );
  XOR U7656 ( .A(DB[1243]), .B(DB[1236]), .Z(n4581) );
  AND U7657 ( .A(n1342), .B(n4582), .Z(n4580) );
  XOR U7658 ( .A(n4583), .B(n4584), .Z(n4582) );
  XOR U7659 ( .A(DB[1236]), .B(DB[1229]), .Z(n4584) );
  AND U7660 ( .A(n1346), .B(n4585), .Z(n4583) );
  XOR U7661 ( .A(n4586), .B(n4587), .Z(n4585) );
  XOR U7662 ( .A(DB[1229]), .B(DB[1222]), .Z(n4587) );
  AND U7663 ( .A(n1350), .B(n4588), .Z(n4586) );
  XOR U7664 ( .A(n4589), .B(n4590), .Z(n4588) );
  XOR U7665 ( .A(DB[1222]), .B(DB[1215]), .Z(n4590) );
  AND U7666 ( .A(n1354), .B(n4591), .Z(n4589) );
  XOR U7667 ( .A(n4592), .B(n4593), .Z(n4591) );
  XOR U7668 ( .A(DB[1215]), .B(DB[1208]), .Z(n4593) );
  AND U7669 ( .A(n1358), .B(n4594), .Z(n4592) );
  XOR U7670 ( .A(n4595), .B(n4596), .Z(n4594) );
  XOR U7671 ( .A(DB[1208]), .B(DB[1201]), .Z(n4596) );
  AND U7672 ( .A(n1362), .B(n4597), .Z(n4595) );
  XOR U7673 ( .A(n4598), .B(n4599), .Z(n4597) );
  XOR U7674 ( .A(DB[1201]), .B(DB[1194]), .Z(n4599) );
  AND U7675 ( .A(n1366), .B(n4600), .Z(n4598) );
  XOR U7676 ( .A(n4601), .B(n4602), .Z(n4600) );
  XOR U7677 ( .A(DB[1194]), .B(DB[1187]), .Z(n4602) );
  AND U7678 ( .A(n1370), .B(n4603), .Z(n4601) );
  XOR U7679 ( .A(n4604), .B(n4605), .Z(n4603) );
  XOR U7680 ( .A(DB[1187]), .B(DB[1180]), .Z(n4605) );
  AND U7681 ( .A(n1374), .B(n4606), .Z(n4604) );
  XOR U7682 ( .A(n4607), .B(n4608), .Z(n4606) );
  XOR U7683 ( .A(DB[1180]), .B(DB[1173]), .Z(n4608) );
  AND U7684 ( .A(n1378), .B(n4609), .Z(n4607) );
  XOR U7685 ( .A(n4610), .B(n4611), .Z(n4609) );
  XOR U7686 ( .A(DB[1173]), .B(DB[1166]), .Z(n4611) );
  AND U7687 ( .A(n1382), .B(n4612), .Z(n4610) );
  XOR U7688 ( .A(n4613), .B(n4614), .Z(n4612) );
  XOR U7689 ( .A(DB[1166]), .B(DB[1159]), .Z(n4614) );
  AND U7690 ( .A(n1386), .B(n4615), .Z(n4613) );
  XOR U7691 ( .A(n4616), .B(n4617), .Z(n4615) );
  XOR U7692 ( .A(DB[1159]), .B(DB[1152]), .Z(n4617) );
  AND U7693 ( .A(n1390), .B(n4618), .Z(n4616) );
  XOR U7694 ( .A(n4619), .B(n4620), .Z(n4618) );
  XOR U7695 ( .A(DB[1152]), .B(DB[1145]), .Z(n4620) );
  AND U7696 ( .A(n1394), .B(n4621), .Z(n4619) );
  XOR U7697 ( .A(n4622), .B(n4623), .Z(n4621) );
  XOR U7698 ( .A(DB[1145]), .B(DB[1138]), .Z(n4623) );
  AND U7699 ( .A(n1398), .B(n4624), .Z(n4622) );
  XOR U7700 ( .A(n4625), .B(n4626), .Z(n4624) );
  XOR U7701 ( .A(DB[1138]), .B(DB[1131]), .Z(n4626) );
  AND U7702 ( .A(n1402), .B(n4627), .Z(n4625) );
  XOR U7703 ( .A(n4628), .B(n4629), .Z(n4627) );
  XOR U7704 ( .A(DB[1131]), .B(DB[1124]), .Z(n4629) );
  AND U7705 ( .A(n1406), .B(n4630), .Z(n4628) );
  XOR U7706 ( .A(n4631), .B(n4632), .Z(n4630) );
  XOR U7707 ( .A(DB[1124]), .B(DB[1117]), .Z(n4632) );
  AND U7708 ( .A(n1410), .B(n4633), .Z(n4631) );
  XOR U7709 ( .A(n4634), .B(n4635), .Z(n4633) );
  XOR U7710 ( .A(DB[1117]), .B(DB[1110]), .Z(n4635) );
  AND U7711 ( .A(n1414), .B(n4636), .Z(n4634) );
  XOR U7712 ( .A(n4637), .B(n4638), .Z(n4636) );
  XOR U7713 ( .A(DB[1110]), .B(DB[1103]), .Z(n4638) );
  AND U7714 ( .A(n1418), .B(n4639), .Z(n4637) );
  XOR U7715 ( .A(n4640), .B(n4641), .Z(n4639) );
  XOR U7716 ( .A(DB[1103]), .B(DB[1096]), .Z(n4641) );
  AND U7717 ( .A(n1422), .B(n4642), .Z(n4640) );
  XOR U7718 ( .A(n4643), .B(n4644), .Z(n4642) );
  XOR U7719 ( .A(DB[1096]), .B(DB[1089]), .Z(n4644) );
  AND U7720 ( .A(n1426), .B(n4645), .Z(n4643) );
  XOR U7721 ( .A(n4646), .B(n4647), .Z(n4645) );
  XOR U7722 ( .A(DB[1089]), .B(DB[1082]), .Z(n4647) );
  AND U7723 ( .A(n1430), .B(n4648), .Z(n4646) );
  XOR U7724 ( .A(n4649), .B(n4650), .Z(n4648) );
  XOR U7725 ( .A(DB[1082]), .B(DB[1075]), .Z(n4650) );
  AND U7726 ( .A(n1434), .B(n4651), .Z(n4649) );
  XOR U7727 ( .A(n4652), .B(n4653), .Z(n4651) );
  XOR U7728 ( .A(DB[1075]), .B(DB[1068]), .Z(n4653) );
  AND U7729 ( .A(n1438), .B(n4654), .Z(n4652) );
  XOR U7730 ( .A(n4655), .B(n4656), .Z(n4654) );
  XOR U7731 ( .A(DB[1068]), .B(DB[1061]), .Z(n4656) );
  AND U7732 ( .A(n1442), .B(n4657), .Z(n4655) );
  XOR U7733 ( .A(n4658), .B(n4659), .Z(n4657) );
  XOR U7734 ( .A(DB[1061]), .B(DB[1054]), .Z(n4659) );
  AND U7735 ( .A(n1446), .B(n4660), .Z(n4658) );
  XOR U7736 ( .A(n4661), .B(n4662), .Z(n4660) );
  XOR U7737 ( .A(DB[1054]), .B(DB[1047]), .Z(n4662) );
  AND U7738 ( .A(n1450), .B(n4663), .Z(n4661) );
  XOR U7739 ( .A(n4664), .B(n4665), .Z(n4663) );
  XOR U7740 ( .A(DB[1047]), .B(DB[1040]), .Z(n4665) );
  AND U7741 ( .A(n1454), .B(n4666), .Z(n4664) );
  XOR U7742 ( .A(n4667), .B(n4668), .Z(n4666) );
  XOR U7743 ( .A(DB[1040]), .B(DB[1033]), .Z(n4668) );
  AND U7744 ( .A(n1458), .B(n4669), .Z(n4667) );
  XOR U7745 ( .A(n4670), .B(n4671), .Z(n4669) );
  XOR U7746 ( .A(DB[1033]), .B(DB[1026]), .Z(n4671) );
  AND U7747 ( .A(n1462), .B(n4672), .Z(n4670) );
  XOR U7748 ( .A(n4673), .B(n4674), .Z(n4672) );
  XOR U7749 ( .A(DB[1026]), .B(DB[1019]), .Z(n4674) );
  AND U7750 ( .A(n1466), .B(n4675), .Z(n4673) );
  XOR U7751 ( .A(n4676), .B(n4677), .Z(n4675) );
  XOR U7752 ( .A(DB[1019]), .B(DB[1012]), .Z(n4677) );
  AND U7753 ( .A(n1470), .B(n4678), .Z(n4676) );
  XOR U7754 ( .A(n4679), .B(n4680), .Z(n4678) );
  XOR U7755 ( .A(DB[1012]), .B(DB[1005]), .Z(n4680) );
  AND U7756 ( .A(n1474), .B(n4681), .Z(n4679) );
  XOR U7757 ( .A(n4682), .B(n4683), .Z(n4681) );
  XOR U7758 ( .A(DB[998]), .B(DB[1005]), .Z(n4683) );
  AND U7759 ( .A(n1478), .B(n4684), .Z(n4682) );
  XOR U7760 ( .A(n4685), .B(n4686), .Z(n4684) );
  XOR U7761 ( .A(DB[998]), .B(DB[991]), .Z(n4686) );
  AND U7762 ( .A(n1482), .B(n4687), .Z(n4685) );
  XOR U7763 ( .A(n4688), .B(n4689), .Z(n4687) );
  XOR U7764 ( .A(DB[991]), .B(DB[984]), .Z(n4689) );
  AND U7765 ( .A(n1486), .B(n4690), .Z(n4688) );
  XOR U7766 ( .A(n4691), .B(n4692), .Z(n4690) );
  XOR U7767 ( .A(DB[984]), .B(DB[977]), .Z(n4692) );
  AND U7768 ( .A(n1490), .B(n4693), .Z(n4691) );
  XOR U7769 ( .A(n4694), .B(n4695), .Z(n4693) );
  XOR U7770 ( .A(DB[977]), .B(DB[970]), .Z(n4695) );
  AND U7771 ( .A(n1494), .B(n4696), .Z(n4694) );
  XOR U7772 ( .A(n4697), .B(n4698), .Z(n4696) );
  XOR U7773 ( .A(DB[970]), .B(DB[963]), .Z(n4698) );
  AND U7774 ( .A(n1498), .B(n4699), .Z(n4697) );
  XOR U7775 ( .A(n4700), .B(n4701), .Z(n4699) );
  XOR U7776 ( .A(DB[963]), .B(DB[956]), .Z(n4701) );
  AND U7777 ( .A(n1502), .B(n4702), .Z(n4700) );
  XOR U7778 ( .A(n4703), .B(n4704), .Z(n4702) );
  XOR U7779 ( .A(DB[956]), .B(DB[949]), .Z(n4704) );
  AND U7780 ( .A(n1506), .B(n4705), .Z(n4703) );
  XOR U7781 ( .A(n4706), .B(n4707), .Z(n4705) );
  XOR U7782 ( .A(DB[949]), .B(DB[942]), .Z(n4707) );
  AND U7783 ( .A(n1510), .B(n4708), .Z(n4706) );
  XOR U7784 ( .A(n4709), .B(n4710), .Z(n4708) );
  XOR U7785 ( .A(DB[942]), .B(DB[935]), .Z(n4710) );
  AND U7786 ( .A(n1514), .B(n4711), .Z(n4709) );
  XOR U7787 ( .A(n4712), .B(n4713), .Z(n4711) );
  XOR U7788 ( .A(DB[935]), .B(DB[928]), .Z(n4713) );
  AND U7789 ( .A(n1518), .B(n4714), .Z(n4712) );
  XOR U7790 ( .A(n4715), .B(n4716), .Z(n4714) );
  XOR U7791 ( .A(DB[928]), .B(DB[921]), .Z(n4716) );
  AND U7792 ( .A(n1522), .B(n4717), .Z(n4715) );
  XOR U7793 ( .A(n4718), .B(n4719), .Z(n4717) );
  XOR U7794 ( .A(DB[921]), .B(DB[914]), .Z(n4719) );
  AND U7795 ( .A(n1526), .B(n4720), .Z(n4718) );
  XOR U7796 ( .A(n4721), .B(n4722), .Z(n4720) );
  XOR U7797 ( .A(DB[914]), .B(DB[907]), .Z(n4722) );
  AND U7798 ( .A(n1530), .B(n4723), .Z(n4721) );
  XOR U7799 ( .A(n4724), .B(n4725), .Z(n4723) );
  XOR U7800 ( .A(DB[907]), .B(DB[900]), .Z(n4725) );
  AND U7801 ( .A(n1534), .B(n4726), .Z(n4724) );
  XOR U7802 ( .A(n4727), .B(n4728), .Z(n4726) );
  XOR U7803 ( .A(DB[900]), .B(DB[893]), .Z(n4728) );
  AND U7804 ( .A(n1538), .B(n4729), .Z(n4727) );
  XOR U7805 ( .A(n4730), .B(n4731), .Z(n4729) );
  XOR U7806 ( .A(DB[893]), .B(DB[886]), .Z(n4731) );
  AND U7807 ( .A(n1542), .B(n4732), .Z(n4730) );
  XOR U7808 ( .A(n4733), .B(n4734), .Z(n4732) );
  XOR U7809 ( .A(DB[886]), .B(DB[879]), .Z(n4734) );
  AND U7810 ( .A(n1546), .B(n4735), .Z(n4733) );
  XOR U7811 ( .A(n4736), .B(n4737), .Z(n4735) );
  XOR U7812 ( .A(DB[879]), .B(DB[872]), .Z(n4737) );
  AND U7813 ( .A(n1550), .B(n4738), .Z(n4736) );
  XOR U7814 ( .A(n4739), .B(n4740), .Z(n4738) );
  XOR U7815 ( .A(DB[872]), .B(DB[865]), .Z(n4740) );
  AND U7816 ( .A(n1554), .B(n4741), .Z(n4739) );
  XOR U7817 ( .A(n4742), .B(n4743), .Z(n4741) );
  XOR U7818 ( .A(DB[865]), .B(DB[858]), .Z(n4743) );
  AND U7819 ( .A(n1558), .B(n4744), .Z(n4742) );
  XOR U7820 ( .A(n4745), .B(n4746), .Z(n4744) );
  XOR U7821 ( .A(DB[858]), .B(DB[851]), .Z(n4746) );
  AND U7822 ( .A(n1562), .B(n4747), .Z(n4745) );
  XOR U7823 ( .A(n4748), .B(n4749), .Z(n4747) );
  XOR U7824 ( .A(DB[851]), .B(DB[844]), .Z(n4749) );
  AND U7825 ( .A(n1566), .B(n4750), .Z(n4748) );
  XOR U7826 ( .A(n4751), .B(n4752), .Z(n4750) );
  XOR U7827 ( .A(DB[844]), .B(DB[837]), .Z(n4752) );
  AND U7828 ( .A(n1570), .B(n4753), .Z(n4751) );
  XOR U7829 ( .A(n4754), .B(n4755), .Z(n4753) );
  XOR U7830 ( .A(DB[837]), .B(DB[830]), .Z(n4755) );
  AND U7831 ( .A(n1574), .B(n4756), .Z(n4754) );
  XOR U7832 ( .A(n4757), .B(n4758), .Z(n4756) );
  XOR U7833 ( .A(DB[830]), .B(DB[823]), .Z(n4758) );
  AND U7834 ( .A(n1578), .B(n4759), .Z(n4757) );
  XOR U7835 ( .A(n4760), .B(n4761), .Z(n4759) );
  XOR U7836 ( .A(DB[823]), .B(DB[816]), .Z(n4761) );
  AND U7837 ( .A(n1582), .B(n4762), .Z(n4760) );
  XOR U7838 ( .A(n4763), .B(n4764), .Z(n4762) );
  XOR U7839 ( .A(DB[816]), .B(DB[809]), .Z(n4764) );
  AND U7840 ( .A(n1586), .B(n4765), .Z(n4763) );
  XOR U7841 ( .A(n4766), .B(n4767), .Z(n4765) );
  XOR U7842 ( .A(DB[809]), .B(DB[802]), .Z(n4767) );
  AND U7843 ( .A(n1590), .B(n4768), .Z(n4766) );
  XOR U7844 ( .A(n4769), .B(n4770), .Z(n4768) );
  XOR U7845 ( .A(DB[802]), .B(DB[795]), .Z(n4770) );
  AND U7846 ( .A(n1594), .B(n4771), .Z(n4769) );
  XOR U7847 ( .A(n4772), .B(n4773), .Z(n4771) );
  XOR U7848 ( .A(DB[795]), .B(DB[788]), .Z(n4773) );
  AND U7849 ( .A(n1598), .B(n4774), .Z(n4772) );
  XOR U7850 ( .A(n4775), .B(n4776), .Z(n4774) );
  XOR U7851 ( .A(DB[788]), .B(DB[781]), .Z(n4776) );
  AND U7852 ( .A(n1602), .B(n4777), .Z(n4775) );
  XOR U7853 ( .A(n4778), .B(n4779), .Z(n4777) );
  XOR U7854 ( .A(DB[781]), .B(DB[774]), .Z(n4779) );
  AND U7855 ( .A(n1606), .B(n4780), .Z(n4778) );
  XOR U7856 ( .A(n4781), .B(n4782), .Z(n4780) );
  XOR U7857 ( .A(DB[774]), .B(DB[767]), .Z(n4782) );
  AND U7858 ( .A(n1610), .B(n4783), .Z(n4781) );
  XOR U7859 ( .A(n4784), .B(n4785), .Z(n4783) );
  XOR U7860 ( .A(DB[767]), .B(DB[760]), .Z(n4785) );
  AND U7861 ( .A(n1614), .B(n4786), .Z(n4784) );
  XOR U7862 ( .A(n4787), .B(n4788), .Z(n4786) );
  XOR U7863 ( .A(DB[760]), .B(DB[753]), .Z(n4788) );
  AND U7864 ( .A(n1618), .B(n4789), .Z(n4787) );
  XOR U7865 ( .A(n4790), .B(n4791), .Z(n4789) );
  XOR U7866 ( .A(DB[753]), .B(DB[746]), .Z(n4791) );
  AND U7867 ( .A(n1622), .B(n4792), .Z(n4790) );
  XOR U7868 ( .A(n4793), .B(n4794), .Z(n4792) );
  XOR U7869 ( .A(DB[746]), .B(DB[739]), .Z(n4794) );
  AND U7870 ( .A(n1626), .B(n4795), .Z(n4793) );
  XOR U7871 ( .A(n4796), .B(n4797), .Z(n4795) );
  XOR U7872 ( .A(DB[739]), .B(DB[732]), .Z(n4797) );
  AND U7873 ( .A(n1630), .B(n4798), .Z(n4796) );
  XOR U7874 ( .A(n4799), .B(n4800), .Z(n4798) );
  XOR U7875 ( .A(DB[732]), .B(DB[725]), .Z(n4800) );
  AND U7876 ( .A(n1634), .B(n4801), .Z(n4799) );
  XOR U7877 ( .A(n4802), .B(n4803), .Z(n4801) );
  XOR U7878 ( .A(DB[725]), .B(DB[718]), .Z(n4803) );
  AND U7879 ( .A(n1638), .B(n4804), .Z(n4802) );
  XOR U7880 ( .A(n4805), .B(n4806), .Z(n4804) );
  XOR U7881 ( .A(DB[718]), .B(DB[711]), .Z(n4806) );
  AND U7882 ( .A(n1642), .B(n4807), .Z(n4805) );
  XOR U7883 ( .A(n4808), .B(n4809), .Z(n4807) );
  XOR U7884 ( .A(DB[711]), .B(DB[704]), .Z(n4809) );
  AND U7885 ( .A(n1646), .B(n4810), .Z(n4808) );
  XOR U7886 ( .A(n4811), .B(n4812), .Z(n4810) );
  XOR U7887 ( .A(DB[704]), .B(DB[697]), .Z(n4812) );
  AND U7888 ( .A(n1650), .B(n4813), .Z(n4811) );
  XOR U7889 ( .A(n4814), .B(n4815), .Z(n4813) );
  XOR U7890 ( .A(DB[697]), .B(DB[690]), .Z(n4815) );
  AND U7891 ( .A(n1654), .B(n4816), .Z(n4814) );
  XOR U7892 ( .A(n4817), .B(n4818), .Z(n4816) );
  XOR U7893 ( .A(DB[690]), .B(DB[683]), .Z(n4818) );
  AND U7894 ( .A(n1658), .B(n4819), .Z(n4817) );
  XOR U7895 ( .A(n4820), .B(n4821), .Z(n4819) );
  XOR U7896 ( .A(DB[683]), .B(DB[676]), .Z(n4821) );
  AND U7897 ( .A(n1662), .B(n4822), .Z(n4820) );
  XOR U7898 ( .A(n4823), .B(n4824), .Z(n4822) );
  XOR U7899 ( .A(DB[676]), .B(DB[669]), .Z(n4824) );
  AND U7900 ( .A(n1666), .B(n4825), .Z(n4823) );
  XOR U7901 ( .A(n4826), .B(n4827), .Z(n4825) );
  XOR U7902 ( .A(DB[669]), .B(DB[662]), .Z(n4827) );
  AND U7903 ( .A(n1670), .B(n4828), .Z(n4826) );
  XOR U7904 ( .A(n4829), .B(n4830), .Z(n4828) );
  XOR U7905 ( .A(DB[662]), .B(DB[655]), .Z(n4830) );
  AND U7906 ( .A(n1674), .B(n4831), .Z(n4829) );
  XOR U7907 ( .A(n4832), .B(n4833), .Z(n4831) );
  XOR U7908 ( .A(DB[655]), .B(DB[648]), .Z(n4833) );
  AND U7909 ( .A(n1678), .B(n4834), .Z(n4832) );
  XOR U7910 ( .A(n4835), .B(n4836), .Z(n4834) );
  XOR U7911 ( .A(DB[648]), .B(DB[641]), .Z(n4836) );
  AND U7912 ( .A(n1682), .B(n4837), .Z(n4835) );
  XOR U7913 ( .A(n4838), .B(n4839), .Z(n4837) );
  XOR U7914 ( .A(DB[641]), .B(DB[634]), .Z(n4839) );
  AND U7915 ( .A(n1686), .B(n4840), .Z(n4838) );
  XOR U7916 ( .A(n4841), .B(n4842), .Z(n4840) );
  XOR U7917 ( .A(DB[634]), .B(DB[627]), .Z(n4842) );
  AND U7918 ( .A(n1690), .B(n4843), .Z(n4841) );
  XOR U7919 ( .A(n4844), .B(n4845), .Z(n4843) );
  XOR U7920 ( .A(DB[627]), .B(DB[620]), .Z(n4845) );
  AND U7921 ( .A(n1694), .B(n4846), .Z(n4844) );
  XOR U7922 ( .A(n4847), .B(n4848), .Z(n4846) );
  XOR U7923 ( .A(DB[620]), .B(DB[613]), .Z(n4848) );
  AND U7924 ( .A(n1698), .B(n4849), .Z(n4847) );
  XOR U7925 ( .A(n4850), .B(n4851), .Z(n4849) );
  XOR U7926 ( .A(DB[613]), .B(DB[606]), .Z(n4851) );
  AND U7927 ( .A(n1702), .B(n4852), .Z(n4850) );
  XOR U7928 ( .A(n4853), .B(n4854), .Z(n4852) );
  XOR U7929 ( .A(DB[606]), .B(DB[599]), .Z(n4854) );
  AND U7930 ( .A(n1706), .B(n4855), .Z(n4853) );
  XOR U7931 ( .A(n4856), .B(n4857), .Z(n4855) );
  XOR U7932 ( .A(DB[599]), .B(DB[592]), .Z(n4857) );
  AND U7933 ( .A(n1710), .B(n4858), .Z(n4856) );
  XOR U7934 ( .A(n4859), .B(n4860), .Z(n4858) );
  XOR U7935 ( .A(DB[592]), .B(DB[585]), .Z(n4860) );
  AND U7936 ( .A(n1714), .B(n4861), .Z(n4859) );
  XOR U7937 ( .A(n4862), .B(n4863), .Z(n4861) );
  XOR U7938 ( .A(DB[585]), .B(DB[578]), .Z(n4863) );
  AND U7939 ( .A(n1718), .B(n4864), .Z(n4862) );
  XOR U7940 ( .A(n4865), .B(n4866), .Z(n4864) );
  XOR U7941 ( .A(DB[578]), .B(DB[571]), .Z(n4866) );
  AND U7942 ( .A(n1722), .B(n4867), .Z(n4865) );
  XOR U7943 ( .A(n4868), .B(n4869), .Z(n4867) );
  XOR U7944 ( .A(DB[571]), .B(DB[564]), .Z(n4869) );
  AND U7945 ( .A(n1726), .B(n4870), .Z(n4868) );
  XOR U7946 ( .A(n4871), .B(n4872), .Z(n4870) );
  XOR U7947 ( .A(DB[564]), .B(DB[557]), .Z(n4872) );
  AND U7948 ( .A(n1730), .B(n4873), .Z(n4871) );
  XOR U7949 ( .A(n4874), .B(n4875), .Z(n4873) );
  XOR U7950 ( .A(DB[557]), .B(DB[550]), .Z(n4875) );
  AND U7951 ( .A(n1734), .B(n4876), .Z(n4874) );
  XOR U7952 ( .A(n4877), .B(n4878), .Z(n4876) );
  XOR U7953 ( .A(DB[550]), .B(DB[543]), .Z(n4878) );
  AND U7954 ( .A(n1738), .B(n4879), .Z(n4877) );
  XOR U7955 ( .A(n4880), .B(n4881), .Z(n4879) );
  XOR U7956 ( .A(DB[543]), .B(DB[536]), .Z(n4881) );
  AND U7957 ( .A(n1742), .B(n4882), .Z(n4880) );
  XOR U7958 ( .A(n4883), .B(n4884), .Z(n4882) );
  XOR U7959 ( .A(DB[536]), .B(DB[529]), .Z(n4884) );
  AND U7960 ( .A(n1746), .B(n4885), .Z(n4883) );
  XOR U7961 ( .A(n4886), .B(n4887), .Z(n4885) );
  XOR U7962 ( .A(DB[529]), .B(DB[522]), .Z(n4887) );
  AND U7963 ( .A(n1750), .B(n4888), .Z(n4886) );
  XOR U7964 ( .A(n4889), .B(n4890), .Z(n4888) );
  XOR U7965 ( .A(DB[522]), .B(DB[515]), .Z(n4890) );
  AND U7966 ( .A(n1754), .B(n4891), .Z(n4889) );
  XOR U7967 ( .A(n4892), .B(n4893), .Z(n4891) );
  XOR U7968 ( .A(DB[515]), .B(DB[508]), .Z(n4893) );
  AND U7969 ( .A(n1758), .B(n4894), .Z(n4892) );
  XOR U7970 ( .A(n4895), .B(n4896), .Z(n4894) );
  XOR U7971 ( .A(DB[508]), .B(DB[501]), .Z(n4896) );
  AND U7972 ( .A(n1762), .B(n4897), .Z(n4895) );
  XOR U7973 ( .A(n4898), .B(n4899), .Z(n4897) );
  XOR U7974 ( .A(DB[501]), .B(DB[494]), .Z(n4899) );
  AND U7975 ( .A(n1766), .B(n4900), .Z(n4898) );
  XOR U7976 ( .A(n4901), .B(n4902), .Z(n4900) );
  XOR U7977 ( .A(DB[494]), .B(DB[487]), .Z(n4902) );
  AND U7978 ( .A(n1770), .B(n4903), .Z(n4901) );
  XOR U7979 ( .A(n4904), .B(n4905), .Z(n4903) );
  XOR U7980 ( .A(DB[487]), .B(DB[480]), .Z(n4905) );
  AND U7981 ( .A(n1774), .B(n4906), .Z(n4904) );
  XOR U7982 ( .A(n4907), .B(n4908), .Z(n4906) );
  XOR U7983 ( .A(DB[480]), .B(DB[473]), .Z(n4908) );
  AND U7984 ( .A(n1778), .B(n4909), .Z(n4907) );
  XOR U7985 ( .A(n4910), .B(n4911), .Z(n4909) );
  XOR U7986 ( .A(DB[473]), .B(DB[466]), .Z(n4911) );
  AND U7987 ( .A(n1782), .B(n4912), .Z(n4910) );
  XOR U7988 ( .A(n4913), .B(n4914), .Z(n4912) );
  XOR U7989 ( .A(DB[466]), .B(DB[459]), .Z(n4914) );
  AND U7990 ( .A(n1786), .B(n4915), .Z(n4913) );
  XOR U7991 ( .A(n4916), .B(n4917), .Z(n4915) );
  XOR U7992 ( .A(DB[459]), .B(DB[452]), .Z(n4917) );
  AND U7993 ( .A(n1790), .B(n4918), .Z(n4916) );
  XOR U7994 ( .A(n4919), .B(n4920), .Z(n4918) );
  XOR U7995 ( .A(DB[452]), .B(DB[445]), .Z(n4920) );
  AND U7996 ( .A(n1794), .B(n4921), .Z(n4919) );
  XOR U7997 ( .A(n4922), .B(n4923), .Z(n4921) );
  XOR U7998 ( .A(DB[445]), .B(DB[438]), .Z(n4923) );
  AND U7999 ( .A(n1798), .B(n4924), .Z(n4922) );
  XOR U8000 ( .A(n4925), .B(n4926), .Z(n4924) );
  XOR U8001 ( .A(DB[438]), .B(DB[431]), .Z(n4926) );
  AND U8002 ( .A(n1802), .B(n4927), .Z(n4925) );
  XOR U8003 ( .A(n4928), .B(n4929), .Z(n4927) );
  XOR U8004 ( .A(DB[431]), .B(DB[424]), .Z(n4929) );
  AND U8005 ( .A(n1806), .B(n4930), .Z(n4928) );
  XOR U8006 ( .A(n4931), .B(n4932), .Z(n4930) );
  XOR U8007 ( .A(DB[424]), .B(DB[417]), .Z(n4932) );
  AND U8008 ( .A(n1810), .B(n4933), .Z(n4931) );
  XOR U8009 ( .A(n4934), .B(n4935), .Z(n4933) );
  XOR U8010 ( .A(DB[417]), .B(DB[410]), .Z(n4935) );
  AND U8011 ( .A(n1814), .B(n4936), .Z(n4934) );
  XOR U8012 ( .A(n4937), .B(n4938), .Z(n4936) );
  XOR U8013 ( .A(DB[410]), .B(DB[403]), .Z(n4938) );
  AND U8014 ( .A(n1818), .B(n4939), .Z(n4937) );
  XOR U8015 ( .A(n4940), .B(n4941), .Z(n4939) );
  XOR U8016 ( .A(DB[403]), .B(DB[396]), .Z(n4941) );
  AND U8017 ( .A(n1822), .B(n4942), .Z(n4940) );
  XOR U8018 ( .A(n4943), .B(n4944), .Z(n4942) );
  XOR U8019 ( .A(DB[396]), .B(DB[389]), .Z(n4944) );
  AND U8020 ( .A(n1826), .B(n4945), .Z(n4943) );
  XOR U8021 ( .A(n4946), .B(n4947), .Z(n4945) );
  XOR U8022 ( .A(DB[389]), .B(DB[382]), .Z(n4947) );
  AND U8023 ( .A(n1830), .B(n4948), .Z(n4946) );
  XOR U8024 ( .A(n4949), .B(n4950), .Z(n4948) );
  XOR U8025 ( .A(DB[382]), .B(DB[375]), .Z(n4950) );
  AND U8026 ( .A(n1834), .B(n4951), .Z(n4949) );
  XOR U8027 ( .A(n4952), .B(n4953), .Z(n4951) );
  XOR U8028 ( .A(DB[375]), .B(DB[368]), .Z(n4953) );
  AND U8029 ( .A(n1838), .B(n4954), .Z(n4952) );
  XOR U8030 ( .A(n4955), .B(n4956), .Z(n4954) );
  XOR U8031 ( .A(DB[368]), .B(DB[361]), .Z(n4956) );
  AND U8032 ( .A(n1842), .B(n4957), .Z(n4955) );
  XOR U8033 ( .A(n4958), .B(n4959), .Z(n4957) );
  XOR U8034 ( .A(DB[361]), .B(DB[354]), .Z(n4959) );
  AND U8035 ( .A(n1846), .B(n4960), .Z(n4958) );
  XOR U8036 ( .A(n4961), .B(n4962), .Z(n4960) );
  XOR U8037 ( .A(DB[354]), .B(DB[347]), .Z(n4962) );
  AND U8038 ( .A(n1850), .B(n4963), .Z(n4961) );
  XOR U8039 ( .A(n4964), .B(n4965), .Z(n4963) );
  XOR U8040 ( .A(DB[347]), .B(DB[340]), .Z(n4965) );
  AND U8041 ( .A(n1854), .B(n4966), .Z(n4964) );
  XOR U8042 ( .A(n4967), .B(n4968), .Z(n4966) );
  XOR U8043 ( .A(DB[340]), .B(DB[333]), .Z(n4968) );
  AND U8044 ( .A(n1858), .B(n4969), .Z(n4967) );
  XOR U8045 ( .A(n4970), .B(n4971), .Z(n4969) );
  XOR U8046 ( .A(DB[333]), .B(DB[326]), .Z(n4971) );
  AND U8047 ( .A(n1862), .B(n4972), .Z(n4970) );
  XOR U8048 ( .A(n4973), .B(n4974), .Z(n4972) );
  XOR U8049 ( .A(DB[326]), .B(DB[319]), .Z(n4974) );
  AND U8050 ( .A(n1866), .B(n4975), .Z(n4973) );
  XOR U8051 ( .A(n4976), .B(n4977), .Z(n4975) );
  XOR U8052 ( .A(DB[319]), .B(DB[312]), .Z(n4977) );
  AND U8053 ( .A(n1870), .B(n4978), .Z(n4976) );
  XOR U8054 ( .A(n4979), .B(n4980), .Z(n4978) );
  XOR U8055 ( .A(DB[312]), .B(DB[305]), .Z(n4980) );
  AND U8056 ( .A(n1874), .B(n4981), .Z(n4979) );
  XOR U8057 ( .A(n4982), .B(n4983), .Z(n4981) );
  XOR U8058 ( .A(DB[305]), .B(DB[298]), .Z(n4983) );
  AND U8059 ( .A(n1878), .B(n4984), .Z(n4982) );
  XOR U8060 ( .A(n4985), .B(n4986), .Z(n4984) );
  XOR U8061 ( .A(DB[298]), .B(DB[291]), .Z(n4986) );
  AND U8062 ( .A(n1882), .B(n4987), .Z(n4985) );
  XOR U8063 ( .A(n4988), .B(n4989), .Z(n4987) );
  XOR U8064 ( .A(DB[291]), .B(DB[284]), .Z(n4989) );
  AND U8065 ( .A(n1886), .B(n4990), .Z(n4988) );
  XOR U8066 ( .A(n4991), .B(n4992), .Z(n4990) );
  XOR U8067 ( .A(DB[284]), .B(DB[277]), .Z(n4992) );
  AND U8068 ( .A(n1890), .B(n4993), .Z(n4991) );
  XOR U8069 ( .A(n4994), .B(n4995), .Z(n4993) );
  XOR U8070 ( .A(DB[277]), .B(DB[270]), .Z(n4995) );
  AND U8071 ( .A(n1894), .B(n4996), .Z(n4994) );
  XOR U8072 ( .A(n4997), .B(n4998), .Z(n4996) );
  XOR U8073 ( .A(DB[270]), .B(DB[263]), .Z(n4998) );
  AND U8074 ( .A(n1898), .B(n4999), .Z(n4997) );
  XOR U8075 ( .A(n5000), .B(n5001), .Z(n4999) );
  XOR U8076 ( .A(DB[263]), .B(DB[256]), .Z(n5001) );
  AND U8077 ( .A(n1902), .B(n5002), .Z(n5000) );
  XOR U8078 ( .A(n5003), .B(n5004), .Z(n5002) );
  XOR U8079 ( .A(DB[256]), .B(DB[249]), .Z(n5004) );
  AND U8080 ( .A(n1906), .B(n5005), .Z(n5003) );
  XOR U8081 ( .A(n5006), .B(n5007), .Z(n5005) );
  XOR U8082 ( .A(DB[249]), .B(DB[242]), .Z(n5007) );
  AND U8083 ( .A(n1910), .B(n5008), .Z(n5006) );
  XOR U8084 ( .A(n5009), .B(n5010), .Z(n5008) );
  XOR U8085 ( .A(DB[242]), .B(DB[235]), .Z(n5010) );
  AND U8086 ( .A(n1914), .B(n5011), .Z(n5009) );
  XOR U8087 ( .A(n5012), .B(n5013), .Z(n5011) );
  XOR U8088 ( .A(DB[235]), .B(DB[228]), .Z(n5013) );
  AND U8089 ( .A(n1918), .B(n5014), .Z(n5012) );
  XOR U8090 ( .A(n5015), .B(n5016), .Z(n5014) );
  XOR U8091 ( .A(DB[228]), .B(DB[221]), .Z(n5016) );
  AND U8092 ( .A(n1922), .B(n5017), .Z(n5015) );
  XOR U8093 ( .A(n5018), .B(n5019), .Z(n5017) );
  XOR U8094 ( .A(DB[221]), .B(DB[214]), .Z(n5019) );
  AND U8095 ( .A(n1926), .B(n5020), .Z(n5018) );
  XOR U8096 ( .A(n5021), .B(n5022), .Z(n5020) );
  XOR U8097 ( .A(DB[214]), .B(DB[207]), .Z(n5022) );
  AND U8098 ( .A(n1930), .B(n5023), .Z(n5021) );
  XOR U8099 ( .A(n5024), .B(n5025), .Z(n5023) );
  XOR U8100 ( .A(DB[207]), .B(DB[200]), .Z(n5025) );
  AND U8101 ( .A(n1934), .B(n5026), .Z(n5024) );
  XOR U8102 ( .A(n5027), .B(n5028), .Z(n5026) );
  XOR U8103 ( .A(DB[200]), .B(DB[193]), .Z(n5028) );
  AND U8104 ( .A(n1938), .B(n5029), .Z(n5027) );
  XOR U8105 ( .A(n5030), .B(n5031), .Z(n5029) );
  XOR U8106 ( .A(DB[193]), .B(DB[186]), .Z(n5031) );
  AND U8107 ( .A(n1942), .B(n5032), .Z(n5030) );
  XOR U8108 ( .A(n5033), .B(n5034), .Z(n5032) );
  XOR U8109 ( .A(DB[186]), .B(DB[179]), .Z(n5034) );
  AND U8110 ( .A(n1946), .B(n5035), .Z(n5033) );
  XOR U8111 ( .A(n5036), .B(n5037), .Z(n5035) );
  XOR U8112 ( .A(DB[179]), .B(DB[172]), .Z(n5037) );
  AND U8113 ( .A(n1950), .B(n5038), .Z(n5036) );
  XOR U8114 ( .A(n5039), .B(n5040), .Z(n5038) );
  XOR U8115 ( .A(DB[172]), .B(DB[165]), .Z(n5040) );
  AND U8116 ( .A(n1954), .B(n5041), .Z(n5039) );
  XOR U8117 ( .A(n5042), .B(n5043), .Z(n5041) );
  XOR U8118 ( .A(DB[165]), .B(DB[158]), .Z(n5043) );
  AND U8119 ( .A(n1958), .B(n5044), .Z(n5042) );
  XOR U8120 ( .A(n5045), .B(n5046), .Z(n5044) );
  XOR U8121 ( .A(DB[158]), .B(DB[151]), .Z(n5046) );
  AND U8122 ( .A(n1962), .B(n5047), .Z(n5045) );
  XOR U8123 ( .A(n5048), .B(n5049), .Z(n5047) );
  XOR U8124 ( .A(DB[151]), .B(DB[144]), .Z(n5049) );
  AND U8125 ( .A(n1966), .B(n5050), .Z(n5048) );
  XOR U8126 ( .A(n5051), .B(n5052), .Z(n5050) );
  XOR U8127 ( .A(DB[144]), .B(DB[137]), .Z(n5052) );
  AND U8128 ( .A(n1970), .B(n5053), .Z(n5051) );
  XOR U8129 ( .A(n5054), .B(n5055), .Z(n5053) );
  XOR U8130 ( .A(DB[137]), .B(DB[130]), .Z(n5055) );
  AND U8131 ( .A(n1974), .B(n5056), .Z(n5054) );
  XOR U8132 ( .A(n5057), .B(n5058), .Z(n5056) );
  XOR U8133 ( .A(DB[130]), .B(DB[123]), .Z(n5058) );
  AND U8134 ( .A(n1978), .B(n5059), .Z(n5057) );
  XOR U8135 ( .A(n5060), .B(n5061), .Z(n5059) );
  XOR U8136 ( .A(DB[123]), .B(DB[116]), .Z(n5061) );
  AND U8137 ( .A(n1982), .B(n5062), .Z(n5060) );
  XOR U8138 ( .A(n5063), .B(n5064), .Z(n5062) );
  XOR U8139 ( .A(DB[116]), .B(DB[109]), .Z(n5064) );
  AND U8140 ( .A(n1986), .B(n5065), .Z(n5063) );
  XOR U8141 ( .A(n5066), .B(n5067), .Z(n5065) );
  XOR U8142 ( .A(DB[109]), .B(DB[102]), .Z(n5067) );
  AND U8143 ( .A(n1990), .B(n5068), .Z(n5066) );
  XOR U8144 ( .A(n5069), .B(n5070), .Z(n5068) );
  XOR U8145 ( .A(DB[95]), .B(DB[102]), .Z(n5070) );
  AND U8146 ( .A(n1994), .B(n5071), .Z(n5069) );
  XOR U8147 ( .A(n5072), .B(n5073), .Z(n5071) );
  XOR U8148 ( .A(DB[95]), .B(DB[88]), .Z(n5073) );
  AND U8149 ( .A(n1998), .B(n5074), .Z(n5072) );
  XOR U8150 ( .A(n5075), .B(n5076), .Z(n5074) );
  XOR U8151 ( .A(DB[88]), .B(DB[81]), .Z(n5076) );
  AND U8152 ( .A(n2002), .B(n5077), .Z(n5075) );
  XOR U8153 ( .A(n5078), .B(n5079), .Z(n5077) );
  XOR U8154 ( .A(DB[81]), .B(DB[74]), .Z(n5079) );
  AND U8155 ( .A(n2006), .B(n5080), .Z(n5078) );
  XOR U8156 ( .A(n5081), .B(n5082), .Z(n5080) );
  XOR U8157 ( .A(DB[74]), .B(DB[67]), .Z(n5082) );
  AND U8158 ( .A(n2010), .B(n5083), .Z(n5081) );
  XOR U8159 ( .A(n5084), .B(n5085), .Z(n5083) );
  XOR U8160 ( .A(DB[67]), .B(DB[60]), .Z(n5085) );
  AND U8161 ( .A(n2014), .B(n5086), .Z(n5084) );
  XOR U8162 ( .A(n5087), .B(n5088), .Z(n5086) );
  XOR U8163 ( .A(DB[60]), .B(DB[53]), .Z(n5088) );
  AND U8164 ( .A(n2018), .B(n5089), .Z(n5087) );
  XOR U8165 ( .A(n5090), .B(n5091), .Z(n5089) );
  XOR U8166 ( .A(DB[53]), .B(DB[46]), .Z(n5091) );
  AND U8167 ( .A(n2022), .B(n5092), .Z(n5090) );
  XOR U8168 ( .A(n5093), .B(n5094), .Z(n5092) );
  XOR U8169 ( .A(DB[46]), .B(DB[39]), .Z(n5094) );
  AND U8170 ( .A(n2026), .B(n5095), .Z(n5093) );
  XOR U8171 ( .A(n5096), .B(n5097), .Z(n5095) );
  XOR U8172 ( .A(DB[39]), .B(DB[32]), .Z(n5097) );
  AND U8173 ( .A(n2030), .B(n5098), .Z(n5096) );
  XOR U8174 ( .A(n5099), .B(n5100), .Z(n5098) );
  XOR U8175 ( .A(DB[32]), .B(DB[25]), .Z(n5100) );
  AND U8176 ( .A(n2034), .B(n5101), .Z(n5099) );
  XOR U8177 ( .A(n5102), .B(n5103), .Z(n5101) );
  XOR U8178 ( .A(DB[25]), .B(DB[18]), .Z(n5103) );
  AND U8179 ( .A(n2038), .B(n5104), .Z(n5102) );
  XOR U8180 ( .A(n5105), .B(n5106), .Z(n5104) );
  XOR U8181 ( .A(DB[18]), .B(DB[11]), .Z(n5106) );
  AND U8182 ( .A(n2042), .B(n5107), .Z(n5105) );
  XOR U8183 ( .A(DB[4]), .B(DB[11]), .Z(n5107) );
  XOR U8184 ( .A(DB[3580]), .B(n5108), .Z(min_val_out[3]) );
  AND U8185 ( .A(n2), .B(n5109), .Z(n5108) );
  XOR U8186 ( .A(n5110), .B(n5111), .Z(n5109) );
  XOR U8187 ( .A(DB[3580]), .B(DB[3573]), .Z(n5111) );
  AND U8188 ( .A(n6), .B(n5112), .Z(n5110) );
  XOR U8189 ( .A(n5113), .B(n5114), .Z(n5112) );
  XOR U8190 ( .A(DB[3573]), .B(DB[3566]), .Z(n5114) );
  AND U8191 ( .A(n10), .B(n5115), .Z(n5113) );
  XOR U8192 ( .A(n5116), .B(n5117), .Z(n5115) );
  XOR U8193 ( .A(DB[3566]), .B(DB[3559]), .Z(n5117) );
  AND U8194 ( .A(n14), .B(n5118), .Z(n5116) );
  XOR U8195 ( .A(n5119), .B(n5120), .Z(n5118) );
  XOR U8196 ( .A(DB[3559]), .B(DB[3552]), .Z(n5120) );
  AND U8197 ( .A(n18), .B(n5121), .Z(n5119) );
  XOR U8198 ( .A(n5122), .B(n5123), .Z(n5121) );
  XOR U8199 ( .A(DB[3552]), .B(DB[3545]), .Z(n5123) );
  AND U8200 ( .A(n22), .B(n5124), .Z(n5122) );
  XOR U8201 ( .A(n5125), .B(n5126), .Z(n5124) );
  XOR U8202 ( .A(DB[3545]), .B(DB[3538]), .Z(n5126) );
  AND U8203 ( .A(n26), .B(n5127), .Z(n5125) );
  XOR U8204 ( .A(n5128), .B(n5129), .Z(n5127) );
  XOR U8205 ( .A(DB[3538]), .B(DB[3531]), .Z(n5129) );
  AND U8206 ( .A(n30), .B(n5130), .Z(n5128) );
  XOR U8207 ( .A(n5131), .B(n5132), .Z(n5130) );
  XOR U8208 ( .A(DB[3531]), .B(DB[3524]), .Z(n5132) );
  AND U8209 ( .A(n34), .B(n5133), .Z(n5131) );
  XOR U8210 ( .A(n5134), .B(n5135), .Z(n5133) );
  XOR U8211 ( .A(DB[3524]), .B(DB[3517]), .Z(n5135) );
  AND U8212 ( .A(n38), .B(n5136), .Z(n5134) );
  XOR U8213 ( .A(n5137), .B(n5138), .Z(n5136) );
  XOR U8214 ( .A(DB[3517]), .B(DB[3510]), .Z(n5138) );
  AND U8215 ( .A(n42), .B(n5139), .Z(n5137) );
  XOR U8216 ( .A(n5140), .B(n5141), .Z(n5139) );
  XOR U8217 ( .A(DB[3510]), .B(DB[3503]), .Z(n5141) );
  AND U8218 ( .A(n46), .B(n5142), .Z(n5140) );
  XOR U8219 ( .A(n5143), .B(n5144), .Z(n5142) );
  XOR U8220 ( .A(DB[3503]), .B(DB[3496]), .Z(n5144) );
  AND U8221 ( .A(n50), .B(n5145), .Z(n5143) );
  XOR U8222 ( .A(n5146), .B(n5147), .Z(n5145) );
  XOR U8223 ( .A(DB[3496]), .B(DB[3489]), .Z(n5147) );
  AND U8224 ( .A(n54), .B(n5148), .Z(n5146) );
  XOR U8225 ( .A(n5149), .B(n5150), .Z(n5148) );
  XOR U8226 ( .A(DB[3489]), .B(DB[3482]), .Z(n5150) );
  AND U8227 ( .A(n58), .B(n5151), .Z(n5149) );
  XOR U8228 ( .A(n5152), .B(n5153), .Z(n5151) );
  XOR U8229 ( .A(DB[3482]), .B(DB[3475]), .Z(n5153) );
  AND U8230 ( .A(n62), .B(n5154), .Z(n5152) );
  XOR U8231 ( .A(n5155), .B(n5156), .Z(n5154) );
  XOR U8232 ( .A(DB[3475]), .B(DB[3468]), .Z(n5156) );
  AND U8233 ( .A(n66), .B(n5157), .Z(n5155) );
  XOR U8234 ( .A(n5158), .B(n5159), .Z(n5157) );
  XOR U8235 ( .A(DB[3468]), .B(DB[3461]), .Z(n5159) );
  AND U8236 ( .A(n70), .B(n5160), .Z(n5158) );
  XOR U8237 ( .A(n5161), .B(n5162), .Z(n5160) );
  XOR U8238 ( .A(DB[3461]), .B(DB[3454]), .Z(n5162) );
  AND U8239 ( .A(n74), .B(n5163), .Z(n5161) );
  XOR U8240 ( .A(n5164), .B(n5165), .Z(n5163) );
  XOR U8241 ( .A(DB[3454]), .B(DB[3447]), .Z(n5165) );
  AND U8242 ( .A(n78), .B(n5166), .Z(n5164) );
  XOR U8243 ( .A(n5167), .B(n5168), .Z(n5166) );
  XOR U8244 ( .A(DB[3447]), .B(DB[3440]), .Z(n5168) );
  AND U8245 ( .A(n82), .B(n5169), .Z(n5167) );
  XOR U8246 ( .A(n5170), .B(n5171), .Z(n5169) );
  XOR U8247 ( .A(DB[3440]), .B(DB[3433]), .Z(n5171) );
  AND U8248 ( .A(n86), .B(n5172), .Z(n5170) );
  XOR U8249 ( .A(n5173), .B(n5174), .Z(n5172) );
  XOR U8250 ( .A(DB[3433]), .B(DB[3426]), .Z(n5174) );
  AND U8251 ( .A(n90), .B(n5175), .Z(n5173) );
  XOR U8252 ( .A(n5176), .B(n5177), .Z(n5175) );
  XOR U8253 ( .A(DB[3426]), .B(DB[3419]), .Z(n5177) );
  AND U8254 ( .A(n94), .B(n5178), .Z(n5176) );
  XOR U8255 ( .A(n5179), .B(n5180), .Z(n5178) );
  XOR U8256 ( .A(DB[3419]), .B(DB[3412]), .Z(n5180) );
  AND U8257 ( .A(n98), .B(n5181), .Z(n5179) );
  XOR U8258 ( .A(n5182), .B(n5183), .Z(n5181) );
  XOR U8259 ( .A(DB[3412]), .B(DB[3405]), .Z(n5183) );
  AND U8260 ( .A(n102), .B(n5184), .Z(n5182) );
  XOR U8261 ( .A(n5185), .B(n5186), .Z(n5184) );
  XOR U8262 ( .A(DB[3405]), .B(DB[3398]), .Z(n5186) );
  AND U8263 ( .A(n106), .B(n5187), .Z(n5185) );
  XOR U8264 ( .A(n5188), .B(n5189), .Z(n5187) );
  XOR U8265 ( .A(DB[3398]), .B(DB[3391]), .Z(n5189) );
  AND U8266 ( .A(n110), .B(n5190), .Z(n5188) );
  XOR U8267 ( .A(n5191), .B(n5192), .Z(n5190) );
  XOR U8268 ( .A(DB[3391]), .B(DB[3384]), .Z(n5192) );
  AND U8269 ( .A(n114), .B(n5193), .Z(n5191) );
  XOR U8270 ( .A(n5194), .B(n5195), .Z(n5193) );
  XOR U8271 ( .A(DB[3384]), .B(DB[3377]), .Z(n5195) );
  AND U8272 ( .A(n118), .B(n5196), .Z(n5194) );
  XOR U8273 ( .A(n5197), .B(n5198), .Z(n5196) );
  XOR U8274 ( .A(DB[3377]), .B(DB[3370]), .Z(n5198) );
  AND U8275 ( .A(n122), .B(n5199), .Z(n5197) );
  XOR U8276 ( .A(n5200), .B(n5201), .Z(n5199) );
  XOR U8277 ( .A(DB[3370]), .B(DB[3363]), .Z(n5201) );
  AND U8278 ( .A(n126), .B(n5202), .Z(n5200) );
  XOR U8279 ( .A(n5203), .B(n5204), .Z(n5202) );
  XOR U8280 ( .A(DB[3363]), .B(DB[3356]), .Z(n5204) );
  AND U8281 ( .A(n130), .B(n5205), .Z(n5203) );
  XOR U8282 ( .A(n5206), .B(n5207), .Z(n5205) );
  XOR U8283 ( .A(DB[3356]), .B(DB[3349]), .Z(n5207) );
  AND U8284 ( .A(n134), .B(n5208), .Z(n5206) );
  XOR U8285 ( .A(n5209), .B(n5210), .Z(n5208) );
  XOR U8286 ( .A(DB[3349]), .B(DB[3342]), .Z(n5210) );
  AND U8287 ( .A(n138), .B(n5211), .Z(n5209) );
  XOR U8288 ( .A(n5212), .B(n5213), .Z(n5211) );
  XOR U8289 ( .A(DB[3342]), .B(DB[3335]), .Z(n5213) );
  AND U8290 ( .A(n142), .B(n5214), .Z(n5212) );
  XOR U8291 ( .A(n5215), .B(n5216), .Z(n5214) );
  XOR U8292 ( .A(DB[3335]), .B(DB[3328]), .Z(n5216) );
  AND U8293 ( .A(n146), .B(n5217), .Z(n5215) );
  XOR U8294 ( .A(n5218), .B(n5219), .Z(n5217) );
  XOR U8295 ( .A(DB[3328]), .B(DB[3321]), .Z(n5219) );
  AND U8296 ( .A(n150), .B(n5220), .Z(n5218) );
  XOR U8297 ( .A(n5221), .B(n5222), .Z(n5220) );
  XOR U8298 ( .A(DB[3321]), .B(DB[3314]), .Z(n5222) );
  AND U8299 ( .A(n154), .B(n5223), .Z(n5221) );
  XOR U8300 ( .A(n5224), .B(n5225), .Z(n5223) );
  XOR U8301 ( .A(DB[3314]), .B(DB[3307]), .Z(n5225) );
  AND U8302 ( .A(n158), .B(n5226), .Z(n5224) );
  XOR U8303 ( .A(n5227), .B(n5228), .Z(n5226) );
  XOR U8304 ( .A(DB[3307]), .B(DB[3300]), .Z(n5228) );
  AND U8305 ( .A(n162), .B(n5229), .Z(n5227) );
  XOR U8306 ( .A(n5230), .B(n5231), .Z(n5229) );
  XOR U8307 ( .A(DB[3300]), .B(DB[3293]), .Z(n5231) );
  AND U8308 ( .A(n166), .B(n5232), .Z(n5230) );
  XOR U8309 ( .A(n5233), .B(n5234), .Z(n5232) );
  XOR U8310 ( .A(DB[3293]), .B(DB[3286]), .Z(n5234) );
  AND U8311 ( .A(n170), .B(n5235), .Z(n5233) );
  XOR U8312 ( .A(n5236), .B(n5237), .Z(n5235) );
  XOR U8313 ( .A(DB[3286]), .B(DB[3279]), .Z(n5237) );
  AND U8314 ( .A(n174), .B(n5238), .Z(n5236) );
  XOR U8315 ( .A(n5239), .B(n5240), .Z(n5238) );
  XOR U8316 ( .A(DB[3279]), .B(DB[3272]), .Z(n5240) );
  AND U8317 ( .A(n178), .B(n5241), .Z(n5239) );
  XOR U8318 ( .A(n5242), .B(n5243), .Z(n5241) );
  XOR U8319 ( .A(DB[3272]), .B(DB[3265]), .Z(n5243) );
  AND U8320 ( .A(n182), .B(n5244), .Z(n5242) );
  XOR U8321 ( .A(n5245), .B(n5246), .Z(n5244) );
  XOR U8322 ( .A(DB[3265]), .B(DB[3258]), .Z(n5246) );
  AND U8323 ( .A(n186), .B(n5247), .Z(n5245) );
  XOR U8324 ( .A(n5248), .B(n5249), .Z(n5247) );
  XOR U8325 ( .A(DB[3258]), .B(DB[3251]), .Z(n5249) );
  AND U8326 ( .A(n190), .B(n5250), .Z(n5248) );
  XOR U8327 ( .A(n5251), .B(n5252), .Z(n5250) );
  XOR U8328 ( .A(DB[3251]), .B(DB[3244]), .Z(n5252) );
  AND U8329 ( .A(n194), .B(n5253), .Z(n5251) );
  XOR U8330 ( .A(n5254), .B(n5255), .Z(n5253) );
  XOR U8331 ( .A(DB[3244]), .B(DB[3237]), .Z(n5255) );
  AND U8332 ( .A(n198), .B(n5256), .Z(n5254) );
  XOR U8333 ( .A(n5257), .B(n5258), .Z(n5256) );
  XOR U8334 ( .A(DB[3237]), .B(DB[3230]), .Z(n5258) );
  AND U8335 ( .A(n202), .B(n5259), .Z(n5257) );
  XOR U8336 ( .A(n5260), .B(n5261), .Z(n5259) );
  XOR U8337 ( .A(DB[3230]), .B(DB[3223]), .Z(n5261) );
  AND U8338 ( .A(n206), .B(n5262), .Z(n5260) );
  XOR U8339 ( .A(n5263), .B(n5264), .Z(n5262) );
  XOR U8340 ( .A(DB[3223]), .B(DB[3216]), .Z(n5264) );
  AND U8341 ( .A(n210), .B(n5265), .Z(n5263) );
  XOR U8342 ( .A(n5266), .B(n5267), .Z(n5265) );
  XOR U8343 ( .A(DB[3216]), .B(DB[3209]), .Z(n5267) );
  AND U8344 ( .A(n214), .B(n5268), .Z(n5266) );
  XOR U8345 ( .A(n5269), .B(n5270), .Z(n5268) );
  XOR U8346 ( .A(DB[3209]), .B(DB[3202]), .Z(n5270) );
  AND U8347 ( .A(n218), .B(n5271), .Z(n5269) );
  XOR U8348 ( .A(n5272), .B(n5273), .Z(n5271) );
  XOR U8349 ( .A(DB[3202]), .B(DB[3195]), .Z(n5273) );
  AND U8350 ( .A(n222), .B(n5274), .Z(n5272) );
  XOR U8351 ( .A(n5275), .B(n5276), .Z(n5274) );
  XOR U8352 ( .A(DB[3195]), .B(DB[3188]), .Z(n5276) );
  AND U8353 ( .A(n226), .B(n5277), .Z(n5275) );
  XOR U8354 ( .A(n5278), .B(n5279), .Z(n5277) );
  XOR U8355 ( .A(DB[3188]), .B(DB[3181]), .Z(n5279) );
  AND U8356 ( .A(n230), .B(n5280), .Z(n5278) );
  XOR U8357 ( .A(n5281), .B(n5282), .Z(n5280) );
  XOR U8358 ( .A(DB[3181]), .B(DB[3174]), .Z(n5282) );
  AND U8359 ( .A(n234), .B(n5283), .Z(n5281) );
  XOR U8360 ( .A(n5284), .B(n5285), .Z(n5283) );
  XOR U8361 ( .A(DB[3174]), .B(DB[3167]), .Z(n5285) );
  AND U8362 ( .A(n238), .B(n5286), .Z(n5284) );
  XOR U8363 ( .A(n5287), .B(n5288), .Z(n5286) );
  XOR U8364 ( .A(DB[3167]), .B(DB[3160]), .Z(n5288) );
  AND U8365 ( .A(n242), .B(n5289), .Z(n5287) );
  XOR U8366 ( .A(n5290), .B(n5291), .Z(n5289) );
  XOR U8367 ( .A(DB[3160]), .B(DB[3153]), .Z(n5291) );
  AND U8368 ( .A(n246), .B(n5292), .Z(n5290) );
  XOR U8369 ( .A(n5293), .B(n5294), .Z(n5292) );
  XOR U8370 ( .A(DB[3153]), .B(DB[3146]), .Z(n5294) );
  AND U8371 ( .A(n250), .B(n5295), .Z(n5293) );
  XOR U8372 ( .A(n5296), .B(n5297), .Z(n5295) );
  XOR U8373 ( .A(DB[3146]), .B(DB[3139]), .Z(n5297) );
  AND U8374 ( .A(n254), .B(n5298), .Z(n5296) );
  XOR U8375 ( .A(n5299), .B(n5300), .Z(n5298) );
  XOR U8376 ( .A(DB[3139]), .B(DB[3132]), .Z(n5300) );
  AND U8377 ( .A(n258), .B(n5301), .Z(n5299) );
  XOR U8378 ( .A(n5302), .B(n5303), .Z(n5301) );
  XOR U8379 ( .A(DB[3132]), .B(DB[3125]), .Z(n5303) );
  AND U8380 ( .A(n262), .B(n5304), .Z(n5302) );
  XOR U8381 ( .A(n5305), .B(n5306), .Z(n5304) );
  XOR U8382 ( .A(DB[3125]), .B(DB[3118]), .Z(n5306) );
  AND U8383 ( .A(n266), .B(n5307), .Z(n5305) );
  XOR U8384 ( .A(n5308), .B(n5309), .Z(n5307) );
  XOR U8385 ( .A(DB[3118]), .B(DB[3111]), .Z(n5309) );
  AND U8386 ( .A(n270), .B(n5310), .Z(n5308) );
  XOR U8387 ( .A(n5311), .B(n5312), .Z(n5310) );
  XOR U8388 ( .A(DB[3111]), .B(DB[3104]), .Z(n5312) );
  AND U8389 ( .A(n274), .B(n5313), .Z(n5311) );
  XOR U8390 ( .A(n5314), .B(n5315), .Z(n5313) );
  XOR U8391 ( .A(DB[3104]), .B(DB[3097]), .Z(n5315) );
  AND U8392 ( .A(n278), .B(n5316), .Z(n5314) );
  XOR U8393 ( .A(n5317), .B(n5318), .Z(n5316) );
  XOR U8394 ( .A(DB[3097]), .B(DB[3090]), .Z(n5318) );
  AND U8395 ( .A(n282), .B(n5319), .Z(n5317) );
  XOR U8396 ( .A(n5320), .B(n5321), .Z(n5319) );
  XOR U8397 ( .A(DB[3090]), .B(DB[3083]), .Z(n5321) );
  AND U8398 ( .A(n286), .B(n5322), .Z(n5320) );
  XOR U8399 ( .A(n5323), .B(n5324), .Z(n5322) );
  XOR U8400 ( .A(DB[3083]), .B(DB[3076]), .Z(n5324) );
  AND U8401 ( .A(n290), .B(n5325), .Z(n5323) );
  XOR U8402 ( .A(n5326), .B(n5327), .Z(n5325) );
  XOR U8403 ( .A(DB[3076]), .B(DB[3069]), .Z(n5327) );
  AND U8404 ( .A(n294), .B(n5328), .Z(n5326) );
  XOR U8405 ( .A(n5329), .B(n5330), .Z(n5328) );
  XOR U8406 ( .A(DB[3069]), .B(DB[3062]), .Z(n5330) );
  AND U8407 ( .A(n298), .B(n5331), .Z(n5329) );
  XOR U8408 ( .A(n5332), .B(n5333), .Z(n5331) );
  XOR U8409 ( .A(DB[3062]), .B(DB[3055]), .Z(n5333) );
  AND U8410 ( .A(n302), .B(n5334), .Z(n5332) );
  XOR U8411 ( .A(n5335), .B(n5336), .Z(n5334) );
  XOR U8412 ( .A(DB[3055]), .B(DB[3048]), .Z(n5336) );
  AND U8413 ( .A(n306), .B(n5337), .Z(n5335) );
  XOR U8414 ( .A(n5338), .B(n5339), .Z(n5337) );
  XOR U8415 ( .A(DB[3048]), .B(DB[3041]), .Z(n5339) );
  AND U8416 ( .A(n310), .B(n5340), .Z(n5338) );
  XOR U8417 ( .A(n5341), .B(n5342), .Z(n5340) );
  XOR U8418 ( .A(DB[3041]), .B(DB[3034]), .Z(n5342) );
  AND U8419 ( .A(n314), .B(n5343), .Z(n5341) );
  XOR U8420 ( .A(n5344), .B(n5345), .Z(n5343) );
  XOR U8421 ( .A(DB[3034]), .B(DB[3027]), .Z(n5345) );
  AND U8422 ( .A(n318), .B(n5346), .Z(n5344) );
  XOR U8423 ( .A(n5347), .B(n5348), .Z(n5346) );
  XOR U8424 ( .A(DB[3027]), .B(DB[3020]), .Z(n5348) );
  AND U8425 ( .A(n322), .B(n5349), .Z(n5347) );
  XOR U8426 ( .A(n5350), .B(n5351), .Z(n5349) );
  XOR U8427 ( .A(DB[3020]), .B(DB[3013]), .Z(n5351) );
  AND U8428 ( .A(n326), .B(n5352), .Z(n5350) );
  XOR U8429 ( .A(n5353), .B(n5354), .Z(n5352) );
  XOR U8430 ( .A(DB[3013]), .B(DB[3006]), .Z(n5354) );
  AND U8431 ( .A(n330), .B(n5355), .Z(n5353) );
  XOR U8432 ( .A(n5356), .B(n5357), .Z(n5355) );
  XOR U8433 ( .A(DB[3006]), .B(DB[2999]), .Z(n5357) );
  AND U8434 ( .A(n334), .B(n5358), .Z(n5356) );
  XOR U8435 ( .A(n5359), .B(n5360), .Z(n5358) );
  XOR U8436 ( .A(DB[2999]), .B(DB[2992]), .Z(n5360) );
  AND U8437 ( .A(n338), .B(n5361), .Z(n5359) );
  XOR U8438 ( .A(n5362), .B(n5363), .Z(n5361) );
  XOR U8439 ( .A(DB[2992]), .B(DB[2985]), .Z(n5363) );
  AND U8440 ( .A(n342), .B(n5364), .Z(n5362) );
  XOR U8441 ( .A(n5365), .B(n5366), .Z(n5364) );
  XOR U8442 ( .A(DB[2985]), .B(DB[2978]), .Z(n5366) );
  AND U8443 ( .A(n346), .B(n5367), .Z(n5365) );
  XOR U8444 ( .A(n5368), .B(n5369), .Z(n5367) );
  XOR U8445 ( .A(DB[2978]), .B(DB[2971]), .Z(n5369) );
  AND U8446 ( .A(n350), .B(n5370), .Z(n5368) );
  XOR U8447 ( .A(n5371), .B(n5372), .Z(n5370) );
  XOR U8448 ( .A(DB[2971]), .B(DB[2964]), .Z(n5372) );
  AND U8449 ( .A(n354), .B(n5373), .Z(n5371) );
  XOR U8450 ( .A(n5374), .B(n5375), .Z(n5373) );
  XOR U8451 ( .A(DB[2964]), .B(DB[2957]), .Z(n5375) );
  AND U8452 ( .A(n358), .B(n5376), .Z(n5374) );
  XOR U8453 ( .A(n5377), .B(n5378), .Z(n5376) );
  XOR U8454 ( .A(DB[2957]), .B(DB[2950]), .Z(n5378) );
  AND U8455 ( .A(n362), .B(n5379), .Z(n5377) );
  XOR U8456 ( .A(n5380), .B(n5381), .Z(n5379) );
  XOR U8457 ( .A(DB[2950]), .B(DB[2943]), .Z(n5381) );
  AND U8458 ( .A(n366), .B(n5382), .Z(n5380) );
  XOR U8459 ( .A(n5383), .B(n5384), .Z(n5382) );
  XOR U8460 ( .A(DB[2943]), .B(DB[2936]), .Z(n5384) );
  AND U8461 ( .A(n370), .B(n5385), .Z(n5383) );
  XOR U8462 ( .A(n5386), .B(n5387), .Z(n5385) );
  XOR U8463 ( .A(DB[2936]), .B(DB[2929]), .Z(n5387) );
  AND U8464 ( .A(n374), .B(n5388), .Z(n5386) );
  XOR U8465 ( .A(n5389), .B(n5390), .Z(n5388) );
  XOR U8466 ( .A(DB[2929]), .B(DB[2922]), .Z(n5390) );
  AND U8467 ( .A(n378), .B(n5391), .Z(n5389) );
  XOR U8468 ( .A(n5392), .B(n5393), .Z(n5391) );
  XOR U8469 ( .A(DB[2922]), .B(DB[2915]), .Z(n5393) );
  AND U8470 ( .A(n382), .B(n5394), .Z(n5392) );
  XOR U8471 ( .A(n5395), .B(n5396), .Z(n5394) );
  XOR U8472 ( .A(DB[2915]), .B(DB[2908]), .Z(n5396) );
  AND U8473 ( .A(n386), .B(n5397), .Z(n5395) );
  XOR U8474 ( .A(n5398), .B(n5399), .Z(n5397) );
  XOR U8475 ( .A(DB[2908]), .B(DB[2901]), .Z(n5399) );
  AND U8476 ( .A(n390), .B(n5400), .Z(n5398) );
  XOR U8477 ( .A(n5401), .B(n5402), .Z(n5400) );
  XOR U8478 ( .A(DB[2901]), .B(DB[2894]), .Z(n5402) );
  AND U8479 ( .A(n394), .B(n5403), .Z(n5401) );
  XOR U8480 ( .A(n5404), .B(n5405), .Z(n5403) );
  XOR U8481 ( .A(DB[2894]), .B(DB[2887]), .Z(n5405) );
  AND U8482 ( .A(n398), .B(n5406), .Z(n5404) );
  XOR U8483 ( .A(n5407), .B(n5408), .Z(n5406) );
  XOR U8484 ( .A(DB[2887]), .B(DB[2880]), .Z(n5408) );
  AND U8485 ( .A(n402), .B(n5409), .Z(n5407) );
  XOR U8486 ( .A(n5410), .B(n5411), .Z(n5409) );
  XOR U8487 ( .A(DB[2880]), .B(DB[2873]), .Z(n5411) );
  AND U8488 ( .A(n406), .B(n5412), .Z(n5410) );
  XOR U8489 ( .A(n5413), .B(n5414), .Z(n5412) );
  XOR U8490 ( .A(DB[2873]), .B(DB[2866]), .Z(n5414) );
  AND U8491 ( .A(n410), .B(n5415), .Z(n5413) );
  XOR U8492 ( .A(n5416), .B(n5417), .Z(n5415) );
  XOR U8493 ( .A(DB[2866]), .B(DB[2859]), .Z(n5417) );
  AND U8494 ( .A(n414), .B(n5418), .Z(n5416) );
  XOR U8495 ( .A(n5419), .B(n5420), .Z(n5418) );
  XOR U8496 ( .A(DB[2859]), .B(DB[2852]), .Z(n5420) );
  AND U8497 ( .A(n418), .B(n5421), .Z(n5419) );
  XOR U8498 ( .A(n5422), .B(n5423), .Z(n5421) );
  XOR U8499 ( .A(DB[2852]), .B(DB[2845]), .Z(n5423) );
  AND U8500 ( .A(n422), .B(n5424), .Z(n5422) );
  XOR U8501 ( .A(n5425), .B(n5426), .Z(n5424) );
  XOR U8502 ( .A(DB[2845]), .B(DB[2838]), .Z(n5426) );
  AND U8503 ( .A(n426), .B(n5427), .Z(n5425) );
  XOR U8504 ( .A(n5428), .B(n5429), .Z(n5427) );
  XOR U8505 ( .A(DB[2838]), .B(DB[2831]), .Z(n5429) );
  AND U8506 ( .A(n430), .B(n5430), .Z(n5428) );
  XOR U8507 ( .A(n5431), .B(n5432), .Z(n5430) );
  XOR U8508 ( .A(DB[2831]), .B(DB[2824]), .Z(n5432) );
  AND U8509 ( .A(n434), .B(n5433), .Z(n5431) );
  XOR U8510 ( .A(n5434), .B(n5435), .Z(n5433) );
  XOR U8511 ( .A(DB[2824]), .B(DB[2817]), .Z(n5435) );
  AND U8512 ( .A(n438), .B(n5436), .Z(n5434) );
  XOR U8513 ( .A(n5437), .B(n5438), .Z(n5436) );
  XOR U8514 ( .A(DB[2817]), .B(DB[2810]), .Z(n5438) );
  AND U8515 ( .A(n442), .B(n5439), .Z(n5437) );
  XOR U8516 ( .A(n5440), .B(n5441), .Z(n5439) );
  XOR U8517 ( .A(DB[2810]), .B(DB[2803]), .Z(n5441) );
  AND U8518 ( .A(n446), .B(n5442), .Z(n5440) );
  XOR U8519 ( .A(n5443), .B(n5444), .Z(n5442) );
  XOR U8520 ( .A(DB[2803]), .B(DB[2796]), .Z(n5444) );
  AND U8521 ( .A(n450), .B(n5445), .Z(n5443) );
  XOR U8522 ( .A(n5446), .B(n5447), .Z(n5445) );
  XOR U8523 ( .A(DB[2796]), .B(DB[2789]), .Z(n5447) );
  AND U8524 ( .A(n454), .B(n5448), .Z(n5446) );
  XOR U8525 ( .A(n5449), .B(n5450), .Z(n5448) );
  XOR U8526 ( .A(DB[2789]), .B(DB[2782]), .Z(n5450) );
  AND U8527 ( .A(n458), .B(n5451), .Z(n5449) );
  XOR U8528 ( .A(n5452), .B(n5453), .Z(n5451) );
  XOR U8529 ( .A(DB[2782]), .B(DB[2775]), .Z(n5453) );
  AND U8530 ( .A(n462), .B(n5454), .Z(n5452) );
  XOR U8531 ( .A(n5455), .B(n5456), .Z(n5454) );
  XOR U8532 ( .A(DB[2775]), .B(DB[2768]), .Z(n5456) );
  AND U8533 ( .A(n466), .B(n5457), .Z(n5455) );
  XOR U8534 ( .A(n5458), .B(n5459), .Z(n5457) );
  XOR U8535 ( .A(DB[2768]), .B(DB[2761]), .Z(n5459) );
  AND U8536 ( .A(n470), .B(n5460), .Z(n5458) );
  XOR U8537 ( .A(n5461), .B(n5462), .Z(n5460) );
  XOR U8538 ( .A(DB[2761]), .B(DB[2754]), .Z(n5462) );
  AND U8539 ( .A(n474), .B(n5463), .Z(n5461) );
  XOR U8540 ( .A(n5464), .B(n5465), .Z(n5463) );
  XOR U8541 ( .A(DB[2754]), .B(DB[2747]), .Z(n5465) );
  AND U8542 ( .A(n478), .B(n5466), .Z(n5464) );
  XOR U8543 ( .A(n5467), .B(n5468), .Z(n5466) );
  XOR U8544 ( .A(DB[2747]), .B(DB[2740]), .Z(n5468) );
  AND U8545 ( .A(n482), .B(n5469), .Z(n5467) );
  XOR U8546 ( .A(n5470), .B(n5471), .Z(n5469) );
  XOR U8547 ( .A(DB[2740]), .B(DB[2733]), .Z(n5471) );
  AND U8548 ( .A(n486), .B(n5472), .Z(n5470) );
  XOR U8549 ( .A(n5473), .B(n5474), .Z(n5472) );
  XOR U8550 ( .A(DB[2733]), .B(DB[2726]), .Z(n5474) );
  AND U8551 ( .A(n490), .B(n5475), .Z(n5473) );
  XOR U8552 ( .A(n5476), .B(n5477), .Z(n5475) );
  XOR U8553 ( .A(DB[2726]), .B(DB[2719]), .Z(n5477) );
  AND U8554 ( .A(n494), .B(n5478), .Z(n5476) );
  XOR U8555 ( .A(n5479), .B(n5480), .Z(n5478) );
  XOR U8556 ( .A(DB[2719]), .B(DB[2712]), .Z(n5480) );
  AND U8557 ( .A(n498), .B(n5481), .Z(n5479) );
  XOR U8558 ( .A(n5482), .B(n5483), .Z(n5481) );
  XOR U8559 ( .A(DB[2712]), .B(DB[2705]), .Z(n5483) );
  AND U8560 ( .A(n502), .B(n5484), .Z(n5482) );
  XOR U8561 ( .A(n5485), .B(n5486), .Z(n5484) );
  XOR U8562 ( .A(DB[2705]), .B(DB[2698]), .Z(n5486) );
  AND U8563 ( .A(n506), .B(n5487), .Z(n5485) );
  XOR U8564 ( .A(n5488), .B(n5489), .Z(n5487) );
  XOR U8565 ( .A(DB[2698]), .B(DB[2691]), .Z(n5489) );
  AND U8566 ( .A(n510), .B(n5490), .Z(n5488) );
  XOR U8567 ( .A(n5491), .B(n5492), .Z(n5490) );
  XOR U8568 ( .A(DB[2691]), .B(DB[2684]), .Z(n5492) );
  AND U8569 ( .A(n514), .B(n5493), .Z(n5491) );
  XOR U8570 ( .A(n5494), .B(n5495), .Z(n5493) );
  XOR U8571 ( .A(DB[2684]), .B(DB[2677]), .Z(n5495) );
  AND U8572 ( .A(n518), .B(n5496), .Z(n5494) );
  XOR U8573 ( .A(n5497), .B(n5498), .Z(n5496) );
  XOR U8574 ( .A(DB[2677]), .B(DB[2670]), .Z(n5498) );
  AND U8575 ( .A(n522), .B(n5499), .Z(n5497) );
  XOR U8576 ( .A(n5500), .B(n5501), .Z(n5499) );
  XOR U8577 ( .A(DB[2670]), .B(DB[2663]), .Z(n5501) );
  AND U8578 ( .A(n526), .B(n5502), .Z(n5500) );
  XOR U8579 ( .A(n5503), .B(n5504), .Z(n5502) );
  XOR U8580 ( .A(DB[2663]), .B(DB[2656]), .Z(n5504) );
  AND U8581 ( .A(n530), .B(n5505), .Z(n5503) );
  XOR U8582 ( .A(n5506), .B(n5507), .Z(n5505) );
  XOR U8583 ( .A(DB[2656]), .B(DB[2649]), .Z(n5507) );
  AND U8584 ( .A(n534), .B(n5508), .Z(n5506) );
  XOR U8585 ( .A(n5509), .B(n5510), .Z(n5508) );
  XOR U8586 ( .A(DB[2649]), .B(DB[2642]), .Z(n5510) );
  AND U8587 ( .A(n538), .B(n5511), .Z(n5509) );
  XOR U8588 ( .A(n5512), .B(n5513), .Z(n5511) );
  XOR U8589 ( .A(DB[2642]), .B(DB[2635]), .Z(n5513) );
  AND U8590 ( .A(n542), .B(n5514), .Z(n5512) );
  XOR U8591 ( .A(n5515), .B(n5516), .Z(n5514) );
  XOR U8592 ( .A(DB[2635]), .B(DB[2628]), .Z(n5516) );
  AND U8593 ( .A(n546), .B(n5517), .Z(n5515) );
  XOR U8594 ( .A(n5518), .B(n5519), .Z(n5517) );
  XOR U8595 ( .A(DB[2628]), .B(DB[2621]), .Z(n5519) );
  AND U8596 ( .A(n550), .B(n5520), .Z(n5518) );
  XOR U8597 ( .A(n5521), .B(n5522), .Z(n5520) );
  XOR U8598 ( .A(DB[2621]), .B(DB[2614]), .Z(n5522) );
  AND U8599 ( .A(n554), .B(n5523), .Z(n5521) );
  XOR U8600 ( .A(n5524), .B(n5525), .Z(n5523) );
  XOR U8601 ( .A(DB[2614]), .B(DB[2607]), .Z(n5525) );
  AND U8602 ( .A(n558), .B(n5526), .Z(n5524) );
  XOR U8603 ( .A(n5527), .B(n5528), .Z(n5526) );
  XOR U8604 ( .A(DB[2607]), .B(DB[2600]), .Z(n5528) );
  AND U8605 ( .A(n562), .B(n5529), .Z(n5527) );
  XOR U8606 ( .A(n5530), .B(n5531), .Z(n5529) );
  XOR U8607 ( .A(DB[2600]), .B(DB[2593]), .Z(n5531) );
  AND U8608 ( .A(n566), .B(n5532), .Z(n5530) );
  XOR U8609 ( .A(n5533), .B(n5534), .Z(n5532) );
  XOR U8610 ( .A(DB[2593]), .B(DB[2586]), .Z(n5534) );
  AND U8611 ( .A(n570), .B(n5535), .Z(n5533) );
  XOR U8612 ( .A(n5536), .B(n5537), .Z(n5535) );
  XOR U8613 ( .A(DB[2586]), .B(DB[2579]), .Z(n5537) );
  AND U8614 ( .A(n574), .B(n5538), .Z(n5536) );
  XOR U8615 ( .A(n5539), .B(n5540), .Z(n5538) );
  XOR U8616 ( .A(DB[2579]), .B(DB[2572]), .Z(n5540) );
  AND U8617 ( .A(n578), .B(n5541), .Z(n5539) );
  XOR U8618 ( .A(n5542), .B(n5543), .Z(n5541) );
  XOR U8619 ( .A(DB[2572]), .B(DB[2565]), .Z(n5543) );
  AND U8620 ( .A(n582), .B(n5544), .Z(n5542) );
  XOR U8621 ( .A(n5545), .B(n5546), .Z(n5544) );
  XOR U8622 ( .A(DB[2565]), .B(DB[2558]), .Z(n5546) );
  AND U8623 ( .A(n586), .B(n5547), .Z(n5545) );
  XOR U8624 ( .A(n5548), .B(n5549), .Z(n5547) );
  XOR U8625 ( .A(DB[2558]), .B(DB[2551]), .Z(n5549) );
  AND U8626 ( .A(n590), .B(n5550), .Z(n5548) );
  XOR U8627 ( .A(n5551), .B(n5552), .Z(n5550) );
  XOR U8628 ( .A(DB[2551]), .B(DB[2544]), .Z(n5552) );
  AND U8629 ( .A(n594), .B(n5553), .Z(n5551) );
  XOR U8630 ( .A(n5554), .B(n5555), .Z(n5553) );
  XOR U8631 ( .A(DB[2544]), .B(DB[2537]), .Z(n5555) );
  AND U8632 ( .A(n598), .B(n5556), .Z(n5554) );
  XOR U8633 ( .A(n5557), .B(n5558), .Z(n5556) );
  XOR U8634 ( .A(DB[2537]), .B(DB[2530]), .Z(n5558) );
  AND U8635 ( .A(n602), .B(n5559), .Z(n5557) );
  XOR U8636 ( .A(n5560), .B(n5561), .Z(n5559) );
  XOR U8637 ( .A(DB[2530]), .B(DB[2523]), .Z(n5561) );
  AND U8638 ( .A(n606), .B(n5562), .Z(n5560) );
  XOR U8639 ( .A(n5563), .B(n5564), .Z(n5562) );
  XOR U8640 ( .A(DB[2523]), .B(DB[2516]), .Z(n5564) );
  AND U8641 ( .A(n610), .B(n5565), .Z(n5563) );
  XOR U8642 ( .A(n5566), .B(n5567), .Z(n5565) );
  XOR U8643 ( .A(DB[2516]), .B(DB[2509]), .Z(n5567) );
  AND U8644 ( .A(n614), .B(n5568), .Z(n5566) );
  XOR U8645 ( .A(n5569), .B(n5570), .Z(n5568) );
  XOR U8646 ( .A(DB[2509]), .B(DB[2502]), .Z(n5570) );
  AND U8647 ( .A(n618), .B(n5571), .Z(n5569) );
  XOR U8648 ( .A(n5572), .B(n5573), .Z(n5571) );
  XOR U8649 ( .A(DB[2502]), .B(DB[2495]), .Z(n5573) );
  AND U8650 ( .A(n622), .B(n5574), .Z(n5572) );
  XOR U8651 ( .A(n5575), .B(n5576), .Z(n5574) );
  XOR U8652 ( .A(DB[2495]), .B(DB[2488]), .Z(n5576) );
  AND U8653 ( .A(n626), .B(n5577), .Z(n5575) );
  XOR U8654 ( .A(n5578), .B(n5579), .Z(n5577) );
  XOR U8655 ( .A(DB[2488]), .B(DB[2481]), .Z(n5579) );
  AND U8656 ( .A(n630), .B(n5580), .Z(n5578) );
  XOR U8657 ( .A(n5581), .B(n5582), .Z(n5580) );
  XOR U8658 ( .A(DB[2481]), .B(DB[2474]), .Z(n5582) );
  AND U8659 ( .A(n634), .B(n5583), .Z(n5581) );
  XOR U8660 ( .A(n5584), .B(n5585), .Z(n5583) );
  XOR U8661 ( .A(DB[2474]), .B(DB[2467]), .Z(n5585) );
  AND U8662 ( .A(n638), .B(n5586), .Z(n5584) );
  XOR U8663 ( .A(n5587), .B(n5588), .Z(n5586) );
  XOR U8664 ( .A(DB[2467]), .B(DB[2460]), .Z(n5588) );
  AND U8665 ( .A(n642), .B(n5589), .Z(n5587) );
  XOR U8666 ( .A(n5590), .B(n5591), .Z(n5589) );
  XOR U8667 ( .A(DB[2460]), .B(DB[2453]), .Z(n5591) );
  AND U8668 ( .A(n646), .B(n5592), .Z(n5590) );
  XOR U8669 ( .A(n5593), .B(n5594), .Z(n5592) );
  XOR U8670 ( .A(DB[2453]), .B(DB[2446]), .Z(n5594) );
  AND U8671 ( .A(n650), .B(n5595), .Z(n5593) );
  XOR U8672 ( .A(n5596), .B(n5597), .Z(n5595) );
  XOR U8673 ( .A(DB[2446]), .B(DB[2439]), .Z(n5597) );
  AND U8674 ( .A(n654), .B(n5598), .Z(n5596) );
  XOR U8675 ( .A(n5599), .B(n5600), .Z(n5598) );
  XOR U8676 ( .A(DB[2439]), .B(DB[2432]), .Z(n5600) );
  AND U8677 ( .A(n658), .B(n5601), .Z(n5599) );
  XOR U8678 ( .A(n5602), .B(n5603), .Z(n5601) );
  XOR U8679 ( .A(DB[2432]), .B(DB[2425]), .Z(n5603) );
  AND U8680 ( .A(n662), .B(n5604), .Z(n5602) );
  XOR U8681 ( .A(n5605), .B(n5606), .Z(n5604) );
  XOR U8682 ( .A(DB[2425]), .B(DB[2418]), .Z(n5606) );
  AND U8683 ( .A(n666), .B(n5607), .Z(n5605) );
  XOR U8684 ( .A(n5608), .B(n5609), .Z(n5607) );
  XOR U8685 ( .A(DB[2418]), .B(DB[2411]), .Z(n5609) );
  AND U8686 ( .A(n670), .B(n5610), .Z(n5608) );
  XOR U8687 ( .A(n5611), .B(n5612), .Z(n5610) );
  XOR U8688 ( .A(DB[2411]), .B(DB[2404]), .Z(n5612) );
  AND U8689 ( .A(n674), .B(n5613), .Z(n5611) );
  XOR U8690 ( .A(n5614), .B(n5615), .Z(n5613) );
  XOR U8691 ( .A(DB[2404]), .B(DB[2397]), .Z(n5615) );
  AND U8692 ( .A(n678), .B(n5616), .Z(n5614) );
  XOR U8693 ( .A(n5617), .B(n5618), .Z(n5616) );
  XOR U8694 ( .A(DB[2397]), .B(DB[2390]), .Z(n5618) );
  AND U8695 ( .A(n682), .B(n5619), .Z(n5617) );
  XOR U8696 ( .A(n5620), .B(n5621), .Z(n5619) );
  XOR U8697 ( .A(DB[2390]), .B(DB[2383]), .Z(n5621) );
  AND U8698 ( .A(n686), .B(n5622), .Z(n5620) );
  XOR U8699 ( .A(n5623), .B(n5624), .Z(n5622) );
  XOR U8700 ( .A(DB[2383]), .B(DB[2376]), .Z(n5624) );
  AND U8701 ( .A(n690), .B(n5625), .Z(n5623) );
  XOR U8702 ( .A(n5626), .B(n5627), .Z(n5625) );
  XOR U8703 ( .A(DB[2376]), .B(DB[2369]), .Z(n5627) );
  AND U8704 ( .A(n694), .B(n5628), .Z(n5626) );
  XOR U8705 ( .A(n5629), .B(n5630), .Z(n5628) );
  XOR U8706 ( .A(DB[2369]), .B(DB[2362]), .Z(n5630) );
  AND U8707 ( .A(n698), .B(n5631), .Z(n5629) );
  XOR U8708 ( .A(n5632), .B(n5633), .Z(n5631) );
  XOR U8709 ( .A(DB[2362]), .B(DB[2355]), .Z(n5633) );
  AND U8710 ( .A(n702), .B(n5634), .Z(n5632) );
  XOR U8711 ( .A(n5635), .B(n5636), .Z(n5634) );
  XOR U8712 ( .A(DB[2355]), .B(DB[2348]), .Z(n5636) );
  AND U8713 ( .A(n706), .B(n5637), .Z(n5635) );
  XOR U8714 ( .A(n5638), .B(n5639), .Z(n5637) );
  XOR U8715 ( .A(DB[2348]), .B(DB[2341]), .Z(n5639) );
  AND U8716 ( .A(n710), .B(n5640), .Z(n5638) );
  XOR U8717 ( .A(n5641), .B(n5642), .Z(n5640) );
  XOR U8718 ( .A(DB[2341]), .B(DB[2334]), .Z(n5642) );
  AND U8719 ( .A(n714), .B(n5643), .Z(n5641) );
  XOR U8720 ( .A(n5644), .B(n5645), .Z(n5643) );
  XOR U8721 ( .A(DB[2334]), .B(DB[2327]), .Z(n5645) );
  AND U8722 ( .A(n718), .B(n5646), .Z(n5644) );
  XOR U8723 ( .A(n5647), .B(n5648), .Z(n5646) );
  XOR U8724 ( .A(DB[2327]), .B(DB[2320]), .Z(n5648) );
  AND U8725 ( .A(n722), .B(n5649), .Z(n5647) );
  XOR U8726 ( .A(n5650), .B(n5651), .Z(n5649) );
  XOR U8727 ( .A(DB[2320]), .B(DB[2313]), .Z(n5651) );
  AND U8728 ( .A(n726), .B(n5652), .Z(n5650) );
  XOR U8729 ( .A(n5653), .B(n5654), .Z(n5652) );
  XOR U8730 ( .A(DB[2313]), .B(DB[2306]), .Z(n5654) );
  AND U8731 ( .A(n730), .B(n5655), .Z(n5653) );
  XOR U8732 ( .A(n5656), .B(n5657), .Z(n5655) );
  XOR U8733 ( .A(DB[2306]), .B(DB[2299]), .Z(n5657) );
  AND U8734 ( .A(n734), .B(n5658), .Z(n5656) );
  XOR U8735 ( .A(n5659), .B(n5660), .Z(n5658) );
  XOR U8736 ( .A(DB[2299]), .B(DB[2292]), .Z(n5660) );
  AND U8737 ( .A(n738), .B(n5661), .Z(n5659) );
  XOR U8738 ( .A(n5662), .B(n5663), .Z(n5661) );
  XOR U8739 ( .A(DB[2292]), .B(DB[2285]), .Z(n5663) );
  AND U8740 ( .A(n742), .B(n5664), .Z(n5662) );
  XOR U8741 ( .A(n5665), .B(n5666), .Z(n5664) );
  XOR U8742 ( .A(DB[2285]), .B(DB[2278]), .Z(n5666) );
  AND U8743 ( .A(n746), .B(n5667), .Z(n5665) );
  XOR U8744 ( .A(n5668), .B(n5669), .Z(n5667) );
  XOR U8745 ( .A(DB[2278]), .B(DB[2271]), .Z(n5669) );
  AND U8746 ( .A(n750), .B(n5670), .Z(n5668) );
  XOR U8747 ( .A(n5671), .B(n5672), .Z(n5670) );
  XOR U8748 ( .A(DB[2271]), .B(DB[2264]), .Z(n5672) );
  AND U8749 ( .A(n754), .B(n5673), .Z(n5671) );
  XOR U8750 ( .A(n5674), .B(n5675), .Z(n5673) );
  XOR U8751 ( .A(DB[2264]), .B(DB[2257]), .Z(n5675) );
  AND U8752 ( .A(n758), .B(n5676), .Z(n5674) );
  XOR U8753 ( .A(n5677), .B(n5678), .Z(n5676) );
  XOR U8754 ( .A(DB[2257]), .B(DB[2250]), .Z(n5678) );
  AND U8755 ( .A(n762), .B(n5679), .Z(n5677) );
  XOR U8756 ( .A(n5680), .B(n5681), .Z(n5679) );
  XOR U8757 ( .A(DB[2250]), .B(DB[2243]), .Z(n5681) );
  AND U8758 ( .A(n766), .B(n5682), .Z(n5680) );
  XOR U8759 ( .A(n5683), .B(n5684), .Z(n5682) );
  XOR U8760 ( .A(DB[2243]), .B(DB[2236]), .Z(n5684) );
  AND U8761 ( .A(n770), .B(n5685), .Z(n5683) );
  XOR U8762 ( .A(n5686), .B(n5687), .Z(n5685) );
  XOR U8763 ( .A(DB[2236]), .B(DB[2229]), .Z(n5687) );
  AND U8764 ( .A(n774), .B(n5688), .Z(n5686) );
  XOR U8765 ( .A(n5689), .B(n5690), .Z(n5688) );
  XOR U8766 ( .A(DB[2229]), .B(DB[2222]), .Z(n5690) );
  AND U8767 ( .A(n778), .B(n5691), .Z(n5689) );
  XOR U8768 ( .A(n5692), .B(n5693), .Z(n5691) );
  XOR U8769 ( .A(DB[2222]), .B(DB[2215]), .Z(n5693) );
  AND U8770 ( .A(n782), .B(n5694), .Z(n5692) );
  XOR U8771 ( .A(n5695), .B(n5696), .Z(n5694) );
  XOR U8772 ( .A(DB[2215]), .B(DB[2208]), .Z(n5696) );
  AND U8773 ( .A(n786), .B(n5697), .Z(n5695) );
  XOR U8774 ( .A(n5698), .B(n5699), .Z(n5697) );
  XOR U8775 ( .A(DB[2208]), .B(DB[2201]), .Z(n5699) );
  AND U8776 ( .A(n790), .B(n5700), .Z(n5698) );
  XOR U8777 ( .A(n5701), .B(n5702), .Z(n5700) );
  XOR U8778 ( .A(DB[2201]), .B(DB[2194]), .Z(n5702) );
  AND U8779 ( .A(n794), .B(n5703), .Z(n5701) );
  XOR U8780 ( .A(n5704), .B(n5705), .Z(n5703) );
  XOR U8781 ( .A(DB[2194]), .B(DB[2187]), .Z(n5705) );
  AND U8782 ( .A(n798), .B(n5706), .Z(n5704) );
  XOR U8783 ( .A(n5707), .B(n5708), .Z(n5706) );
  XOR U8784 ( .A(DB[2187]), .B(DB[2180]), .Z(n5708) );
  AND U8785 ( .A(n802), .B(n5709), .Z(n5707) );
  XOR U8786 ( .A(n5710), .B(n5711), .Z(n5709) );
  XOR U8787 ( .A(DB[2180]), .B(DB[2173]), .Z(n5711) );
  AND U8788 ( .A(n806), .B(n5712), .Z(n5710) );
  XOR U8789 ( .A(n5713), .B(n5714), .Z(n5712) );
  XOR U8790 ( .A(DB[2173]), .B(DB[2166]), .Z(n5714) );
  AND U8791 ( .A(n810), .B(n5715), .Z(n5713) );
  XOR U8792 ( .A(n5716), .B(n5717), .Z(n5715) );
  XOR U8793 ( .A(DB[2166]), .B(DB[2159]), .Z(n5717) );
  AND U8794 ( .A(n814), .B(n5718), .Z(n5716) );
  XOR U8795 ( .A(n5719), .B(n5720), .Z(n5718) );
  XOR U8796 ( .A(DB[2159]), .B(DB[2152]), .Z(n5720) );
  AND U8797 ( .A(n818), .B(n5721), .Z(n5719) );
  XOR U8798 ( .A(n5722), .B(n5723), .Z(n5721) );
  XOR U8799 ( .A(DB[2152]), .B(DB[2145]), .Z(n5723) );
  AND U8800 ( .A(n822), .B(n5724), .Z(n5722) );
  XOR U8801 ( .A(n5725), .B(n5726), .Z(n5724) );
  XOR U8802 ( .A(DB[2145]), .B(DB[2138]), .Z(n5726) );
  AND U8803 ( .A(n826), .B(n5727), .Z(n5725) );
  XOR U8804 ( .A(n5728), .B(n5729), .Z(n5727) );
  XOR U8805 ( .A(DB[2138]), .B(DB[2131]), .Z(n5729) );
  AND U8806 ( .A(n830), .B(n5730), .Z(n5728) );
  XOR U8807 ( .A(n5731), .B(n5732), .Z(n5730) );
  XOR U8808 ( .A(DB[2131]), .B(DB[2124]), .Z(n5732) );
  AND U8809 ( .A(n834), .B(n5733), .Z(n5731) );
  XOR U8810 ( .A(n5734), .B(n5735), .Z(n5733) );
  XOR U8811 ( .A(DB[2124]), .B(DB[2117]), .Z(n5735) );
  AND U8812 ( .A(n838), .B(n5736), .Z(n5734) );
  XOR U8813 ( .A(n5737), .B(n5738), .Z(n5736) );
  XOR U8814 ( .A(DB[2117]), .B(DB[2110]), .Z(n5738) );
  AND U8815 ( .A(n842), .B(n5739), .Z(n5737) );
  XOR U8816 ( .A(n5740), .B(n5741), .Z(n5739) );
  XOR U8817 ( .A(DB[2110]), .B(DB[2103]), .Z(n5741) );
  AND U8818 ( .A(n846), .B(n5742), .Z(n5740) );
  XOR U8819 ( .A(n5743), .B(n5744), .Z(n5742) );
  XOR U8820 ( .A(DB[2103]), .B(DB[2096]), .Z(n5744) );
  AND U8821 ( .A(n850), .B(n5745), .Z(n5743) );
  XOR U8822 ( .A(n5746), .B(n5747), .Z(n5745) );
  XOR U8823 ( .A(DB[2096]), .B(DB[2089]), .Z(n5747) );
  AND U8824 ( .A(n854), .B(n5748), .Z(n5746) );
  XOR U8825 ( .A(n5749), .B(n5750), .Z(n5748) );
  XOR U8826 ( .A(DB[2089]), .B(DB[2082]), .Z(n5750) );
  AND U8827 ( .A(n858), .B(n5751), .Z(n5749) );
  XOR U8828 ( .A(n5752), .B(n5753), .Z(n5751) );
  XOR U8829 ( .A(DB[2082]), .B(DB[2075]), .Z(n5753) );
  AND U8830 ( .A(n862), .B(n5754), .Z(n5752) );
  XOR U8831 ( .A(n5755), .B(n5756), .Z(n5754) );
  XOR U8832 ( .A(DB[2075]), .B(DB[2068]), .Z(n5756) );
  AND U8833 ( .A(n866), .B(n5757), .Z(n5755) );
  XOR U8834 ( .A(n5758), .B(n5759), .Z(n5757) );
  XOR U8835 ( .A(DB[2068]), .B(DB[2061]), .Z(n5759) );
  AND U8836 ( .A(n870), .B(n5760), .Z(n5758) );
  XOR U8837 ( .A(n5761), .B(n5762), .Z(n5760) );
  XOR U8838 ( .A(DB[2061]), .B(DB[2054]), .Z(n5762) );
  AND U8839 ( .A(n874), .B(n5763), .Z(n5761) );
  XOR U8840 ( .A(n5764), .B(n5765), .Z(n5763) );
  XOR U8841 ( .A(DB[2054]), .B(DB[2047]), .Z(n5765) );
  AND U8842 ( .A(n878), .B(n5766), .Z(n5764) );
  XOR U8843 ( .A(n5767), .B(n5768), .Z(n5766) );
  XOR U8844 ( .A(DB[2047]), .B(DB[2040]), .Z(n5768) );
  AND U8845 ( .A(n882), .B(n5769), .Z(n5767) );
  XOR U8846 ( .A(n5770), .B(n5771), .Z(n5769) );
  XOR U8847 ( .A(DB[2040]), .B(DB[2033]), .Z(n5771) );
  AND U8848 ( .A(n886), .B(n5772), .Z(n5770) );
  XOR U8849 ( .A(n5773), .B(n5774), .Z(n5772) );
  XOR U8850 ( .A(DB[2033]), .B(DB[2026]), .Z(n5774) );
  AND U8851 ( .A(n890), .B(n5775), .Z(n5773) );
  XOR U8852 ( .A(n5776), .B(n5777), .Z(n5775) );
  XOR U8853 ( .A(DB[2026]), .B(DB[2019]), .Z(n5777) );
  AND U8854 ( .A(n894), .B(n5778), .Z(n5776) );
  XOR U8855 ( .A(n5779), .B(n5780), .Z(n5778) );
  XOR U8856 ( .A(DB[2019]), .B(DB[2012]), .Z(n5780) );
  AND U8857 ( .A(n898), .B(n5781), .Z(n5779) );
  XOR U8858 ( .A(n5782), .B(n5783), .Z(n5781) );
  XOR U8859 ( .A(DB[2012]), .B(DB[2005]), .Z(n5783) );
  AND U8860 ( .A(n902), .B(n5784), .Z(n5782) );
  XOR U8861 ( .A(n5785), .B(n5786), .Z(n5784) );
  XOR U8862 ( .A(DB[2005]), .B(DB[1998]), .Z(n5786) );
  AND U8863 ( .A(n906), .B(n5787), .Z(n5785) );
  XOR U8864 ( .A(n5788), .B(n5789), .Z(n5787) );
  XOR U8865 ( .A(DB[1998]), .B(DB[1991]), .Z(n5789) );
  AND U8866 ( .A(n910), .B(n5790), .Z(n5788) );
  XOR U8867 ( .A(n5791), .B(n5792), .Z(n5790) );
  XOR U8868 ( .A(DB[1991]), .B(DB[1984]), .Z(n5792) );
  AND U8869 ( .A(n914), .B(n5793), .Z(n5791) );
  XOR U8870 ( .A(n5794), .B(n5795), .Z(n5793) );
  XOR U8871 ( .A(DB[1984]), .B(DB[1977]), .Z(n5795) );
  AND U8872 ( .A(n918), .B(n5796), .Z(n5794) );
  XOR U8873 ( .A(n5797), .B(n5798), .Z(n5796) );
  XOR U8874 ( .A(DB[1977]), .B(DB[1970]), .Z(n5798) );
  AND U8875 ( .A(n922), .B(n5799), .Z(n5797) );
  XOR U8876 ( .A(n5800), .B(n5801), .Z(n5799) );
  XOR U8877 ( .A(DB[1970]), .B(DB[1963]), .Z(n5801) );
  AND U8878 ( .A(n926), .B(n5802), .Z(n5800) );
  XOR U8879 ( .A(n5803), .B(n5804), .Z(n5802) );
  XOR U8880 ( .A(DB[1963]), .B(DB[1956]), .Z(n5804) );
  AND U8881 ( .A(n930), .B(n5805), .Z(n5803) );
  XOR U8882 ( .A(n5806), .B(n5807), .Z(n5805) );
  XOR U8883 ( .A(DB[1956]), .B(DB[1949]), .Z(n5807) );
  AND U8884 ( .A(n934), .B(n5808), .Z(n5806) );
  XOR U8885 ( .A(n5809), .B(n5810), .Z(n5808) );
  XOR U8886 ( .A(DB[1949]), .B(DB[1942]), .Z(n5810) );
  AND U8887 ( .A(n938), .B(n5811), .Z(n5809) );
  XOR U8888 ( .A(n5812), .B(n5813), .Z(n5811) );
  XOR U8889 ( .A(DB[1942]), .B(DB[1935]), .Z(n5813) );
  AND U8890 ( .A(n942), .B(n5814), .Z(n5812) );
  XOR U8891 ( .A(n5815), .B(n5816), .Z(n5814) );
  XOR U8892 ( .A(DB[1935]), .B(DB[1928]), .Z(n5816) );
  AND U8893 ( .A(n946), .B(n5817), .Z(n5815) );
  XOR U8894 ( .A(n5818), .B(n5819), .Z(n5817) );
  XOR U8895 ( .A(DB[1928]), .B(DB[1921]), .Z(n5819) );
  AND U8896 ( .A(n950), .B(n5820), .Z(n5818) );
  XOR U8897 ( .A(n5821), .B(n5822), .Z(n5820) );
  XOR U8898 ( .A(DB[1921]), .B(DB[1914]), .Z(n5822) );
  AND U8899 ( .A(n954), .B(n5823), .Z(n5821) );
  XOR U8900 ( .A(n5824), .B(n5825), .Z(n5823) );
  XOR U8901 ( .A(DB[1914]), .B(DB[1907]), .Z(n5825) );
  AND U8902 ( .A(n958), .B(n5826), .Z(n5824) );
  XOR U8903 ( .A(n5827), .B(n5828), .Z(n5826) );
  XOR U8904 ( .A(DB[1907]), .B(DB[1900]), .Z(n5828) );
  AND U8905 ( .A(n962), .B(n5829), .Z(n5827) );
  XOR U8906 ( .A(n5830), .B(n5831), .Z(n5829) );
  XOR U8907 ( .A(DB[1900]), .B(DB[1893]), .Z(n5831) );
  AND U8908 ( .A(n966), .B(n5832), .Z(n5830) );
  XOR U8909 ( .A(n5833), .B(n5834), .Z(n5832) );
  XOR U8910 ( .A(DB[1893]), .B(DB[1886]), .Z(n5834) );
  AND U8911 ( .A(n970), .B(n5835), .Z(n5833) );
  XOR U8912 ( .A(n5836), .B(n5837), .Z(n5835) );
  XOR U8913 ( .A(DB[1886]), .B(DB[1879]), .Z(n5837) );
  AND U8914 ( .A(n974), .B(n5838), .Z(n5836) );
  XOR U8915 ( .A(n5839), .B(n5840), .Z(n5838) );
  XOR U8916 ( .A(DB[1879]), .B(DB[1872]), .Z(n5840) );
  AND U8917 ( .A(n978), .B(n5841), .Z(n5839) );
  XOR U8918 ( .A(n5842), .B(n5843), .Z(n5841) );
  XOR U8919 ( .A(DB[1872]), .B(DB[1865]), .Z(n5843) );
  AND U8920 ( .A(n982), .B(n5844), .Z(n5842) );
  XOR U8921 ( .A(n5845), .B(n5846), .Z(n5844) );
  XOR U8922 ( .A(DB[1865]), .B(DB[1858]), .Z(n5846) );
  AND U8923 ( .A(n986), .B(n5847), .Z(n5845) );
  XOR U8924 ( .A(n5848), .B(n5849), .Z(n5847) );
  XOR U8925 ( .A(DB[1858]), .B(DB[1851]), .Z(n5849) );
  AND U8926 ( .A(n990), .B(n5850), .Z(n5848) );
  XOR U8927 ( .A(n5851), .B(n5852), .Z(n5850) );
  XOR U8928 ( .A(DB[1851]), .B(DB[1844]), .Z(n5852) );
  AND U8929 ( .A(n994), .B(n5853), .Z(n5851) );
  XOR U8930 ( .A(n5854), .B(n5855), .Z(n5853) );
  XOR U8931 ( .A(DB[1844]), .B(DB[1837]), .Z(n5855) );
  AND U8932 ( .A(n998), .B(n5856), .Z(n5854) );
  XOR U8933 ( .A(n5857), .B(n5858), .Z(n5856) );
  XOR U8934 ( .A(DB[1837]), .B(DB[1830]), .Z(n5858) );
  AND U8935 ( .A(n1002), .B(n5859), .Z(n5857) );
  XOR U8936 ( .A(n5860), .B(n5861), .Z(n5859) );
  XOR U8937 ( .A(DB[1830]), .B(DB[1823]), .Z(n5861) );
  AND U8938 ( .A(n1006), .B(n5862), .Z(n5860) );
  XOR U8939 ( .A(n5863), .B(n5864), .Z(n5862) );
  XOR U8940 ( .A(DB[1823]), .B(DB[1816]), .Z(n5864) );
  AND U8941 ( .A(n1010), .B(n5865), .Z(n5863) );
  XOR U8942 ( .A(n5866), .B(n5867), .Z(n5865) );
  XOR U8943 ( .A(DB[1816]), .B(DB[1809]), .Z(n5867) );
  AND U8944 ( .A(n1014), .B(n5868), .Z(n5866) );
  XOR U8945 ( .A(n5869), .B(n5870), .Z(n5868) );
  XOR U8946 ( .A(DB[1809]), .B(DB[1802]), .Z(n5870) );
  AND U8947 ( .A(n1018), .B(n5871), .Z(n5869) );
  XOR U8948 ( .A(n5872), .B(n5873), .Z(n5871) );
  XOR U8949 ( .A(DB[1802]), .B(DB[1795]), .Z(n5873) );
  AND U8950 ( .A(n1022), .B(n5874), .Z(n5872) );
  XOR U8951 ( .A(n5875), .B(n5876), .Z(n5874) );
  XOR U8952 ( .A(DB[1795]), .B(DB[1788]), .Z(n5876) );
  AND U8953 ( .A(n1026), .B(n5877), .Z(n5875) );
  XOR U8954 ( .A(n5878), .B(n5879), .Z(n5877) );
  XOR U8955 ( .A(DB[1788]), .B(DB[1781]), .Z(n5879) );
  AND U8956 ( .A(n1030), .B(n5880), .Z(n5878) );
  XOR U8957 ( .A(n5881), .B(n5882), .Z(n5880) );
  XOR U8958 ( .A(DB[1781]), .B(DB[1774]), .Z(n5882) );
  AND U8959 ( .A(n1034), .B(n5883), .Z(n5881) );
  XOR U8960 ( .A(n5884), .B(n5885), .Z(n5883) );
  XOR U8961 ( .A(DB[1774]), .B(DB[1767]), .Z(n5885) );
  AND U8962 ( .A(n1038), .B(n5886), .Z(n5884) );
  XOR U8963 ( .A(n5887), .B(n5888), .Z(n5886) );
  XOR U8964 ( .A(DB[1767]), .B(DB[1760]), .Z(n5888) );
  AND U8965 ( .A(n1042), .B(n5889), .Z(n5887) );
  XOR U8966 ( .A(n5890), .B(n5891), .Z(n5889) );
  XOR U8967 ( .A(DB[1760]), .B(DB[1753]), .Z(n5891) );
  AND U8968 ( .A(n1046), .B(n5892), .Z(n5890) );
  XOR U8969 ( .A(n5893), .B(n5894), .Z(n5892) );
  XOR U8970 ( .A(DB[1753]), .B(DB[1746]), .Z(n5894) );
  AND U8971 ( .A(n1050), .B(n5895), .Z(n5893) );
  XOR U8972 ( .A(n5896), .B(n5897), .Z(n5895) );
  XOR U8973 ( .A(DB[1746]), .B(DB[1739]), .Z(n5897) );
  AND U8974 ( .A(n1054), .B(n5898), .Z(n5896) );
  XOR U8975 ( .A(n5899), .B(n5900), .Z(n5898) );
  XOR U8976 ( .A(DB[1739]), .B(DB[1732]), .Z(n5900) );
  AND U8977 ( .A(n1058), .B(n5901), .Z(n5899) );
  XOR U8978 ( .A(n5902), .B(n5903), .Z(n5901) );
  XOR U8979 ( .A(DB[1732]), .B(DB[1725]), .Z(n5903) );
  AND U8980 ( .A(n1062), .B(n5904), .Z(n5902) );
  XOR U8981 ( .A(n5905), .B(n5906), .Z(n5904) );
  XOR U8982 ( .A(DB[1725]), .B(DB[1718]), .Z(n5906) );
  AND U8983 ( .A(n1066), .B(n5907), .Z(n5905) );
  XOR U8984 ( .A(n5908), .B(n5909), .Z(n5907) );
  XOR U8985 ( .A(DB[1718]), .B(DB[1711]), .Z(n5909) );
  AND U8986 ( .A(n1070), .B(n5910), .Z(n5908) );
  XOR U8987 ( .A(n5911), .B(n5912), .Z(n5910) );
  XOR U8988 ( .A(DB[1711]), .B(DB[1704]), .Z(n5912) );
  AND U8989 ( .A(n1074), .B(n5913), .Z(n5911) );
  XOR U8990 ( .A(n5914), .B(n5915), .Z(n5913) );
  XOR U8991 ( .A(DB[1704]), .B(DB[1697]), .Z(n5915) );
  AND U8992 ( .A(n1078), .B(n5916), .Z(n5914) );
  XOR U8993 ( .A(n5917), .B(n5918), .Z(n5916) );
  XOR U8994 ( .A(DB[1697]), .B(DB[1690]), .Z(n5918) );
  AND U8995 ( .A(n1082), .B(n5919), .Z(n5917) );
  XOR U8996 ( .A(n5920), .B(n5921), .Z(n5919) );
  XOR U8997 ( .A(DB[1690]), .B(DB[1683]), .Z(n5921) );
  AND U8998 ( .A(n1086), .B(n5922), .Z(n5920) );
  XOR U8999 ( .A(n5923), .B(n5924), .Z(n5922) );
  XOR U9000 ( .A(DB[1683]), .B(DB[1676]), .Z(n5924) );
  AND U9001 ( .A(n1090), .B(n5925), .Z(n5923) );
  XOR U9002 ( .A(n5926), .B(n5927), .Z(n5925) );
  XOR U9003 ( .A(DB[1676]), .B(DB[1669]), .Z(n5927) );
  AND U9004 ( .A(n1094), .B(n5928), .Z(n5926) );
  XOR U9005 ( .A(n5929), .B(n5930), .Z(n5928) );
  XOR U9006 ( .A(DB[1669]), .B(DB[1662]), .Z(n5930) );
  AND U9007 ( .A(n1098), .B(n5931), .Z(n5929) );
  XOR U9008 ( .A(n5932), .B(n5933), .Z(n5931) );
  XOR U9009 ( .A(DB[1662]), .B(DB[1655]), .Z(n5933) );
  AND U9010 ( .A(n1102), .B(n5934), .Z(n5932) );
  XOR U9011 ( .A(n5935), .B(n5936), .Z(n5934) );
  XOR U9012 ( .A(DB[1655]), .B(DB[1648]), .Z(n5936) );
  AND U9013 ( .A(n1106), .B(n5937), .Z(n5935) );
  XOR U9014 ( .A(n5938), .B(n5939), .Z(n5937) );
  XOR U9015 ( .A(DB[1648]), .B(DB[1641]), .Z(n5939) );
  AND U9016 ( .A(n1110), .B(n5940), .Z(n5938) );
  XOR U9017 ( .A(n5941), .B(n5942), .Z(n5940) );
  XOR U9018 ( .A(DB[1641]), .B(DB[1634]), .Z(n5942) );
  AND U9019 ( .A(n1114), .B(n5943), .Z(n5941) );
  XOR U9020 ( .A(n5944), .B(n5945), .Z(n5943) );
  XOR U9021 ( .A(DB[1634]), .B(DB[1627]), .Z(n5945) );
  AND U9022 ( .A(n1118), .B(n5946), .Z(n5944) );
  XOR U9023 ( .A(n5947), .B(n5948), .Z(n5946) );
  XOR U9024 ( .A(DB[1627]), .B(DB[1620]), .Z(n5948) );
  AND U9025 ( .A(n1122), .B(n5949), .Z(n5947) );
  XOR U9026 ( .A(n5950), .B(n5951), .Z(n5949) );
  XOR U9027 ( .A(DB[1620]), .B(DB[1613]), .Z(n5951) );
  AND U9028 ( .A(n1126), .B(n5952), .Z(n5950) );
  XOR U9029 ( .A(n5953), .B(n5954), .Z(n5952) );
  XOR U9030 ( .A(DB[1613]), .B(DB[1606]), .Z(n5954) );
  AND U9031 ( .A(n1130), .B(n5955), .Z(n5953) );
  XOR U9032 ( .A(n5956), .B(n5957), .Z(n5955) );
  XOR U9033 ( .A(DB[1606]), .B(DB[1599]), .Z(n5957) );
  AND U9034 ( .A(n1134), .B(n5958), .Z(n5956) );
  XOR U9035 ( .A(n5959), .B(n5960), .Z(n5958) );
  XOR U9036 ( .A(DB[1599]), .B(DB[1592]), .Z(n5960) );
  AND U9037 ( .A(n1138), .B(n5961), .Z(n5959) );
  XOR U9038 ( .A(n5962), .B(n5963), .Z(n5961) );
  XOR U9039 ( .A(DB[1592]), .B(DB[1585]), .Z(n5963) );
  AND U9040 ( .A(n1142), .B(n5964), .Z(n5962) );
  XOR U9041 ( .A(n5965), .B(n5966), .Z(n5964) );
  XOR U9042 ( .A(DB[1585]), .B(DB[1578]), .Z(n5966) );
  AND U9043 ( .A(n1146), .B(n5967), .Z(n5965) );
  XOR U9044 ( .A(n5968), .B(n5969), .Z(n5967) );
  XOR U9045 ( .A(DB[1578]), .B(DB[1571]), .Z(n5969) );
  AND U9046 ( .A(n1150), .B(n5970), .Z(n5968) );
  XOR U9047 ( .A(n5971), .B(n5972), .Z(n5970) );
  XOR U9048 ( .A(DB[1571]), .B(DB[1564]), .Z(n5972) );
  AND U9049 ( .A(n1154), .B(n5973), .Z(n5971) );
  XOR U9050 ( .A(n5974), .B(n5975), .Z(n5973) );
  XOR U9051 ( .A(DB[1564]), .B(DB[1557]), .Z(n5975) );
  AND U9052 ( .A(n1158), .B(n5976), .Z(n5974) );
  XOR U9053 ( .A(n5977), .B(n5978), .Z(n5976) );
  XOR U9054 ( .A(DB[1557]), .B(DB[1550]), .Z(n5978) );
  AND U9055 ( .A(n1162), .B(n5979), .Z(n5977) );
  XOR U9056 ( .A(n5980), .B(n5981), .Z(n5979) );
  XOR U9057 ( .A(DB[1550]), .B(DB[1543]), .Z(n5981) );
  AND U9058 ( .A(n1166), .B(n5982), .Z(n5980) );
  XOR U9059 ( .A(n5983), .B(n5984), .Z(n5982) );
  XOR U9060 ( .A(DB[1543]), .B(DB[1536]), .Z(n5984) );
  AND U9061 ( .A(n1170), .B(n5985), .Z(n5983) );
  XOR U9062 ( .A(n5986), .B(n5987), .Z(n5985) );
  XOR U9063 ( .A(DB[1536]), .B(DB[1529]), .Z(n5987) );
  AND U9064 ( .A(n1174), .B(n5988), .Z(n5986) );
  XOR U9065 ( .A(n5989), .B(n5990), .Z(n5988) );
  XOR U9066 ( .A(DB[1529]), .B(DB[1522]), .Z(n5990) );
  AND U9067 ( .A(n1178), .B(n5991), .Z(n5989) );
  XOR U9068 ( .A(n5992), .B(n5993), .Z(n5991) );
  XOR U9069 ( .A(DB[1522]), .B(DB[1515]), .Z(n5993) );
  AND U9070 ( .A(n1182), .B(n5994), .Z(n5992) );
  XOR U9071 ( .A(n5995), .B(n5996), .Z(n5994) );
  XOR U9072 ( .A(DB[1515]), .B(DB[1508]), .Z(n5996) );
  AND U9073 ( .A(n1186), .B(n5997), .Z(n5995) );
  XOR U9074 ( .A(n5998), .B(n5999), .Z(n5997) );
  XOR U9075 ( .A(DB[1508]), .B(DB[1501]), .Z(n5999) );
  AND U9076 ( .A(n1190), .B(n6000), .Z(n5998) );
  XOR U9077 ( .A(n6001), .B(n6002), .Z(n6000) );
  XOR U9078 ( .A(DB[1501]), .B(DB[1494]), .Z(n6002) );
  AND U9079 ( .A(n1194), .B(n6003), .Z(n6001) );
  XOR U9080 ( .A(n6004), .B(n6005), .Z(n6003) );
  XOR U9081 ( .A(DB[1494]), .B(DB[1487]), .Z(n6005) );
  AND U9082 ( .A(n1198), .B(n6006), .Z(n6004) );
  XOR U9083 ( .A(n6007), .B(n6008), .Z(n6006) );
  XOR U9084 ( .A(DB[1487]), .B(DB[1480]), .Z(n6008) );
  AND U9085 ( .A(n1202), .B(n6009), .Z(n6007) );
  XOR U9086 ( .A(n6010), .B(n6011), .Z(n6009) );
  XOR U9087 ( .A(DB[1480]), .B(DB[1473]), .Z(n6011) );
  AND U9088 ( .A(n1206), .B(n6012), .Z(n6010) );
  XOR U9089 ( .A(n6013), .B(n6014), .Z(n6012) );
  XOR U9090 ( .A(DB[1473]), .B(DB[1466]), .Z(n6014) );
  AND U9091 ( .A(n1210), .B(n6015), .Z(n6013) );
  XOR U9092 ( .A(n6016), .B(n6017), .Z(n6015) );
  XOR U9093 ( .A(DB[1466]), .B(DB[1459]), .Z(n6017) );
  AND U9094 ( .A(n1214), .B(n6018), .Z(n6016) );
  XOR U9095 ( .A(n6019), .B(n6020), .Z(n6018) );
  XOR U9096 ( .A(DB[1459]), .B(DB[1452]), .Z(n6020) );
  AND U9097 ( .A(n1218), .B(n6021), .Z(n6019) );
  XOR U9098 ( .A(n6022), .B(n6023), .Z(n6021) );
  XOR U9099 ( .A(DB[1452]), .B(DB[1445]), .Z(n6023) );
  AND U9100 ( .A(n1222), .B(n6024), .Z(n6022) );
  XOR U9101 ( .A(n6025), .B(n6026), .Z(n6024) );
  XOR U9102 ( .A(DB[1445]), .B(DB[1438]), .Z(n6026) );
  AND U9103 ( .A(n1226), .B(n6027), .Z(n6025) );
  XOR U9104 ( .A(n6028), .B(n6029), .Z(n6027) );
  XOR U9105 ( .A(DB[1438]), .B(DB[1431]), .Z(n6029) );
  AND U9106 ( .A(n1230), .B(n6030), .Z(n6028) );
  XOR U9107 ( .A(n6031), .B(n6032), .Z(n6030) );
  XOR U9108 ( .A(DB[1431]), .B(DB[1424]), .Z(n6032) );
  AND U9109 ( .A(n1234), .B(n6033), .Z(n6031) );
  XOR U9110 ( .A(n6034), .B(n6035), .Z(n6033) );
  XOR U9111 ( .A(DB[1424]), .B(DB[1417]), .Z(n6035) );
  AND U9112 ( .A(n1238), .B(n6036), .Z(n6034) );
  XOR U9113 ( .A(n6037), .B(n6038), .Z(n6036) );
  XOR U9114 ( .A(DB[1417]), .B(DB[1410]), .Z(n6038) );
  AND U9115 ( .A(n1242), .B(n6039), .Z(n6037) );
  XOR U9116 ( .A(n6040), .B(n6041), .Z(n6039) );
  XOR U9117 ( .A(DB[1410]), .B(DB[1403]), .Z(n6041) );
  AND U9118 ( .A(n1246), .B(n6042), .Z(n6040) );
  XOR U9119 ( .A(n6043), .B(n6044), .Z(n6042) );
  XOR U9120 ( .A(DB[1403]), .B(DB[1396]), .Z(n6044) );
  AND U9121 ( .A(n1250), .B(n6045), .Z(n6043) );
  XOR U9122 ( .A(n6046), .B(n6047), .Z(n6045) );
  XOR U9123 ( .A(DB[1396]), .B(DB[1389]), .Z(n6047) );
  AND U9124 ( .A(n1254), .B(n6048), .Z(n6046) );
  XOR U9125 ( .A(n6049), .B(n6050), .Z(n6048) );
  XOR U9126 ( .A(DB[1389]), .B(DB[1382]), .Z(n6050) );
  AND U9127 ( .A(n1258), .B(n6051), .Z(n6049) );
  XOR U9128 ( .A(n6052), .B(n6053), .Z(n6051) );
  XOR U9129 ( .A(DB[1382]), .B(DB[1375]), .Z(n6053) );
  AND U9130 ( .A(n1262), .B(n6054), .Z(n6052) );
  XOR U9131 ( .A(n6055), .B(n6056), .Z(n6054) );
  XOR U9132 ( .A(DB[1375]), .B(DB[1368]), .Z(n6056) );
  AND U9133 ( .A(n1266), .B(n6057), .Z(n6055) );
  XOR U9134 ( .A(n6058), .B(n6059), .Z(n6057) );
  XOR U9135 ( .A(DB[1368]), .B(DB[1361]), .Z(n6059) );
  AND U9136 ( .A(n1270), .B(n6060), .Z(n6058) );
  XOR U9137 ( .A(n6061), .B(n6062), .Z(n6060) );
  XOR U9138 ( .A(DB[1361]), .B(DB[1354]), .Z(n6062) );
  AND U9139 ( .A(n1274), .B(n6063), .Z(n6061) );
  XOR U9140 ( .A(n6064), .B(n6065), .Z(n6063) );
  XOR U9141 ( .A(DB[1354]), .B(DB[1347]), .Z(n6065) );
  AND U9142 ( .A(n1278), .B(n6066), .Z(n6064) );
  XOR U9143 ( .A(n6067), .B(n6068), .Z(n6066) );
  XOR U9144 ( .A(DB[1347]), .B(DB[1340]), .Z(n6068) );
  AND U9145 ( .A(n1282), .B(n6069), .Z(n6067) );
  XOR U9146 ( .A(n6070), .B(n6071), .Z(n6069) );
  XOR U9147 ( .A(DB[1340]), .B(DB[1333]), .Z(n6071) );
  AND U9148 ( .A(n1286), .B(n6072), .Z(n6070) );
  XOR U9149 ( .A(n6073), .B(n6074), .Z(n6072) );
  XOR U9150 ( .A(DB[1333]), .B(DB[1326]), .Z(n6074) );
  AND U9151 ( .A(n1290), .B(n6075), .Z(n6073) );
  XOR U9152 ( .A(n6076), .B(n6077), .Z(n6075) );
  XOR U9153 ( .A(DB[1326]), .B(DB[1319]), .Z(n6077) );
  AND U9154 ( .A(n1294), .B(n6078), .Z(n6076) );
  XOR U9155 ( .A(n6079), .B(n6080), .Z(n6078) );
  XOR U9156 ( .A(DB[1319]), .B(DB[1312]), .Z(n6080) );
  AND U9157 ( .A(n1298), .B(n6081), .Z(n6079) );
  XOR U9158 ( .A(n6082), .B(n6083), .Z(n6081) );
  XOR U9159 ( .A(DB[1312]), .B(DB[1305]), .Z(n6083) );
  AND U9160 ( .A(n1302), .B(n6084), .Z(n6082) );
  XOR U9161 ( .A(n6085), .B(n6086), .Z(n6084) );
  XOR U9162 ( .A(DB[1305]), .B(DB[1298]), .Z(n6086) );
  AND U9163 ( .A(n1306), .B(n6087), .Z(n6085) );
  XOR U9164 ( .A(n6088), .B(n6089), .Z(n6087) );
  XOR U9165 ( .A(DB[1298]), .B(DB[1291]), .Z(n6089) );
  AND U9166 ( .A(n1310), .B(n6090), .Z(n6088) );
  XOR U9167 ( .A(n6091), .B(n6092), .Z(n6090) );
  XOR U9168 ( .A(DB[1291]), .B(DB[1284]), .Z(n6092) );
  AND U9169 ( .A(n1314), .B(n6093), .Z(n6091) );
  XOR U9170 ( .A(n6094), .B(n6095), .Z(n6093) );
  XOR U9171 ( .A(DB[1284]), .B(DB[1277]), .Z(n6095) );
  AND U9172 ( .A(n1318), .B(n6096), .Z(n6094) );
  XOR U9173 ( .A(n6097), .B(n6098), .Z(n6096) );
  XOR U9174 ( .A(DB[1277]), .B(DB[1270]), .Z(n6098) );
  AND U9175 ( .A(n1322), .B(n6099), .Z(n6097) );
  XOR U9176 ( .A(n6100), .B(n6101), .Z(n6099) );
  XOR U9177 ( .A(DB[1270]), .B(DB[1263]), .Z(n6101) );
  AND U9178 ( .A(n1326), .B(n6102), .Z(n6100) );
  XOR U9179 ( .A(n6103), .B(n6104), .Z(n6102) );
  XOR U9180 ( .A(DB[1263]), .B(DB[1256]), .Z(n6104) );
  AND U9181 ( .A(n1330), .B(n6105), .Z(n6103) );
  XOR U9182 ( .A(n6106), .B(n6107), .Z(n6105) );
  XOR U9183 ( .A(DB[1256]), .B(DB[1249]), .Z(n6107) );
  AND U9184 ( .A(n1334), .B(n6108), .Z(n6106) );
  XOR U9185 ( .A(n6109), .B(n6110), .Z(n6108) );
  XOR U9186 ( .A(DB[1249]), .B(DB[1242]), .Z(n6110) );
  AND U9187 ( .A(n1338), .B(n6111), .Z(n6109) );
  XOR U9188 ( .A(n6112), .B(n6113), .Z(n6111) );
  XOR U9189 ( .A(DB[1242]), .B(DB[1235]), .Z(n6113) );
  AND U9190 ( .A(n1342), .B(n6114), .Z(n6112) );
  XOR U9191 ( .A(n6115), .B(n6116), .Z(n6114) );
  XOR U9192 ( .A(DB[1235]), .B(DB[1228]), .Z(n6116) );
  AND U9193 ( .A(n1346), .B(n6117), .Z(n6115) );
  XOR U9194 ( .A(n6118), .B(n6119), .Z(n6117) );
  XOR U9195 ( .A(DB[1228]), .B(DB[1221]), .Z(n6119) );
  AND U9196 ( .A(n1350), .B(n6120), .Z(n6118) );
  XOR U9197 ( .A(n6121), .B(n6122), .Z(n6120) );
  XOR U9198 ( .A(DB[1221]), .B(DB[1214]), .Z(n6122) );
  AND U9199 ( .A(n1354), .B(n6123), .Z(n6121) );
  XOR U9200 ( .A(n6124), .B(n6125), .Z(n6123) );
  XOR U9201 ( .A(DB[1214]), .B(DB[1207]), .Z(n6125) );
  AND U9202 ( .A(n1358), .B(n6126), .Z(n6124) );
  XOR U9203 ( .A(n6127), .B(n6128), .Z(n6126) );
  XOR U9204 ( .A(DB[1207]), .B(DB[1200]), .Z(n6128) );
  AND U9205 ( .A(n1362), .B(n6129), .Z(n6127) );
  XOR U9206 ( .A(n6130), .B(n6131), .Z(n6129) );
  XOR U9207 ( .A(DB[1200]), .B(DB[1193]), .Z(n6131) );
  AND U9208 ( .A(n1366), .B(n6132), .Z(n6130) );
  XOR U9209 ( .A(n6133), .B(n6134), .Z(n6132) );
  XOR U9210 ( .A(DB[1193]), .B(DB[1186]), .Z(n6134) );
  AND U9211 ( .A(n1370), .B(n6135), .Z(n6133) );
  XOR U9212 ( .A(n6136), .B(n6137), .Z(n6135) );
  XOR U9213 ( .A(DB[1186]), .B(DB[1179]), .Z(n6137) );
  AND U9214 ( .A(n1374), .B(n6138), .Z(n6136) );
  XOR U9215 ( .A(n6139), .B(n6140), .Z(n6138) );
  XOR U9216 ( .A(DB[1179]), .B(DB[1172]), .Z(n6140) );
  AND U9217 ( .A(n1378), .B(n6141), .Z(n6139) );
  XOR U9218 ( .A(n6142), .B(n6143), .Z(n6141) );
  XOR U9219 ( .A(DB[1172]), .B(DB[1165]), .Z(n6143) );
  AND U9220 ( .A(n1382), .B(n6144), .Z(n6142) );
  XOR U9221 ( .A(n6145), .B(n6146), .Z(n6144) );
  XOR U9222 ( .A(DB[1165]), .B(DB[1158]), .Z(n6146) );
  AND U9223 ( .A(n1386), .B(n6147), .Z(n6145) );
  XOR U9224 ( .A(n6148), .B(n6149), .Z(n6147) );
  XOR U9225 ( .A(DB[1158]), .B(DB[1151]), .Z(n6149) );
  AND U9226 ( .A(n1390), .B(n6150), .Z(n6148) );
  XOR U9227 ( .A(n6151), .B(n6152), .Z(n6150) );
  XOR U9228 ( .A(DB[1151]), .B(DB[1144]), .Z(n6152) );
  AND U9229 ( .A(n1394), .B(n6153), .Z(n6151) );
  XOR U9230 ( .A(n6154), .B(n6155), .Z(n6153) );
  XOR U9231 ( .A(DB[1144]), .B(DB[1137]), .Z(n6155) );
  AND U9232 ( .A(n1398), .B(n6156), .Z(n6154) );
  XOR U9233 ( .A(n6157), .B(n6158), .Z(n6156) );
  XOR U9234 ( .A(DB[1137]), .B(DB[1130]), .Z(n6158) );
  AND U9235 ( .A(n1402), .B(n6159), .Z(n6157) );
  XOR U9236 ( .A(n6160), .B(n6161), .Z(n6159) );
  XOR U9237 ( .A(DB[1130]), .B(DB[1123]), .Z(n6161) );
  AND U9238 ( .A(n1406), .B(n6162), .Z(n6160) );
  XOR U9239 ( .A(n6163), .B(n6164), .Z(n6162) );
  XOR U9240 ( .A(DB[1123]), .B(DB[1116]), .Z(n6164) );
  AND U9241 ( .A(n1410), .B(n6165), .Z(n6163) );
  XOR U9242 ( .A(n6166), .B(n6167), .Z(n6165) );
  XOR U9243 ( .A(DB[1116]), .B(DB[1109]), .Z(n6167) );
  AND U9244 ( .A(n1414), .B(n6168), .Z(n6166) );
  XOR U9245 ( .A(n6169), .B(n6170), .Z(n6168) );
  XOR U9246 ( .A(DB[1109]), .B(DB[1102]), .Z(n6170) );
  AND U9247 ( .A(n1418), .B(n6171), .Z(n6169) );
  XOR U9248 ( .A(n6172), .B(n6173), .Z(n6171) );
  XOR U9249 ( .A(DB[1102]), .B(DB[1095]), .Z(n6173) );
  AND U9250 ( .A(n1422), .B(n6174), .Z(n6172) );
  XOR U9251 ( .A(n6175), .B(n6176), .Z(n6174) );
  XOR U9252 ( .A(DB[1095]), .B(DB[1088]), .Z(n6176) );
  AND U9253 ( .A(n1426), .B(n6177), .Z(n6175) );
  XOR U9254 ( .A(n6178), .B(n6179), .Z(n6177) );
  XOR U9255 ( .A(DB[1088]), .B(DB[1081]), .Z(n6179) );
  AND U9256 ( .A(n1430), .B(n6180), .Z(n6178) );
  XOR U9257 ( .A(n6181), .B(n6182), .Z(n6180) );
  XOR U9258 ( .A(DB[1081]), .B(DB[1074]), .Z(n6182) );
  AND U9259 ( .A(n1434), .B(n6183), .Z(n6181) );
  XOR U9260 ( .A(n6184), .B(n6185), .Z(n6183) );
  XOR U9261 ( .A(DB[1074]), .B(DB[1067]), .Z(n6185) );
  AND U9262 ( .A(n1438), .B(n6186), .Z(n6184) );
  XOR U9263 ( .A(n6187), .B(n6188), .Z(n6186) );
  XOR U9264 ( .A(DB[1067]), .B(DB[1060]), .Z(n6188) );
  AND U9265 ( .A(n1442), .B(n6189), .Z(n6187) );
  XOR U9266 ( .A(n6190), .B(n6191), .Z(n6189) );
  XOR U9267 ( .A(DB[1060]), .B(DB[1053]), .Z(n6191) );
  AND U9268 ( .A(n1446), .B(n6192), .Z(n6190) );
  XOR U9269 ( .A(n6193), .B(n6194), .Z(n6192) );
  XOR U9270 ( .A(DB[1053]), .B(DB[1046]), .Z(n6194) );
  AND U9271 ( .A(n1450), .B(n6195), .Z(n6193) );
  XOR U9272 ( .A(n6196), .B(n6197), .Z(n6195) );
  XOR U9273 ( .A(DB[1046]), .B(DB[1039]), .Z(n6197) );
  AND U9274 ( .A(n1454), .B(n6198), .Z(n6196) );
  XOR U9275 ( .A(n6199), .B(n6200), .Z(n6198) );
  XOR U9276 ( .A(DB[1039]), .B(DB[1032]), .Z(n6200) );
  AND U9277 ( .A(n1458), .B(n6201), .Z(n6199) );
  XOR U9278 ( .A(n6202), .B(n6203), .Z(n6201) );
  XOR U9279 ( .A(DB[1032]), .B(DB[1025]), .Z(n6203) );
  AND U9280 ( .A(n1462), .B(n6204), .Z(n6202) );
  XOR U9281 ( .A(n6205), .B(n6206), .Z(n6204) );
  XOR U9282 ( .A(DB[1025]), .B(DB[1018]), .Z(n6206) );
  AND U9283 ( .A(n1466), .B(n6207), .Z(n6205) );
  XOR U9284 ( .A(n6208), .B(n6209), .Z(n6207) );
  XOR U9285 ( .A(DB[1018]), .B(DB[1011]), .Z(n6209) );
  AND U9286 ( .A(n1470), .B(n6210), .Z(n6208) );
  XOR U9287 ( .A(n6211), .B(n6212), .Z(n6210) );
  XOR U9288 ( .A(DB[1011]), .B(DB[1004]), .Z(n6212) );
  AND U9289 ( .A(n1474), .B(n6213), .Z(n6211) );
  XOR U9290 ( .A(n6214), .B(n6215), .Z(n6213) );
  XOR U9291 ( .A(DB[997]), .B(DB[1004]), .Z(n6215) );
  AND U9292 ( .A(n1478), .B(n6216), .Z(n6214) );
  XOR U9293 ( .A(n6217), .B(n6218), .Z(n6216) );
  XOR U9294 ( .A(DB[997]), .B(DB[990]), .Z(n6218) );
  AND U9295 ( .A(n1482), .B(n6219), .Z(n6217) );
  XOR U9296 ( .A(n6220), .B(n6221), .Z(n6219) );
  XOR U9297 ( .A(DB[990]), .B(DB[983]), .Z(n6221) );
  AND U9298 ( .A(n1486), .B(n6222), .Z(n6220) );
  XOR U9299 ( .A(n6223), .B(n6224), .Z(n6222) );
  XOR U9300 ( .A(DB[983]), .B(DB[976]), .Z(n6224) );
  AND U9301 ( .A(n1490), .B(n6225), .Z(n6223) );
  XOR U9302 ( .A(n6226), .B(n6227), .Z(n6225) );
  XOR U9303 ( .A(DB[976]), .B(DB[969]), .Z(n6227) );
  AND U9304 ( .A(n1494), .B(n6228), .Z(n6226) );
  XOR U9305 ( .A(n6229), .B(n6230), .Z(n6228) );
  XOR U9306 ( .A(DB[969]), .B(DB[962]), .Z(n6230) );
  AND U9307 ( .A(n1498), .B(n6231), .Z(n6229) );
  XOR U9308 ( .A(n6232), .B(n6233), .Z(n6231) );
  XOR U9309 ( .A(DB[962]), .B(DB[955]), .Z(n6233) );
  AND U9310 ( .A(n1502), .B(n6234), .Z(n6232) );
  XOR U9311 ( .A(n6235), .B(n6236), .Z(n6234) );
  XOR U9312 ( .A(DB[955]), .B(DB[948]), .Z(n6236) );
  AND U9313 ( .A(n1506), .B(n6237), .Z(n6235) );
  XOR U9314 ( .A(n6238), .B(n6239), .Z(n6237) );
  XOR U9315 ( .A(DB[948]), .B(DB[941]), .Z(n6239) );
  AND U9316 ( .A(n1510), .B(n6240), .Z(n6238) );
  XOR U9317 ( .A(n6241), .B(n6242), .Z(n6240) );
  XOR U9318 ( .A(DB[941]), .B(DB[934]), .Z(n6242) );
  AND U9319 ( .A(n1514), .B(n6243), .Z(n6241) );
  XOR U9320 ( .A(n6244), .B(n6245), .Z(n6243) );
  XOR U9321 ( .A(DB[934]), .B(DB[927]), .Z(n6245) );
  AND U9322 ( .A(n1518), .B(n6246), .Z(n6244) );
  XOR U9323 ( .A(n6247), .B(n6248), .Z(n6246) );
  XOR U9324 ( .A(DB[927]), .B(DB[920]), .Z(n6248) );
  AND U9325 ( .A(n1522), .B(n6249), .Z(n6247) );
  XOR U9326 ( .A(n6250), .B(n6251), .Z(n6249) );
  XOR U9327 ( .A(DB[920]), .B(DB[913]), .Z(n6251) );
  AND U9328 ( .A(n1526), .B(n6252), .Z(n6250) );
  XOR U9329 ( .A(n6253), .B(n6254), .Z(n6252) );
  XOR U9330 ( .A(DB[913]), .B(DB[906]), .Z(n6254) );
  AND U9331 ( .A(n1530), .B(n6255), .Z(n6253) );
  XOR U9332 ( .A(n6256), .B(n6257), .Z(n6255) );
  XOR U9333 ( .A(DB[906]), .B(DB[899]), .Z(n6257) );
  AND U9334 ( .A(n1534), .B(n6258), .Z(n6256) );
  XOR U9335 ( .A(n6259), .B(n6260), .Z(n6258) );
  XOR U9336 ( .A(DB[899]), .B(DB[892]), .Z(n6260) );
  AND U9337 ( .A(n1538), .B(n6261), .Z(n6259) );
  XOR U9338 ( .A(n6262), .B(n6263), .Z(n6261) );
  XOR U9339 ( .A(DB[892]), .B(DB[885]), .Z(n6263) );
  AND U9340 ( .A(n1542), .B(n6264), .Z(n6262) );
  XOR U9341 ( .A(n6265), .B(n6266), .Z(n6264) );
  XOR U9342 ( .A(DB[885]), .B(DB[878]), .Z(n6266) );
  AND U9343 ( .A(n1546), .B(n6267), .Z(n6265) );
  XOR U9344 ( .A(n6268), .B(n6269), .Z(n6267) );
  XOR U9345 ( .A(DB[878]), .B(DB[871]), .Z(n6269) );
  AND U9346 ( .A(n1550), .B(n6270), .Z(n6268) );
  XOR U9347 ( .A(n6271), .B(n6272), .Z(n6270) );
  XOR U9348 ( .A(DB[871]), .B(DB[864]), .Z(n6272) );
  AND U9349 ( .A(n1554), .B(n6273), .Z(n6271) );
  XOR U9350 ( .A(n6274), .B(n6275), .Z(n6273) );
  XOR U9351 ( .A(DB[864]), .B(DB[857]), .Z(n6275) );
  AND U9352 ( .A(n1558), .B(n6276), .Z(n6274) );
  XOR U9353 ( .A(n6277), .B(n6278), .Z(n6276) );
  XOR U9354 ( .A(DB[857]), .B(DB[850]), .Z(n6278) );
  AND U9355 ( .A(n1562), .B(n6279), .Z(n6277) );
  XOR U9356 ( .A(n6280), .B(n6281), .Z(n6279) );
  XOR U9357 ( .A(DB[850]), .B(DB[843]), .Z(n6281) );
  AND U9358 ( .A(n1566), .B(n6282), .Z(n6280) );
  XOR U9359 ( .A(n6283), .B(n6284), .Z(n6282) );
  XOR U9360 ( .A(DB[843]), .B(DB[836]), .Z(n6284) );
  AND U9361 ( .A(n1570), .B(n6285), .Z(n6283) );
  XOR U9362 ( .A(n6286), .B(n6287), .Z(n6285) );
  XOR U9363 ( .A(DB[836]), .B(DB[829]), .Z(n6287) );
  AND U9364 ( .A(n1574), .B(n6288), .Z(n6286) );
  XOR U9365 ( .A(n6289), .B(n6290), .Z(n6288) );
  XOR U9366 ( .A(DB[829]), .B(DB[822]), .Z(n6290) );
  AND U9367 ( .A(n1578), .B(n6291), .Z(n6289) );
  XOR U9368 ( .A(n6292), .B(n6293), .Z(n6291) );
  XOR U9369 ( .A(DB[822]), .B(DB[815]), .Z(n6293) );
  AND U9370 ( .A(n1582), .B(n6294), .Z(n6292) );
  XOR U9371 ( .A(n6295), .B(n6296), .Z(n6294) );
  XOR U9372 ( .A(DB[815]), .B(DB[808]), .Z(n6296) );
  AND U9373 ( .A(n1586), .B(n6297), .Z(n6295) );
  XOR U9374 ( .A(n6298), .B(n6299), .Z(n6297) );
  XOR U9375 ( .A(DB[808]), .B(DB[801]), .Z(n6299) );
  AND U9376 ( .A(n1590), .B(n6300), .Z(n6298) );
  XOR U9377 ( .A(n6301), .B(n6302), .Z(n6300) );
  XOR U9378 ( .A(DB[801]), .B(DB[794]), .Z(n6302) );
  AND U9379 ( .A(n1594), .B(n6303), .Z(n6301) );
  XOR U9380 ( .A(n6304), .B(n6305), .Z(n6303) );
  XOR U9381 ( .A(DB[794]), .B(DB[787]), .Z(n6305) );
  AND U9382 ( .A(n1598), .B(n6306), .Z(n6304) );
  XOR U9383 ( .A(n6307), .B(n6308), .Z(n6306) );
  XOR U9384 ( .A(DB[787]), .B(DB[780]), .Z(n6308) );
  AND U9385 ( .A(n1602), .B(n6309), .Z(n6307) );
  XOR U9386 ( .A(n6310), .B(n6311), .Z(n6309) );
  XOR U9387 ( .A(DB[780]), .B(DB[773]), .Z(n6311) );
  AND U9388 ( .A(n1606), .B(n6312), .Z(n6310) );
  XOR U9389 ( .A(n6313), .B(n6314), .Z(n6312) );
  XOR U9390 ( .A(DB[773]), .B(DB[766]), .Z(n6314) );
  AND U9391 ( .A(n1610), .B(n6315), .Z(n6313) );
  XOR U9392 ( .A(n6316), .B(n6317), .Z(n6315) );
  XOR U9393 ( .A(DB[766]), .B(DB[759]), .Z(n6317) );
  AND U9394 ( .A(n1614), .B(n6318), .Z(n6316) );
  XOR U9395 ( .A(n6319), .B(n6320), .Z(n6318) );
  XOR U9396 ( .A(DB[759]), .B(DB[752]), .Z(n6320) );
  AND U9397 ( .A(n1618), .B(n6321), .Z(n6319) );
  XOR U9398 ( .A(n6322), .B(n6323), .Z(n6321) );
  XOR U9399 ( .A(DB[752]), .B(DB[745]), .Z(n6323) );
  AND U9400 ( .A(n1622), .B(n6324), .Z(n6322) );
  XOR U9401 ( .A(n6325), .B(n6326), .Z(n6324) );
  XOR U9402 ( .A(DB[745]), .B(DB[738]), .Z(n6326) );
  AND U9403 ( .A(n1626), .B(n6327), .Z(n6325) );
  XOR U9404 ( .A(n6328), .B(n6329), .Z(n6327) );
  XOR U9405 ( .A(DB[738]), .B(DB[731]), .Z(n6329) );
  AND U9406 ( .A(n1630), .B(n6330), .Z(n6328) );
  XOR U9407 ( .A(n6331), .B(n6332), .Z(n6330) );
  XOR U9408 ( .A(DB[731]), .B(DB[724]), .Z(n6332) );
  AND U9409 ( .A(n1634), .B(n6333), .Z(n6331) );
  XOR U9410 ( .A(n6334), .B(n6335), .Z(n6333) );
  XOR U9411 ( .A(DB[724]), .B(DB[717]), .Z(n6335) );
  AND U9412 ( .A(n1638), .B(n6336), .Z(n6334) );
  XOR U9413 ( .A(n6337), .B(n6338), .Z(n6336) );
  XOR U9414 ( .A(DB[717]), .B(DB[710]), .Z(n6338) );
  AND U9415 ( .A(n1642), .B(n6339), .Z(n6337) );
  XOR U9416 ( .A(n6340), .B(n6341), .Z(n6339) );
  XOR U9417 ( .A(DB[710]), .B(DB[703]), .Z(n6341) );
  AND U9418 ( .A(n1646), .B(n6342), .Z(n6340) );
  XOR U9419 ( .A(n6343), .B(n6344), .Z(n6342) );
  XOR U9420 ( .A(DB[703]), .B(DB[696]), .Z(n6344) );
  AND U9421 ( .A(n1650), .B(n6345), .Z(n6343) );
  XOR U9422 ( .A(n6346), .B(n6347), .Z(n6345) );
  XOR U9423 ( .A(DB[696]), .B(DB[689]), .Z(n6347) );
  AND U9424 ( .A(n1654), .B(n6348), .Z(n6346) );
  XOR U9425 ( .A(n6349), .B(n6350), .Z(n6348) );
  XOR U9426 ( .A(DB[689]), .B(DB[682]), .Z(n6350) );
  AND U9427 ( .A(n1658), .B(n6351), .Z(n6349) );
  XOR U9428 ( .A(n6352), .B(n6353), .Z(n6351) );
  XOR U9429 ( .A(DB[682]), .B(DB[675]), .Z(n6353) );
  AND U9430 ( .A(n1662), .B(n6354), .Z(n6352) );
  XOR U9431 ( .A(n6355), .B(n6356), .Z(n6354) );
  XOR U9432 ( .A(DB[675]), .B(DB[668]), .Z(n6356) );
  AND U9433 ( .A(n1666), .B(n6357), .Z(n6355) );
  XOR U9434 ( .A(n6358), .B(n6359), .Z(n6357) );
  XOR U9435 ( .A(DB[668]), .B(DB[661]), .Z(n6359) );
  AND U9436 ( .A(n1670), .B(n6360), .Z(n6358) );
  XOR U9437 ( .A(n6361), .B(n6362), .Z(n6360) );
  XOR U9438 ( .A(DB[661]), .B(DB[654]), .Z(n6362) );
  AND U9439 ( .A(n1674), .B(n6363), .Z(n6361) );
  XOR U9440 ( .A(n6364), .B(n6365), .Z(n6363) );
  XOR U9441 ( .A(DB[654]), .B(DB[647]), .Z(n6365) );
  AND U9442 ( .A(n1678), .B(n6366), .Z(n6364) );
  XOR U9443 ( .A(n6367), .B(n6368), .Z(n6366) );
  XOR U9444 ( .A(DB[647]), .B(DB[640]), .Z(n6368) );
  AND U9445 ( .A(n1682), .B(n6369), .Z(n6367) );
  XOR U9446 ( .A(n6370), .B(n6371), .Z(n6369) );
  XOR U9447 ( .A(DB[640]), .B(DB[633]), .Z(n6371) );
  AND U9448 ( .A(n1686), .B(n6372), .Z(n6370) );
  XOR U9449 ( .A(n6373), .B(n6374), .Z(n6372) );
  XOR U9450 ( .A(DB[633]), .B(DB[626]), .Z(n6374) );
  AND U9451 ( .A(n1690), .B(n6375), .Z(n6373) );
  XOR U9452 ( .A(n6376), .B(n6377), .Z(n6375) );
  XOR U9453 ( .A(DB[626]), .B(DB[619]), .Z(n6377) );
  AND U9454 ( .A(n1694), .B(n6378), .Z(n6376) );
  XOR U9455 ( .A(n6379), .B(n6380), .Z(n6378) );
  XOR U9456 ( .A(DB[619]), .B(DB[612]), .Z(n6380) );
  AND U9457 ( .A(n1698), .B(n6381), .Z(n6379) );
  XOR U9458 ( .A(n6382), .B(n6383), .Z(n6381) );
  XOR U9459 ( .A(DB[612]), .B(DB[605]), .Z(n6383) );
  AND U9460 ( .A(n1702), .B(n6384), .Z(n6382) );
  XOR U9461 ( .A(n6385), .B(n6386), .Z(n6384) );
  XOR U9462 ( .A(DB[605]), .B(DB[598]), .Z(n6386) );
  AND U9463 ( .A(n1706), .B(n6387), .Z(n6385) );
  XOR U9464 ( .A(n6388), .B(n6389), .Z(n6387) );
  XOR U9465 ( .A(DB[598]), .B(DB[591]), .Z(n6389) );
  AND U9466 ( .A(n1710), .B(n6390), .Z(n6388) );
  XOR U9467 ( .A(n6391), .B(n6392), .Z(n6390) );
  XOR U9468 ( .A(DB[591]), .B(DB[584]), .Z(n6392) );
  AND U9469 ( .A(n1714), .B(n6393), .Z(n6391) );
  XOR U9470 ( .A(n6394), .B(n6395), .Z(n6393) );
  XOR U9471 ( .A(DB[584]), .B(DB[577]), .Z(n6395) );
  AND U9472 ( .A(n1718), .B(n6396), .Z(n6394) );
  XOR U9473 ( .A(n6397), .B(n6398), .Z(n6396) );
  XOR U9474 ( .A(DB[577]), .B(DB[570]), .Z(n6398) );
  AND U9475 ( .A(n1722), .B(n6399), .Z(n6397) );
  XOR U9476 ( .A(n6400), .B(n6401), .Z(n6399) );
  XOR U9477 ( .A(DB[570]), .B(DB[563]), .Z(n6401) );
  AND U9478 ( .A(n1726), .B(n6402), .Z(n6400) );
  XOR U9479 ( .A(n6403), .B(n6404), .Z(n6402) );
  XOR U9480 ( .A(DB[563]), .B(DB[556]), .Z(n6404) );
  AND U9481 ( .A(n1730), .B(n6405), .Z(n6403) );
  XOR U9482 ( .A(n6406), .B(n6407), .Z(n6405) );
  XOR U9483 ( .A(DB[556]), .B(DB[549]), .Z(n6407) );
  AND U9484 ( .A(n1734), .B(n6408), .Z(n6406) );
  XOR U9485 ( .A(n6409), .B(n6410), .Z(n6408) );
  XOR U9486 ( .A(DB[549]), .B(DB[542]), .Z(n6410) );
  AND U9487 ( .A(n1738), .B(n6411), .Z(n6409) );
  XOR U9488 ( .A(n6412), .B(n6413), .Z(n6411) );
  XOR U9489 ( .A(DB[542]), .B(DB[535]), .Z(n6413) );
  AND U9490 ( .A(n1742), .B(n6414), .Z(n6412) );
  XOR U9491 ( .A(n6415), .B(n6416), .Z(n6414) );
  XOR U9492 ( .A(DB[535]), .B(DB[528]), .Z(n6416) );
  AND U9493 ( .A(n1746), .B(n6417), .Z(n6415) );
  XOR U9494 ( .A(n6418), .B(n6419), .Z(n6417) );
  XOR U9495 ( .A(DB[528]), .B(DB[521]), .Z(n6419) );
  AND U9496 ( .A(n1750), .B(n6420), .Z(n6418) );
  XOR U9497 ( .A(n6421), .B(n6422), .Z(n6420) );
  XOR U9498 ( .A(DB[521]), .B(DB[514]), .Z(n6422) );
  AND U9499 ( .A(n1754), .B(n6423), .Z(n6421) );
  XOR U9500 ( .A(n6424), .B(n6425), .Z(n6423) );
  XOR U9501 ( .A(DB[514]), .B(DB[507]), .Z(n6425) );
  AND U9502 ( .A(n1758), .B(n6426), .Z(n6424) );
  XOR U9503 ( .A(n6427), .B(n6428), .Z(n6426) );
  XOR U9504 ( .A(DB[507]), .B(DB[500]), .Z(n6428) );
  AND U9505 ( .A(n1762), .B(n6429), .Z(n6427) );
  XOR U9506 ( .A(n6430), .B(n6431), .Z(n6429) );
  XOR U9507 ( .A(DB[500]), .B(DB[493]), .Z(n6431) );
  AND U9508 ( .A(n1766), .B(n6432), .Z(n6430) );
  XOR U9509 ( .A(n6433), .B(n6434), .Z(n6432) );
  XOR U9510 ( .A(DB[493]), .B(DB[486]), .Z(n6434) );
  AND U9511 ( .A(n1770), .B(n6435), .Z(n6433) );
  XOR U9512 ( .A(n6436), .B(n6437), .Z(n6435) );
  XOR U9513 ( .A(DB[486]), .B(DB[479]), .Z(n6437) );
  AND U9514 ( .A(n1774), .B(n6438), .Z(n6436) );
  XOR U9515 ( .A(n6439), .B(n6440), .Z(n6438) );
  XOR U9516 ( .A(DB[479]), .B(DB[472]), .Z(n6440) );
  AND U9517 ( .A(n1778), .B(n6441), .Z(n6439) );
  XOR U9518 ( .A(n6442), .B(n6443), .Z(n6441) );
  XOR U9519 ( .A(DB[472]), .B(DB[465]), .Z(n6443) );
  AND U9520 ( .A(n1782), .B(n6444), .Z(n6442) );
  XOR U9521 ( .A(n6445), .B(n6446), .Z(n6444) );
  XOR U9522 ( .A(DB[465]), .B(DB[458]), .Z(n6446) );
  AND U9523 ( .A(n1786), .B(n6447), .Z(n6445) );
  XOR U9524 ( .A(n6448), .B(n6449), .Z(n6447) );
  XOR U9525 ( .A(DB[458]), .B(DB[451]), .Z(n6449) );
  AND U9526 ( .A(n1790), .B(n6450), .Z(n6448) );
  XOR U9527 ( .A(n6451), .B(n6452), .Z(n6450) );
  XOR U9528 ( .A(DB[451]), .B(DB[444]), .Z(n6452) );
  AND U9529 ( .A(n1794), .B(n6453), .Z(n6451) );
  XOR U9530 ( .A(n6454), .B(n6455), .Z(n6453) );
  XOR U9531 ( .A(DB[444]), .B(DB[437]), .Z(n6455) );
  AND U9532 ( .A(n1798), .B(n6456), .Z(n6454) );
  XOR U9533 ( .A(n6457), .B(n6458), .Z(n6456) );
  XOR U9534 ( .A(DB[437]), .B(DB[430]), .Z(n6458) );
  AND U9535 ( .A(n1802), .B(n6459), .Z(n6457) );
  XOR U9536 ( .A(n6460), .B(n6461), .Z(n6459) );
  XOR U9537 ( .A(DB[430]), .B(DB[423]), .Z(n6461) );
  AND U9538 ( .A(n1806), .B(n6462), .Z(n6460) );
  XOR U9539 ( .A(n6463), .B(n6464), .Z(n6462) );
  XOR U9540 ( .A(DB[423]), .B(DB[416]), .Z(n6464) );
  AND U9541 ( .A(n1810), .B(n6465), .Z(n6463) );
  XOR U9542 ( .A(n6466), .B(n6467), .Z(n6465) );
  XOR U9543 ( .A(DB[416]), .B(DB[409]), .Z(n6467) );
  AND U9544 ( .A(n1814), .B(n6468), .Z(n6466) );
  XOR U9545 ( .A(n6469), .B(n6470), .Z(n6468) );
  XOR U9546 ( .A(DB[409]), .B(DB[402]), .Z(n6470) );
  AND U9547 ( .A(n1818), .B(n6471), .Z(n6469) );
  XOR U9548 ( .A(n6472), .B(n6473), .Z(n6471) );
  XOR U9549 ( .A(DB[402]), .B(DB[395]), .Z(n6473) );
  AND U9550 ( .A(n1822), .B(n6474), .Z(n6472) );
  XOR U9551 ( .A(n6475), .B(n6476), .Z(n6474) );
  XOR U9552 ( .A(DB[395]), .B(DB[388]), .Z(n6476) );
  AND U9553 ( .A(n1826), .B(n6477), .Z(n6475) );
  XOR U9554 ( .A(n6478), .B(n6479), .Z(n6477) );
  XOR U9555 ( .A(DB[388]), .B(DB[381]), .Z(n6479) );
  AND U9556 ( .A(n1830), .B(n6480), .Z(n6478) );
  XOR U9557 ( .A(n6481), .B(n6482), .Z(n6480) );
  XOR U9558 ( .A(DB[381]), .B(DB[374]), .Z(n6482) );
  AND U9559 ( .A(n1834), .B(n6483), .Z(n6481) );
  XOR U9560 ( .A(n6484), .B(n6485), .Z(n6483) );
  XOR U9561 ( .A(DB[374]), .B(DB[367]), .Z(n6485) );
  AND U9562 ( .A(n1838), .B(n6486), .Z(n6484) );
  XOR U9563 ( .A(n6487), .B(n6488), .Z(n6486) );
  XOR U9564 ( .A(DB[367]), .B(DB[360]), .Z(n6488) );
  AND U9565 ( .A(n1842), .B(n6489), .Z(n6487) );
  XOR U9566 ( .A(n6490), .B(n6491), .Z(n6489) );
  XOR U9567 ( .A(DB[360]), .B(DB[353]), .Z(n6491) );
  AND U9568 ( .A(n1846), .B(n6492), .Z(n6490) );
  XOR U9569 ( .A(n6493), .B(n6494), .Z(n6492) );
  XOR U9570 ( .A(DB[353]), .B(DB[346]), .Z(n6494) );
  AND U9571 ( .A(n1850), .B(n6495), .Z(n6493) );
  XOR U9572 ( .A(n6496), .B(n6497), .Z(n6495) );
  XOR U9573 ( .A(DB[346]), .B(DB[339]), .Z(n6497) );
  AND U9574 ( .A(n1854), .B(n6498), .Z(n6496) );
  XOR U9575 ( .A(n6499), .B(n6500), .Z(n6498) );
  XOR U9576 ( .A(DB[339]), .B(DB[332]), .Z(n6500) );
  AND U9577 ( .A(n1858), .B(n6501), .Z(n6499) );
  XOR U9578 ( .A(n6502), .B(n6503), .Z(n6501) );
  XOR U9579 ( .A(DB[332]), .B(DB[325]), .Z(n6503) );
  AND U9580 ( .A(n1862), .B(n6504), .Z(n6502) );
  XOR U9581 ( .A(n6505), .B(n6506), .Z(n6504) );
  XOR U9582 ( .A(DB[325]), .B(DB[318]), .Z(n6506) );
  AND U9583 ( .A(n1866), .B(n6507), .Z(n6505) );
  XOR U9584 ( .A(n6508), .B(n6509), .Z(n6507) );
  XOR U9585 ( .A(DB[318]), .B(DB[311]), .Z(n6509) );
  AND U9586 ( .A(n1870), .B(n6510), .Z(n6508) );
  XOR U9587 ( .A(n6511), .B(n6512), .Z(n6510) );
  XOR U9588 ( .A(DB[311]), .B(DB[304]), .Z(n6512) );
  AND U9589 ( .A(n1874), .B(n6513), .Z(n6511) );
  XOR U9590 ( .A(n6514), .B(n6515), .Z(n6513) );
  XOR U9591 ( .A(DB[304]), .B(DB[297]), .Z(n6515) );
  AND U9592 ( .A(n1878), .B(n6516), .Z(n6514) );
  XOR U9593 ( .A(n6517), .B(n6518), .Z(n6516) );
  XOR U9594 ( .A(DB[297]), .B(DB[290]), .Z(n6518) );
  AND U9595 ( .A(n1882), .B(n6519), .Z(n6517) );
  XOR U9596 ( .A(n6520), .B(n6521), .Z(n6519) );
  XOR U9597 ( .A(DB[290]), .B(DB[283]), .Z(n6521) );
  AND U9598 ( .A(n1886), .B(n6522), .Z(n6520) );
  XOR U9599 ( .A(n6523), .B(n6524), .Z(n6522) );
  XOR U9600 ( .A(DB[283]), .B(DB[276]), .Z(n6524) );
  AND U9601 ( .A(n1890), .B(n6525), .Z(n6523) );
  XOR U9602 ( .A(n6526), .B(n6527), .Z(n6525) );
  XOR U9603 ( .A(DB[276]), .B(DB[269]), .Z(n6527) );
  AND U9604 ( .A(n1894), .B(n6528), .Z(n6526) );
  XOR U9605 ( .A(n6529), .B(n6530), .Z(n6528) );
  XOR U9606 ( .A(DB[269]), .B(DB[262]), .Z(n6530) );
  AND U9607 ( .A(n1898), .B(n6531), .Z(n6529) );
  XOR U9608 ( .A(n6532), .B(n6533), .Z(n6531) );
  XOR U9609 ( .A(DB[262]), .B(DB[255]), .Z(n6533) );
  AND U9610 ( .A(n1902), .B(n6534), .Z(n6532) );
  XOR U9611 ( .A(n6535), .B(n6536), .Z(n6534) );
  XOR U9612 ( .A(DB[255]), .B(DB[248]), .Z(n6536) );
  AND U9613 ( .A(n1906), .B(n6537), .Z(n6535) );
  XOR U9614 ( .A(n6538), .B(n6539), .Z(n6537) );
  XOR U9615 ( .A(DB[248]), .B(DB[241]), .Z(n6539) );
  AND U9616 ( .A(n1910), .B(n6540), .Z(n6538) );
  XOR U9617 ( .A(n6541), .B(n6542), .Z(n6540) );
  XOR U9618 ( .A(DB[241]), .B(DB[234]), .Z(n6542) );
  AND U9619 ( .A(n1914), .B(n6543), .Z(n6541) );
  XOR U9620 ( .A(n6544), .B(n6545), .Z(n6543) );
  XOR U9621 ( .A(DB[234]), .B(DB[227]), .Z(n6545) );
  AND U9622 ( .A(n1918), .B(n6546), .Z(n6544) );
  XOR U9623 ( .A(n6547), .B(n6548), .Z(n6546) );
  XOR U9624 ( .A(DB[227]), .B(DB[220]), .Z(n6548) );
  AND U9625 ( .A(n1922), .B(n6549), .Z(n6547) );
  XOR U9626 ( .A(n6550), .B(n6551), .Z(n6549) );
  XOR U9627 ( .A(DB[220]), .B(DB[213]), .Z(n6551) );
  AND U9628 ( .A(n1926), .B(n6552), .Z(n6550) );
  XOR U9629 ( .A(n6553), .B(n6554), .Z(n6552) );
  XOR U9630 ( .A(DB[213]), .B(DB[206]), .Z(n6554) );
  AND U9631 ( .A(n1930), .B(n6555), .Z(n6553) );
  XOR U9632 ( .A(n6556), .B(n6557), .Z(n6555) );
  XOR U9633 ( .A(DB[206]), .B(DB[199]), .Z(n6557) );
  AND U9634 ( .A(n1934), .B(n6558), .Z(n6556) );
  XOR U9635 ( .A(n6559), .B(n6560), .Z(n6558) );
  XOR U9636 ( .A(DB[199]), .B(DB[192]), .Z(n6560) );
  AND U9637 ( .A(n1938), .B(n6561), .Z(n6559) );
  XOR U9638 ( .A(n6562), .B(n6563), .Z(n6561) );
  XOR U9639 ( .A(DB[192]), .B(DB[185]), .Z(n6563) );
  AND U9640 ( .A(n1942), .B(n6564), .Z(n6562) );
  XOR U9641 ( .A(n6565), .B(n6566), .Z(n6564) );
  XOR U9642 ( .A(DB[185]), .B(DB[178]), .Z(n6566) );
  AND U9643 ( .A(n1946), .B(n6567), .Z(n6565) );
  XOR U9644 ( .A(n6568), .B(n6569), .Z(n6567) );
  XOR U9645 ( .A(DB[178]), .B(DB[171]), .Z(n6569) );
  AND U9646 ( .A(n1950), .B(n6570), .Z(n6568) );
  XOR U9647 ( .A(n6571), .B(n6572), .Z(n6570) );
  XOR U9648 ( .A(DB[171]), .B(DB[164]), .Z(n6572) );
  AND U9649 ( .A(n1954), .B(n6573), .Z(n6571) );
  XOR U9650 ( .A(n6574), .B(n6575), .Z(n6573) );
  XOR U9651 ( .A(DB[164]), .B(DB[157]), .Z(n6575) );
  AND U9652 ( .A(n1958), .B(n6576), .Z(n6574) );
  XOR U9653 ( .A(n6577), .B(n6578), .Z(n6576) );
  XOR U9654 ( .A(DB[157]), .B(DB[150]), .Z(n6578) );
  AND U9655 ( .A(n1962), .B(n6579), .Z(n6577) );
  XOR U9656 ( .A(n6580), .B(n6581), .Z(n6579) );
  XOR U9657 ( .A(DB[150]), .B(DB[143]), .Z(n6581) );
  AND U9658 ( .A(n1966), .B(n6582), .Z(n6580) );
  XOR U9659 ( .A(n6583), .B(n6584), .Z(n6582) );
  XOR U9660 ( .A(DB[143]), .B(DB[136]), .Z(n6584) );
  AND U9661 ( .A(n1970), .B(n6585), .Z(n6583) );
  XOR U9662 ( .A(n6586), .B(n6587), .Z(n6585) );
  XOR U9663 ( .A(DB[136]), .B(DB[129]), .Z(n6587) );
  AND U9664 ( .A(n1974), .B(n6588), .Z(n6586) );
  XOR U9665 ( .A(n6589), .B(n6590), .Z(n6588) );
  XOR U9666 ( .A(DB[129]), .B(DB[122]), .Z(n6590) );
  AND U9667 ( .A(n1978), .B(n6591), .Z(n6589) );
  XOR U9668 ( .A(n6592), .B(n6593), .Z(n6591) );
  XOR U9669 ( .A(DB[122]), .B(DB[115]), .Z(n6593) );
  AND U9670 ( .A(n1982), .B(n6594), .Z(n6592) );
  XOR U9671 ( .A(n6595), .B(n6596), .Z(n6594) );
  XOR U9672 ( .A(DB[115]), .B(DB[108]), .Z(n6596) );
  AND U9673 ( .A(n1986), .B(n6597), .Z(n6595) );
  XOR U9674 ( .A(n6598), .B(n6599), .Z(n6597) );
  XOR U9675 ( .A(DB[108]), .B(DB[101]), .Z(n6599) );
  AND U9676 ( .A(n1990), .B(n6600), .Z(n6598) );
  XOR U9677 ( .A(n6601), .B(n6602), .Z(n6600) );
  XOR U9678 ( .A(DB[94]), .B(DB[101]), .Z(n6602) );
  AND U9679 ( .A(n1994), .B(n6603), .Z(n6601) );
  XOR U9680 ( .A(n6604), .B(n6605), .Z(n6603) );
  XOR U9681 ( .A(DB[94]), .B(DB[87]), .Z(n6605) );
  AND U9682 ( .A(n1998), .B(n6606), .Z(n6604) );
  XOR U9683 ( .A(n6607), .B(n6608), .Z(n6606) );
  XOR U9684 ( .A(DB[87]), .B(DB[80]), .Z(n6608) );
  AND U9685 ( .A(n2002), .B(n6609), .Z(n6607) );
  XOR U9686 ( .A(n6610), .B(n6611), .Z(n6609) );
  XOR U9687 ( .A(DB[80]), .B(DB[73]), .Z(n6611) );
  AND U9688 ( .A(n2006), .B(n6612), .Z(n6610) );
  XOR U9689 ( .A(n6613), .B(n6614), .Z(n6612) );
  XOR U9690 ( .A(DB[73]), .B(DB[66]), .Z(n6614) );
  AND U9691 ( .A(n2010), .B(n6615), .Z(n6613) );
  XOR U9692 ( .A(n6616), .B(n6617), .Z(n6615) );
  XOR U9693 ( .A(DB[66]), .B(DB[59]), .Z(n6617) );
  AND U9694 ( .A(n2014), .B(n6618), .Z(n6616) );
  XOR U9695 ( .A(n6619), .B(n6620), .Z(n6618) );
  XOR U9696 ( .A(DB[59]), .B(DB[52]), .Z(n6620) );
  AND U9697 ( .A(n2018), .B(n6621), .Z(n6619) );
  XOR U9698 ( .A(n6622), .B(n6623), .Z(n6621) );
  XOR U9699 ( .A(DB[52]), .B(DB[45]), .Z(n6623) );
  AND U9700 ( .A(n2022), .B(n6624), .Z(n6622) );
  XOR U9701 ( .A(n6625), .B(n6626), .Z(n6624) );
  XOR U9702 ( .A(DB[45]), .B(DB[38]), .Z(n6626) );
  AND U9703 ( .A(n2026), .B(n6627), .Z(n6625) );
  XOR U9704 ( .A(n6628), .B(n6629), .Z(n6627) );
  XOR U9705 ( .A(DB[38]), .B(DB[31]), .Z(n6629) );
  AND U9706 ( .A(n2030), .B(n6630), .Z(n6628) );
  XOR U9707 ( .A(n6631), .B(n6632), .Z(n6630) );
  XOR U9708 ( .A(DB[31]), .B(DB[24]), .Z(n6632) );
  AND U9709 ( .A(n2034), .B(n6633), .Z(n6631) );
  XOR U9710 ( .A(n6634), .B(n6635), .Z(n6633) );
  XOR U9711 ( .A(DB[24]), .B(DB[17]), .Z(n6635) );
  AND U9712 ( .A(n2038), .B(n6636), .Z(n6634) );
  XOR U9713 ( .A(n6637), .B(n6638), .Z(n6636) );
  XOR U9714 ( .A(DB[17]), .B(DB[10]), .Z(n6638) );
  AND U9715 ( .A(n2042), .B(n6639), .Z(n6637) );
  XOR U9716 ( .A(DB[3]), .B(DB[10]), .Z(n6639) );
  XOR U9717 ( .A(DB[3579]), .B(n6640), .Z(min_val_out[2]) );
  AND U9718 ( .A(n2), .B(n6641), .Z(n6640) );
  XOR U9719 ( .A(n6642), .B(n6643), .Z(n6641) );
  XOR U9720 ( .A(DB[3579]), .B(DB[3572]), .Z(n6643) );
  AND U9721 ( .A(n6), .B(n6644), .Z(n6642) );
  XOR U9722 ( .A(n6645), .B(n6646), .Z(n6644) );
  XOR U9723 ( .A(DB[3572]), .B(DB[3565]), .Z(n6646) );
  AND U9724 ( .A(n10), .B(n6647), .Z(n6645) );
  XOR U9725 ( .A(n6648), .B(n6649), .Z(n6647) );
  XOR U9726 ( .A(DB[3565]), .B(DB[3558]), .Z(n6649) );
  AND U9727 ( .A(n14), .B(n6650), .Z(n6648) );
  XOR U9728 ( .A(n6651), .B(n6652), .Z(n6650) );
  XOR U9729 ( .A(DB[3558]), .B(DB[3551]), .Z(n6652) );
  AND U9730 ( .A(n18), .B(n6653), .Z(n6651) );
  XOR U9731 ( .A(n6654), .B(n6655), .Z(n6653) );
  XOR U9732 ( .A(DB[3551]), .B(DB[3544]), .Z(n6655) );
  AND U9733 ( .A(n22), .B(n6656), .Z(n6654) );
  XOR U9734 ( .A(n6657), .B(n6658), .Z(n6656) );
  XOR U9735 ( .A(DB[3544]), .B(DB[3537]), .Z(n6658) );
  AND U9736 ( .A(n26), .B(n6659), .Z(n6657) );
  XOR U9737 ( .A(n6660), .B(n6661), .Z(n6659) );
  XOR U9738 ( .A(DB[3537]), .B(DB[3530]), .Z(n6661) );
  AND U9739 ( .A(n30), .B(n6662), .Z(n6660) );
  XOR U9740 ( .A(n6663), .B(n6664), .Z(n6662) );
  XOR U9741 ( .A(DB[3530]), .B(DB[3523]), .Z(n6664) );
  AND U9742 ( .A(n34), .B(n6665), .Z(n6663) );
  XOR U9743 ( .A(n6666), .B(n6667), .Z(n6665) );
  XOR U9744 ( .A(DB[3523]), .B(DB[3516]), .Z(n6667) );
  AND U9745 ( .A(n38), .B(n6668), .Z(n6666) );
  XOR U9746 ( .A(n6669), .B(n6670), .Z(n6668) );
  XOR U9747 ( .A(DB[3516]), .B(DB[3509]), .Z(n6670) );
  AND U9748 ( .A(n42), .B(n6671), .Z(n6669) );
  XOR U9749 ( .A(n6672), .B(n6673), .Z(n6671) );
  XOR U9750 ( .A(DB[3509]), .B(DB[3502]), .Z(n6673) );
  AND U9751 ( .A(n46), .B(n6674), .Z(n6672) );
  XOR U9752 ( .A(n6675), .B(n6676), .Z(n6674) );
  XOR U9753 ( .A(DB[3502]), .B(DB[3495]), .Z(n6676) );
  AND U9754 ( .A(n50), .B(n6677), .Z(n6675) );
  XOR U9755 ( .A(n6678), .B(n6679), .Z(n6677) );
  XOR U9756 ( .A(DB[3495]), .B(DB[3488]), .Z(n6679) );
  AND U9757 ( .A(n54), .B(n6680), .Z(n6678) );
  XOR U9758 ( .A(n6681), .B(n6682), .Z(n6680) );
  XOR U9759 ( .A(DB[3488]), .B(DB[3481]), .Z(n6682) );
  AND U9760 ( .A(n58), .B(n6683), .Z(n6681) );
  XOR U9761 ( .A(n6684), .B(n6685), .Z(n6683) );
  XOR U9762 ( .A(DB[3481]), .B(DB[3474]), .Z(n6685) );
  AND U9763 ( .A(n62), .B(n6686), .Z(n6684) );
  XOR U9764 ( .A(n6687), .B(n6688), .Z(n6686) );
  XOR U9765 ( .A(DB[3474]), .B(DB[3467]), .Z(n6688) );
  AND U9766 ( .A(n66), .B(n6689), .Z(n6687) );
  XOR U9767 ( .A(n6690), .B(n6691), .Z(n6689) );
  XOR U9768 ( .A(DB[3467]), .B(DB[3460]), .Z(n6691) );
  AND U9769 ( .A(n70), .B(n6692), .Z(n6690) );
  XOR U9770 ( .A(n6693), .B(n6694), .Z(n6692) );
  XOR U9771 ( .A(DB[3460]), .B(DB[3453]), .Z(n6694) );
  AND U9772 ( .A(n74), .B(n6695), .Z(n6693) );
  XOR U9773 ( .A(n6696), .B(n6697), .Z(n6695) );
  XOR U9774 ( .A(DB[3453]), .B(DB[3446]), .Z(n6697) );
  AND U9775 ( .A(n78), .B(n6698), .Z(n6696) );
  XOR U9776 ( .A(n6699), .B(n6700), .Z(n6698) );
  XOR U9777 ( .A(DB[3446]), .B(DB[3439]), .Z(n6700) );
  AND U9778 ( .A(n82), .B(n6701), .Z(n6699) );
  XOR U9779 ( .A(n6702), .B(n6703), .Z(n6701) );
  XOR U9780 ( .A(DB[3439]), .B(DB[3432]), .Z(n6703) );
  AND U9781 ( .A(n86), .B(n6704), .Z(n6702) );
  XOR U9782 ( .A(n6705), .B(n6706), .Z(n6704) );
  XOR U9783 ( .A(DB[3432]), .B(DB[3425]), .Z(n6706) );
  AND U9784 ( .A(n90), .B(n6707), .Z(n6705) );
  XOR U9785 ( .A(n6708), .B(n6709), .Z(n6707) );
  XOR U9786 ( .A(DB[3425]), .B(DB[3418]), .Z(n6709) );
  AND U9787 ( .A(n94), .B(n6710), .Z(n6708) );
  XOR U9788 ( .A(n6711), .B(n6712), .Z(n6710) );
  XOR U9789 ( .A(DB[3418]), .B(DB[3411]), .Z(n6712) );
  AND U9790 ( .A(n98), .B(n6713), .Z(n6711) );
  XOR U9791 ( .A(n6714), .B(n6715), .Z(n6713) );
  XOR U9792 ( .A(DB[3411]), .B(DB[3404]), .Z(n6715) );
  AND U9793 ( .A(n102), .B(n6716), .Z(n6714) );
  XOR U9794 ( .A(n6717), .B(n6718), .Z(n6716) );
  XOR U9795 ( .A(DB[3404]), .B(DB[3397]), .Z(n6718) );
  AND U9796 ( .A(n106), .B(n6719), .Z(n6717) );
  XOR U9797 ( .A(n6720), .B(n6721), .Z(n6719) );
  XOR U9798 ( .A(DB[3397]), .B(DB[3390]), .Z(n6721) );
  AND U9799 ( .A(n110), .B(n6722), .Z(n6720) );
  XOR U9800 ( .A(n6723), .B(n6724), .Z(n6722) );
  XOR U9801 ( .A(DB[3390]), .B(DB[3383]), .Z(n6724) );
  AND U9802 ( .A(n114), .B(n6725), .Z(n6723) );
  XOR U9803 ( .A(n6726), .B(n6727), .Z(n6725) );
  XOR U9804 ( .A(DB[3383]), .B(DB[3376]), .Z(n6727) );
  AND U9805 ( .A(n118), .B(n6728), .Z(n6726) );
  XOR U9806 ( .A(n6729), .B(n6730), .Z(n6728) );
  XOR U9807 ( .A(DB[3376]), .B(DB[3369]), .Z(n6730) );
  AND U9808 ( .A(n122), .B(n6731), .Z(n6729) );
  XOR U9809 ( .A(n6732), .B(n6733), .Z(n6731) );
  XOR U9810 ( .A(DB[3369]), .B(DB[3362]), .Z(n6733) );
  AND U9811 ( .A(n126), .B(n6734), .Z(n6732) );
  XOR U9812 ( .A(n6735), .B(n6736), .Z(n6734) );
  XOR U9813 ( .A(DB[3362]), .B(DB[3355]), .Z(n6736) );
  AND U9814 ( .A(n130), .B(n6737), .Z(n6735) );
  XOR U9815 ( .A(n6738), .B(n6739), .Z(n6737) );
  XOR U9816 ( .A(DB[3355]), .B(DB[3348]), .Z(n6739) );
  AND U9817 ( .A(n134), .B(n6740), .Z(n6738) );
  XOR U9818 ( .A(n6741), .B(n6742), .Z(n6740) );
  XOR U9819 ( .A(DB[3348]), .B(DB[3341]), .Z(n6742) );
  AND U9820 ( .A(n138), .B(n6743), .Z(n6741) );
  XOR U9821 ( .A(n6744), .B(n6745), .Z(n6743) );
  XOR U9822 ( .A(DB[3341]), .B(DB[3334]), .Z(n6745) );
  AND U9823 ( .A(n142), .B(n6746), .Z(n6744) );
  XOR U9824 ( .A(n6747), .B(n6748), .Z(n6746) );
  XOR U9825 ( .A(DB[3334]), .B(DB[3327]), .Z(n6748) );
  AND U9826 ( .A(n146), .B(n6749), .Z(n6747) );
  XOR U9827 ( .A(n6750), .B(n6751), .Z(n6749) );
  XOR U9828 ( .A(DB[3327]), .B(DB[3320]), .Z(n6751) );
  AND U9829 ( .A(n150), .B(n6752), .Z(n6750) );
  XOR U9830 ( .A(n6753), .B(n6754), .Z(n6752) );
  XOR U9831 ( .A(DB[3320]), .B(DB[3313]), .Z(n6754) );
  AND U9832 ( .A(n154), .B(n6755), .Z(n6753) );
  XOR U9833 ( .A(n6756), .B(n6757), .Z(n6755) );
  XOR U9834 ( .A(DB[3313]), .B(DB[3306]), .Z(n6757) );
  AND U9835 ( .A(n158), .B(n6758), .Z(n6756) );
  XOR U9836 ( .A(n6759), .B(n6760), .Z(n6758) );
  XOR U9837 ( .A(DB[3306]), .B(DB[3299]), .Z(n6760) );
  AND U9838 ( .A(n162), .B(n6761), .Z(n6759) );
  XOR U9839 ( .A(n6762), .B(n6763), .Z(n6761) );
  XOR U9840 ( .A(DB[3299]), .B(DB[3292]), .Z(n6763) );
  AND U9841 ( .A(n166), .B(n6764), .Z(n6762) );
  XOR U9842 ( .A(n6765), .B(n6766), .Z(n6764) );
  XOR U9843 ( .A(DB[3292]), .B(DB[3285]), .Z(n6766) );
  AND U9844 ( .A(n170), .B(n6767), .Z(n6765) );
  XOR U9845 ( .A(n6768), .B(n6769), .Z(n6767) );
  XOR U9846 ( .A(DB[3285]), .B(DB[3278]), .Z(n6769) );
  AND U9847 ( .A(n174), .B(n6770), .Z(n6768) );
  XOR U9848 ( .A(n6771), .B(n6772), .Z(n6770) );
  XOR U9849 ( .A(DB[3278]), .B(DB[3271]), .Z(n6772) );
  AND U9850 ( .A(n178), .B(n6773), .Z(n6771) );
  XOR U9851 ( .A(n6774), .B(n6775), .Z(n6773) );
  XOR U9852 ( .A(DB[3271]), .B(DB[3264]), .Z(n6775) );
  AND U9853 ( .A(n182), .B(n6776), .Z(n6774) );
  XOR U9854 ( .A(n6777), .B(n6778), .Z(n6776) );
  XOR U9855 ( .A(DB[3264]), .B(DB[3257]), .Z(n6778) );
  AND U9856 ( .A(n186), .B(n6779), .Z(n6777) );
  XOR U9857 ( .A(n6780), .B(n6781), .Z(n6779) );
  XOR U9858 ( .A(DB[3257]), .B(DB[3250]), .Z(n6781) );
  AND U9859 ( .A(n190), .B(n6782), .Z(n6780) );
  XOR U9860 ( .A(n6783), .B(n6784), .Z(n6782) );
  XOR U9861 ( .A(DB[3250]), .B(DB[3243]), .Z(n6784) );
  AND U9862 ( .A(n194), .B(n6785), .Z(n6783) );
  XOR U9863 ( .A(n6786), .B(n6787), .Z(n6785) );
  XOR U9864 ( .A(DB[3243]), .B(DB[3236]), .Z(n6787) );
  AND U9865 ( .A(n198), .B(n6788), .Z(n6786) );
  XOR U9866 ( .A(n6789), .B(n6790), .Z(n6788) );
  XOR U9867 ( .A(DB[3236]), .B(DB[3229]), .Z(n6790) );
  AND U9868 ( .A(n202), .B(n6791), .Z(n6789) );
  XOR U9869 ( .A(n6792), .B(n6793), .Z(n6791) );
  XOR U9870 ( .A(DB[3229]), .B(DB[3222]), .Z(n6793) );
  AND U9871 ( .A(n206), .B(n6794), .Z(n6792) );
  XOR U9872 ( .A(n6795), .B(n6796), .Z(n6794) );
  XOR U9873 ( .A(DB[3222]), .B(DB[3215]), .Z(n6796) );
  AND U9874 ( .A(n210), .B(n6797), .Z(n6795) );
  XOR U9875 ( .A(n6798), .B(n6799), .Z(n6797) );
  XOR U9876 ( .A(DB[3215]), .B(DB[3208]), .Z(n6799) );
  AND U9877 ( .A(n214), .B(n6800), .Z(n6798) );
  XOR U9878 ( .A(n6801), .B(n6802), .Z(n6800) );
  XOR U9879 ( .A(DB[3208]), .B(DB[3201]), .Z(n6802) );
  AND U9880 ( .A(n218), .B(n6803), .Z(n6801) );
  XOR U9881 ( .A(n6804), .B(n6805), .Z(n6803) );
  XOR U9882 ( .A(DB[3201]), .B(DB[3194]), .Z(n6805) );
  AND U9883 ( .A(n222), .B(n6806), .Z(n6804) );
  XOR U9884 ( .A(n6807), .B(n6808), .Z(n6806) );
  XOR U9885 ( .A(DB[3194]), .B(DB[3187]), .Z(n6808) );
  AND U9886 ( .A(n226), .B(n6809), .Z(n6807) );
  XOR U9887 ( .A(n6810), .B(n6811), .Z(n6809) );
  XOR U9888 ( .A(DB[3187]), .B(DB[3180]), .Z(n6811) );
  AND U9889 ( .A(n230), .B(n6812), .Z(n6810) );
  XOR U9890 ( .A(n6813), .B(n6814), .Z(n6812) );
  XOR U9891 ( .A(DB[3180]), .B(DB[3173]), .Z(n6814) );
  AND U9892 ( .A(n234), .B(n6815), .Z(n6813) );
  XOR U9893 ( .A(n6816), .B(n6817), .Z(n6815) );
  XOR U9894 ( .A(DB[3173]), .B(DB[3166]), .Z(n6817) );
  AND U9895 ( .A(n238), .B(n6818), .Z(n6816) );
  XOR U9896 ( .A(n6819), .B(n6820), .Z(n6818) );
  XOR U9897 ( .A(DB[3166]), .B(DB[3159]), .Z(n6820) );
  AND U9898 ( .A(n242), .B(n6821), .Z(n6819) );
  XOR U9899 ( .A(n6822), .B(n6823), .Z(n6821) );
  XOR U9900 ( .A(DB[3159]), .B(DB[3152]), .Z(n6823) );
  AND U9901 ( .A(n246), .B(n6824), .Z(n6822) );
  XOR U9902 ( .A(n6825), .B(n6826), .Z(n6824) );
  XOR U9903 ( .A(DB[3152]), .B(DB[3145]), .Z(n6826) );
  AND U9904 ( .A(n250), .B(n6827), .Z(n6825) );
  XOR U9905 ( .A(n6828), .B(n6829), .Z(n6827) );
  XOR U9906 ( .A(DB[3145]), .B(DB[3138]), .Z(n6829) );
  AND U9907 ( .A(n254), .B(n6830), .Z(n6828) );
  XOR U9908 ( .A(n6831), .B(n6832), .Z(n6830) );
  XOR U9909 ( .A(DB[3138]), .B(DB[3131]), .Z(n6832) );
  AND U9910 ( .A(n258), .B(n6833), .Z(n6831) );
  XOR U9911 ( .A(n6834), .B(n6835), .Z(n6833) );
  XOR U9912 ( .A(DB[3131]), .B(DB[3124]), .Z(n6835) );
  AND U9913 ( .A(n262), .B(n6836), .Z(n6834) );
  XOR U9914 ( .A(n6837), .B(n6838), .Z(n6836) );
  XOR U9915 ( .A(DB[3124]), .B(DB[3117]), .Z(n6838) );
  AND U9916 ( .A(n266), .B(n6839), .Z(n6837) );
  XOR U9917 ( .A(n6840), .B(n6841), .Z(n6839) );
  XOR U9918 ( .A(DB[3117]), .B(DB[3110]), .Z(n6841) );
  AND U9919 ( .A(n270), .B(n6842), .Z(n6840) );
  XOR U9920 ( .A(n6843), .B(n6844), .Z(n6842) );
  XOR U9921 ( .A(DB[3110]), .B(DB[3103]), .Z(n6844) );
  AND U9922 ( .A(n274), .B(n6845), .Z(n6843) );
  XOR U9923 ( .A(n6846), .B(n6847), .Z(n6845) );
  XOR U9924 ( .A(DB[3103]), .B(DB[3096]), .Z(n6847) );
  AND U9925 ( .A(n278), .B(n6848), .Z(n6846) );
  XOR U9926 ( .A(n6849), .B(n6850), .Z(n6848) );
  XOR U9927 ( .A(DB[3096]), .B(DB[3089]), .Z(n6850) );
  AND U9928 ( .A(n282), .B(n6851), .Z(n6849) );
  XOR U9929 ( .A(n6852), .B(n6853), .Z(n6851) );
  XOR U9930 ( .A(DB[3089]), .B(DB[3082]), .Z(n6853) );
  AND U9931 ( .A(n286), .B(n6854), .Z(n6852) );
  XOR U9932 ( .A(n6855), .B(n6856), .Z(n6854) );
  XOR U9933 ( .A(DB[3082]), .B(DB[3075]), .Z(n6856) );
  AND U9934 ( .A(n290), .B(n6857), .Z(n6855) );
  XOR U9935 ( .A(n6858), .B(n6859), .Z(n6857) );
  XOR U9936 ( .A(DB[3075]), .B(DB[3068]), .Z(n6859) );
  AND U9937 ( .A(n294), .B(n6860), .Z(n6858) );
  XOR U9938 ( .A(n6861), .B(n6862), .Z(n6860) );
  XOR U9939 ( .A(DB[3068]), .B(DB[3061]), .Z(n6862) );
  AND U9940 ( .A(n298), .B(n6863), .Z(n6861) );
  XOR U9941 ( .A(n6864), .B(n6865), .Z(n6863) );
  XOR U9942 ( .A(DB[3061]), .B(DB[3054]), .Z(n6865) );
  AND U9943 ( .A(n302), .B(n6866), .Z(n6864) );
  XOR U9944 ( .A(n6867), .B(n6868), .Z(n6866) );
  XOR U9945 ( .A(DB[3054]), .B(DB[3047]), .Z(n6868) );
  AND U9946 ( .A(n306), .B(n6869), .Z(n6867) );
  XOR U9947 ( .A(n6870), .B(n6871), .Z(n6869) );
  XOR U9948 ( .A(DB[3047]), .B(DB[3040]), .Z(n6871) );
  AND U9949 ( .A(n310), .B(n6872), .Z(n6870) );
  XOR U9950 ( .A(n6873), .B(n6874), .Z(n6872) );
  XOR U9951 ( .A(DB[3040]), .B(DB[3033]), .Z(n6874) );
  AND U9952 ( .A(n314), .B(n6875), .Z(n6873) );
  XOR U9953 ( .A(n6876), .B(n6877), .Z(n6875) );
  XOR U9954 ( .A(DB[3033]), .B(DB[3026]), .Z(n6877) );
  AND U9955 ( .A(n318), .B(n6878), .Z(n6876) );
  XOR U9956 ( .A(n6879), .B(n6880), .Z(n6878) );
  XOR U9957 ( .A(DB[3026]), .B(DB[3019]), .Z(n6880) );
  AND U9958 ( .A(n322), .B(n6881), .Z(n6879) );
  XOR U9959 ( .A(n6882), .B(n6883), .Z(n6881) );
  XOR U9960 ( .A(DB[3019]), .B(DB[3012]), .Z(n6883) );
  AND U9961 ( .A(n326), .B(n6884), .Z(n6882) );
  XOR U9962 ( .A(n6885), .B(n6886), .Z(n6884) );
  XOR U9963 ( .A(DB[3012]), .B(DB[3005]), .Z(n6886) );
  AND U9964 ( .A(n330), .B(n6887), .Z(n6885) );
  XOR U9965 ( .A(n6888), .B(n6889), .Z(n6887) );
  XOR U9966 ( .A(DB[3005]), .B(DB[2998]), .Z(n6889) );
  AND U9967 ( .A(n334), .B(n6890), .Z(n6888) );
  XOR U9968 ( .A(n6891), .B(n6892), .Z(n6890) );
  XOR U9969 ( .A(DB[2998]), .B(DB[2991]), .Z(n6892) );
  AND U9970 ( .A(n338), .B(n6893), .Z(n6891) );
  XOR U9971 ( .A(n6894), .B(n6895), .Z(n6893) );
  XOR U9972 ( .A(DB[2991]), .B(DB[2984]), .Z(n6895) );
  AND U9973 ( .A(n342), .B(n6896), .Z(n6894) );
  XOR U9974 ( .A(n6897), .B(n6898), .Z(n6896) );
  XOR U9975 ( .A(DB[2984]), .B(DB[2977]), .Z(n6898) );
  AND U9976 ( .A(n346), .B(n6899), .Z(n6897) );
  XOR U9977 ( .A(n6900), .B(n6901), .Z(n6899) );
  XOR U9978 ( .A(DB[2977]), .B(DB[2970]), .Z(n6901) );
  AND U9979 ( .A(n350), .B(n6902), .Z(n6900) );
  XOR U9980 ( .A(n6903), .B(n6904), .Z(n6902) );
  XOR U9981 ( .A(DB[2970]), .B(DB[2963]), .Z(n6904) );
  AND U9982 ( .A(n354), .B(n6905), .Z(n6903) );
  XOR U9983 ( .A(n6906), .B(n6907), .Z(n6905) );
  XOR U9984 ( .A(DB[2963]), .B(DB[2956]), .Z(n6907) );
  AND U9985 ( .A(n358), .B(n6908), .Z(n6906) );
  XOR U9986 ( .A(n6909), .B(n6910), .Z(n6908) );
  XOR U9987 ( .A(DB[2956]), .B(DB[2949]), .Z(n6910) );
  AND U9988 ( .A(n362), .B(n6911), .Z(n6909) );
  XOR U9989 ( .A(n6912), .B(n6913), .Z(n6911) );
  XOR U9990 ( .A(DB[2949]), .B(DB[2942]), .Z(n6913) );
  AND U9991 ( .A(n366), .B(n6914), .Z(n6912) );
  XOR U9992 ( .A(n6915), .B(n6916), .Z(n6914) );
  XOR U9993 ( .A(DB[2942]), .B(DB[2935]), .Z(n6916) );
  AND U9994 ( .A(n370), .B(n6917), .Z(n6915) );
  XOR U9995 ( .A(n6918), .B(n6919), .Z(n6917) );
  XOR U9996 ( .A(DB[2935]), .B(DB[2928]), .Z(n6919) );
  AND U9997 ( .A(n374), .B(n6920), .Z(n6918) );
  XOR U9998 ( .A(n6921), .B(n6922), .Z(n6920) );
  XOR U9999 ( .A(DB[2928]), .B(DB[2921]), .Z(n6922) );
  AND U10000 ( .A(n378), .B(n6923), .Z(n6921) );
  XOR U10001 ( .A(n6924), .B(n6925), .Z(n6923) );
  XOR U10002 ( .A(DB[2921]), .B(DB[2914]), .Z(n6925) );
  AND U10003 ( .A(n382), .B(n6926), .Z(n6924) );
  XOR U10004 ( .A(n6927), .B(n6928), .Z(n6926) );
  XOR U10005 ( .A(DB[2914]), .B(DB[2907]), .Z(n6928) );
  AND U10006 ( .A(n386), .B(n6929), .Z(n6927) );
  XOR U10007 ( .A(n6930), .B(n6931), .Z(n6929) );
  XOR U10008 ( .A(DB[2907]), .B(DB[2900]), .Z(n6931) );
  AND U10009 ( .A(n390), .B(n6932), .Z(n6930) );
  XOR U10010 ( .A(n6933), .B(n6934), .Z(n6932) );
  XOR U10011 ( .A(DB[2900]), .B(DB[2893]), .Z(n6934) );
  AND U10012 ( .A(n394), .B(n6935), .Z(n6933) );
  XOR U10013 ( .A(n6936), .B(n6937), .Z(n6935) );
  XOR U10014 ( .A(DB[2893]), .B(DB[2886]), .Z(n6937) );
  AND U10015 ( .A(n398), .B(n6938), .Z(n6936) );
  XOR U10016 ( .A(n6939), .B(n6940), .Z(n6938) );
  XOR U10017 ( .A(DB[2886]), .B(DB[2879]), .Z(n6940) );
  AND U10018 ( .A(n402), .B(n6941), .Z(n6939) );
  XOR U10019 ( .A(n6942), .B(n6943), .Z(n6941) );
  XOR U10020 ( .A(DB[2879]), .B(DB[2872]), .Z(n6943) );
  AND U10021 ( .A(n406), .B(n6944), .Z(n6942) );
  XOR U10022 ( .A(n6945), .B(n6946), .Z(n6944) );
  XOR U10023 ( .A(DB[2872]), .B(DB[2865]), .Z(n6946) );
  AND U10024 ( .A(n410), .B(n6947), .Z(n6945) );
  XOR U10025 ( .A(n6948), .B(n6949), .Z(n6947) );
  XOR U10026 ( .A(DB[2865]), .B(DB[2858]), .Z(n6949) );
  AND U10027 ( .A(n414), .B(n6950), .Z(n6948) );
  XOR U10028 ( .A(n6951), .B(n6952), .Z(n6950) );
  XOR U10029 ( .A(DB[2858]), .B(DB[2851]), .Z(n6952) );
  AND U10030 ( .A(n418), .B(n6953), .Z(n6951) );
  XOR U10031 ( .A(n6954), .B(n6955), .Z(n6953) );
  XOR U10032 ( .A(DB[2851]), .B(DB[2844]), .Z(n6955) );
  AND U10033 ( .A(n422), .B(n6956), .Z(n6954) );
  XOR U10034 ( .A(n6957), .B(n6958), .Z(n6956) );
  XOR U10035 ( .A(DB[2844]), .B(DB[2837]), .Z(n6958) );
  AND U10036 ( .A(n426), .B(n6959), .Z(n6957) );
  XOR U10037 ( .A(n6960), .B(n6961), .Z(n6959) );
  XOR U10038 ( .A(DB[2837]), .B(DB[2830]), .Z(n6961) );
  AND U10039 ( .A(n430), .B(n6962), .Z(n6960) );
  XOR U10040 ( .A(n6963), .B(n6964), .Z(n6962) );
  XOR U10041 ( .A(DB[2830]), .B(DB[2823]), .Z(n6964) );
  AND U10042 ( .A(n434), .B(n6965), .Z(n6963) );
  XOR U10043 ( .A(n6966), .B(n6967), .Z(n6965) );
  XOR U10044 ( .A(DB[2823]), .B(DB[2816]), .Z(n6967) );
  AND U10045 ( .A(n438), .B(n6968), .Z(n6966) );
  XOR U10046 ( .A(n6969), .B(n6970), .Z(n6968) );
  XOR U10047 ( .A(DB[2816]), .B(DB[2809]), .Z(n6970) );
  AND U10048 ( .A(n442), .B(n6971), .Z(n6969) );
  XOR U10049 ( .A(n6972), .B(n6973), .Z(n6971) );
  XOR U10050 ( .A(DB[2809]), .B(DB[2802]), .Z(n6973) );
  AND U10051 ( .A(n446), .B(n6974), .Z(n6972) );
  XOR U10052 ( .A(n6975), .B(n6976), .Z(n6974) );
  XOR U10053 ( .A(DB[2802]), .B(DB[2795]), .Z(n6976) );
  AND U10054 ( .A(n450), .B(n6977), .Z(n6975) );
  XOR U10055 ( .A(n6978), .B(n6979), .Z(n6977) );
  XOR U10056 ( .A(DB[2795]), .B(DB[2788]), .Z(n6979) );
  AND U10057 ( .A(n454), .B(n6980), .Z(n6978) );
  XOR U10058 ( .A(n6981), .B(n6982), .Z(n6980) );
  XOR U10059 ( .A(DB[2788]), .B(DB[2781]), .Z(n6982) );
  AND U10060 ( .A(n458), .B(n6983), .Z(n6981) );
  XOR U10061 ( .A(n6984), .B(n6985), .Z(n6983) );
  XOR U10062 ( .A(DB[2781]), .B(DB[2774]), .Z(n6985) );
  AND U10063 ( .A(n462), .B(n6986), .Z(n6984) );
  XOR U10064 ( .A(n6987), .B(n6988), .Z(n6986) );
  XOR U10065 ( .A(DB[2774]), .B(DB[2767]), .Z(n6988) );
  AND U10066 ( .A(n466), .B(n6989), .Z(n6987) );
  XOR U10067 ( .A(n6990), .B(n6991), .Z(n6989) );
  XOR U10068 ( .A(DB[2767]), .B(DB[2760]), .Z(n6991) );
  AND U10069 ( .A(n470), .B(n6992), .Z(n6990) );
  XOR U10070 ( .A(n6993), .B(n6994), .Z(n6992) );
  XOR U10071 ( .A(DB[2760]), .B(DB[2753]), .Z(n6994) );
  AND U10072 ( .A(n474), .B(n6995), .Z(n6993) );
  XOR U10073 ( .A(n6996), .B(n6997), .Z(n6995) );
  XOR U10074 ( .A(DB[2753]), .B(DB[2746]), .Z(n6997) );
  AND U10075 ( .A(n478), .B(n6998), .Z(n6996) );
  XOR U10076 ( .A(n6999), .B(n7000), .Z(n6998) );
  XOR U10077 ( .A(DB[2746]), .B(DB[2739]), .Z(n7000) );
  AND U10078 ( .A(n482), .B(n7001), .Z(n6999) );
  XOR U10079 ( .A(n7002), .B(n7003), .Z(n7001) );
  XOR U10080 ( .A(DB[2739]), .B(DB[2732]), .Z(n7003) );
  AND U10081 ( .A(n486), .B(n7004), .Z(n7002) );
  XOR U10082 ( .A(n7005), .B(n7006), .Z(n7004) );
  XOR U10083 ( .A(DB[2732]), .B(DB[2725]), .Z(n7006) );
  AND U10084 ( .A(n490), .B(n7007), .Z(n7005) );
  XOR U10085 ( .A(n7008), .B(n7009), .Z(n7007) );
  XOR U10086 ( .A(DB[2725]), .B(DB[2718]), .Z(n7009) );
  AND U10087 ( .A(n494), .B(n7010), .Z(n7008) );
  XOR U10088 ( .A(n7011), .B(n7012), .Z(n7010) );
  XOR U10089 ( .A(DB[2718]), .B(DB[2711]), .Z(n7012) );
  AND U10090 ( .A(n498), .B(n7013), .Z(n7011) );
  XOR U10091 ( .A(n7014), .B(n7015), .Z(n7013) );
  XOR U10092 ( .A(DB[2711]), .B(DB[2704]), .Z(n7015) );
  AND U10093 ( .A(n502), .B(n7016), .Z(n7014) );
  XOR U10094 ( .A(n7017), .B(n7018), .Z(n7016) );
  XOR U10095 ( .A(DB[2704]), .B(DB[2697]), .Z(n7018) );
  AND U10096 ( .A(n506), .B(n7019), .Z(n7017) );
  XOR U10097 ( .A(n7020), .B(n7021), .Z(n7019) );
  XOR U10098 ( .A(DB[2697]), .B(DB[2690]), .Z(n7021) );
  AND U10099 ( .A(n510), .B(n7022), .Z(n7020) );
  XOR U10100 ( .A(n7023), .B(n7024), .Z(n7022) );
  XOR U10101 ( .A(DB[2690]), .B(DB[2683]), .Z(n7024) );
  AND U10102 ( .A(n514), .B(n7025), .Z(n7023) );
  XOR U10103 ( .A(n7026), .B(n7027), .Z(n7025) );
  XOR U10104 ( .A(DB[2683]), .B(DB[2676]), .Z(n7027) );
  AND U10105 ( .A(n518), .B(n7028), .Z(n7026) );
  XOR U10106 ( .A(n7029), .B(n7030), .Z(n7028) );
  XOR U10107 ( .A(DB[2676]), .B(DB[2669]), .Z(n7030) );
  AND U10108 ( .A(n522), .B(n7031), .Z(n7029) );
  XOR U10109 ( .A(n7032), .B(n7033), .Z(n7031) );
  XOR U10110 ( .A(DB[2669]), .B(DB[2662]), .Z(n7033) );
  AND U10111 ( .A(n526), .B(n7034), .Z(n7032) );
  XOR U10112 ( .A(n7035), .B(n7036), .Z(n7034) );
  XOR U10113 ( .A(DB[2662]), .B(DB[2655]), .Z(n7036) );
  AND U10114 ( .A(n530), .B(n7037), .Z(n7035) );
  XOR U10115 ( .A(n7038), .B(n7039), .Z(n7037) );
  XOR U10116 ( .A(DB[2655]), .B(DB[2648]), .Z(n7039) );
  AND U10117 ( .A(n534), .B(n7040), .Z(n7038) );
  XOR U10118 ( .A(n7041), .B(n7042), .Z(n7040) );
  XOR U10119 ( .A(DB[2648]), .B(DB[2641]), .Z(n7042) );
  AND U10120 ( .A(n538), .B(n7043), .Z(n7041) );
  XOR U10121 ( .A(n7044), .B(n7045), .Z(n7043) );
  XOR U10122 ( .A(DB[2641]), .B(DB[2634]), .Z(n7045) );
  AND U10123 ( .A(n542), .B(n7046), .Z(n7044) );
  XOR U10124 ( .A(n7047), .B(n7048), .Z(n7046) );
  XOR U10125 ( .A(DB[2634]), .B(DB[2627]), .Z(n7048) );
  AND U10126 ( .A(n546), .B(n7049), .Z(n7047) );
  XOR U10127 ( .A(n7050), .B(n7051), .Z(n7049) );
  XOR U10128 ( .A(DB[2627]), .B(DB[2620]), .Z(n7051) );
  AND U10129 ( .A(n550), .B(n7052), .Z(n7050) );
  XOR U10130 ( .A(n7053), .B(n7054), .Z(n7052) );
  XOR U10131 ( .A(DB[2620]), .B(DB[2613]), .Z(n7054) );
  AND U10132 ( .A(n554), .B(n7055), .Z(n7053) );
  XOR U10133 ( .A(n7056), .B(n7057), .Z(n7055) );
  XOR U10134 ( .A(DB[2613]), .B(DB[2606]), .Z(n7057) );
  AND U10135 ( .A(n558), .B(n7058), .Z(n7056) );
  XOR U10136 ( .A(n7059), .B(n7060), .Z(n7058) );
  XOR U10137 ( .A(DB[2606]), .B(DB[2599]), .Z(n7060) );
  AND U10138 ( .A(n562), .B(n7061), .Z(n7059) );
  XOR U10139 ( .A(n7062), .B(n7063), .Z(n7061) );
  XOR U10140 ( .A(DB[2599]), .B(DB[2592]), .Z(n7063) );
  AND U10141 ( .A(n566), .B(n7064), .Z(n7062) );
  XOR U10142 ( .A(n7065), .B(n7066), .Z(n7064) );
  XOR U10143 ( .A(DB[2592]), .B(DB[2585]), .Z(n7066) );
  AND U10144 ( .A(n570), .B(n7067), .Z(n7065) );
  XOR U10145 ( .A(n7068), .B(n7069), .Z(n7067) );
  XOR U10146 ( .A(DB[2585]), .B(DB[2578]), .Z(n7069) );
  AND U10147 ( .A(n574), .B(n7070), .Z(n7068) );
  XOR U10148 ( .A(n7071), .B(n7072), .Z(n7070) );
  XOR U10149 ( .A(DB[2578]), .B(DB[2571]), .Z(n7072) );
  AND U10150 ( .A(n578), .B(n7073), .Z(n7071) );
  XOR U10151 ( .A(n7074), .B(n7075), .Z(n7073) );
  XOR U10152 ( .A(DB[2571]), .B(DB[2564]), .Z(n7075) );
  AND U10153 ( .A(n582), .B(n7076), .Z(n7074) );
  XOR U10154 ( .A(n7077), .B(n7078), .Z(n7076) );
  XOR U10155 ( .A(DB[2564]), .B(DB[2557]), .Z(n7078) );
  AND U10156 ( .A(n586), .B(n7079), .Z(n7077) );
  XOR U10157 ( .A(n7080), .B(n7081), .Z(n7079) );
  XOR U10158 ( .A(DB[2557]), .B(DB[2550]), .Z(n7081) );
  AND U10159 ( .A(n590), .B(n7082), .Z(n7080) );
  XOR U10160 ( .A(n7083), .B(n7084), .Z(n7082) );
  XOR U10161 ( .A(DB[2550]), .B(DB[2543]), .Z(n7084) );
  AND U10162 ( .A(n594), .B(n7085), .Z(n7083) );
  XOR U10163 ( .A(n7086), .B(n7087), .Z(n7085) );
  XOR U10164 ( .A(DB[2543]), .B(DB[2536]), .Z(n7087) );
  AND U10165 ( .A(n598), .B(n7088), .Z(n7086) );
  XOR U10166 ( .A(n7089), .B(n7090), .Z(n7088) );
  XOR U10167 ( .A(DB[2536]), .B(DB[2529]), .Z(n7090) );
  AND U10168 ( .A(n602), .B(n7091), .Z(n7089) );
  XOR U10169 ( .A(n7092), .B(n7093), .Z(n7091) );
  XOR U10170 ( .A(DB[2529]), .B(DB[2522]), .Z(n7093) );
  AND U10171 ( .A(n606), .B(n7094), .Z(n7092) );
  XOR U10172 ( .A(n7095), .B(n7096), .Z(n7094) );
  XOR U10173 ( .A(DB[2522]), .B(DB[2515]), .Z(n7096) );
  AND U10174 ( .A(n610), .B(n7097), .Z(n7095) );
  XOR U10175 ( .A(n7098), .B(n7099), .Z(n7097) );
  XOR U10176 ( .A(DB[2515]), .B(DB[2508]), .Z(n7099) );
  AND U10177 ( .A(n614), .B(n7100), .Z(n7098) );
  XOR U10178 ( .A(n7101), .B(n7102), .Z(n7100) );
  XOR U10179 ( .A(DB[2508]), .B(DB[2501]), .Z(n7102) );
  AND U10180 ( .A(n618), .B(n7103), .Z(n7101) );
  XOR U10181 ( .A(n7104), .B(n7105), .Z(n7103) );
  XOR U10182 ( .A(DB[2501]), .B(DB[2494]), .Z(n7105) );
  AND U10183 ( .A(n622), .B(n7106), .Z(n7104) );
  XOR U10184 ( .A(n7107), .B(n7108), .Z(n7106) );
  XOR U10185 ( .A(DB[2494]), .B(DB[2487]), .Z(n7108) );
  AND U10186 ( .A(n626), .B(n7109), .Z(n7107) );
  XOR U10187 ( .A(n7110), .B(n7111), .Z(n7109) );
  XOR U10188 ( .A(DB[2487]), .B(DB[2480]), .Z(n7111) );
  AND U10189 ( .A(n630), .B(n7112), .Z(n7110) );
  XOR U10190 ( .A(n7113), .B(n7114), .Z(n7112) );
  XOR U10191 ( .A(DB[2480]), .B(DB[2473]), .Z(n7114) );
  AND U10192 ( .A(n634), .B(n7115), .Z(n7113) );
  XOR U10193 ( .A(n7116), .B(n7117), .Z(n7115) );
  XOR U10194 ( .A(DB[2473]), .B(DB[2466]), .Z(n7117) );
  AND U10195 ( .A(n638), .B(n7118), .Z(n7116) );
  XOR U10196 ( .A(n7119), .B(n7120), .Z(n7118) );
  XOR U10197 ( .A(DB[2466]), .B(DB[2459]), .Z(n7120) );
  AND U10198 ( .A(n642), .B(n7121), .Z(n7119) );
  XOR U10199 ( .A(n7122), .B(n7123), .Z(n7121) );
  XOR U10200 ( .A(DB[2459]), .B(DB[2452]), .Z(n7123) );
  AND U10201 ( .A(n646), .B(n7124), .Z(n7122) );
  XOR U10202 ( .A(n7125), .B(n7126), .Z(n7124) );
  XOR U10203 ( .A(DB[2452]), .B(DB[2445]), .Z(n7126) );
  AND U10204 ( .A(n650), .B(n7127), .Z(n7125) );
  XOR U10205 ( .A(n7128), .B(n7129), .Z(n7127) );
  XOR U10206 ( .A(DB[2445]), .B(DB[2438]), .Z(n7129) );
  AND U10207 ( .A(n654), .B(n7130), .Z(n7128) );
  XOR U10208 ( .A(n7131), .B(n7132), .Z(n7130) );
  XOR U10209 ( .A(DB[2438]), .B(DB[2431]), .Z(n7132) );
  AND U10210 ( .A(n658), .B(n7133), .Z(n7131) );
  XOR U10211 ( .A(n7134), .B(n7135), .Z(n7133) );
  XOR U10212 ( .A(DB[2431]), .B(DB[2424]), .Z(n7135) );
  AND U10213 ( .A(n662), .B(n7136), .Z(n7134) );
  XOR U10214 ( .A(n7137), .B(n7138), .Z(n7136) );
  XOR U10215 ( .A(DB[2424]), .B(DB[2417]), .Z(n7138) );
  AND U10216 ( .A(n666), .B(n7139), .Z(n7137) );
  XOR U10217 ( .A(n7140), .B(n7141), .Z(n7139) );
  XOR U10218 ( .A(DB[2417]), .B(DB[2410]), .Z(n7141) );
  AND U10219 ( .A(n670), .B(n7142), .Z(n7140) );
  XOR U10220 ( .A(n7143), .B(n7144), .Z(n7142) );
  XOR U10221 ( .A(DB[2410]), .B(DB[2403]), .Z(n7144) );
  AND U10222 ( .A(n674), .B(n7145), .Z(n7143) );
  XOR U10223 ( .A(n7146), .B(n7147), .Z(n7145) );
  XOR U10224 ( .A(DB[2403]), .B(DB[2396]), .Z(n7147) );
  AND U10225 ( .A(n678), .B(n7148), .Z(n7146) );
  XOR U10226 ( .A(n7149), .B(n7150), .Z(n7148) );
  XOR U10227 ( .A(DB[2396]), .B(DB[2389]), .Z(n7150) );
  AND U10228 ( .A(n682), .B(n7151), .Z(n7149) );
  XOR U10229 ( .A(n7152), .B(n7153), .Z(n7151) );
  XOR U10230 ( .A(DB[2389]), .B(DB[2382]), .Z(n7153) );
  AND U10231 ( .A(n686), .B(n7154), .Z(n7152) );
  XOR U10232 ( .A(n7155), .B(n7156), .Z(n7154) );
  XOR U10233 ( .A(DB[2382]), .B(DB[2375]), .Z(n7156) );
  AND U10234 ( .A(n690), .B(n7157), .Z(n7155) );
  XOR U10235 ( .A(n7158), .B(n7159), .Z(n7157) );
  XOR U10236 ( .A(DB[2375]), .B(DB[2368]), .Z(n7159) );
  AND U10237 ( .A(n694), .B(n7160), .Z(n7158) );
  XOR U10238 ( .A(n7161), .B(n7162), .Z(n7160) );
  XOR U10239 ( .A(DB[2368]), .B(DB[2361]), .Z(n7162) );
  AND U10240 ( .A(n698), .B(n7163), .Z(n7161) );
  XOR U10241 ( .A(n7164), .B(n7165), .Z(n7163) );
  XOR U10242 ( .A(DB[2361]), .B(DB[2354]), .Z(n7165) );
  AND U10243 ( .A(n702), .B(n7166), .Z(n7164) );
  XOR U10244 ( .A(n7167), .B(n7168), .Z(n7166) );
  XOR U10245 ( .A(DB[2354]), .B(DB[2347]), .Z(n7168) );
  AND U10246 ( .A(n706), .B(n7169), .Z(n7167) );
  XOR U10247 ( .A(n7170), .B(n7171), .Z(n7169) );
  XOR U10248 ( .A(DB[2347]), .B(DB[2340]), .Z(n7171) );
  AND U10249 ( .A(n710), .B(n7172), .Z(n7170) );
  XOR U10250 ( .A(n7173), .B(n7174), .Z(n7172) );
  XOR U10251 ( .A(DB[2340]), .B(DB[2333]), .Z(n7174) );
  AND U10252 ( .A(n714), .B(n7175), .Z(n7173) );
  XOR U10253 ( .A(n7176), .B(n7177), .Z(n7175) );
  XOR U10254 ( .A(DB[2333]), .B(DB[2326]), .Z(n7177) );
  AND U10255 ( .A(n718), .B(n7178), .Z(n7176) );
  XOR U10256 ( .A(n7179), .B(n7180), .Z(n7178) );
  XOR U10257 ( .A(DB[2326]), .B(DB[2319]), .Z(n7180) );
  AND U10258 ( .A(n722), .B(n7181), .Z(n7179) );
  XOR U10259 ( .A(n7182), .B(n7183), .Z(n7181) );
  XOR U10260 ( .A(DB[2319]), .B(DB[2312]), .Z(n7183) );
  AND U10261 ( .A(n726), .B(n7184), .Z(n7182) );
  XOR U10262 ( .A(n7185), .B(n7186), .Z(n7184) );
  XOR U10263 ( .A(DB[2312]), .B(DB[2305]), .Z(n7186) );
  AND U10264 ( .A(n730), .B(n7187), .Z(n7185) );
  XOR U10265 ( .A(n7188), .B(n7189), .Z(n7187) );
  XOR U10266 ( .A(DB[2305]), .B(DB[2298]), .Z(n7189) );
  AND U10267 ( .A(n734), .B(n7190), .Z(n7188) );
  XOR U10268 ( .A(n7191), .B(n7192), .Z(n7190) );
  XOR U10269 ( .A(DB[2298]), .B(DB[2291]), .Z(n7192) );
  AND U10270 ( .A(n738), .B(n7193), .Z(n7191) );
  XOR U10271 ( .A(n7194), .B(n7195), .Z(n7193) );
  XOR U10272 ( .A(DB[2291]), .B(DB[2284]), .Z(n7195) );
  AND U10273 ( .A(n742), .B(n7196), .Z(n7194) );
  XOR U10274 ( .A(n7197), .B(n7198), .Z(n7196) );
  XOR U10275 ( .A(DB[2284]), .B(DB[2277]), .Z(n7198) );
  AND U10276 ( .A(n746), .B(n7199), .Z(n7197) );
  XOR U10277 ( .A(n7200), .B(n7201), .Z(n7199) );
  XOR U10278 ( .A(DB[2277]), .B(DB[2270]), .Z(n7201) );
  AND U10279 ( .A(n750), .B(n7202), .Z(n7200) );
  XOR U10280 ( .A(n7203), .B(n7204), .Z(n7202) );
  XOR U10281 ( .A(DB[2270]), .B(DB[2263]), .Z(n7204) );
  AND U10282 ( .A(n754), .B(n7205), .Z(n7203) );
  XOR U10283 ( .A(n7206), .B(n7207), .Z(n7205) );
  XOR U10284 ( .A(DB[2263]), .B(DB[2256]), .Z(n7207) );
  AND U10285 ( .A(n758), .B(n7208), .Z(n7206) );
  XOR U10286 ( .A(n7209), .B(n7210), .Z(n7208) );
  XOR U10287 ( .A(DB[2256]), .B(DB[2249]), .Z(n7210) );
  AND U10288 ( .A(n762), .B(n7211), .Z(n7209) );
  XOR U10289 ( .A(n7212), .B(n7213), .Z(n7211) );
  XOR U10290 ( .A(DB[2249]), .B(DB[2242]), .Z(n7213) );
  AND U10291 ( .A(n766), .B(n7214), .Z(n7212) );
  XOR U10292 ( .A(n7215), .B(n7216), .Z(n7214) );
  XOR U10293 ( .A(DB[2242]), .B(DB[2235]), .Z(n7216) );
  AND U10294 ( .A(n770), .B(n7217), .Z(n7215) );
  XOR U10295 ( .A(n7218), .B(n7219), .Z(n7217) );
  XOR U10296 ( .A(DB[2235]), .B(DB[2228]), .Z(n7219) );
  AND U10297 ( .A(n774), .B(n7220), .Z(n7218) );
  XOR U10298 ( .A(n7221), .B(n7222), .Z(n7220) );
  XOR U10299 ( .A(DB[2228]), .B(DB[2221]), .Z(n7222) );
  AND U10300 ( .A(n778), .B(n7223), .Z(n7221) );
  XOR U10301 ( .A(n7224), .B(n7225), .Z(n7223) );
  XOR U10302 ( .A(DB[2221]), .B(DB[2214]), .Z(n7225) );
  AND U10303 ( .A(n782), .B(n7226), .Z(n7224) );
  XOR U10304 ( .A(n7227), .B(n7228), .Z(n7226) );
  XOR U10305 ( .A(DB[2214]), .B(DB[2207]), .Z(n7228) );
  AND U10306 ( .A(n786), .B(n7229), .Z(n7227) );
  XOR U10307 ( .A(n7230), .B(n7231), .Z(n7229) );
  XOR U10308 ( .A(DB[2207]), .B(DB[2200]), .Z(n7231) );
  AND U10309 ( .A(n790), .B(n7232), .Z(n7230) );
  XOR U10310 ( .A(n7233), .B(n7234), .Z(n7232) );
  XOR U10311 ( .A(DB[2200]), .B(DB[2193]), .Z(n7234) );
  AND U10312 ( .A(n794), .B(n7235), .Z(n7233) );
  XOR U10313 ( .A(n7236), .B(n7237), .Z(n7235) );
  XOR U10314 ( .A(DB[2193]), .B(DB[2186]), .Z(n7237) );
  AND U10315 ( .A(n798), .B(n7238), .Z(n7236) );
  XOR U10316 ( .A(n7239), .B(n7240), .Z(n7238) );
  XOR U10317 ( .A(DB[2186]), .B(DB[2179]), .Z(n7240) );
  AND U10318 ( .A(n802), .B(n7241), .Z(n7239) );
  XOR U10319 ( .A(n7242), .B(n7243), .Z(n7241) );
  XOR U10320 ( .A(DB[2179]), .B(DB[2172]), .Z(n7243) );
  AND U10321 ( .A(n806), .B(n7244), .Z(n7242) );
  XOR U10322 ( .A(n7245), .B(n7246), .Z(n7244) );
  XOR U10323 ( .A(DB[2172]), .B(DB[2165]), .Z(n7246) );
  AND U10324 ( .A(n810), .B(n7247), .Z(n7245) );
  XOR U10325 ( .A(n7248), .B(n7249), .Z(n7247) );
  XOR U10326 ( .A(DB[2165]), .B(DB[2158]), .Z(n7249) );
  AND U10327 ( .A(n814), .B(n7250), .Z(n7248) );
  XOR U10328 ( .A(n7251), .B(n7252), .Z(n7250) );
  XOR U10329 ( .A(DB[2158]), .B(DB[2151]), .Z(n7252) );
  AND U10330 ( .A(n818), .B(n7253), .Z(n7251) );
  XOR U10331 ( .A(n7254), .B(n7255), .Z(n7253) );
  XOR U10332 ( .A(DB[2151]), .B(DB[2144]), .Z(n7255) );
  AND U10333 ( .A(n822), .B(n7256), .Z(n7254) );
  XOR U10334 ( .A(n7257), .B(n7258), .Z(n7256) );
  XOR U10335 ( .A(DB[2144]), .B(DB[2137]), .Z(n7258) );
  AND U10336 ( .A(n826), .B(n7259), .Z(n7257) );
  XOR U10337 ( .A(n7260), .B(n7261), .Z(n7259) );
  XOR U10338 ( .A(DB[2137]), .B(DB[2130]), .Z(n7261) );
  AND U10339 ( .A(n830), .B(n7262), .Z(n7260) );
  XOR U10340 ( .A(n7263), .B(n7264), .Z(n7262) );
  XOR U10341 ( .A(DB[2130]), .B(DB[2123]), .Z(n7264) );
  AND U10342 ( .A(n834), .B(n7265), .Z(n7263) );
  XOR U10343 ( .A(n7266), .B(n7267), .Z(n7265) );
  XOR U10344 ( .A(DB[2123]), .B(DB[2116]), .Z(n7267) );
  AND U10345 ( .A(n838), .B(n7268), .Z(n7266) );
  XOR U10346 ( .A(n7269), .B(n7270), .Z(n7268) );
  XOR U10347 ( .A(DB[2116]), .B(DB[2109]), .Z(n7270) );
  AND U10348 ( .A(n842), .B(n7271), .Z(n7269) );
  XOR U10349 ( .A(n7272), .B(n7273), .Z(n7271) );
  XOR U10350 ( .A(DB[2109]), .B(DB[2102]), .Z(n7273) );
  AND U10351 ( .A(n846), .B(n7274), .Z(n7272) );
  XOR U10352 ( .A(n7275), .B(n7276), .Z(n7274) );
  XOR U10353 ( .A(DB[2102]), .B(DB[2095]), .Z(n7276) );
  AND U10354 ( .A(n850), .B(n7277), .Z(n7275) );
  XOR U10355 ( .A(n7278), .B(n7279), .Z(n7277) );
  XOR U10356 ( .A(DB[2095]), .B(DB[2088]), .Z(n7279) );
  AND U10357 ( .A(n854), .B(n7280), .Z(n7278) );
  XOR U10358 ( .A(n7281), .B(n7282), .Z(n7280) );
  XOR U10359 ( .A(DB[2088]), .B(DB[2081]), .Z(n7282) );
  AND U10360 ( .A(n858), .B(n7283), .Z(n7281) );
  XOR U10361 ( .A(n7284), .B(n7285), .Z(n7283) );
  XOR U10362 ( .A(DB[2081]), .B(DB[2074]), .Z(n7285) );
  AND U10363 ( .A(n862), .B(n7286), .Z(n7284) );
  XOR U10364 ( .A(n7287), .B(n7288), .Z(n7286) );
  XOR U10365 ( .A(DB[2074]), .B(DB[2067]), .Z(n7288) );
  AND U10366 ( .A(n866), .B(n7289), .Z(n7287) );
  XOR U10367 ( .A(n7290), .B(n7291), .Z(n7289) );
  XOR U10368 ( .A(DB[2067]), .B(DB[2060]), .Z(n7291) );
  AND U10369 ( .A(n870), .B(n7292), .Z(n7290) );
  XOR U10370 ( .A(n7293), .B(n7294), .Z(n7292) );
  XOR U10371 ( .A(DB[2060]), .B(DB[2053]), .Z(n7294) );
  AND U10372 ( .A(n874), .B(n7295), .Z(n7293) );
  XOR U10373 ( .A(n7296), .B(n7297), .Z(n7295) );
  XOR U10374 ( .A(DB[2053]), .B(DB[2046]), .Z(n7297) );
  AND U10375 ( .A(n878), .B(n7298), .Z(n7296) );
  XOR U10376 ( .A(n7299), .B(n7300), .Z(n7298) );
  XOR U10377 ( .A(DB[2046]), .B(DB[2039]), .Z(n7300) );
  AND U10378 ( .A(n882), .B(n7301), .Z(n7299) );
  XOR U10379 ( .A(n7302), .B(n7303), .Z(n7301) );
  XOR U10380 ( .A(DB[2039]), .B(DB[2032]), .Z(n7303) );
  AND U10381 ( .A(n886), .B(n7304), .Z(n7302) );
  XOR U10382 ( .A(n7305), .B(n7306), .Z(n7304) );
  XOR U10383 ( .A(DB[2032]), .B(DB[2025]), .Z(n7306) );
  AND U10384 ( .A(n890), .B(n7307), .Z(n7305) );
  XOR U10385 ( .A(n7308), .B(n7309), .Z(n7307) );
  XOR U10386 ( .A(DB[2025]), .B(DB[2018]), .Z(n7309) );
  AND U10387 ( .A(n894), .B(n7310), .Z(n7308) );
  XOR U10388 ( .A(n7311), .B(n7312), .Z(n7310) );
  XOR U10389 ( .A(DB[2018]), .B(DB[2011]), .Z(n7312) );
  AND U10390 ( .A(n898), .B(n7313), .Z(n7311) );
  XOR U10391 ( .A(n7314), .B(n7315), .Z(n7313) );
  XOR U10392 ( .A(DB[2011]), .B(DB[2004]), .Z(n7315) );
  AND U10393 ( .A(n902), .B(n7316), .Z(n7314) );
  XOR U10394 ( .A(n7317), .B(n7318), .Z(n7316) );
  XOR U10395 ( .A(DB[2004]), .B(DB[1997]), .Z(n7318) );
  AND U10396 ( .A(n906), .B(n7319), .Z(n7317) );
  XOR U10397 ( .A(n7320), .B(n7321), .Z(n7319) );
  XOR U10398 ( .A(DB[1997]), .B(DB[1990]), .Z(n7321) );
  AND U10399 ( .A(n910), .B(n7322), .Z(n7320) );
  XOR U10400 ( .A(n7323), .B(n7324), .Z(n7322) );
  XOR U10401 ( .A(DB[1990]), .B(DB[1983]), .Z(n7324) );
  AND U10402 ( .A(n914), .B(n7325), .Z(n7323) );
  XOR U10403 ( .A(n7326), .B(n7327), .Z(n7325) );
  XOR U10404 ( .A(DB[1983]), .B(DB[1976]), .Z(n7327) );
  AND U10405 ( .A(n918), .B(n7328), .Z(n7326) );
  XOR U10406 ( .A(n7329), .B(n7330), .Z(n7328) );
  XOR U10407 ( .A(DB[1976]), .B(DB[1969]), .Z(n7330) );
  AND U10408 ( .A(n922), .B(n7331), .Z(n7329) );
  XOR U10409 ( .A(n7332), .B(n7333), .Z(n7331) );
  XOR U10410 ( .A(DB[1969]), .B(DB[1962]), .Z(n7333) );
  AND U10411 ( .A(n926), .B(n7334), .Z(n7332) );
  XOR U10412 ( .A(n7335), .B(n7336), .Z(n7334) );
  XOR U10413 ( .A(DB[1962]), .B(DB[1955]), .Z(n7336) );
  AND U10414 ( .A(n930), .B(n7337), .Z(n7335) );
  XOR U10415 ( .A(n7338), .B(n7339), .Z(n7337) );
  XOR U10416 ( .A(DB[1955]), .B(DB[1948]), .Z(n7339) );
  AND U10417 ( .A(n934), .B(n7340), .Z(n7338) );
  XOR U10418 ( .A(n7341), .B(n7342), .Z(n7340) );
  XOR U10419 ( .A(DB[1948]), .B(DB[1941]), .Z(n7342) );
  AND U10420 ( .A(n938), .B(n7343), .Z(n7341) );
  XOR U10421 ( .A(n7344), .B(n7345), .Z(n7343) );
  XOR U10422 ( .A(DB[1941]), .B(DB[1934]), .Z(n7345) );
  AND U10423 ( .A(n942), .B(n7346), .Z(n7344) );
  XOR U10424 ( .A(n7347), .B(n7348), .Z(n7346) );
  XOR U10425 ( .A(DB[1934]), .B(DB[1927]), .Z(n7348) );
  AND U10426 ( .A(n946), .B(n7349), .Z(n7347) );
  XOR U10427 ( .A(n7350), .B(n7351), .Z(n7349) );
  XOR U10428 ( .A(DB[1927]), .B(DB[1920]), .Z(n7351) );
  AND U10429 ( .A(n950), .B(n7352), .Z(n7350) );
  XOR U10430 ( .A(n7353), .B(n7354), .Z(n7352) );
  XOR U10431 ( .A(DB[1920]), .B(DB[1913]), .Z(n7354) );
  AND U10432 ( .A(n954), .B(n7355), .Z(n7353) );
  XOR U10433 ( .A(n7356), .B(n7357), .Z(n7355) );
  XOR U10434 ( .A(DB[1913]), .B(DB[1906]), .Z(n7357) );
  AND U10435 ( .A(n958), .B(n7358), .Z(n7356) );
  XOR U10436 ( .A(n7359), .B(n7360), .Z(n7358) );
  XOR U10437 ( .A(DB[1906]), .B(DB[1899]), .Z(n7360) );
  AND U10438 ( .A(n962), .B(n7361), .Z(n7359) );
  XOR U10439 ( .A(n7362), .B(n7363), .Z(n7361) );
  XOR U10440 ( .A(DB[1899]), .B(DB[1892]), .Z(n7363) );
  AND U10441 ( .A(n966), .B(n7364), .Z(n7362) );
  XOR U10442 ( .A(n7365), .B(n7366), .Z(n7364) );
  XOR U10443 ( .A(DB[1892]), .B(DB[1885]), .Z(n7366) );
  AND U10444 ( .A(n970), .B(n7367), .Z(n7365) );
  XOR U10445 ( .A(n7368), .B(n7369), .Z(n7367) );
  XOR U10446 ( .A(DB[1885]), .B(DB[1878]), .Z(n7369) );
  AND U10447 ( .A(n974), .B(n7370), .Z(n7368) );
  XOR U10448 ( .A(n7371), .B(n7372), .Z(n7370) );
  XOR U10449 ( .A(DB[1878]), .B(DB[1871]), .Z(n7372) );
  AND U10450 ( .A(n978), .B(n7373), .Z(n7371) );
  XOR U10451 ( .A(n7374), .B(n7375), .Z(n7373) );
  XOR U10452 ( .A(DB[1871]), .B(DB[1864]), .Z(n7375) );
  AND U10453 ( .A(n982), .B(n7376), .Z(n7374) );
  XOR U10454 ( .A(n7377), .B(n7378), .Z(n7376) );
  XOR U10455 ( .A(DB[1864]), .B(DB[1857]), .Z(n7378) );
  AND U10456 ( .A(n986), .B(n7379), .Z(n7377) );
  XOR U10457 ( .A(n7380), .B(n7381), .Z(n7379) );
  XOR U10458 ( .A(DB[1857]), .B(DB[1850]), .Z(n7381) );
  AND U10459 ( .A(n990), .B(n7382), .Z(n7380) );
  XOR U10460 ( .A(n7383), .B(n7384), .Z(n7382) );
  XOR U10461 ( .A(DB[1850]), .B(DB[1843]), .Z(n7384) );
  AND U10462 ( .A(n994), .B(n7385), .Z(n7383) );
  XOR U10463 ( .A(n7386), .B(n7387), .Z(n7385) );
  XOR U10464 ( .A(DB[1843]), .B(DB[1836]), .Z(n7387) );
  AND U10465 ( .A(n998), .B(n7388), .Z(n7386) );
  XOR U10466 ( .A(n7389), .B(n7390), .Z(n7388) );
  XOR U10467 ( .A(DB[1836]), .B(DB[1829]), .Z(n7390) );
  AND U10468 ( .A(n1002), .B(n7391), .Z(n7389) );
  XOR U10469 ( .A(n7392), .B(n7393), .Z(n7391) );
  XOR U10470 ( .A(DB[1829]), .B(DB[1822]), .Z(n7393) );
  AND U10471 ( .A(n1006), .B(n7394), .Z(n7392) );
  XOR U10472 ( .A(n7395), .B(n7396), .Z(n7394) );
  XOR U10473 ( .A(DB[1822]), .B(DB[1815]), .Z(n7396) );
  AND U10474 ( .A(n1010), .B(n7397), .Z(n7395) );
  XOR U10475 ( .A(n7398), .B(n7399), .Z(n7397) );
  XOR U10476 ( .A(DB[1815]), .B(DB[1808]), .Z(n7399) );
  AND U10477 ( .A(n1014), .B(n7400), .Z(n7398) );
  XOR U10478 ( .A(n7401), .B(n7402), .Z(n7400) );
  XOR U10479 ( .A(DB[1808]), .B(DB[1801]), .Z(n7402) );
  AND U10480 ( .A(n1018), .B(n7403), .Z(n7401) );
  XOR U10481 ( .A(n7404), .B(n7405), .Z(n7403) );
  XOR U10482 ( .A(DB[1801]), .B(DB[1794]), .Z(n7405) );
  AND U10483 ( .A(n1022), .B(n7406), .Z(n7404) );
  XOR U10484 ( .A(n7407), .B(n7408), .Z(n7406) );
  XOR U10485 ( .A(DB[1794]), .B(DB[1787]), .Z(n7408) );
  AND U10486 ( .A(n1026), .B(n7409), .Z(n7407) );
  XOR U10487 ( .A(n7410), .B(n7411), .Z(n7409) );
  XOR U10488 ( .A(DB[1787]), .B(DB[1780]), .Z(n7411) );
  AND U10489 ( .A(n1030), .B(n7412), .Z(n7410) );
  XOR U10490 ( .A(n7413), .B(n7414), .Z(n7412) );
  XOR U10491 ( .A(DB[1780]), .B(DB[1773]), .Z(n7414) );
  AND U10492 ( .A(n1034), .B(n7415), .Z(n7413) );
  XOR U10493 ( .A(n7416), .B(n7417), .Z(n7415) );
  XOR U10494 ( .A(DB[1773]), .B(DB[1766]), .Z(n7417) );
  AND U10495 ( .A(n1038), .B(n7418), .Z(n7416) );
  XOR U10496 ( .A(n7419), .B(n7420), .Z(n7418) );
  XOR U10497 ( .A(DB[1766]), .B(DB[1759]), .Z(n7420) );
  AND U10498 ( .A(n1042), .B(n7421), .Z(n7419) );
  XOR U10499 ( .A(n7422), .B(n7423), .Z(n7421) );
  XOR U10500 ( .A(DB[1759]), .B(DB[1752]), .Z(n7423) );
  AND U10501 ( .A(n1046), .B(n7424), .Z(n7422) );
  XOR U10502 ( .A(n7425), .B(n7426), .Z(n7424) );
  XOR U10503 ( .A(DB[1752]), .B(DB[1745]), .Z(n7426) );
  AND U10504 ( .A(n1050), .B(n7427), .Z(n7425) );
  XOR U10505 ( .A(n7428), .B(n7429), .Z(n7427) );
  XOR U10506 ( .A(DB[1745]), .B(DB[1738]), .Z(n7429) );
  AND U10507 ( .A(n1054), .B(n7430), .Z(n7428) );
  XOR U10508 ( .A(n7431), .B(n7432), .Z(n7430) );
  XOR U10509 ( .A(DB[1738]), .B(DB[1731]), .Z(n7432) );
  AND U10510 ( .A(n1058), .B(n7433), .Z(n7431) );
  XOR U10511 ( .A(n7434), .B(n7435), .Z(n7433) );
  XOR U10512 ( .A(DB[1731]), .B(DB[1724]), .Z(n7435) );
  AND U10513 ( .A(n1062), .B(n7436), .Z(n7434) );
  XOR U10514 ( .A(n7437), .B(n7438), .Z(n7436) );
  XOR U10515 ( .A(DB[1724]), .B(DB[1717]), .Z(n7438) );
  AND U10516 ( .A(n1066), .B(n7439), .Z(n7437) );
  XOR U10517 ( .A(n7440), .B(n7441), .Z(n7439) );
  XOR U10518 ( .A(DB[1717]), .B(DB[1710]), .Z(n7441) );
  AND U10519 ( .A(n1070), .B(n7442), .Z(n7440) );
  XOR U10520 ( .A(n7443), .B(n7444), .Z(n7442) );
  XOR U10521 ( .A(DB[1710]), .B(DB[1703]), .Z(n7444) );
  AND U10522 ( .A(n1074), .B(n7445), .Z(n7443) );
  XOR U10523 ( .A(n7446), .B(n7447), .Z(n7445) );
  XOR U10524 ( .A(DB[1703]), .B(DB[1696]), .Z(n7447) );
  AND U10525 ( .A(n1078), .B(n7448), .Z(n7446) );
  XOR U10526 ( .A(n7449), .B(n7450), .Z(n7448) );
  XOR U10527 ( .A(DB[1696]), .B(DB[1689]), .Z(n7450) );
  AND U10528 ( .A(n1082), .B(n7451), .Z(n7449) );
  XOR U10529 ( .A(n7452), .B(n7453), .Z(n7451) );
  XOR U10530 ( .A(DB[1689]), .B(DB[1682]), .Z(n7453) );
  AND U10531 ( .A(n1086), .B(n7454), .Z(n7452) );
  XOR U10532 ( .A(n7455), .B(n7456), .Z(n7454) );
  XOR U10533 ( .A(DB[1682]), .B(DB[1675]), .Z(n7456) );
  AND U10534 ( .A(n1090), .B(n7457), .Z(n7455) );
  XOR U10535 ( .A(n7458), .B(n7459), .Z(n7457) );
  XOR U10536 ( .A(DB[1675]), .B(DB[1668]), .Z(n7459) );
  AND U10537 ( .A(n1094), .B(n7460), .Z(n7458) );
  XOR U10538 ( .A(n7461), .B(n7462), .Z(n7460) );
  XOR U10539 ( .A(DB[1668]), .B(DB[1661]), .Z(n7462) );
  AND U10540 ( .A(n1098), .B(n7463), .Z(n7461) );
  XOR U10541 ( .A(n7464), .B(n7465), .Z(n7463) );
  XOR U10542 ( .A(DB[1661]), .B(DB[1654]), .Z(n7465) );
  AND U10543 ( .A(n1102), .B(n7466), .Z(n7464) );
  XOR U10544 ( .A(n7467), .B(n7468), .Z(n7466) );
  XOR U10545 ( .A(DB[1654]), .B(DB[1647]), .Z(n7468) );
  AND U10546 ( .A(n1106), .B(n7469), .Z(n7467) );
  XOR U10547 ( .A(n7470), .B(n7471), .Z(n7469) );
  XOR U10548 ( .A(DB[1647]), .B(DB[1640]), .Z(n7471) );
  AND U10549 ( .A(n1110), .B(n7472), .Z(n7470) );
  XOR U10550 ( .A(n7473), .B(n7474), .Z(n7472) );
  XOR U10551 ( .A(DB[1640]), .B(DB[1633]), .Z(n7474) );
  AND U10552 ( .A(n1114), .B(n7475), .Z(n7473) );
  XOR U10553 ( .A(n7476), .B(n7477), .Z(n7475) );
  XOR U10554 ( .A(DB[1633]), .B(DB[1626]), .Z(n7477) );
  AND U10555 ( .A(n1118), .B(n7478), .Z(n7476) );
  XOR U10556 ( .A(n7479), .B(n7480), .Z(n7478) );
  XOR U10557 ( .A(DB[1626]), .B(DB[1619]), .Z(n7480) );
  AND U10558 ( .A(n1122), .B(n7481), .Z(n7479) );
  XOR U10559 ( .A(n7482), .B(n7483), .Z(n7481) );
  XOR U10560 ( .A(DB[1619]), .B(DB[1612]), .Z(n7483) );
  AND U10561 ( .A(n1126), .B(n7484), .Z(n7482) );
  XOR U10562 ( .A(n7485), .B(n7486), .Z(n7484) );
  XOR U10563 ( .A(DB[1612]), .B(DB[1605]), .Z(n7486) );
  AND U10564 ( .A(n1130), .B(n7487), .Z(n7485) );
  XOR U10565 ( .A(n7488), .B(n7489), .Z(n7487) );
  XOR U10566 ( .A(DB[1605]), .B(DB[1598]), .Z(n7489) );
  AND U10567 ( .A(n1134), .B(n7490), .Z(n7488) );
  XOR U10568 ( .A(n7491), .B(n7492), .Z(n7490) );
  XOR U10569 ( .A(DB[1598]), .B(DB[1591]), .Z(n7492) );
  AND U10570 ( .A(n1138), .B(n7493), .Z(n7491) );
  XOR U10571 ( .A(n7494), .B(n7495), .Z(n7493) );
  XOR U10572 ( .A(DB[1591]), .B(DB[1584]), .Z(n7495) );
  AND U10573 ( .A(n1142), .B(n7496), .Z(n7494) );
  XOR U10574 ( .A(n7497), .B(n7498), .Z(n7496) );
  XOR U10575 ( .A(DB[1584]), .B(DB[1577]), .Z(n7498) );
  AND U10576 ( .A(n1146), .B(n7499), .Z(n7497) );
  XOR U10577 ( .A(n7500), .B(n7501), .Z(n7499) );
  XOR U10578 ( .A(DB[1577]), .B(DB[1570]), .Z(n7501) );
  AND U10579 ( .A(n1150), .B(n7502), .Z(n7500) );
  XOR U10580 ( .A(n7503), .B(n7504), .Z(n7502) );
  XOR U10581 ( .A(DB[1570]), .B(DB[1563]), .Z(n7504) );
  AND U10582 ( .A(n1154), .B(n7505), .Z(n7503) );
  XOR U10583 ( .A(n7506), .B(n7507), .Z(n7505) );
  XOR U10584 ( .A(DB[1563]), .B(DB[1556]), .Z(n7507) );
  AND U10585 ( .A(n1158), .B(n7508), .Z(n7506) );
  XOR U10586 ( .A(n7509), .B(n7510), .Z(n7508) );
  XOR U10587 ( .A(DB[1556]), .B(DB[1549]), .Z(n7510) );
  AND U10588 ( .A(n1162), .B(n7511), .Z(n7509) );
  XOR U10589 ( .A(n7512), .B(n7513), .Z(n7511) );
  XOR U10590 ( .A(DB[1549]), .B(DB[1542]), .Z(n7513) );
  AND U10591 ( .A(n1166), .B(n7514), .Z(n7512) );
  XOR U10592 ( .A(n7515), .B(n7516), .Z(n7514) );
  XOR U10593 ( .A(DB[1542]), .B(DB[1535]), .Z(n7516) );
  AND U10594 ( .A(n1170), .B(n7517), .Z(n7515) );
  XOR U10595 ( .A(n7518), .B(n7519), .Z(n7517) );
  XOR U10596 ( .A(DB[1535]), .B(DB[1528]), .Z(n7519) );
  AND U10597 ( .A(n1174), .B(n7520), .Z(n7518) );
  XOR U10598 ( .A(n7521), .B(n7522), .Z(n7520) );
  XOR U10599 ( .A(DB[1528]), .B(DB[1521]), .Z(n7522) );
  AND U10600 ( .A(n1178), .B(n7523), .Z(n7521) );
  XOR U10601 ( .A(n7524), .B(n7525), .Z(n7523) );
  XOR U10602 ( .A(DB[1521]), .B(DB[1514]), .Z(n7525) );
  AND U10603 ( .A(n1182), .B(n7526), .Z(n7524) );
  XOR U10604 ( .A(n7527), .B(n7528), .Z(n7526) );
  XOR U10605 ( .A(DB[1514]), .B(DB[1507]), .Z(n7528) );
  AND U10606 ( .A(n1186), .B(n7529), .Z(n7527) );
  XOR U10607 ( .A(n7530), .B(n7531), .Z(n7529) );
  XOR U10608 ( .A(DB[1507]), .B(DB[1500]), .Z(n7531) );
  AND U10609 ( .A(n1190), .B(n7532), .Z(n7530) );
  XOR U10610 ( .A(n7533), .B(n7534), .Z(n7532) );
  XOR U10611 ( .A(DB[1500]), .B(DB[1493]), .Z(n7534) );
  AND U10612 ( .A(n1194), .B(n7535), .Z(n7533) );
  XOR U10613 ( .A(n7536), .B(n7537), .Z(n7535) );
  XOR U10614 ( .A(DB[1493]), .B(DB[1486]), .Z(n7537) );
  AND U10615 ( .A(n1198), .B(n7538), .Z(n7536) );
  XOR U10616 ( .A(n7539), .B(n7540), .Z(n7538) );
  XOR U10617 ( .A(DB[1486]), .B(DB[1479]), .Z(n7540) );
  AND U10618 ( .A(n1202), .B(n7541), .Z(n7539) );
  XOR U10619 ( .A(n7542), .B(n7543), .Z(n7541) );
  XOR U10620 ( .A(DB[1479]), .B(DB[1472]), .Z(n7543) );
  AND U10621 ( .A(n1206), .B(n7544), .Z(n7542) );
  XOR U10622 ( .A(n7545), .B(n7546), .Z(n7544) );
  XOR U10623 ( .A(DB[1472]), .B(DB[1465]), .Z(n7546) );
  AND U10624 ( .A(n1210), .B(n7547), .Z(n7545) );
  XOR U10625 ( .A(n7548), .B(n7549), .Z(n7547) );
  XOR U10626 ( .A(DB[1465]), .B(DB[1458]), .Z(n7549) );
  AND U10627 ( .A(n1214), .B(n7550), .Z(n7548) );
  XOR U10628 ( .A(n7551), .B(n7552), .Z(n7550) );
  XOR U10629 ( .A(DB[1458]), .B(DB[1451]), .Z(n7552) );
  AND U10630 ( .A(n1218), .B(n7553), .Z(n7551) );
  XOR U10631 ( .A(n7554), .B(n7555), .Z(n7553) );
  XOR U10632 ( .A(DB[1451]), .B(DB[1444]), .Z(n7555) );
  AND U10633 ( .A(n1222), .B(n7556), .Z(n7554) );
  XOR U10634 ( .A(n7557), .B(n7558), .Z(n7556) );
  XOR U10635 ( .A(DB[1444]), .B(DB[1437]), .Z(n7558) );
  AND U10636 ( .A(n1226), .B(n7559), .Z(n7557) );
  XOR U10637 ( .A(n7560), .B(n7561), .Z(n7559) );
  XOR U10638 ( .A(DB[1437]), .B(DB[1430]), .Z(n7561) );
  AND U10639 ( .A(n1230), .B(n7562), .Z(n7560) );
  XOR U10640 ( .A(n7563), .B(n7564), .Z(n7562) );
  XOR U10641 ( .A(DB[1430]), .B(DB[1423]), .Z(n7564) );
  AND U10642 ( .A(n1234), .B(n7565), .Z(n7563) );
  XOR U10643 ( .A(n7566), .B(n7567), .Z(n7565) );
  XOR U10644 ( .A(DB[1423]), .B(DB[1416]), .Z(n7567) );
  AND U10645 ( .A(n1238), .B(n7568), .Z(n7566) );
  XOR U10646 ( .A(n7569), .B(n7570), .Z(n7568) );
  XOR U10647 ( .A(DB[1416]), .B(DB[1409]), .Z(n7570) );
  AND U10648 ( .A(n1242), .B(n7571), .Z(n7569) );
  XOR U10649 ( .A(n7572), .B(n7573), .Z(n7571) );
  XOR U10650 ( .A(DB[1409]), .B(DB[1402]), .Z(n7573) );
  AND U10651 ( .A(n1246), .B(n7574), .Z(n7572) );
  XOR U10652 ( .A(n7575), .B(n7576), .Z(n7574) );
  XOR U10653 ( .A(DB[1402]), .B(DB[1395]), .Z(n7576) );
  AND U10654 ( .A(n1250), .B(n7577), .Z(n7575) );
  XOR U10655 ( .A(n7578), .B(n7579), .Z(n7577) );
  XOR U10656 ( .A(DB[1395]), .B(DB[1388]), .Z(n7579) );
  AND U10657 ( .A(n1254), .B(n7580), .Z(n7578) );
  XOR U10658 ( .A(n7581), .B(n7582), .Z(n7580) );
  XOR U10659 ( .A(DB[1388]), .B(DB[1381]), .Z(n7582) );
  AND U10660 ( .A(n1258), .B(n7583), .Z(n7581) );
  XOR U10661 ( .A(n7584), .B(n7585), .Z(n7583) );
  XOR U10662 ( .A(DB[1381]), .B(DB[1374]), .Z(n7585) );
  AND U10663 ( .A(n1262), .B(n7586), .Z(n7584) );
  XOR U10664 ( .A(n7587), .B(n7588), .Z(n7586) );
  XOR U10665 ( .A(DB[1374]), .B(DB[1367]), .Z(n7588) );
  AND U10666 ( .A(n1266), .B(n7589), .Z(n7587) );
  XOR U10667 ( .A(n7590), .B(n7591), .Z(n7589) );
  XOR U10668 ( .A(DB[1367]), .B(DB[1360]), .Z(n7591) );
  AND U10669 ( .A(n1270), .B(n7592), .Z(n7590) );
  XOR U10670 ( .A(n7593), .B(n7594), .Z(n7592) );
  XOR U10671 ( .A(DB[1360]), .B(DB[1353]), .Z(n7594) );
  AND U10672 ( .A(n1274), .B(n7595), .Z(n7593) );
  XOR U10673 ( .A(n7596), .B(n7597), .Z(n7595) );
  XOR U10674 ( .A(DB[1353]), .B(DB[1346]), .Z(n7597) );
  AND U10675 ( .A(n1278), .B(n7598), .Z(n7596) );
  XOR U10676 ( .A(n7599), .B(n7600), .Z(n7598) );
  XOR U10677 ( .A(DB[1346]), .B(DB[1339]), .Z(n7600) );
  AND U10678 ( .A(n1282), .B(n7601), .Z(n7599) );
  XOR U10679 ( .A(n7602), .B(n7603), .Z(n7601) );
  XOR U10680 ( .A(DB[1339]), .B(DB[1332]), .Z(n7603) );
  AND U10681 ( .A(n1286), .B(n7604), .Z(n7602) );
  XOR U10682 ( .A(n7605), .B(n7606), .Z(n7604) );
  XOR U10683 ( .A(DB[1332]), .B(DB[1325]), .Z(n7606) );
  AND U10684 ( .A(n1290), .B(n7607), .Z(n7605) );
  XOR U10685 ( .A(n7608), .B(n7609), .Z(n7607) );
  XOR U10686 ( .A(DB[1325]), .B(DB[1318]), .Z(n7609) );
  AND U10687 ( .A(n1294), .B(n7610), .Z(n7608) );
  XOR U10688 ( .A(n7611), .B(n7612), .Z(n7610) );
  XOR U10689 ( .A(DB[1318]), .B(DB[1311]), .Z(n7612) );
  AND U10690 ( .A(n1298), .B(n7613), .Z(n7611) );
  XOR U10691 ( .A(n7614), .B(n7615), .Z(n7613) );
  XOR U10692 ( .A(DB[1311]), .B(DB[1304]), .Z(n7615) );
  AND U10693 ( .A(n1302), .B(n7616), .Z(n7614) );
  XOR U10694 ( .A(n7617), .B(n7618), .Z(n7616) );
  XOR U10695 ( .A(DB[1304]), .B(DB[1297]), .Z(n7618) );
  AND U10696 ( .A(n1306), .B(n7619), .Z(n7617) );
  XOR U10697 ( .A(n7620), .B(n7621), .Z(n7619) );
  XOR U10698 ( .A(DB[1297]), .B(DB[1290]), .Z(n7621) );
  AND U10699 ( .A(n1310), .B(n7622), .Z(n7620) );
  XOR U10700 ( .A(n7623), .B(n7624), .Z(n7622) );
  XOR U10701 ( .A(DB[1290]), .B(DB[1283]), .Z(n7624) );
  AND U10702 ( .A(n1314), .B(n7625), .Z(n7623) );
  XOR U10703 ( .A(n7626), .B(n7627), .Z(n7625) );
  XOR U10704 ( .A(DB[1283]), .B(DB[1276]), .Z(n7627) );
  AND U10705 ( .A(n1318), .B(n7628), .Z(n7626) );
  XOR U10706 ( .A(n7629), .B(n7630), .Z(n7628) );
  XOR U10707 ( .A(DB[1276]), .B(DB[1269]), .Z(n7630) );
  AND U10708 ( .A(n1322), .B(n7631), .Z(n7629) );
  XOR U10709 ( .A(n7632), .B(n7633), .Z(n7631) );
  XOR U10710 ( .A(DB[1269]), .B(DB[1262]), .Z(n7633) );
  AND U10711 ( .A(n1326), .B(n7634), .Z(n7632) );
  XOR U10712 ( .A(n7635), .B(n7636), .Z(n7634) );
  XOR U10713 ( .A(DB[1262]), .B(DB[1255]), .Z(n7636) );
  AND U10714 ( .A(n1330), .B(n7637), .Z(n7635) );
  XOR U10715 ( .A(n7638), .B(n7639), .Z(n7637) );
  XOR U10716 ( .A(DB[1255]), .B(DB[1248]), .Z(n7639) );
  AND U10717 ( .A(n1334), .B(n7640), .Z(n7638) );
  XOR U10718 ( .A(n7641), .B(n7642), .Z(n7640) );
  XOR U10719 ( .A(DB[1248]), .B(DB[1241]), .Z(n7642) );
  AND U10720 ( .A(n1338), .B(n7643), .Z(n7641) );
  XOR U10721 ( .A(n7644), .B(n7645), .Z(n7643) );
  XOR U10722 ( .A(DB[1241]), .B(DB[1234]), .Z(n7645) );
  AND U10723 ( .A(n1342), .B(n7646), .Z(n7644) );
  XOR U10724 ( .A(n7647), .B(n7648), .Z(n7646) );
  XOR U10725 ( .A(DB[1234]), .B(DB[1227]), .Z(n7648) );
  AND U10726 ( .A(n1346), .B(n7649), .Z(n7647) );
  XOR U10727 ( .A(n7650), .B(n7651), .Z(n7649) );
  XOR U10728 ( .A(DB[1227]), .B(DB[1220]), .Z(n7651) );
  AND U10729 ( .A(n1350), .B(n7652), .Z(n7650) );
  XOR U10730 ( .A(n7653), .B(n7654), .Z(n7652) );
  XOR U10731 ( .A(DB[1220]), .B(DB[1213]), .Z(n7654) );
  AND U10732 ( .A(n1354), .B(n7655), .Z(n7653) );
  XOR U10733 ( .A(n7656), .B(n7657), .Z(n7655) );
  XOR U10734 ( .A(DB[1213]), .B(DB[1206]), .Z(n7657) );
  AND U10735 ( .A(n1358), .B(n7658), .Z(n7656) );
  XOR U10736 ( .A(n7659), .B(n7660), .Z(n7658) );
  XOR U10737 ( .A(DB[1206]), .B(DB[1199]), .Z(n7660) );
  AND U10738 ( .A(n1362), .B(n7661), .Z(n7659) );
  XOR U10739 ( .A(n7662), .B(n7663), .Z(n7661) );
  XOR U10740 ( .A(DB[1199]), .B(DB[1192]), .Z(n7663) );
  AND U10741 ( .A(n1366), .B(n7664), .Z(n7662) );
  XOR U10742 ( .A(n7665), .B(n7666), .Z(n7664) );
  XOR U10743 ( .A(DB[1192]), .B(DB[1185]), .Z(n7666) );
  AND U10744 ( .A(n1370), .B(n7667), .Z(n7665) );
  XOR U10745 ( .A(n7668), .B(n7669), .Z(n7667) );
  XOR U10746 ( .A(DB[1185]), .B(DB[1178]), .Z(n7669) );
  AND U10747 ( .A(n1374), .B(n7670), .Z(n7668) );
  XOR U10748 ( .A(n7671), .B(n7672), .Z(n7670) );
  XOR U10749 ( .A(DB[1178]), .B(DB[1171]), .Z(n7672) );
  AND U10750 ( .A(n1378), .B(n7673), .Z(n7671) );
  XOR U10751 ( .A(n7674), .B(n7675), .Z(n7673) );
  XOR U10752 ( .A(DB[1171]), .B(DB[1164]), .Z(n7675) );
  AND U10753 ( .A(n1382), .B(n7676), .Z(n7674) );
  XOR U10754 ( .A(n7677), .B(n7678), .Z(n7676) );
  XOR U10755 ( .A(DB[1164]), .B(DB[1157]), .Z(n7678) );
  AND U10756 ( .A(n1386), .B(n7679), .Z(n7677) );
  XOR U10757 ( .A(n7680), .B(n7681), .Z(n7679) );
  XOR U10758 ( .A(DB[1157]), .B(DB[1150]), .Z(n7681) );
  AND U10759 ( .A(n1390), .B(n7682), .Z(n7680) );
  XOR U10760 ( .A(n7683), .B(n7684), .Z(n7682) );
  XOR U10761 ( .A(DB[1150]), .B(DB[1143]), .Z(n7684) );
  AND U10762 ( .A(n1394), .B(n7685), .Z(n7683) );
  XOR U10763 ( .A(n7686), .B(n7687), .Z(n7685) );
  XOR U10764 ( .A(DB[1143]), .B(DB[1136]), .Z(n7687) );
  AND U10765 ( .A(n1398), .B(n7688), .Z(n7686) );
  XOR U10766 ( .A(n7689), .B(n7690), .Z(n7688) );
  XOR U10767 ( .A(DB[1136]), .B(DB[1129]), .Z(n7690) );
  AND U10768 ( .A(n1402), .B(n7691), .Z(n7689) );
  XOR U10769 ( .A(n7692), .B(n7693), .Z(n7691) );
  XOR U10770 ( .A(DB[1129]), .B(DB[1122]), .Z(n7693) );
  AND U10771 ( .A(n1406), .B(n7694), .Z(n7692) );
  XOR U10772 ( .A(n7695), .B(n7696), .Z(n7694) );
  XOR U10773 ( .A(DB[1122]), .B(DB[1115]), .Z(n7696) );
  AND U10774 ( .A(n1410), .B(n7697), .Z(n7695) );
  XOR U10775 ( .A(n7698), .B(n7699), .Z(n7697) );
  XOR U10776 ( .A(DB[1115]), .B(DB[1108]), .Z(n7699) );
  AND U10777 ( .A(n1414), .B(n7700), .Z(n7698) );
  XOR U10778 ( .A(n7701), .B(n7702), .Z(n7700) );
  XOR U10779 ( .A(DB[1108]), .B(DB[1101]), .Z(n7702) );
  AND U10780 ( .A(n1418), .B(n7703), .Z(n7701) );
  XOR U10781 ( .A(n7704), .B(n7705), .Z(n7703) );
  XOR U10782 ( .A(DB[1101]), .B(DB[1094]), .Z(n7705) );
  AND U10783 ( .A(n1422), .B(n7706), .Z(n7704) );
  XOR U10784 ( .A(n7707), .B(n7708), .Z(n7706) );
  XOR U10785 ( .A(DB[1094]), .B(DB[1087]), .Z(n7708) );
  AND U10786 ( .A(n1426), .B(n7709), .Z(n7707) );
  XOR U10787 ( .A(n7710), .B(n7711), .Z(n7709) );
  XOR U10788 ( .A(DB[1087]), .B(DB[1080]), .Z(n7711) );
  AND U10789 ( .A(n1430), .B(n7712), .Z(n7710) );
  XOR U10790 ( .A(n7713), .B(n7714), .Z(n7712) );
  XOR U10791 ( .A(DB[1080]), .B(DB[1073]), .Z(n7714) );
  AND U10792 ( .A(n1434), .B(n7715), .Z(n7713) );
  XOR U10793 ( .A(n7716), .B(n7717), .Z(n7715) );
  XOR U10794 ( .A(DB[1073]), .B(DB[1066]), .Z(n7717) );
  AND U10795 ( .A(n1438), .B(n7718), .Z(n7716) );
  XOR U10796 ( .A(n7719), .B(n7720), .Z(n7718) );
  XOR U10797 ( .A(DB[1066]), .B(DB[1059]), .Z(n7720) );
  AND U10798 ( .A(n1442), .B(n7721), .Z(n7719) );
  XOR U10799 ( .A(n7722), .B(n7723), .Z(n7721) );
  XOR U10800 ( .A(DB[1059]), .B(DB[1052]), .Z(n7723) );
  AND U10801 ( .A(n1446), .B(n7724), .Z(n7722) );
  XOR U10802 ( .A(n7725), .B(n7726), .Z(n7724) );
  XOR U10803 ( .A(DB[1052]), .B(DB[1045]), .Z(n7726) );
  AND U10804 ( .A(n1450), .B(n7727), .Z(n7725) );
  XOR U10805 ( .A(n7728), .B(n7729), .Z(n7727) );
  XOR U10806 ( .A(DB[1045]), .B(DB[1038]), .Z(n7729) );
  AND U10807 ( .A(n1454), .B(n7730), .Z(n7728) );
  XOR U10808 ( .A(n7731), .B(n7732), .Z(n7730) );
  XOR U10809 ( .A(DB[1038]), .B(DB[1031]), .Z(n7732) );
  AND U10810 ( .A(n1458), .B(n7733), .Z(n7731) );
  XOR U10811 ( .A(n7734), .B(n7735), .Z(n7733) );
  XOR U10812 ( .A(DB[1031]), .B(DB[1024]), .Z(n7735) );
  AND U10813 ( .A(n1462), .B(n7736), .Z(n7734) );
  XOR U10814 ( .A(n7737), .B(n7738), .Z(n7736) );
  XOR U10815 ( .A(DB[1024]), .B(DB[1017]), .Z(n7738) );
  AND U10816 ( .A(n1466), .B(n7739), .Z(n7737) );
  XOR U10817 ( .A(n7740), .B(n7741), .Z(n7739) );
  XOR U10818 ( .A(DB[1017]), .B(DB[1010]), .Z(n7741) );
  AND U10819 ( .A(n1470), .B(n7742), .Z(n7740) );
  XOR U10820 ( .A(n7743), .B(n7744), .Z(n7742) );
  XOR U10821 ( .A(DB[1010]), .B(DB[1003]), .Z(n7744) );
  AND U10822 ( .A(n1474), .B(n7745), .Z(n7743) );
  XOR U10823 ( .A(n7746), .B(n7747), .Z(n7745) );
  XOR U10824 ( .A(DB[996]), .B(DB[1003]), .Z(n7747) );
  AND U10825 ( .A(n1478), .B(n7748), .Z(n7746) );
  XOR U10826 ( .A(n7749), .B(n7750), .Z(n7748) );
  XOR U10827 ( .A(DB[996]), .B(DB[989]), .Z(n7750) );
  AND U10828 ( .A(n1482), .B(n7751), .Z(n7749) );
  XOR U10829 ( .A(n7752), .B(n7753), .Z(n7751) );
  XOR U10830 ( .A(DB[989]), .B(DB[982]), .Z(n7753) );
  AND U10831 ( .A(n1486), .B(n7754), .Z(n7752) );
  XOR U10832 ( .A(n7755), .B(n7756), .Z(n7754) );
  XOR U10833 ( .A(DB[982]), .B(DB[975]), .Z(n7756) );
  AND U10834 ( .A(n1490), .B(n7757), .Z(n7755) );
  XOR U10835 ( .A(n7758), .B(n7759), .Z(n7757) );
  XOR U10836 ( .A(DB[975]), .B(DB[968]), .Z(n7759) );
  AND U10837 ( .A(n1494), .B(n7760), .Z(n7758) );
  XOR U10838 ( .A(n7761), .B(n7762), .Z(n7760) );
  XOR U10839 ( .A(DB[968]), .B(DB[961]), .Z(n7762) );
  AND U10840 ( .A(n1498), .B(n7763), .Z(n7761) );
  XOR U10841 ( .A(n7764), .B(n7765), .Z(n7763) );
  XOR U10842 ( .A(DB[961]), .B(DB[954]), .Z(n7765) );
  AND U10843 ( .A(n1502), .B(n7766), .Z(n7764) );
  XOR U10844 ( .A(n7767), .B(n7768), .Z(n7766) );
  XOR U10845 ( .A(DB[954]), .B(DB[947]), .Z(n7768) );
  AND U10846 ( .A(n1506), .B(n7769), .Z(n7767) );
  XOR U10847 ( .A(n7770), .B(n7771), .Z(n7769) );
  XOR U10848 ( .A(DB[947]), .B(DB[940]), .Z(n7771) );
  AND U10849 ( .A(n1510), .B(n7772), .Z(n7770) );
  XOR U10850 ( .A(n7773), .B(n7774), .Z(n7772) );
  XOR U10851 ( .A(DB[940]), .B(DB[933]), .Z(n7774) );
  AND U10852 ( .A(n1514), .B(n7775), .Z(n7773) );
  XOR U10853 ( .A(n7776), .B(n7777), .Z(n7775) );
  XOR U10854 ( .A(DB[933]), .B(DB[926]), .Z(n7777) );
  AND U10855 ( .A(n1518), .B(n7778), .Z(n7776) );
  XOR U10856 ( .A(n7779), .B(n7780), .Z(n7778) );
  XOR U10857 ( .A(DB[926]), .B(DB[919]), .Z(n7780) );
  AND U10858 ( .A(n1522), .B(n7781), .Z(n7779) );
  XOR U10859 ( .A(n7782), .B(n7783), .Z(n7781) );
  XOR U10860 ( .A(DB[919]), .B(DB[912]), .Z(n7783) );
  AND U10861 ( .A(n1526), .B(n7784), .Z(n7782) );
  XOR U10862 ( .A(n7785), .B(n7786), .Z(n7784) );
  XOR U10863 ( .A(DB[912]), .B(DB[905]), .Z(n7786) );
  AND U10864 ( .A(n1530), .B(n7787), .Z(n7785) );
  XOR U10865 ( .A(n7788), .B(n7789), .Z(n7787) );
  XOR U10866 ( .A(DB[905]), .B(DB[898]), .Z(n7789) );
  AND U10867 ( .A(n1534), .B(n7790), .Z(n7788) );
  XOR U10868 ( .A(n7791), .B(n7792), .Z(n7790) );
  XOR U10869 ( .A(DB[898]), .B(DB[891]), .Z(n7792) );
  AND U10870 ( .A(n1538), .B(n7793), .Z(n7791) );
  XOR U10871 ( .A(n7794), .B(n7795), .Z(n7793) );
  XOR U10872 ( .A(DB[891]), .B(DB[884]), .Z(n7795) );
  AND U10873 ( .A(n1542), .B(n7796), .Z(n7794) );
  XOR U10874 ( .A(n7797), .B(n7798), .Z(n7796) );
  XOR U10875 ( .A(DB[884]), .B(DB[877]), .Z(n7798) );
  AND U10876 ( .A(n1546), .B(n7799), .Z(n7797) );
  XOR U10877 ( .A(n7800), .B(n7801), .Z(n7799) );
  XOR U10878 ( .A(DB[877]), .B(DB[870]), .Z(n7801) );
  AND U10879 ( .A(n1550), .B(n7802), .Z(n7800) );
  XOR U10880 ( .A(n7803), .B(n7804), .Z(n7802) );
  XOR U10881 ( .A(DB[870]), .B(DB[863]), .Z(n7804) );
  AND U10882 ( .A(n1554), .B(n7805), .Z(n7803) );
  XOR U10883 ( .A(n7806), .B(n7807), .Z(n7805) );
  XOR U10884 ( .A(DB[863]), .B(DB[856]), .Z(n7807) );
  AND U10885 ( .A(n1558), .B(n7808), .Z(n7806) );
  XOR U10886 ( .A(n7809), .B(n7810), .Z(n7808) );
  XOR U10887 ( .A(DB[856]), .B(DB[849]), .Z(n7810) );
  AND U10888 ( .A(n1562), .B(n7811), .Z(n7809) );
  XOR U10889 ( .A(n7812), .B(n7813), .Z(n7811) );
  XOR U10890 ( .A(DB[849]), .B(DB[842]), .Z(n7813) );
  AND U10891 ( .A(n1566), .B(n7814), .Z(n7812) );
  XOR U10892 ( .A(n7815), .B(n7816), .Z(n7814) );
  XOR U10893 ( .A(DB[842]), .B(DB[835]), .Z(n7816) );
  AND U10894 ( .A(n1570), .B(n7817), .Z(n7815) );
  XOR U10895 ( .A(n7818), .B(n7819), .Z(n7817) );
  XOR U10896 ( .A(DB[835]), .B(DB[828]), .Z(n7819) );
  AND U10897 ( .A(n1574), .B(n7820), .Z(n7818) );
  XOR U10898 ( .A(n7821), .B(n7822), .Z(n7820) );
  XOR U10899 ( .A(DB[828]), .B(DB[821]), .Z(n7822) );
  AND U10900 ( .A(n1578), .B(n7823), .Z(n7821) );
  XOR U10901 ( .A(n7824), .B(n7825), .Z(n7823) );
  XOR U10902 ( .A(DB[821]), .B(DB[814]), .Z(n7825) );
  AND U10903 ( .A(n1582), .B(n7826), .Z(n7824) );
  XOR U10904 ( .A(n7827), .B(n7828), .Z(n7826) );
  XOR U10905 ( .A(DB[814]), .B(DB[807]), .Z(n7828) );
  AND U10906 ( .A(n1586), .B(n7829), .Z(n7827) );
  XOR U10907 ( .A(n7830), .B(n7831), .Z(n7829) );
  XOR U10908 ( .A(DB[807]), .B(DB[800]), .Z(n7831) );
  AND U10909 ( .A(n1590), .B(n7832), .Z(n7830) );
  XOR U10910 ( .A(n7833), .B(n7834), .Z(n7832) );
  XOR U10911 ( .A(DB[800]), .B(DB[793]), .Z(n7834) );
  AND U10912 ( .A(n1594), .B(n7835), .Z(n7833) );
  XOR U10913 ( .A(n7836), .B(n7837), .Z(n7835) );
  XOR U10914 ( .A(DB[793]), .B(DB[786]), .Z(n7837) );
  AND U10915 ( .A(n1598), .B(n7838), .Z(n7836) );
  XOR U10916 ( .A(n7839), .B(n7840), .Z(n7838) );
  XOR U10917 ( .A(DB[786]), .B(DB[779]), .Z(n7840) );
  AND U10918 ( .A(n1602), .B(n7841), .Z(n7839) );
  XOR U10919 ( .A(n7842), .B(n7843), .Z(n7841) );
  XOR U10920 ( .A(DB[779]), .B(DB[772]), .Z(n7843) );
  AND U10921 ( .A(n1606), .B(n7844), .Z(n7842) );
  XOR U10922 ( .A(n7845), .B(n7846), .Z(n7844) );
  XOR U10923 ( .A(DB[772]), .B(DB[765]), .Z(n7846) );
  AND U10924 ( .A(n1610), .B(n7847), .Z(n7845) );
  XOR U10925 ( .A(n7848), .B(n7849), .Z(n7847) );
  XOR U10926 ( .A(DB[765]), .B(DB[758]), .Z(n7849) );
  AND U10927 ( .A(n1614), .B(n7850), .Z(n7848) );
  XOR U10928 ( .A(n7851), .B(n7852), .Z(n7850) );
  XOR U10929 ( .A(DB[758]), .B(DB[751]), .Z(n7852) );
  AND U10930 ( .A(n1618), .B(n7853), .Z(n7851) );
  XOR U10931 ( .A(n7854), .B(n7855), .Z(n7853) );
  XOR U10932 ( .A(DB[751]), .B(DB[744]), .Z(n7855) );
  AND U10933 ( .A(n1622), .B(n7856), .Z(n7854) );
  XOR U10934 ( .A(n7857), .B(n7858), .Z(n7856) );
  XOR U10935 ( .A(DB[744]), .B(DB[737]), .Z(n7858) );
  AND U10936 ( .A(n1626), .B(n7859), .Z(n7857) );
  XOR U10937 ( .A(n7860), .B(n7861), .Z(n7859) );
  XOR U10938 ( .A(DB[737]), .B(DB[730]), .Z(n7861) );
  AND U10939 ( .A(n1630), .B(n7862), .Z(n7860) );
  XOR U10940 ( .A(n7863), .B(n7864), .Z(n7862) );
  XOR U10941 ( .A(DB[730]), .B(DB[723]), .Z(n7864) );
  AND U10942 ( .A(n1634), .B(n7865), .Z(n7863) );
  XOR U10943 ( .A(n7866), .B(n7867), .Z(n7865) );
  XOR U10944 ( .A(DB[723]), .B(DB[716]), .Z(n7867) );
  AND U10945 ( .A(n1638), .B(n7868), .Z(n7866) );
  XOR U10946 ( .A(n7869), .B(n7870), .Z(n7868) );
  XOR U10947 ( .A(DB[716]), .B(DB[709]), .Z(n7870) );
  AND U10948 ( .A(n1642), .B(n7871), .Z(n7869) );
  XOR U10949 ( .A(n7872), .B(n7873), .Z(n7871) );
  XOR U10950 ( .A(DB[709]), .B(DB[702]), .Z(n7873) );
  AND U10951 ( .A(n1646), .B(n7874), .Z(n7872) );
  XOR U10952 ( .A(n7875), .B(n7876), .Z(n7874) );
  XOR U10953 ( .A(DB[702]), .B(DB[695]), .Z(n7876) );
  AND U10954 ( .A(n1650), .B(n7877), .Z(n7875) );
  XOR U10955 ( .A(n7878), .B(n7879), .Z(n7877) );
  XOR U10956 ( .A(DB[695]), .B(DB[688]), .Z(n7879) );
  AND U10957 ( .A(n1654), .B(n7880), .Z(n7878) );
  XOR U10958 ( .A(n7881), .B(n7882), .Z(n7880) );
  XOR U10959 ( .A(DB[688]), .B(DB[681]), .Z(n7882) );
  AND U10960 ( .A(n1658), .B(n7883), .Z(n7881) );
  XOR U10961 ( .A(n7884), .B(n7885), .Z(n7883) );
  XOR U10962 ( .A(DB[681]), .B(DB[674]), .Z(n7885) );
  AND U10963 ( .A(n1662), .B(n7886), .Z(n7884) );
  XOR U10964 ( .A(n7887), .B(n7888), .Z(n7886) );
  XOR U10965 ( .A(DB[674]), .B(DB[667]), .Z(n7888) );
  AND U10966 ( .A(n1666), .B(n7889), .Z(n7887) );
  XOR U10967 ( .A(n7890), .B(n7891), .Z(n7889) );
  XOR U10968 ( .A(DB[667]), .B(DB[660]), .Z(n7891) );
  AND U10969 ( .A(n1670), .B(n7892), .Z(n7890) );
  XOR U10970 ( .A(n7893), .B(n7894), .Z(n7892) );
  XOR U10971 ( .A(DB[660]), .B(DB[653]), .Z(n7894) );
  AND U10972 ( .A(n1674), .B(n7895), .Z(n7893) );
  XOR U10973 ( .A(n7896), .B(n7897), .Z(n7895) );
  XOR U10974 ( .A(DB[653]), .B(DB[646]), .Z(n7897) );
  AND U10975 ( .A(n1678), .B(n7898), .Z(n7896) );
  XOR U10976 ( .A(n7899), .B(n7900), .Z(n7898) );
  XOR U10977 ( .A(DB[646]), .B(DB[639]), .Z(n7900) );
  AND U10978 ( .A(n1682), .B(n7901), .Z(n7899) );
  XOR U10979 ( .A(n7902), .B(n7903), .Z(n7901) );
  XOR U10980 ( .A(DB[639]), .B(DB[632]), .Z(n7903) );
  AND U10981 ( .A(n1686), .B(n7904), .Z(n7902) );
  XOR U10982 ( .A(n7905), .B(n7906), .Z(n7904) );
  XOR U10983 ( .A(DB[632]), .B(DB[625]), .Z(n7906) );
  AND U10984 ( .A(n1690), .B(n7907), .Z(n7905) );
  XOR U10985 ( .A(n7908), .B(n7909), .Z(n7907) );
  XOR U10986 ( .A(DB[625]), .B(DB[618]), .Z(n7909) );
  AND U10987 ( .A(n1694), .B(n7910), .Z(n7908) );
  XOR U10988 ( .A(n7911), .B(n7912), .Z(n7910) );
  XOR U10989 ( .A(DB[618]), .B(DB[611]), .Z(n7912) );
  AND U10990 ( .A(n1698), .B(n7913), .Z(n7911) );
  XOR U10991 ( .A(n7914), .B(n7915), .Z(n7913) );
  XOR U10992 ( .A(DB[611]), .B(DB[604]), .Z(n7915) );
  AND U10993 ( .A(n1702), .B(n7916), .Z(n7914) );
  XOR U10994 ( .A(n7917), .B(n7918), .Z(n7916) );
  XOR U10995 ( .A(DB[604]), .B(DB[597]), .Z(n7918) );
  AND U10996 ( .A(n1706), .B(n7919), .Z(n7917) );
  XOR U10997 ( .A(n7920), .B(n7921), .Z(n7919) );
  XOR U10998 ( .A(DB[597]), .B(DB[590]), .Z(n7921) );
  AND U10999 ( .A(n1710), .B(n7922), .Z(n7920) );
  XOR U11000 ( .A(n7923), .B(n7924), .Z(n7922) );
  XOR U11001 ( .A(DB[590]), .B(DB[583]), .Z(n7924) );
  AND U11002 ( .A(n1714), .B(n7925), .Z(n7923) );
  XOR U11003 ( .A(n7926), .B(n7927), .Z(n7925) );
  XOR U11004 ( .A(DB[583]), .B(DB[576]), .Z(n7927) );
  AND U11005 ( .A(n1718), .B(n7928), .Z(n7926) );
  XOR U11006 ( .A(n7929), .B(n7930), .Z(n7928) );
  XOR U11007 ( .A(DB[576]), .B(DB[569]), .Z(n7930) );
  AND U11008 ( .A(n1722), .B(n7931), .Z(n7929) );
  XOR U11009 ( .A(n7932), .B(n7933), .Z(n7931) );
  XOR U11010 ( .A(DB[569]), .B(DB[562]), .Z(n7933) );
  AND U11011 ( .A(n1726), .B(n7934), .Z(n7932) );
  XOR U11012 ( .A(n7935), .B(n7936), .Z(n7934) );
  XOR U11013 ( .A(DB[562]), .B(DB[555]), .Z(n7936) );
  AND U11014 ( .A(n1730), .B(n7937), .Z(n7935) );
  XOR U11015 ( .A(n7938), .B(n7939), .Z(n7937) );
  XOR U11016 ( .A(DB[555]), .B(DB[548]), .Z(n7939) );
  AND U11017 ( .A(n1734), .B(n7940), .Z(n7938) );
  XOR U11018 ( .A(n7941), .B(n7942), .Z(n7940) );
  XOR U11019 ( .A(DB[548]), .B(DB[541]), .Z(n7942) );
  AND U11020 ( .A(n1738), .B(n7943), .Z(n7941) );
  XOR U11021 ( .A(n7944), .B(n7945), .Z(n7943) );
  XOR U11022 ( .A(DB[541]), .B(DB[534]), .Z(n7945) );
  AND U11023 ( .A(n1742), .B(n7946), .Z(n7944) );
  XOR U11024 ( .A(n7947), .B(n7948), .Z(n7946) );
  XOR U11025 ( .A(DB[534]), .B(DB[527]), .Z(n7948) );
  AND U11026 ( .A(n1746), .B(n7949), .Z(n7947) );
  XOR U11027 ( .A(n7950), .B(n7951), .Z(n7949) );
  XOR U11028 ( .A(DB[527]), .B(DB[520]), .Z(n7951) );
  AND U11029 ( .A(n1750), .B(n7952), .Z(n7950) );
  XOR U11030 ( .A(n7953), .B(n7954), .Z(n7952) );
  XOR U11031 ( .A(DB[520]), .B(DB[513]), .Z(n7954) );
  AND U11032 ( .A(n1754), .B(n7955), .Z(n7953) );
  XOR U11033 ( .A(n7956), .B(n7957), .Z(n7955) );
  XOR U11034 ( .A(DB[513]), .B(DB[506]), .Z(n7957) );
  AND U11035 ( .A(n1758), .B(n7958), .Z(n7956) );
  XOR U11036 ( .A(n7959), .B(n7960), .Z(n7958) );
  XOR U11037 ( .A(DB[506]), .B(DB[499]), .Z(n7960) );
  AND U11038 ( .A(n1762), .B(n7961), .Z(n7959) );
  XOR U11039 ( .A(n7962), .B(n7963), .Z(n7961) );
  XOR U11040 ( .A(DB[499]), .B(DB[492]), .Z(n7963) );
  AND U11041 ( .A(n1766), .B(n7964), .Z(n7962) );
  XOR U11042 ( .A(n7965), .B(n7966), .Z(n7964) );
  XOR U11043 ( .A(DB[492]), .B(DB[485]), .Z(n7966) );
  AND U11044 ( .A(n1770), .B(n7967), .Z(n7965) );
  XOR U11045 ( .A(n7968), .B(n7969), .Z(n7967) );
  XOR U11046 ( .A(DB[485]), .B(DB[478]), .Z(n7969) );
  AND U11047 ( .A(n1774), .B(n7970), .Z(n7968) );
  XOR U11048 ( .A(n7971), .B(n7972), .Z(n7970) );
  XOR U11049 ( .A(DB[478]), .B(DB[471]), .Z(n7972) );
  AND U11050 ( .A(n1778), .B(n7973), .Z(n7971) );
  XOR U11051 ( .A(n7974), .B(n7975), .Z(n7973) );
  XOR U11052 ( .A(DB[471]), .B(DB[464]), .Z(n7975) );
  AND U11053 ( .A(n1782), .B(n7976), .Z(n7974) );
  XOR U11054 ( .A(n7977), .B(n7978), .Z(n7976) );
  XOR U11055 ( .A(DB[464]), .B(DB[457]), .Z(n7978) );
  AND U11056 ( .A(n1786), .B(n7979), .Z(n7977) );
  XOR U11057 ( .A(n7980), .B(n7981), .Z(n7979) );
  XOR U11058 ( .A(DB[457]), .B(DB[450]), .Z(n7981) );
  AND U11059 ( .A(n1790), .B(n7982), .Z(n7980) );
  XOR U11060 ( .A(n7983), .B(n7984), .Z(n7982) );
  XOR U11061 ( .A(DB[450]), .B(DB[443]), .Z(n7984) );
  AND U11062 ( .A(n1794), .B(n7985), .Z(n7983) );
  XOR U11063 ( .A(n7986), .B(n7987), .Z(n7985) );
  XOR U11064 ( .A(DB[443]), .B(DB[436]), .Z(n7987) );
  AND U11065 ( .A(n1798), .B(n7988), .Z(n7986) );
  XOR U11066 ( .A(n7989), .B(n7990), .Z(n7988) );
  XOR U11067 ( .A(DB[436]), .B(DB[429]), .Z(n7990) );
  AND U11068 ( .A(n1802), .B(n7991), .Z(n7989) );
  XOR U11069 ( .A(n7992), .B(n7993), .Z(n7991) );
  XOR U11070 ( .A(DB[429]), .B(DB[422]), .Z(n7993) );
  AND U11071 ( .A(n1806), .B(n7994), .Z(n7992) );
  XOR U11072 ( .A(n7995), .B(n7996), .Z(n7994) );
  XOR U11073 ( .A(DB[422]), .B(DB[415]), .Z(n7996) );
  AND U11074 ( .A(n1810), .B(n7997), .Z(n7995) );
  XOR U11075 ( .A(n7998), .B(n7999), .Z(n7997) );
  XOR U11076 ( .A(DB[415]), .B(DB[408]), .Z(n7999) );
  AND U11077 ( .A(n1814), .B(n8000), .Z(n7998) );
  XOR U11078 ( .A(n8001), .B(n8002), .Z(n8000) );
  XOR U11079 ( .A(DB[408]), .B(DB[401]), .Z(n8002) );
  AND U11080 ( .A(n1818), .B(n8003), .Z(n8001) );
  XOR U11081 ( .A(n8004), .B(n8005), .Z(n8003) );
  XOR U11082 ( .A(DB[401]), .B(DB[394]), .Z(n8005) );
  AND U11083 ( .A(n1822), .B(n8006), .Z(n8004) );
  XOR U11084 ( .A(n8007), .B(n8008), .Z(n8006) );
  XOR U11085 ( .A(DB[394]), .B(DB[387]), .Z(n8008) );
  AND U11086 ( .A(n1826), .B(n8009), .Z(n8007) );
  XOR U11087 ( .A(n8010), .B(n8011), .Z(n8009) );
  XOR U11088 ( .A(DB[387]), .B(DB[380]), .Z(n8011) );
  AND U11089 ( .A(n1830), .B(n8012), .Z(n8010) );
  XOR U11090 ( .A(n8013), .B(n8014), .Z(n8012) );
  XOR U11091 ( .A(DB[380]), .B(DB[373]), .Z(n8014) );
  AND U11092 ( .A(n1834), .B(n8015), .Z(n8013) );
  XOR U11093 ( .A(n8016), .B(n8017), .Z(n8015) );
  XOR U11094 ( .A(DB[373]), .B(DB[366]), .Z(n8017) );
  AND U11095 ( .A(n1838), .B(n8018), .Z(n8016) );
  XOR U11096 ( .A(n8019), .B(n8020), .Z(n8018) );
  XOR U11097 ( .A(DB[366]), .B(DB[359]), .Z(n8020) );
  AND U11098 ( .A(n1842), .B(n8021), .Z(n8019) );
  XOR U11099 ( .A(n8022), .B(n8023), .Z(n8021) );
  XOR U11100 ( .A(DB[359]), .B(DB[352]), .Z(n8023) );
  AND U11101 ( .A(n1846), .B(n8024), .Z(n8022) );
  XOR U11102 ( .A(n8025), .B(n8026), .Z(n8024) );
  XOR U11103 ( .A(DB[352]), .B(DB[345]), .Z(n8026) );
  AND U11104 ( .A(n1850), .B(n8027), .Z(n8025) );
  XOR U11105 ( .A(n8028), .B(n8029), .Z(n8027) );
  XOR U11106 ( .A(DB[345]), .B(DB[338]), .Z(n8029) );
  AND U11107 ( .A(n1854), .B(n8030), .Z(n8028) );
  XOR U11108 ( .A(n8031), .B(n8032), .Z(n8030) );
  XOR U11109 ( .A(DB[338]), .B(DB[331]), .Z(n8032) );
  AND U11110 ( .A(n1858), .B(n8033), .Z(n8031) );
  XOR U11111 ( .A(n8034), .B(n8035), .Z(n8033) );
  XOR U11112 ( .A(DB[331]), .B(DB[324]), .Z(n8035) );
  AND U11113 ( .A(n1862), .B(n8036), .Z(n8034) );
  XOR U11114 ( .A(n8037), .B(n8038), .Z(n8036) );
  XOR U11115 ( .A(DB[324]), .B(DB[317]), .Z(n8038) );
  AND U11116 ( .A(n1866), .B(n8039), .Z(n8037) );
  XOR U11117 ( .A(n8040), .B(n8041), .Z(n8039) );
  XOR U11118 ( .A(DB[317]), .B(DB[310]), .Z(n8041) );
  AND U11119 ( .A(n1870), .B(n8042), .Z(n8040) );
  XOR U11120 ( .A(n8043), .B(n8044), .Z(n8042) );
  XOR U11121 ( .A(DB[310]), .B(DB[303]), .Z(n8044) );
  AND U11122 ( .A(n1874), .B(n8045), .Z(n8043) );
  XOR U11123 ( .A(n8046), .B(n8047), .Z(n8045) );
  XOR U11124 ( .A(DB[303]), .B(DB[296]), .Z(n8047) );
  AND U11125 ( .A(n1878), .B(n8048), .Z(n8046) );
  XOR U11126 ( .A(n8049), .B(n8050), .Z(n8048) );
  XOR U11127 ( .A(DB[296]), .B(DB[289]), .Z(n8050) );
  AND U11128 ( .A(n1882), .B(n8051), .Z(n8049) );
  XOR U11129 ( .A(n8052), .B(n8053), .Z(n8051) );
  XOR U11130 ( .A(DB[289]), .B(DB[282]), .Z(n8053) );
  AND U11131 ( .A(n1886), .B(n8054), .Z(n8052) );
  XOR U11132 ( .A(n8055), .B(n8056), .Z(n8054) );
  XOR U11133 ( .A(DB[282]), .B(DB[275]), .Z(n8056) );
  AND U11134 ( .A(n1890), .B(n8057), .Z(n8055) );
  XOR U11135 ( .A(n8058), .B(n8059), .Z(n8057) );
  XOR U11136 ( .A(DB[275]), .B(DB[268]), .Z(n8059) );
  AND U11137 ( .A(n1894), .B(n8060), .Z(n8058) );
  XOR U11138 ( .A(n8061), .B(n8062), .Z(n8060) );
  XOR U11139 ( .A(DB[268]), .B(DB[261]), .Z(n8062) );
  AND U11140 ( .A(n1898), .B(n8063), .Z(n8061) );
  XOR U11141 ( .A(n8064), .B(n8065), .Z(n8063) );
  XOR U11142 ( .A(DB[261]), .B(DB[254]), .Z(n8065) );
  AND U11143 ( .A(n1902), .B(n8066), .Z(n8064) );
  XOR U11144 ( .A(n8067), .B(n8068), .Z(n8066) );
  XOR U11145 ( .A(DB[254]), .B(DB[247]), .Z(n8068) );
  AND U11146 ( .A(n1906), .B(n8069), .Z(n8067) );
  XOR U11147 ( .A(n8070), .B(n8071), .Z(n8069) );
  XOR U11148 ( .A(DB[247]), .B(DB[240]), .Z(n8071) );
  AND U11149 ( .A(n1910), .B(n8072), .Z(n8070) );
  XOR U11150 ( .A(n8073), .B(n8074), .Z(n8072) );
  XOR U11151 ( .A(DB[240]), .B(DB[233]), .Z(n8074) );
  AND U11152 ( .A(n1914), .B(n8075), .Z(n8073) );
  XOR U11153 ( .A(n8076), .B(n8077), .Z(n8075) );
  XOR U11154 ( .A(DB[233]), .B(DB[226]), .Z(n8077) );
  AND U11155 ( .A(n1918), .B(n8078), .Z(n8076) );
  XOR U11156 ( .A(n8079), .B(n8080), .Z(n8078) );
  XOR U11157 ( .A(DB[226]), .B(DB[219]), .Z(n8080) );
  AND U11158 ( .A(n1922), .B(n8081), .Z(n8079) );
  XOR U11159 ( .A(n8082), .B(n8083), .Z(n8081) );
  XOR U11160 ( .A(DB[219]), .B(DB[212]), .Z(n8083) );
  AND U11161 ( .A(n1926), .B(n8084), .Z(n8082) );
  XOR U11162 ( .A(n8085), .B(n8086), .Z(n8084) );
  XOR U11163 ( .A(DB[212]), .B(DB[205]), .Z(n8086) );
  AND U11164 ( .A(n1930), .B(n8087), .Z(n8085) );
  XOR U11165 ( .A(n8088), .B(n8089), .Z(n8087) );
  XOR U11166 ( .A(DB[205]), .B(DB[198]), .Z(n8089) );
  AND U11167 ( .A(n1934), .B(n8090), .Z(n8088) );
  XOR U11168 ( .A(n8091), .B(n8092), .Z(n8090) );
  XOR U11169 ( .A(DB[198]), .B(DB[191]), .Z(n8092) );
  AND U11170 ( .A(n1938), .B(n8093), .Z(n8091) );
  XOR U11171 ( .A(n8094), .B(n8095), .Z(n8093) );
  XOR U11172 ( .A(DB[191]), .B(DB[184]), .Z(n8095) );
  AND U11173 ( .A(n1942), .B(n8096), .Z(n8094) );
  XOR U11174 ( .A(n8097), .B(n8098), .Z(n8096) );
  XOR U11175 ( .A(DB[184]), .B(DB[177]), .Z(n8098) );
  AND U11176 ( .A(n1946), .B(n8099), .Z(n8097) );
  XOR U11177 ( .A(n8100), .B(n8101), .Z(n8099) );
  XOR U11178 ( .A(DB[177]), .B(DB[170]), .Z(n8101) );
  AND U11179 ( .A(n1950), .B(n8102), .Z(n8100) );
  XOR U11180 ( .A(n8103), .B(n8104), .Z(n8102) );
  XOR U11181 ( .A(DB[170]), .B(DB[163]), .Z(n8104) );
  AND U11182 ( .A(n1954), .B(n8105), .Z(n8103) );
  XOR U11183 ( .A(n8106), .B(n8107), .Z(n8105) );
  XOR U11184 ( .A(DB[163]), .B(DB[156]), .Z(n8107) );
  AND U11185 ( .A(n1958), .B(n8108), .Z(n8106) );
  XOR U11186 ( .A(n8109), .B(n8110), .Z(n8108) );
  XOR U11187 ( .A(DB[156]), .B(DB[149]), .Z(n8110) );
  AND U11188 ( .A(n1962), .B(n8111), .Z(n8109) );
  XOR U11189 ( .A(n8112), .B(n8113), .Z(n8111) );
  XOR U11190 ( .A(DB[149]), .B(DB[142]), .Z(n8113) );
  AND U11191 ( .A(n1966), .B(n8114), .Z(n8112) );
  XOR U11192 ( .A(n8115), .B(n8116), .Z(n8114) );
  XOR U11193 ( .A(DB[142]), .B(DB[135]), .Z(n8116) );
  AND U11194 ( .A(n1970), .B(n8117), .Z(n8115) );
  XOR U11195 ( .A(n8118), .B(n8119), .Z(n8117) );
  XOR U11196 ( .A(DB[135]), .B(DB[128]), .Z(n8119) );
  AND U11197 ( .A(n1974), .B(n8120), .Z(n8118) );
  XOR U11198 ( .A(n8121), .B(n8122), .Z(n8120) );
  XOR U11199 ( .A(DB[128]), .B(DB[121]), .Z(n8122) );
  AND U11200 ( .A(n1978), .B(n8123), .Z(n8121) );
  XOR U11201 ( .A(n8124), .B(n8125), .Z(n8123) );
  XOR U11202 ( .A(DB[121]), .B(DB[114]), .Z(n8125) );
  AND U11203 ( .A(n1982), .B(n8126), .Z(n8124) );
  XOR U11204 ( .A(n8127), .B(n8128), .Z(n8126) );
  XOR U11205 ( .A(DB[114]), .B(DB[107]), .Z(n8128) );
  AND U11206 ( .A(n1986), .B(n8129), .Z(n8127) );
  XOR U11207 ( .A(n8130), .B(n8131), .Z(n8129) );
  XOR U11208 ( .A(DB[107]), .B(DB[100]), .Z(n8131) );
  AND U11209 ( .A(n1990), .B(n8132), .Z(n8130) );
  XOR U11210 ( .A(n8133), .B(n8134), .Z(n8132) );
  XOR U11211 ( .A(DB[93]), .B(DB[100]), .Z(n8134) );
  AND U11212 ( .A(n1994), .B(n8135), .Z(n8133) );
  XOR U11213 ( .A(n8136), .B(n8137), .Z(n8135) );
  XOR U11214 ( .A(DB[93]), .B(DB[86]), .Z(n8137) );
  AND U11215 ( .A(n1998), .B(n8138), .Z(n8136) );
  XOR U11216 ( .A(n8139), .B(n8140), .Z(n8138) );
  XOR U11217 ( .A(DB[86]), .B(DB[79]), .Z(n8140) );
  AND U11218 ( .A(n2002), .B(n8141), .Z(n8139) );
  XOR U11219 ( .A(n8142), .B(n8143), .Z(n8141) );
  XOR U11220 ( .A(DB[79]), .B(DB[72]), .Z(n8143) );
  AND U11221 ( .A(n2006), .B(n8144), .Z(n8142) );
  XOR U11222 ( .A(n8145), .B(n8146), .Z(n8144) );
  XOR U11223 ( .A(DB[72]), .B(DB[65]), .Z(n8146) );
  AND U11224 ( .A(n2010), .B(n8147), .Z(n8145) );
  XOR U11225 ( .A(n8148), .B(n8149), .Z(n8147) );
  XOR U11226 ( .A(DB[65]), .B(DB[58]), .Z(n8149) );
  AND U11227 ( .A(n2014), .B(n8150), .Z(n8148) );
  XOR U11228 ( .A(n8151), .B(n8152), .Z(n8150) );
  XOR U11229 ( .A(DB[58]), .B(DB[51]), .Z(n8152) );
  AND U11230 ( .A(n2018), .B(n8153), .Z(n8151) );
  XOR U11231 ( .A(n8154), .B(n8155), .Z(n8153) );
  XOR U11232 ( .A(DB[51]), .B(DB[44]), .Z(n8155) );
  AND U11233 ( .A(n2022), .B(n8156), .Z(n8154) );
  XOR U11234 ( .A(n8157), .B(n8158), .Z(n8156) );
  XOR U11235 ( .A(DB[44]), .B(DB[37]), .Z(n8158) );
  AND U11236 ( .A(n2026), .B(n8159), .Z(n8157) );
  XOR U11237 ( .A(n8160), .B(n8161), .Z(n8159) );
  XOR U11238 ( .A(DB[37]), .B(DB[30]), .Z(n8161) );
  AND U11239 ( .A(n2030), .B(n8162), .Z(n8160) );
  XOR U11240 ( .A(n8163), .B(n8164), .Z(n8162) );
  XOR U11241 ( .A(DB[30]), .B(DB[23]), .Z(n8164) );
  AND U11242 ( .A(n2034), .B(n8165), .Z(n8163) );
  XOR U11243 ( .A(n8166), .B(n8167), .Z(n8165) );
  XOR U11244 ( .A(DB[23]), .B(DB[16]), .Z(n8167) );
  AND U11245 ( .A(n2038), .B(n8168), .Z(n8166) );
  XOR U11246 ( .A(n8169), .B(n8170), .Z(n8168) );
  XOR U11247 ( .A(DB[9]), .B(DB[16]), .Z(n8170) );
  AND U11248 ( .A(n2042), .B(n8171), .Z(n8169) );
  XOR U11249 ( .A(DB[9]), .B(DB[2]), .Z(n8171) );
  XOR U11250 ( .A(DB[3578]), .B(n8172), .Z(min_val_out[1]) );
  AND U11251 ( .A(n2), .B(n8173), .Z(n8172) );
  XOR U11252 ( .A(n8174), .B(n8175), .Z(n8173) );
  XOR U11253 ( .A(DB[3578]), .B(DB[3571]), .Z(n8175) );
  AND U11254 ( .A(n6), .B(n8176), .Z(n8174) );
  XOR U11255 ( .A(n8177), .B(n8178), .Z(n8176) );
  XOR U11256 ( .A(DB[3571]), .B(DB[3564]), .Z(n8178) );
  AND U11257 ( .A(n10), .B(n8179), .Z(n8177) );
  XOR U11258 ( .A(n8180), .B(n8181), .Z(n8179) );
  XOR U11259 ( .A(DB[3564]), .B(DB[3557]), .Z(n8181) );
  AND U11260 ( .A(n14), .B(n8182), .Z(n8180) );
  XOR U11261 ( .A(n8183), .B(n8184), .Z(n8182) );
  XOR U11262 ( .A(DB[3557]), .B(DB[3550]), .Z(n8184) );
  AND U11263 ( .A(n18), .B(n8185), .Z(n8183) );
  XOR U11264 ( .A(n8186), .B(n8187), .Z(n8185) );
  XOR U11265 ( .A(DB[3550]), .B(DB[3543]), .Z(n8187) );
  AND U11266 ( .A(n22), .B(n8188), .Z(n8186) );
  XOR U11267 ( .A(n8189), .B(n8190), .Z(n8188) );
  XOR U11268 ( .A(DB[3543]), .B(DB[3536]), .Z(n8190) );
  AND U11269 ( .A(n26), .B(n8191), .Z(n8189) );
  XOR U11270 ( .A(n8192), .B(n8193), .Z(n8191) );
  XOR U11271 ( .A(DB[3536]), .B(DB[3529]), .Z(n8193) );
  AND U11272 ( .A(n30), .B(n8194), .Z(n8192) );
  XOR U11273 ( .A(n8195), .B(n8196), .Z(n8194) );
  XOR U11274 ( .A(DB[3529]), .B(DB[3522]), .Z(n8196) );
  AND U11275 ( .A(n34), .B(n8197), .Z(n8195) );
  XOR U11276 ( .A(n8198), .B(n8199), .Z(n8197) );
  XOR U11277 ( .A(DB[3522]), .B(DB[3515]), .Z(n8199) );
  AND U11278 ( .A(n38), .B(n8200), .Z(n8198) );
  XOR U11279 ( .A(n8201), .B(n8202), .Z(n8200) );
  XOR U11280 ( .A(DB[3515]), .B(DB[3508]), .Z(n8202) );
  AND U11281 ( .A(n42), .B(n8203), .Z(n8201) );
  XOR U11282 ( .A(n8204), .B(n8205), .Z(n8203) );
  XOR U11283 ( .A(DB[3508]), .B(DB[3501]), .Z(n8205) );
  AND U11284 ( .A(n46), .B(n8206), .Z(n8204) );
  XOR U11285 ( .A(n8207), .B(n8208), .Z(n8206) );
  XOR U11286 ( .A(DB[3501]), .B(DB[3494]), .Z(n8208) );
  AND U11287 ( .A(n50), .B(n8209), .Z(n8207) );
  XOR U11288 ( .A(n8210), .B(n8211), .Z(n8209) );
  XOR U11289 ( .A(DB[3494]), .B(DB[3487]), .Z(n8211) );
  AND U11290 ( .A(n54), .B(n8212), .Z(n8210) );
  XOR U11291 ( .A(n8213), .B(n8214), .Z(n8212) );
  XOR U11292 ( .A(DB[3487]), .B(DB[3480]), .Z(n8214) );
  AND U11293 ( .A(n58), .B(n8215), .Z(n8213) );
  XOR U11294 ( .A(n8216), .B(n8217), .Z(n8215) );
  XOR U11295 ( .A(DB[3480]), .B(DB[3473]), .Z(n8217) );
  AND U11296 ( .A(n62), .B(n8218), .Z(n8216) );
  XOR U11297 ( .A(n8219), .B(n8220), .Z(n8218) );
  XOR U11298 ( .A(DB[3473]), .B(DB[3466]), .Z(n8220) );
  AND U11299 ( .A(n66), .B(n8221), .Z(n8219) );
  XOR U11300 ( .A(n8222), .B(n8223), .Z(n8221) );
  XOR U11301 ( .A(DB[3466]), .B(DB[3459]), .Z(n8223) );
  AND U11302 ( .A(n70), .B(n8224), .Z(n8222) );
  XOR U11303 ( .A(n8225), .B(n8226), .Z(n8224) );
  XOR U11304 ( .A(DB[3459]), .B(DB[3452]), .Z(n8226) );
  AND U11305 ( .A(n74), .B(n8227), .Z(n8225) );
  XOR U11306 ( .A(n8228), .B(n8229), .Z(n8227) );
  XOR U11307 ( .A(DB[3452]), .B(DB[3445]), .Z(n8229) );
  AND U11308 ( .A(n78), .B(n8230), .Z(n8228) );
  XOR U11309 ( .A(n8231), .B(n8232), .Z(n8230) );
  XOR U11310 ( .A(DB[3445]), .B(DB[3438]), .Z(n8232) );
  AND U11311 ( .A(n82), .B(n8233), .Z(n8231) );
  XOR U11312 ( .A(n8234), .B(n8235), .Z(n8233) );
  XOR U11313 ( .A(DB[3438]), .B(DB[3431]), .Z(n8235) );
  AND U11314 ( .A(n86), .B(n8236), .Z(n8234) );
  XOR U11315 ( .A(n8237), .B(n8238), .Z(n8236) );
  XOR U11316 ( .A(DB[3431]), .B(DB[3424]), .Z(n8238) );
  AND U11317 ( .A(n90), .B(n8239), .Z(n8237) );
  XOR U11318 ( .A(n8240), .B(n8241), .Z(n8239) );
  XOR U11319 ( .A(DB[3424]), .B(DB[3417]), .Z(n8241) );
  AND U11320 ( .A(n94), .B(n8242), .Z(n8240) );
  XOR U11321 ( .A(n8243), .B(n8244), .Z(n8242) );
  XOR U11322 ( .A(DB[3417]), .B(DB[3410]), .Z(n8244) );
  AND U11323 ( .A(n98), .B(n8245), .Z(n8243) );
  XOR U11324 ( .A(n8246), .B(n8247), .Z(n8245) );
  XOR U11325 ( .A(DB[3410]), .B(DB[3403]), .Z(n8247) );
  AND U11326 ( .A(n102), .B(n8248), .Z(n8246) );
  XOR U11327 ( .A(n8249), .B(n8250), .Z(n8248) );
  XOR U11328 ( .A(DB[3403]), .B(DB[3396]), .Z(n8250) );
  AND U11329 ( .A(n106), .B(n8251), .Z(n8249) );
  XOR U11330 ( .A(n8252), .B(n8253), .Z(n8251) );
  XOR U11331 ( .A(DB[3396]), .B(DB[3389]), .Z(n8253) );
  AND U11332 ( .A(n110), .B(n8254), .Z(n8252) );
  XOR U11333 ( .A(n8255), .B(n8256), .Z(n8254) );
  XOR U11334 ( .A(DB[3389]), .B(DB[3382]), .Z(n8256) );
  AND U11335 ( .A(n114), .B(n8257), .Z(n8255) );
  XOR U11336 ( .A(n8258), .B(n8259), .Z(n8257) );
  XOR U11337 ( .A(DB[3382]), .B(DB[3375]), .Z(n8259) );
  AND U11338 ( .A(n118), .B(n8260), .Z(n8258) );
  XOR U11339 ( .A(n8261), .B(n8262), .Z(n8260) );
  XOR U11340 ( .A(DB[3375]), .B(DB[3368]), .Z(n8262) );
  AND U11341 ( .A(n122), .B(n8263), .Z(n8261) );
  XOR U11342 ( .A(n8264), .B(n8265), .Z(n8263) );
  XOR U11343 ( .A(DB[3368]), .B(DB[3361]), .Z(n8265) );
  AND U11344 ( .A(n126), .B(n8266), .Z(n8264) );
  XOR U11345 ( .A(n8267), .B(n8268), .Z(n8266) );
  XOR U11346 ( .A(DB[3361]), .B(DB[3354]), .Z(n8268) );
  AND U11347 ( .A(n130), .B(n8269), .Z(n8267) );
  XOR U11348 ( .A(n8270), .B(n8271), .Z(n8269) );
  XOR U11349 ( .A(DB[3354]), .B(DB[3347]), .Z(n8271) );
  AND U11350 ( .A(n134), .B(n8272), .Z(n8270) );
  XOR U11351 ( .A(n8273), .B(n8274), .Z(n8272) );
  XOR U11352 ( .A(DB[3347]), .B(DB[3340]), .Z(n8274) );
  AND U11353 ( .A(n138), .B(n8275), .Z(n8273) );
  XOR U11354 ( .A(n8276), .B(n8277), .Z(n8275) );
  XOR U11355 ( .A(DB[3340]), .B(DB[3333]), .Z(n8277) );
  AND U11356 ( .A(n142), .B(n8278), .Z(n8276) );
  XOR U11357 ( .A(n8279), .B(n8280), .Z(n8278) );
  XOR U11358 ( .A(DB[3333]), .B(DB[3326]), .Z(n8280) );
  AND U11359 ( .A(n146), .B(n8281), .Z(n8279) );
  XOR U11360 ( .A(n8282), .B(n8283), .Z(n8281) );
  XOR U11361 ( .A(DB[3326]), .B(DB[3319]), .Z(n8283) );
  AND U11362 ( .A(n150), .B(n8284), .Z(n8282) );
  XOR U11363 ( .A(n8285), .B(n8286), .Z(n8284) );
  XOR U11364 ( .A(DB[3319]), .B(DB[3312]), .Z(n8286) );
  AND U11365 ( .A(n154), .B(n8287), .Z(n8285) );
  XOR U11366 ( .A(n8288), .B(n8289), .Z(n8287) );
  XOR U11367 ( .A(DB[3312]), .B(DB[3305]), .Z(n8289) );
  AND U11368 ( .A(n158), .B(n8290), .Z(n8288) );
  XOR U11369 ( .A(n8291), .B(n8292), .Z(n8290) );
  XOR U11370 ( .A(DB[3305]), .B(DB[3298]), .Z(n8292) );
  AND U11371 ( .A(n162), .B(n8293), .Z(n8291) );
  XOR U11372 ( .A(n8294), .B(n8295), .Z(n8293) );
  XOR U11373 ( .A(DB[3298]), .B(DB[3291]), .Z(n8295) );
  AND U11374 ( .A(n166), .B(n8296), .Z(n8294) );
  XOR U11375 ( .A(n8297), .B(n8298), .Z(n8296) );
  XOR U11376 ( .A(DB[3291]), .B(DB[3284]), .Z(n8298) );
  AND U11377 ( .A(n170), .B(n8299), .Z(n8297) );
  XOR U11378 ( .A(n8300), .B(n8301), .Z(n8299) );
  XOR U11379 ( .A(DB[3284]), .B(DB[3277]), .Z(n8301) );
  AND U11380 ( .A(n174), .B(n8302), .Z(n8300) );
  XOR U11381 ( .A(n8303), .B(n8304), .Z(n8302) );
  XOR U11382 ( .A(DB[3277]), .B(DB[3270]), .Z(n8304) );
  AND U11383 ( .A(n178), .B(n8305), .Z(n8303) );
  XOR U11384 ( .A(n8306), .B(n8307), .Z(n8305) );
  XOR U11385 ( .A(DB[3270]), .B(DB[3263]), .Z(n8307) );
  AND U11386 ( .A(n182), .B(n8308), .Z(n8306) );
  XOR U11387 ( .A(n8309), .B(n8310), .Z(n8308) );
  XOR U11388 ( .A(DB[3263]), .B(DB[3256]), .Z(n8310) );
  AND U11389 ( .A(n186), .B(n8311), .Z(n8309) );
  XOR U11390 ( .A(n8312), .B(n8313), .Z(n8311) );
  XOR U11391 ( .A(DB[3256]), .B(DB[3249]), .Z(n8313) );
  AND U11392 ( .A(n190), .B(n8314), .Z(n8312) );
  XOR U11393 ( .A(n8315), .B(n8316), .Z(n8314) );
  XOR U11394 ( .A(DB[3249]), .B(DB[3242]), .Z(n8316) );
  AND U11395 ( .A(n194), .B(n8317), .Z(n8315) );
  XOR U11396 ( .A(n8318), .B(n8319), .Z(n8317) );
  XOR U11397 ( .A(DB[3242]), .B(DB[3235]), .Z(n8319) );
  AND U11398 ( .A(n198), .B(n8320), .Z(n8318) );
  XOR U11399 ( .A(n8321), .B(n8322), .Z(n8320) );
  XOR U11400 ( .A(DB[3235]), .B(DB[3228]), .Z(n8322) );
  AND U11401 ( .A(n202), .B(n8323), .Z(n8321) );
  XOR U11402 ( .A(n8324), .B(n8325), .Z(n8323) );
  XOR U11403 ( .A(DB[3228]), .B(DB[3221]), .Z(n8325) );
  AND U11404 ( .A(n206), .B(n8326), .Z(n8324) );
  XOR U11405 ( .A(n8327), .B(n8328), .Z(n8326) );
  XOR U11406 ( .A(DB[3221]), .B(DB[3214]), .Z(n8328) );
  AND U11407 ( .A(n210), .B(n8329), .Z(n8327) );
  XOR U11408 ( .A(n8330), .B(n8331), .Z(n8329) );
  XOR U11409 ( .A(DB[3214]), .B(DB[3207]), .Z(n8331) );
  AND U11410 ( .A(n214), .B(n8332), .Z(n8330) );
  XOR U11411 ( .A(n8333), .B(n8334), .Z(n8332) );
  XOR U11412 ( .A(DB[3207]), .B(DB[3200]), .Z(n8334) );
  AND U11413 ( .A(n218), .B(n8335), .Z(n8333) );
  XOR U11414 ( .A(n8336), .B(n8337), .Z(n8335) );
  XOR U11415 ( .A(DB[3200]), .B(DB[3193]), .Z(n8337) );
  AND U11416 ( .A(n222), .B(n8338), .Z(n8336) );
  XOR U11417 ( .A(n8339), .B(n8340), .Z(n8338) );
  XOR U11418 ( .A(DB[3193]), .B(DB[3186]), .Z(n8340) );
  AND U11419 ( .A(n226), .B(n8341), .Z(n8339) );
  XOR U11420 ( .A(n8342), .B(n8343), .Z(n8341) );
  XOR U11421 ( .A(DB[3186]), .B(DB[3179]), .Z(n8343) );
  AND U11422 ( .A(n230), .B(n8344), .Z(n8342) );
  XOR U11423 ( .A(n8345), .B(n8346), .Z(n8344) );
  XOR U11424 ( .A(DB[3179]), .B(DB[3172]), .Z(n8346) );
  AND U11425 ( .A(n234), .B(n8347), .Z(n8345) );
  XOR U11426 ( .A(n8348), .B(n8349), .Z(n8347) );
  XOR U11427 ( .A(DB[3172]), .B(DB[3165]), .Z(n8349) );
  AND U11428 ( .A(n238), .B(n8350), .Z(n8348) );
  XOR U11429 ( .A(n8351), .B(n8352), .Z(n8350) );
  XOR U11430 ( .A(DB[3165]), .B(DB[3158]), .Z(n8352) );
  AND U11431 ( .A(n242), .B(n8353), .Z(n8351) );
  XOR U11432 ( .A(n8354), .B(n8355), .Z(n8353) );
  XOR U11433 ( .A(DB[3158]), .B(DB[3151]), .Z(n8355) );
  AND U11434 ( .A(n246), .B(n8356), .Z(n8354) );
  XOR U11435 ( .A(n8357), .B(n8358), .Z(n8356) );
  XOR U11436 ( .A(DB[3151]), .B(DB[3144]), .Z(n8358) );
  AND U11437 ( .A(n250), .B(n8359), .Z(n8357) );
  XOR U11438 ( .A(n8360), .B(n8361), .Z(n8359) );
  XOR U11439 ( .A(DB[3144]), .B(DB[3137]), .Z(n8361) );
  AND U11440 ( .A(n254), .B(n8362), .Z(n8360) );
  XOR U11441 ( .A(n8363), .B(n8364), .Z(n8362) );
  XOR U11442 ( .A(DB[3137]), .B(DB[3130]), .Z(n8364) );
  AND U11443 ( .A(n258), .B(n8365), .Z(n8363) );
  XOR U11444 ( .A(n8366), .B(n8367), .Z(n8365) );
  XOR U11445 ( .A(DB[3130]), .B(DB[3123]), .Z(n8367) );
  AND U11446 ( .A(n262), .B(n8368), .Z(n8366) );
  XOR U11447 ( .A(n8369), .B(n8370), .Z(n8368) );
  XOR U11448 ( .A(DB[3123]), .B(DB[3116]), .Z(n8370) );
  AND U11449 ( .A(n266), .B(n8371), .Z(n8369) );
  XOR U11450 ( .A(n8372), .B(n8373), .Z(n8371) );
  XOR U11451 ( .A(DB[3116]), .B(DB[3109]), .Z(n8373) );
  AND U11452 ( .A(n270), .B(n8374), .Z(n8372) );
  XOR U11453 ( .A(n8375), .B(n8376), .Z(n8374) );
  XOR U11454 ( .A(DB[3109]), .B(DB[3102]), .Z(n8376) );
  AND U11455 ( .A(n274), .B(n8377), .Z(n8375) );
  XOR U11456 ( .A(n8378), .B(n8379), .Z(n8377) );
  XOR U11457 ( .A(DB[3102]), .B(DB[3095]), .Z(n8379) );
  AND U11458 ( .A(n278), .B(n8380), .Z(n8378) );
  XOR U11459 ( .A(n8381), .B(n8382), .Z(n8380) );
  XOR U11460 ( .A(DB[3095]), .B(DB[3088]), .Z(n8382) );
  AND U11461 ( .A(n282), .B(n8383), .Z(n8381) );
  XOR U11462 ( .A(n8384), .B(n8385), .Z(n8383) );
  XOR U11463 ( .A(DB[3088]), .B(DB[3081]), .Z(n8385) );
  AND U11464 ( .A(n286), .B(n8386), .Z(n8384) );
  XOR U11465 ( .A(n8387), .B(n8388), .Z(n8386) );
  XOR U11466 ( .A(DB[3081]), .B(DB[3074]), .Z(n8388) );
  AND U11467 ( .A(n290), .B(n8389), .Z(n8387) );
  XOR U11468 ( .A(n8390), .B(n8391), .Z(n8389) );
  XOR U11469 ( .A(DB[3074]), .B(DB[3067]), .Z(n8391) );
  AND U11470 ( .A(n294), .B(n8392), .Z(n8390) );
  XOR U11471 ( .A(n8393), .B(n8394), .Z(n8392) );
  XOR U11472 ( .A(DB[3067]), .B(DB[3060]), .Z(n8394) );
  AND U11473 ( .A(n298), .B(n8395), .Z(n8393) );
  XOR U11474 ( .A(n8396), .B(n8397), .Z(n8395) );
  XOR U11475 ( .A(DB[3060]), .B(DB[3053]), .Z(n8397) );
  AND U11476 ( .A(n302), .B(n8398), .Z(n8396) );
  XOR U11477 ( .A(n8399), .B(n8400), .Z(n8398) );
  XOR U11478 ( .A(DB[3053]), .B(DB[3046]), .Z(n8400) );
  AND U11479 ( .A(n306), .B(n8401), .Z(n8399) );
  XOR U11480 ( .A(n8402), .B(n8403), .Z(n8401) );
  XOR U11481 ( .A(DB[3046]), .B(DB[3039]), .Z(n8403) );
  AND U11482 ( .A(n310), .B(n8404), .Z(n8402) );
  XOR U11483 ( .A(n8405), .B(n8406), .Z(n8404) );
  XOR U11484 ( .A(DB[3039]), .B(DB[3032]), .Z(n8406) );
  AND U11485 ( .A(n314), .B(n8407), .Z(n8405) );
  XOR U11486 ( .A(n8408), .B(n8409), .Z(n8407) );
  XOR U11487 ( .A(DB[3032]), .B(DB[3025]), .Z(n8409) );
  AND U11488 ( .A(n318), .B(n8410), .Z(n8408) );
  XOR U11489 ( .A(n8411), .B(n8412), .Z(n8410) );
  XOR U11490 ( .A(DB[3025]), .B(DB[3018]), .Z(n8412) );
  AND U11491 ( .A(n322), .B(n8413), .Z(n8411) );
  XOR U11492 ( .A(n8414), .B(n8415), .Z(n8413) );
  XOR U11493 ( .A(DB[3018]), .B(DB[3011]), .Z(n8415) );
  AND U11494 ( .A(n326), .B(n8416), .Z(n8414) );
  XOR U11495 ( .A(n8417), .B(n8418), .Z(n8416) );
  XOR U11496 ( .A(DB[3011]), .B(DB[3004]), .Z(n8418) );
  AND U11497 ( .A(n330), .B(n8419), .Z(n8417) );
  XOR U11498 ( .A(n8420), .B(n8421), .Z(n8419) );
  XOR U11499 ( .A(DB[3004]), .B(DB[2997]), .Z(n8421) );
  AND U11500 ( .A(n334), .B(n8422), .Z(n8420) );
  XOR U11501 ( .A(n8423), .B(n8424), .Z(n8422) );
  XOR U11502 ( .A(DB[2997]), .B(DB[2990]), .Z(n8424) );
  AND U11503 ( .A(n338), .B(n8425), .Z(n8423) );
  XOR U11504 ( .A(n8426), .B(n8427), .Z(n8425) );
  XOR U11505 ( .A(DB[2990]), .B(DB[2983]), .Z(n8427) );
  AND U11506 ( .A(n342), .B(n8428), .Z(n8426) );
  XOR U11507 ( .A(n8429), .B(n8430), .Z(n8428) );
  XOR U11508 ( .A(DB[2983]), .B(DB[2976]), .Z(n8430) );
  AND U11509 ( .A(n346), .B(n8431), .Z(n8429) );
  XOR U11510 ( .A(n8432), .B(n8433), .Z(n8431) );
  XOR U11511 ( .A(DB[2976]), .B(DB[2969]), .Z(n8433) );
  AND U11512 ( .A(n350), .B(n8434), .Z(n8432) );
  XOR U11513 ( .A(n8435), .B(n8436), .Z(n8434) );
  XOR U11514 ( .A(DB[2969]), .B(DB[2962]), .Z(n8436) );
  AND U11515 ( .A(n354), .B(n8437), .Z(n8435) );
  XOR U11516 ( .A(n8438), .B(n8439), .Z(n8437) );
  XOR U11517 ( .A(DB[2962]), .B(DB[2955]), .Z(n8439) );
  AND U11518 ( .A(n358), .B(n8440), .Z(n8438) );
  XOR U11519 ( .A(n8441), .B(n8442), .Z(n8440) );
  XOR U11520 ( .A(DB[2955]), .B(DB[2948]), .Z(n8442) );
  AND U11521 ( .A(n362), .B(n8443), .Z(n8441) );
  XOR U11522 ( .A(n8444), .B(n8445), .Z(n8443) );
  XOR U11523 ( .A(DB[2948]), .B(DB[2941]), .Z(n8445) );
  AND U11524 ( .A(n366), .B(n8446), .Z(n8444) );
  XOR U11525 ( .A(n8447), .B(n8448), .Z(n8446) );
  XOR U11526 ( .A(DB[2941]), .B(DB[2934]), .Z(n8448) );
  AND U11527 ( .A(n370), .B(n8449), .Z(n8447) );
  XOR U11528 ( .A(n8450), .B(n8451), .Z(n8449) );
  XOR U11529 ( .A(DB[2934]), .B(DB[2927]), .Z(n8451) );
  AND U11530 ( .A(n374), .B(n8452), .Z(n8450) );
  XOR U11531 ( .A(n8453), .B(n8454), .Z(n8452) );
  XOR U11532 ( .A(DB[2927]), .B(DB[2920]), .Z(n8454) );
  AND U11533 ( .A(n378), .B(n8455), .Z(n8453) );
  XOR U11534 ( .A(n8456), .B(n8457), .Z(n8455) );
  XOR U11535 ( .A(DB[2920]), .B(DB[2913]), .Z(n8457) );
  AND U11536 ( .A(n382), .B(n8458), .Z(n8456) );
  XOR U11537 ( .A(n8459), .B(n8460), .Z(n8458) );
  XOR U11538 ( .A(DB[2913]), .B(DB[2906]), .Z(n8460) );
  AND U11539 ( .A(n386), .B(n8461), .Z(n8459) );
  XOR U11540 ( .A(n8462), .B(n8463), .Z(n8461) );
  XOR U11541 ( .A(DB[2906]), .B(DB[2899]), .Z(n8463) );
  AND U11542 ( .A(n390), .B(n8464), .Z(n8462) );
  XOR U11543 ( .A(n8465), .B(n8466), .Z(n8464) );
  XOR U11544 ( .A(DB[2899]), .B(DB[2892]), .Z(n8466) );
  AND U11545 ( .A(n394), .B(n8467), .Z(n8465) );
  XOR U11546 ( .A(n8468), .B(n8469), .Z(n8467) );
  XOR U11547 ( .A(DB[2892]), .B(DB[2885]), .Z(n8469) );
  AND U11548 ( .A(n398), .B(n8470), .Z(n8468) );
  XOR U11549 ( .A(n8471), .B(n8472), .Z(n8470) );
  XOR U11550 ( .A(DB[2885]), .B(DB[2878]), .Z(n8472) );
  AND U11551 ( .A(n402), .B(n8473), .Z(n8471) );
  XOR U11552 ( .A(n8474), .B(n8475), .Z(n8473) );
  XOR U11553 ( .A(DB[2878]), .B(DB[2871]), .Z(n8475) );
  AND U11554 ( .A(n406), .B(n8476), .Z(n8474) );
  XOR U11555 ( .A(n8477), .B(n8478), .Z(n8476) );
  XOR U11556 ( .A(DB[2871]), .B(DB[2864]), .Z(n8478) );
  AND U11557 ( .A(n410), .B(n8479), .Z(n8477) );
  XOR U11558 ( .A(n8480), .B(n8481), .Z(n8479) );
  XOR U11559 ( .A(DB[2864]), .B(DB[2857]), .Z(n8481) );
  AND U11560 ( .A(n414), .B(n8482), .Z(n8480) );
  XOR U11561 ( .A(n8483), .B(n8484), .Z(n8482) );
  XOR U11562 ( .A(DB[2857]), .B(DB[2850]), .Z(n8484) );
  AND U11563 ( .A(n418), .B(n8485), .Z(n8483) );
  XOR U11564 ( .A(n8486), .B(n8487), .Z(n8485) );
  XOR U11565 ( .A(DB[2850]), .B(DB[2843]), .Z(n8487) );
  AND U11566 ( .A(n422), .B(n8488), .Z(n8486) );
  XOR U11567 ( .A(n8489), .B(n8490), .Z(n8488) );
  XOR U11568 ( .A(DB[2843]), .B(DB[2836]), .Z(n8490) );
  AND U11569 ( .A(n426), .B(n8491), .Z(n8489) );
  XOR U11570 ( .A(n8492), .B(n8493), .Z(n8491) );
  XOR U11571 ( .A(DB[2836]), .B(DB[2829]), .Z(n8493) );
  AND U11572 ( .A(n430), .B(n8494), .Z(n8492) );
  XOR U11573 ( .A(n8495), .B(n8496), .Z(n8494) );
  XOR U11574 ( .A(DB[2829]), .B(DB[2822]), .Z(n8496) );
  AND U11575 ( .A(n434), .B(n8497), .Z(n8495) );
  XOR U11576 ( .A(n8498), .B(n8499), .Z(n8497) );
  XOR U11577 ( .A(DB[2822]), .B(DB[2815]), .Z(n8499) );
  AND U11578 ( .A(n438), .B(n8500), .Z(n8498) );
  XOR U11579 ( .A(n8501), .B(n8502), .Z(n8500) );
  XOR U11580 ( .A(DB[2815]), .B(DB[2808]), .Z(n8502) );
  AND U11581 ( .A(n442), .B(n8503), .Z(n8501) );
  XOR U11582 ( .A(n8504), .B(n8505), .Z(n8503) );
  XOR U11583 ( .A(DB[2808]), .B(DB[2801]), .Z(n8505) );
  AND U11584 ( .A(n446), .B(n8506), .Z(n8504) );
  XOR U11585 ( .A(n8507), .B(n8508), .Z(n8506) );
  XOR U11586 ( .A(DB[2801]), .B(DB[2794]), .Z(n8508) );
  AND U11587 ( .A(n450), .B(n8509), .Z(n8507) );
  XOR U11588 ( .A(n8510), .B(n8511), .Z(n8509) );
  XOR U11589 ( .A(DB[2794]), .B(DB[2787]), .Z(n8511) );
  AND U11590 ( .A(n454), .B(n8512), .Z(n8510) );
  XOR U11591 ( .A(n8513), .B(n8514), .Z(n8512) );
  XOR U11592 ( .A(DB[2787]), .B(DB[2780]), .Z(n8514) );
  AND U11593 ( .A(n458), .B(n8515), .Z(n8513) );
  XOR U11594 ( .A(n8516), .B(n8517), .Z(n8515) );
  XOR U11595 ( .A(DB[2780]), .B(DB[2773]), .Z(n8517) );
  AND U11596 ( .A(n462), .B(n8518), .Z(n8516) );
  XOR U11597 ( .A(n8519), .B(n8520), .Z(n8518) );
  XOR U11598 ( .A(DB[2773]), .B(DB[2766]), .Z(n8520) );
  AND U11599 ( .A(n466), .B(n8521), .Z(n8519) );
  XOR U11600 ( .A(n8522), .B(n8523), .Z(n8521) );
  XOR U11601 ( .A(DB[2766]), .B(DB[2759]), .Z(n8523) );
  AND U11602 ( .A(n470), .B(n8524), .Z(n8522) );
  XOR U11603 ( .A(n8525), .B(n8526), .Z(n8524) );
  XOR U11604 ( .A(DB[2759]), .B(DB[2752]), .Z(n8526) );
  AND U11605 ( .A(n474), .B(n8527), .Z(n8525) );
  XOR U11606 ( .A(n8528), .B(n8529), .Z(n8527) );
  XOR U11607 ( .A(DB[2752]), .B(DB[2745]), .Z(n8529) );
  AND U11608 ( .A(n478), .B(n8530), .Z(n8528) );
  XOR U11609 ( .A(n8531), .B(n8532), .Z(n8530) );
  XOR U11610 ( .A(DB[2745]), .B(DB[2738]), .Z(n8532) );
  AND U11611 ( .A(n482), .B(n8533), .Z(n8531) );
  XOR U11612 ( .A(n8534), .B(n8535), .Z(n8533) );
  XOR U11613 ( .A(DB[2738]), .B(DB[2731]), .Z(n8535) );
  AND U11614 ( .A(n486), .B(n8536), .Z(n8534) );
  XOR U11615 ( .A(n8537), .B(n8538), .Z(n8536) );
  XOR U11616 ( .A(DB[2731]), .B(DB[2724]), .Z(n8538) );
  AND U11617 ( .A(n490), .B(n8539), .Z(n8537) );
  XOR U11618 ( .A(n8540), .B(n8541), .Z(n8539) );
  XOR U11619 ( .A(DB[2724]), .B(DB[2717]), .Z(n8541) );
  AND U11620 ( .A(n494), .B(n8542), .Z(n8540) );
  XOR U11621 ( .A(n8543), .B(n8544), .Z(n8542) );
  XOR U11622 ( .A(DB[2717]), .B(DB[2710]), .Z(n8544) );
  AND U11623 ( .A(n498), .B(n8545), .Z(n8543) );
  XOR U11624 ( .A(n8546), .B(n8547), .Z(n8545) );
  XOR U11625 ( .A(DB[2710]), .B(DB[2703]), .Z(n8547) );
  AND U11626 ( .A(n502), .B(n8548), .Z(n8546) );
  XOR U11627 ( .A(n8549), .B(n8550), .Z(n8548) );
  XOR U11628 ( .A(DB[2703]), .B(DB[2696]), .Z(n8550) );
  AND U11629 ( .A(n506), .B(n8551), .Z(n8549) );
  XOR U11630 ( .A(n8552), .B(n8553), .Z(n8551) );
  XOR U11631 ( .A(DB[2696]), .B(DB[2689]), .Z(n8553) );
  AND U11632 ( .A(n510), .B(n8554), .Z(n8552) );
  XOR U11633 ( .A(n8555), .B(n8556), .Z(n8554) );
  XOR U11634 ( .A(DB[2689]), .B(DB[2682]), .Z(n8556) );
  AND U11635 ( .A(n514), .B(n8557), .Z(n8555) );
  XOR U11636 ( .A(n8558), .B(n8559), .Z(n8557) );
  XOR U11637 ( .A(DB[2682]), .B(DB[2675]), .Z(n8559) );
  AND U11638 ( .A(n518), .B(n8560), .Z(n8558) );
  XOR U11639 ( .A(n8561), .B(n8562), .Z(n8560) );
  XOR U11640 ( .A(DB[2675]), .B(DB[2668]), .Z(n8562) );
  AND U11641 ( .A(n522), .B(n8563), .Z(n8561) );
  XOR U11642 ( .A(n8564), .B(n8565), .Z(n8563) );
  XOR U11643 ( .A(DB[2668]), .B(DB[2661]), .Z(n8565) );
  AND U11644 ( .A(n526), .B(n8566), .Z(n8564) );
  XOR U11645 ( .A(n8567), .B(n8568), .Z(n8566) );
  XOR U11646 ( .A(DB[2661]), .B(DB[2654]), .Z(n8568) );
  AND U11647 ( .A(n530), .B(n8569), .Z(n8567) );
  XOR U11648 ( .A(n8570), .B(n8571), .Z(n8569) );
  XOR U11649 ( .A(DB[2654]), .B(DB[2647]), .Z(n8571) );
  AND U11650 ( .A(n534), .B(n8572), .Z(n8570) );
  XOR U11651 ( .A(n8573), .B(n8574), .Z(n8572) );
  XOR U11652 ( .A(DB[2647]), .B(DB[2640]), .Z(n8574) );
  AND U11653 ( .A(n538), .B(n8575), .Z(n8573) );
  XOR U11654 ( .A(n8576), .B(n8577), .Z(n8575) );
  XOR U11655 ( .A(DB[2640]), .B(DB[2633]), .Z(n8577) );
  AND U11656 ( .A(n542), .B(n8578), .Z(n8576) );
  XOR U11657 ( .A(n8579), .B(n8580), .Z(n8578) );
  XOR U11658 ( .A(DB[2633]), .B(DB[2626]), .Z(n8580) );
  AND U11659 ( .A(n546), .B(n8581), .Z(n8579) );
  XOR U11660 ( .A(n8582), .B(n8583), .Z(n8581) );
  XOR U11661 ( .A(DB[2626]), .B(DB[2619]), .Z(n8583) );
  AND U11662 ( .A(n550), .B(n8584), .Z(n8582) );
  XOR U11663 ( .A(n8585), .B(n8586), .Z(n8584) );
  XOR U11664 ( .A(DB[2619]), .B(DB[2612]), .Z(n8586) );
  AND U11665 ( .A(n554), .B(n8587), .Z(n8585) );
  XOR U11666 ( .A(n8588), .B(n8589), .Z(n8587) );
  XOR U11667 ( .A(DB[2612]), .B(DB[2605]), .Z(n8589) );
  AND U11668 ( .A(n558), .B(n8590), .Z(n8588) );
  XOR U11669 ( .A(n8591), .B(n8592), .Z(n8590) );
  XOR U11670 ( .A(DB[2605]), .B(DB[2598]), .Z(n8592) );
  AND U11671 ( .A(n562), .B(n8593), .Z(n8591) );
  XOR U11672 ( .A(n8594), .B(n8595), .Z(n8593) );
  XOR U11673 ( .A(DB[2598]), .B(DB[2591]), .Z(n8595) );
  AND U11674 ( .A(n566), .B(n8596), .Z(n8594) );
  XOR U11675 ( .A(n8597), .B(n8598), .Z(n8596) );
  XOR U11676 ( .A(DB[2591]), .B(DB[2584]), .Z(n8598) );
  AND U11677 ( .A(n570), .B(n8599), .Z(n8597) );
  XOR U11678 ( .A(n8600), .B(n8601), .Z(n8599) );
  XOR U11679 ( .A(DB[2584]), .B(DB[2577]), .Z(n8601) );
  AND U11680 ( .A(n574), .B(n8602), .Z(n8600) );
  XOR U11681 ( .A(n8603), .B(n8604), .Z(n8602) );
  XOR U11682 ( .A(DB[2577]), .B(DB[2570]), .Z(n8604) );
  AND U11683 ( .A(n578), .B(n8605), .Z(n8603) );
  XOR U11684 ( .A(n8606), .B(n8607), .Z(n8605) );
  XOR U11685 ( .A(DB[2570]), .B(DB[2563]), .Z(n8607) );
  AND U11686 ( .A(n582), .B(n8608), .Z(n8606) );
  XOR U11687 ( .A(n8609), .B(n8610), .Z(n8608) );
  XOR U11688 ( .A(DB[2563]), .B(DB[2556]), .Z(n8610) );
  AND U11689 ( .A(n586), .B(n8611), .Z(n8609) );
  XOR U11690 ( .A(n8612), .B(n8613), .Z(n8611) );
  XOR U11691 ( .A(DB[2556]), .B(DB[2549]), .Z(n8613) );
  AND U11692 ( .A(n590), .B(n8614), .Z(n8612) );
  XOR U11693 ( .A(n8615), .B(n8616), .Z(n8614) );
  XOR U11694 ( .A(DB[2549]), .B(DB[2542]), .Z(n8616) );
  AND U11695 ( .A(n594), .B(n8617), .Z(n8615) );
  XOR U11696 ( .A(n8618), .B(n8619), .Z(n8617) );
  XOR U11697 ( .A(DB[2542]), .B(DB[2535]), .Z(n8619) );
  AND U11698 ( .A(n598), .B(n8620), .Z(n8618) );
  XOR U11699 ( .A(n8621), .B(n8622), .Z(n8620) );
  XOR U11700 ( .A(DB[2535]), .B(DB[2528]), .Z(n8622) );
  AND U11701 ( .A(n602), .B(n8623), .Z(n8621) );
  XOR U11702 ( .A(n8624), .B(n8625), .Z(n8623) );
  XOR U11703 ( .A(DB[2528]), .B(DB[2521]), .Z(n8625) );
  AND U11704 ( .A(n606), .B(n8626), .Z(n8624) );
  XOR U11705 ( .A(n8627), .B(n8628), .Z(n8626) );
  XOR U11706 ( .A(DB[2521]), .B(DB[2514]), .Z(n8628) );
  AND U11707 ( .A(n610), .B(n8629), .Z(n8627) );
  XOR U11708 ( .A(n8630), .B(n8631), .Z(n8629) );
  XOR U11709 ( .A(DB[2514]), .B(DB[2507]), .Z(n8631) );
  AND U11710 ( .A(n614), .B(n8632), .Z(n8630) );
  XOR U11711 ( .A(n8633), .B(n8634), .Z(n8632) );
  XOR U11712 ( .A(DB[2507]), .B(DB[2500]), .Z(n8634) );
  AND U11713 ( .A(n618), .B(n8635), .Z(n8633) );
  XOR U11714 ( .A(n8636), .B(n8637), .Z(n8635) );
  XOR U11715 ( .A(DB[2500]), .B(DB[2493]), .Z(n8637) );
  AND U11716 ( .A(n622), .B(n8638), .Z(n8636) );
  XOR U11717 ( .A(n8639), .B(n8640), .Z(n8638) );
  XOR U11718 ( .A(DB[2493]), .B(DB[2486]), .Z(n8640) );
  AND U11719 ( .A(n626), .B(n8641), .Z(n8639) );
  XOR U11720 ( .A(n8642), .B(n8643), .Z(n8641) );
  XOR U11721 ( .A(DB[2486]), .B(DB[2479]), .Z(n8643) );
  AND U11722 ( .A(n630), .B(n8644), .Z(n8642) );
  XOR U11723 ( .A(n8645), .B(n8646), .Z(n8644) );
  XOR U11724 ( .A(DB[2479]), .B(DB[2472]), .Z(n8646) );
  AND U11725 ( .A(n634), .B(n8647), .Z(n8645) );
  XOR U11726 ( .A(n8648), .B(n8649), .Z(n8647) );
  XOR U11727 ( .A(DB[2472]), .B(DB[2465]), .Z(n8649) );
  AND U11728 ( .A(n638), .B(n8650), .Z(n8648) );
  XOR U11729 ( .A(n8651), .B(n8652), .Z(n8650) );
  XOR U11730 ( .A(DB[2465]), .B(DB[2458]), .Z(n8652) );
  AND U11731 ( .A(n642), .B(n8653), .Z(n8651) );
  XOR U11732 ( .A(n8654), .B(n8655), .Z(n8653) );
  XOR U11733 ( .A(DB[2458]), .B(DB[2451]), .Z(n8655) );
  AND U11734 ( .A(n646), .B(n8656), .Z(n8654) );
  XOR U11735 ( .A(n8657), .B(n8658), .Z(n8656) );
  XOR U11736 ( .A(DB[2451]), .B(DB[2444]), .Z(n8658) );
  AND U11737 ( .A(n650), .B(n8659), .Z(n8657) );
  XOR U11738 ( .A(n8660), .B(n8661), .Z(n8659) );
  XOR U11739 ( .A(DB[2444]), .B(DB[2437]), .Z(n8661) );
  AND U11740 ( .A(n654), .B(n8662), .Z(n8660) );
  XOR U11741 ( .A(n8663), .B(n8664), .Z(n8662) );
  XOR U11742 ( .A(DB[2437]), .B(DB[2430]), .Z(n8664) );
  AND U11743 ( .A(n658), .B(n8665), .Z(n8663) );
  XOR U11744 ( .A(n8666), .B(n8667), .Z(n8665) );
  XOR U11745 ( .A(DB[2430]), .B(DB[2423]), .Z(n8667) );
  AND U11746 ( .A(n662), .B(n8668), .Z(n8666) );
  XOR U11747 ( .A(n8669), .B(n8670), .Z(n8668) );
  XOR U11748 ( .A(DB[2423]), .B(DB[2416]), .Z(n8670) );
  AND U11749 ( .A(n666), .B(n8671), .Z(n8669) );
  XOR U11750 ( .A(n8672), .B(n8673), .Z(n8671) );
  XOR U11751 ( .A(DB[2416]), .B(DB[2409]), .Z(n8673) );
  AND U11752 ( .A(n670), .B(n8674), .Z(n8672) );
  XOR U11753 ( .A(n8675), .B(n8676), .Z(n8674) );
  XOR U11754 ( .A(DB[2409]), .B(DB[2402]), .Z(n8676) );
  AND U11755 ( .A(n674), .B(n8677), .Z(n8675) );
  XOR U11756 ( .A(n8678), .B(n8679), .Z(n8677) );
  XOR U11757 ( .A(DB[2402]), .B(DB[2395]), .Z(n8679) );
  AND U11758 ( .A(n678), .B(n8680), .Z(n8678) );
  XOR U11759 ( .A(n8681), .B(n8682), .Z(n8680) );
  XOR U11760 ( .A(DB[2395]), .B(DB[2388]), .Z(n8682) );
  AND U11761 ( .A(n682), .B(n8683), .Z(n8681) );
  XOR U11762 ( .A(n8684), .B(n8685), .Z(n8683) );
  XOR U11763 ( .A(DB[2388]), .B(DB[2381]), .Z(n8685) );
  AND U11764 ( .A(n686), .B(n8686), .Z(n8684) );
  XOR U11765 ( .A(n8687), .B(n8688), .Z(n8686) );
  XOR U11766 ( .A(DB[2381]), .B(DB[2374]), .Z(n8688) );
  AND U11767 ( .A(n690), .B(n8689), .Z(n8687) );
  XOR U11768 ( .A(n8690), .B(n8691), .Z(n8689) );
  XOR U11769 ( .A(DB[2374]), .B(DB[2367]), .Z(n8691) );
  AND U11770 ( .A(n694), .B(n8692), .Z(n8690) );
  XOR U11771 ( .A(n8693), .B(n8694), .Z(n8692) );
  XOR U11772 ( .A(DB[2367]), .B(DB[2360]), .Z(n8694) );
  AND U11773 ( .A(n698), .B(n8695), .Z(n8693) );
  XOR U11774 ( .A(n8696), .B(n8697), .Z(n8695) );
  XOR U11775 ( .A(DB[2360]), .B(DB[2353]), .Z(n8697) );
  AND U11776 ( .A(n702), .B(n8698), .Z(n8696) );
  XOR U11777 ( .A(n8699), .B(n8700), .Z(n8698) );
  XOR U11778 ( .A(DB[2353]), .B(DB[2346]), .Z(n8700) );
  AND U11779 ( .A(n706), .B(n8701), .Z(n8699) );
  XOR U11780 ( .A(n8702), .B(n8703), .Z(n8701) );
  XOR U11781 ( .A(DB[2346]), .B(DB[2339]), .Z(n8703) );
  AND U11782 ( .A(n710), .B(n8704), .Z(n8702) );
  XOR U11783 ( .A(n8705), .B(n8706), .Z(n8704) );
  XOR U11784 ( .A(DB[2339]), .B(DB[2332]), .Z(n8706) );
  AND U11785 ( .A(n714), .B(n8707), .Z(n8705) );
  XOR U11786 ( .A(n8708), .B(n8709), .Z(n8707) );
  XOR U11787 ( .A(DB[2332]), .B(DB[2325]), .Z(n8709) );
  AND U11788 ( .A(n718), .B(n8710), .Z(n8708) );
  XOR U11789 ( .A(n8711), .B(n8712), .Z(n8710) );
  XOR U11790 ( .A(DB[2325]), .B(DB[2318]), .Z(n8712) );
  AND U11791 ( .A(n722), .B(n8713), .Z(n8711) );
  XOR U11792 ( .A(n8714), .B(n8715), .Z(n8713) );
  XOR U11793 ( .A(DB[2318]), .B(DB[2311]), .Z(n8715) );
  AND U11794 ( .A(n726), .B(n8716), .Z(n8714) );
  XOR U11795 ( .A(n8717), .B(n8718), .Z(n8716) );
  XOR U11796 ( .A(DB[2311]), .B(DB[2304]), .Z(n8718) );
  AND U11797 ( .A(n730), .B(n8719), .Z(n8717) );
  XOR U11798 ( .A(n8720), .B(n8721), .Z(n8719) );
  XOR U11799 ( .A(DB[2304]), .B(DB[2297]), .Z(n8721) );
  AND U11800 ( .A(n734), .B(n8722), .Z(n8720) );
  XOR U11801 ( .A(n8723), .B(n8724), .Z(n8722) );
  XOR U11802 ( .A(DB[2297]), .B(DB[2290]), .Z(n8724) );
  AND U11803 ( .A(n738), .B(n8725), .Z(n8723) );
  XOR U11804 ( .A(n8726), .B(n8727), .Z(n8725) );
  XOR U11805 ( .A(DB[2290]), .B(DB[2283]), .Z(n8727) );
  AND U11806 ( .A(n742), .B(n8728), .Z(n8726) );
  XOR U11807 ( .A(n8729), .B(n8730), .Z(n8728) );
  XOR U11808 ( .A(DB[2283]), .B(DB[2276]), .Z(n8730) );
  AND U11809 ( .A(n746), .B(n8731), .Z(n8729) );
  XOR U11810 ( .A(n8732), .B(n8733), .Z(n8731) );
  XOR U11811 ( .A(DB[2276]), .B(DB[2269]), .Z(n8733) );
  AND U11812 ( .A(n750), .B(n8734), .Z(n8732) );
  XOR U11813 ( .A(n8735), .B(n8736), .Z(n8734) );
  XOR U11814 ( .A(DB[2269]), .B(DB[2262]), .Z(n8736) );
  AND U11815 ( .A(n754), .B(n8737), .Z(n8735) );
  XOR U11816 ( .A(n8738), .B(n8739), .Z(n8737) );
  XOR U11817 ( .A(DB[2262]), .B(DB[2255]), .Z(n8739) );
  AND U11818 ( .A(n758), .B(n8740), .Z(n8738) );
  XOR U11819 ( .A(n8741), .B(n8742), .Z(n8740) );
  XOR U11820 ( .A(DB[2255]), .B(DB[2248]), .Z(n8742) );
  AND U11821 ( .A(n762), .B(n8743), .Z(n8741) );
  XOR U11822 ( .A(n8744), .B(n8745), .Z(n8743) );
  XOR U11823 ( .A(DB[2248]), .B(DB[2241]), .Z(n8745) );
  AND U11824 ( .A(n766), .B(n8746), .Z(n8744) );
  XOR U11825 ( .A(n8747), .B(n8748), .Z(n8746) );
  XOR U11826 ( .A(DB[2241]), .B(DB[2234]), .Z(n8748) );
  AND U11827 ( .A(n770), .B(n8749), .Z(n8747) );
  XOR U11828 ( .A(n8750), .B(n8751), .Z(n8749) );
  XOR U11829 ( .A(DB[2234]), .B(DB[2227]), .Z(n8751) );
  AND U11830 ( .A(n774), .B(n8752), .Z(n8750) );
  XOR U11831 ( .A(n8753), .B(n8754), .Z(n8752) );
  XOR U11832 ( .A(DB[2227]), .B(DB[2220]), .Z(n8754) );
  AND U11833 ( .A(n778), .B(n8755), .Z(n8753) );
  XOR U11834 ( .A(n8756), .B(n8757), .Z(n8755) );
  XOR U11835 ( .A(DB[2220]), .B(DB[2213]), .Z(n8757) );
  AND U11836 ( .A(n782), .B(n8758), .Z(n8756) );
  XOR U11837 ( .A(n8759), .B(n8760), .Z(n8758) );
  XOR U11838 ( .A(DB[2213]), .B(DB[2206]), .Z(n8760) );
  AND U11839 ( .A(n786), .B(n8761), .Z(n8759) );
  XOR U11840 ( .A(n8762), .B(n8763), .Z(n8761) );
  XOR U11841 ( .A(DB[2206]), .B(DB[2199]), .Z(n8763) );
  AND U11842 ( .A(n790), .B(n8764), .Z(n8762) );
  XOR U11843 ( .A(n8765), .B(n8766), .Z(n8764) );
  XOR U11844 ( .A(DB[2199]), .B(DB[2192]), .Z(n8766) );
  AND U11845 ( .A(n794), .B(n8767), .Z(n8765) );
  XOR U11846 ( .A(n8768), .B(n8769), .Z(n8767) );
  XOR U11847 ( .A(DB[2192]), .B(DB[2185]), .Z(n8769) );
  AND U11848 ( .A(n798), .B(n8770), .Z(n8768) );
  XOR U11849 ( .A(n8771), .B(n8772), .Z(n8770) );
  XOR U11850 ( .A(DB[2185]), .B(DB[2178]), .Z(n8772) );
  AND U11851 ( .A(n802), .B(n8773), .Z(n8771) );
  XOR U11852 ( .A(n8774), .B(n8775), .Z(n8773) );
  XOR U11853 ( .A(DB[2178]), .B(DB[2171]), .Z(n8775) );
  AND U11854 ( .A(n806), .B(n8776), .Z(n8774) );
  XOR U11855 ( .A(n8777), .B(n8778), .Z(n8776) );
  XOR U11856 ( .A(DB[2171]), .B(DB[2164]), .Z(n8778) );
  AND U11857 ( .A(n810), .B(n8779), .Z(n8777) );
  XOR U11858 ( .A(n8780), .B(n8781), .Z(n8779) );
  XOR U11859 ( .A(DB[2164]), .B(DB[2157]), .Z(n8781) );
  AND U11860 ( .A(n814), .B(n8782), .Z(n8780) );
  XOR U11861 ( .A(n8783), .B(n8784), .Z(n8782) );
  XOR U11862 ( .A(DB[2157]), .B(DB[2150]), .Z(n8784) );
  AND U11863 ( .A(n818), .B(n8785), .Z(n8783) );
  XOR U11864 ( .A(n8786), .B(n8787), .Z(n8785) );
  XOR U11865 ( .A(DB[2150]), .B(DB[2143]), .Z(n8787) );
  AND U11866 ( .A(n822), .B(n8788), .Z(n8786) );
  XOR U11867 ( .A(n8789), .B(n8790), .Z(n8788) );
  XOR U11868 ( .A(DB[2143]), .B(DB[2136]), .Z(n8790) );
  AND U11869 ( .A(n826), .B(n8791), .Z(n8789) );
  XOR U11870 ( .A(n8792), .B(n8793), .Z(n8791) );
  XOR U11871 ( .A(DB[2136]), .B(DB[2129]), .Z(n8793) );
  AND U11872 ( .A(n830), .B(n8794), .Z(n8792) );
  XOR U11873 ( .A(n8795), .B(n8796), .Z(n8794) );
  XOR U11874 ( .A(DB[2129]), .B(DB[2122]), .Z(n8796) );
  AND U11875 ( .A(n834), .B(n8797), .Z(n8795) );
  XOR U11876 ( .A(n8798), .B(n8799), .Z(n8797) );
  XOR U11877 ( .A(DB[2122]), .B(DB[2115]), .Z(n8799) );
  AND U11878 ( .A(n838), .B(n8800), .Z(n8798) );
  XOR U11879 ( .A(n8801), .B(n8802), .Z(n8800) );
  XOR U11880 ( .A(DB[2115]), .B(DB[2108]), .Z(n8802) );
  AND U11881 ( .A(n842), .B(n8803), .Z(n8801) );
  XOR U11882 ( .A(n8804), .B(n8805), .Z(n8803) );
  XOR U11883 ( .A(DB[2108]), .B(DB[2101]), .Z(n8805) );
  AND U11884 ( .A(n846), .B(n8806), .Z(n8804) );
  XOR U11885 ( .A(n8807), .B(n8808), .Z(n8806) );
  XOR U11886 ( .A(DB[2101]), .B(DB[2094]), .Z(n8808) );
  AND U11887 ( .A(n850), .B(n8809), .Z(n8807) );
  XOR U11888 ( .A(n8810), .B(n8811), .Z(n8809) );
  XOR U11889 ( .A(DB[2094]), .B(DB[2087]), .Z(n8811) );
  AND U11890 ( .A(n854), .B(n8812), .Z(n8810) );
  XOR U11891 ( .A(n8813), .B(n8814), .Z(n8812) );
  XOR U11892 ( .A(DB[2087]), .B(DB[2080]), .Z(n8814) );
  AND U11893 ( .A(n858), .B(n8815), .Z(n8813) );
  XOR U11894 ( .A(n8816), .B(n8817), .Z(n8815) );
  XOR U11895 ( .A(DB[2080]), .B(DB[2073]), .Z(n8817) );
  AND U11896 ( .A(n862), .B(n8818), .Z(n8816) );
  XOR U11897 ( .A(n8819), .B(n8820), .Z(n8818) );
  XOR U11898 ( .A(DB[2073]), .B(DB[2066]), .Z(n8820) );
  AND U11899 ( .A(n866), .B(n8821), .Z(n8819) );
  XOR U11900 ( .A(n8822), .B(n8823), .Z(n8821) );
  XOR U11901 ( .A(DB[2066]), .B(DB[2059]), .Z(n8823) );
  AND U11902 ( .A(n870), .B(n8824), .Z(n8822) );
  XOR U11903 ( .A(n8825), .B(n8826), .Z(n8824) );
  XOR U11904 ( .A(DB[2059]), .B(DB[2052]), .Z(n8826) );
  AND U11905 ( .A(n874), .B(n8827), .Z(n8825) );
  XOR U11906 ( .A(n8828), .B(n8829), .Z(n8827) );
  XOR U11907 ( .A(DB[2052]), .B(DB[2045]), .Z(n8829) );
  AND U11908 ( .A(n878), .B(n8830), .Z(n8828) );
  XOR U11909 ( .A(n8831), .B(n8832), .Z(n8830) );
  XOR U11910 ( .A(DB[2045]), .B(DB[2038]), .Z(n8832) );
  AND U11911 ( .A(n882), .B(n8833), .Z(n8831) );
  XOR U11912 ( .A(n8834), .B(n8835), .Z(n8833) );
  XOR U11913 ( .A(DB[2038]), .B(DB[2031]), .Z(n8835) );
  AND U11914 ( .A(n886), .B(n8836), .Z(n8834) );
  XOR U11915 ( .A(n8837), .B(n8838), .Z(n8836) );
  XOR U11916 ( .A(DB[2031]), .B(DB[2024]), .Z(n8838) );
  AND U11917 ( .A(n890), .B(n8839), .Z(n8837) );
  XOR U11918 ( .A(n8840), .B(n8841), .Z(n8839) );
  XOR U11919 ( .A(DB[2024]), .B(DB[2017]), .Z(n8841) );
  AND U11920 ( .A(n894), .B(n8842), .Z(n8840) );
  XOR U11921 ( .A(n8843), .B(n8844), .Z(n8842) );
  XOR U11922 ( .A(DB[2017]), .B(DB[2010]), .Z(n8844) );
  AND U11923 ( .A(n898), .B(n8845), .Z(n8843) );
  XOR U11924 ( .A(n8846), .B(n8847), .Z(n8845) );
  XOR U11925 ( .A(DB[2010]), .B(DB[2003]), .Z(n8847) );
  AND U11926 ( .A(n902), .B(n8848), .Z(n8846) );
  XOR U11927 ( .A(n8849), .B(n8850), .Z(n8848) );
  XOR U11928 ( .A(DB[2003]), .B(DB[1996]), .Z(n8850) );
  AND U11929 ( .A(n906), .B(n8851), .Z(n8849) );
  XOR U11930 ( .A(n8852), .B(n8853), .Z(n8851) );
  XOR U11931 ( .A(DB[1996]), .B(DB[1989]), .Z(n8853) );
  AND U11932 ( .A(n910), .B(n8854), .Z(n8852) );
  XOR U11933 ( .A(n8855), .B(n8856), .Z(n8854) );
  XOR U11934 ( .A(DB[1989]), .B(DB[1982]), .Z(n8856) );
  AND U11935 ( .A(n914), .B(n8857), .Z(n8855) );
  XOR U11936 ( .A(n8858), .B(n8859), .Z(n8857) );
  XOR U11937 ( .A(DB[1982]), .B(DB[1975]), .Z(n8859) );
  AND U11938 ( .A(n918), .B(n8860), .Z(n8858) );
  XOR U11939 ( .A(n8861), .B(n8862), .Z(n8860) );
  XOR U11940 ( .A(DB[1975]), .B(DB[1968]), .Z(n8862) );
  AND U11941 ( .A(n922), .B(n8863), .Z(n8861) );
  XOR U11942 ( .A(n8864), .B(n8865), .Z(n8863) );
  XOR U11943 ( .A(DB[1968]), .B(DB[1961]), .Z(n8865) );
  AND U11944 ( .A(n926), .B(n8866), .Z(n8864) );
  XOR U11945 ( .A(n8867), .B(n8868), .Z(n8866) );
  XOR U11946 ( .A(DB[1961]), .B(DB[1954]), .Z(n8868) );
  AND U11947 ( .A(n930), .B(n8869), .Z(n8867) );
  XOR U11948 ( .A(n8870), .B(n8871), .Z(n8869) );
  XOR U11949 ( .A(DB[1954]), .B(DB[1947]), .Z(n8871) );
  AND U11950 ( .A(n934), .B(n8872), .Z(n8870) );
  XOR U11951 ( .A(n8873), .B(n8874), .Z(n8872) );
  XOR U11952 ( .A(DB[1947]), .B(DB[1940]), .Z(n8874) );
  AND U11953 ( .A(n938), .B(n8875), .Z(n8873) );
  XOR U11954 ( .A(n8876), .B(n8877), .Z(n8875) );
  XOR U11955 ( .A(DB[1940]), .B(DB[1933]), .Z(n8877) );
  AND U11956 ( .A(n942), .B(n8878), .Z(n8876) );
  XOR U11957 ( .A(n8879), .B(n8880), .Z(n8878) );
  XOR U11958 ( .A(DB[1933]), .B(DB[1926]), .Z(n8880) );
  AND U11959 ( .A(n946), .B(n8881), .Z(n8879) );
  XOR U11960 ( .A(n8882), .B(n8883), .Z(n8881) );
  XOR U11961 ( .A(DB[1926]), .B(DB[1919]), .Z(n8883) );
  AND U11962 ( .A(n950), .B(n8884), .Z(n8882) );
  XOR U11963 ( .A(n8885), .B(n8886), .Z(n8884) );
  XOR U11964 ( .A(DB[1919]), .B(DB[1912]), .Z(n8886) );
  AND U11965 ( .A(n954), .B(n8887), .Z(n8885) );
  XOR U11966 ( .A(n8888), .B(n8889), .Z(n8887) );
  XOR U11967 ( .A(DB[1912]), .B(DB[1905]), .Z(n8889) );
  AND U11968 ( .A(n958), .B(n8890), .Z(n8888) );
  XOR U11969 ( .A(n8891), .B(n8892), .Z(n8890) );
  XOR U11970 ( .A(DB[1905]), .B(DB[1898]), .Z(n8892) );
  AND U11971 ( .A(n962), .B(n8893), .Z(n8891) );
  XOR U11972 ( .A(n8894), .B(n8895), .Z(n8893) );
  XOR U11973 ( .A(DB[1898]), .B(DB[1891]), .Z(n8895) );
  AND U11974 ( .A(n966), .B(n8896), .Z(n8894) );
  XOR U11975 ( .A(n8897), .B(n8898), .Z(n8896) );
  XOR U11976 ( .A(DB[1891]), .B(DB[1884]), .Z(n8898) );
  AND U11977 ( .A(n970), .B(n8899), .Z(n8897) );
  XOR U11978 ( .A(n8900), .B(n8901), .Z(n8899) );
  XOR U11979 ( .A(DB[1884]), .B(DB[1877]), .Z(n8901) );
  AND U11980 ( .A(n974), .B(n8902), .Z(n8900) );
  XOR U11981 ( .A(n8903), .B(n8904), .Z(n8902) );
  XOR U11982 ( .A(DB[1877]), .B(DB[1870]), .Z(n8904) );
  AND U11983 ( .A(n978), .B(n8905), .Z(n8903) );
  XOR U11984 ( .A(n8906), .B(n8907), .Z(n8905) );
  XOR U11985 ( .A(DB[1870]), .B(DB[1863]), .Z(n8907) );
  AND U11986 ( .A(n982), .B(n8908), .Z(n8906) );
  XOR U11987 ( .A(n8909), .B(n8910), .Z(n8908) );
  XOR U11988 ( .A(DB[1863]), .B(DB[1856]), .Z(n8910) );
  AND U11989 ( .A(n986), .B(n8911), .Z(n8909) );
  XOR U11990 ( .A(n8912), .B(n8913), .Z(n8911) );
  XOR U11991 ( .A(DB[1856]), .B(DB[1849]), .Z(n8913) );
  AND U11992 ( .A(n990), .B(n8914), .Z(n8912) );
  XOR U11993 ( .A(n8915), .B(n8916), .Z(n8914) );
  XOR U11994 ( .A(DB[1849]), .B(DB[1842]), .Z(n8916) );
  AND U11995 ( .A(n994), .B(n8917), .Z(n8915) );
  XOR U11996 ( .A(n8918), .B(n8919), .Z(n8917) );
  XOR U11997 ( .A(DB[1842]), .B(DB[1835]), .Z(n8919) );
  AND U11998 ( .A(n998), .B(n8920), .Z(n8918) );
  XOR U11999 ( .A(n8921), .B(n8922), .Z(n8920) );
  XOR U12000 ( .A(DB[1835]), .B(DB[1828]), .Z(n8922) );
  AND U12001 ( .A(n1002), .B(n8923), .Z(n8921) );
  XOR U12002 ( .A(n8924), .B(n8925), .Z(n8923) );
  XOR U12003 ( .A(DB[1828]), .B(DB[1821]), .Z(n8925) );
  AND U12004 ( .A(n1006), .B(n8926), .Z(n8924) );
  XOR U12005 ( .A(n8927), .B(n8928), .Z(n8926) );
  XOR U12006 ( .A(DB[1821]), .B(DB[1814]), .Z(n8928) );
  AND U12007 ( .A(n1010), .B(n8929), .Z(n8927) );
  XOR U12008 ( .A(n8930), .B(n8931), .Z(n8929) );
  XOR U12009 ( .A(DB[1814]), .B(DB[1807]), .Z(n8931) );
  AND U12010 ( .A(n1014), .B(n8932), .Z(n8930) );
  XOR U12011 ( .A(n8933), .B(n8934), .Z(n8932) );
  XOR U12012 ( .A(DB[1807]), .B(DB[1800]), .Z(n8934) );
  AND U12013 ( .A(n1018), .B(n8935), .Z(n8933) );
  XOR U12014 ( .A(n8936), .B(n8937), .Z(n8935) );
  XOR U12015 ( .A(DB[1800]), .B(DB[1793]), .Z(n8937) );
  AND U12016 ( .A(n1022), .B(n8938), .Z(n8936) );
  XOR U12017 ( .A(n8939), .B(n8940), .Z(n8938) );
  XOR U12018 ( .A(DB[1793]), .B(DB[1786]), .Z(n8940) );
  AND U12019 ( .A(n1026), .B(n8941), .Z(n8939) );
  XOR U12020 ( .A(n8942), .B(n8943), .Z(n8941) );
  XOR U12021 ( .A(DB[1786]), .B(DB[1779]), .Z(n8943) );
  AND U12022 ( .A(n1030), .B(n8944), .Z(n8942) );
  XOR U12023 ( .A(n8945), .B(n8946), .Z(n8944) );
  XOR U12024 ( .A(DB[1779]), .B(DB[1772]), .Z(n8946) );
  AND U12025 ( .A(n1034), .B(n8947), .Z(n8945) );
  XOR U12026 ( .A(n8948), .B(n8949), .Z(n8947) );
  XOR U12027 ( .A(DB[1772]), .B(DB[1765]), .Z(n8949) );
  AND U12028 ( .A(n1038), .B(n8950), .Z(n8948) );
  XOR U12029 ( .A(n8951), .B(n8952), .Z(n8950) );
  XOR U12030 ( .A(DB[1765]), .B(DB[1758]), .Z(n8952) );
  AND U12031 ( .A(n1042), .B(n8953), .Z(n8951) );
  XOR U12032 ( .A(n8954), .B(n8955), .Z(n8953) );
  XOR U12033 ( .A(DB[1758]), .B(DB[1751]), .Z(n8955) );
  AND U12034 ( .A(n1046), .B(n8956), .Z(n8954) );
  XOR U12035 ( .A(n8957), .B(n8958), .Z(n8956) );
  XOR U12036 ( .A(DB[1751]), .B(DB[1744]), .Z(n8958) );
  AND U12037 ( .A(n1050), .B(n8959), .Z(n8957) );
  XOR U12038 ( .A(n8960), .B(n8961), .Z(n8959) );
  XOR U12039 ( .A(DB[1744]), .B(DB[1737]), .Z(n8961) );
  AND U12040 ( .A(n1054), .B(n8962), .Z(n8960) );
  XOR U12041 ( .A(n8963), .B(n8964), .Z(n8962) );
  XOR U12042 ( .A(DB[1737]), .B(DB[1730]), .Z(n8964) );
  AND U12043 ( .A(n1058), .B(n8965), .Z(n8963) );
  XOR U12044 ( .A(n8966), .B(n8967), .Z(n8965) );
  XOR U12045 ( .A(DB[1730]), .B(DB[1723]), .Z(n8967) );
  AND U12046 ( .A(n1062), .B(n8968), .Z(n8966) );
  XOR U12047 ( .A(n8969), .B(n8970), .Z(n8968) );
  XOR U12048 ( .A(DB[1723]), .B(DB[1716]), .Z(n8970) );
  AND U12049 ( .A(n1066), .B(n8971), .Z(n8969) );
  XOR U12050 ( .A(n8972), .B(n8973), .Z(n8971) );
  XOR U12051 ( .A(DB[1716]), .B(DB[1709]), .Z(n8973) );
  AND U12052 ( .A(n1070), .B(n8974), .Z(n8972) );
  XOR U12053 ( .A(n8975), .B(n8976), .Z(n8974) );
  XOR U12054 ( .A(DB[1709]), .B(DB[1702]), .Z(n8976) );
  AND U12055 ( .A(n1074), .B(n8977), .Z(n8975) );
  XOR U12056 ( .A(n8978), .B(n8979), .Z(n8977) );
  XOR U12057 ( .A(DB[1702]), .B(DB[1695]), .Z(n8979) );
  AND U12058 ( .A(n1078), .B(n8980), .Z(n8978) );
  XOR U12059 ( .A(n8981), .B(n8982), .Z(n8980) );
  XOR U12060 ( .A(DB[1695]), .B(DB[1688]), .Z(n8982) );
  AND U12061 ( .A(n1082), .B(n8983), .Z(n8981) );
  XOR U12062 ( .A(n8984), .B(n8985), .Z(n8983) );
  XOR U12063 ( .A(DB[1688]), .B(DB[1681]), .Z(n8985) );
  AND U12064 ( .A(n1086), .B(n8986), .Z(n8984) );
  XOR U12065 ( .A(n8987), .B(n8988), .Z(n8986) );
  XOR U12066 ( .A(DB[1681]), .B(DB[1674]), .Z(n8988) );
  AND U12067 ( .A(n1090), .B(n8989), .Z(n8987) );
  XOR U12068 ( .A(n8990), .B(n8991), .Z(n8989) );
  XOR U12069 ( .A(DB[1674]), .B(DB[1667]), .Z(n8991) );
  AND U12070 ( .A(n1094), .B(n8992), .Z(n8990) );
  XOR U12071 ( .A(n8993), .B(n8994), .Z(n8992) );
  XOR U12072 ( .A(DB[1667]), .B(DB[1660]), .Z(n8994) );
  AND U12073 ( .A(n1098), .B(n8995), .Z(n8993) );
  XOR U12074 ( .A(n8996), .B(n8997), .Z(n8995) );
  XOR U12075 ( .A(DB[1660]), .B(DB[1653]), .Z(n8997) );
  AND U12076 ( .A(n1102), .B(n8998), .Z(n8996) );
  XOR U12077 ( .A(n8999), .B(n9000), .Z(n8998) );
  XOR U12078 ( .A(DB[1653]), .B(DB[1646]), .Z(n9000) );
  AND U12079 ( .A(n1106), .B(n9001), .Z(n8999) );
  XOR U12080 ( .A(n9002), .B(n9003), .Z(n9001) );
  XOR U12081 ( .A(DB[1646]), .B(DB[1639]), .Z(n9003) );
  AND U12082 ( .A(n1110), .B(n9004), .Z(n9002) );
  XOR U12083 ( .A(n9005), .B(n9006), .Z(n9004) );
  XOR U12084 ( .A(DB[1639]), .B(DB[1632]), .Z(n9006) );
  AND U12085 ( .A(n1114), .B(n9007), .Z(n9005) );
  XOR U12086 ( .A(n9008), .B(n9009), .Z(n9007) );
  XOR U12087 ( .A(DB[1632]), .B(DB[1625]), .Z(n9009) );
  AND U12088 ( .A(n1118), .B(n9010), .Z(n9008) );
  XOR U12089 ( .A(n9011), .B(n9012), .Z(n9010) );
  XOR U12090 ( .A(DB[1625]), .B(DB[1618]), .Z(n9012) );
  AND U12091 ( .A(n1122), .B(n9013), .Z(n9011) );
  XOR U12092 ( .A(n9014), .B(n9015), .Z(n9013) );
  XOR U12093 ( .A(DB[1618]), .B(DB[1611]), .Z(n9015) );
  AND U12094 ( .A(n1126), .B(n9016), .Z(n9014) );
  XOR U12095 ( .A(n9017), .B(n9018), .Z(n9016) );
  XOR U12096 ( .A(DB[1611]), .B(DB[1604]), .Z(n9018) );
  AND U12097 ( .A(n1130), .B(n9019), .Z(n9017) );
  XOR U12098 ( .A(n9020), .B(n9021), .Z(n9019) );
  XOR U12099 ( .A(DB[1604]), .B(DB[1597]), .Z(n9021) );
  AND U12100 ( .A(n1134), .B(n9022), .Z(n9020) );
  XOR U12101 ( .A(n9023), .B(n9024), .Z(n9022) );
  XOR U12102 ( .A(DB[1597]), .B(DB[1590]), .Z(n9024) );
  AND U12103 ( .A(n1138), .B(n9025), .Z(n9023) );
  XOR U12104 ( .A(n9026), .B(n9027), .Z(n9025) );
  XOR U12105 ( .A(DB[1590]), .B(DB[1583]), .Z(n9027) );
  AND U12106 ( .A(n1142), .B(n9028), .Z(n9026) );
  XOR U12107 ( .A(n9029), .B(n9030), .Z(n9028) );
  XOR U12108 ( .A(DB[1583]), .B(DB[1576]), .Z(n9030) );
  AND U12109 ( .A(n1146), .B(n9031), .Z(n9029) );
  XOR U12110 ( .A(n9032), .B(n9033), .Z(n9031) );
  XOR U12111 ( .A(DB[1576]), .B(DB[1569]), .Z(n9033) );
  AND U12112 ( .A(n1150), .B(n9034), .Z(n9032) );
  XOR U12113 ( .A(n9035), .B(n9036), .Z(n9034) );
  XOR U12114 ( .A(DB[1569]), .B(DB[1562]), .Z(n9036) );
  AND U12115 ( .A(n1154), .B(n9037), .Z(n9035) );
  XOR U12116 ( .A(n9038), .B(n9039), .Z(n9037) );
  XOR U12117 ( .A(DB[1562]), .B(DB[1555]), .Z(n9039) );
  AND U12118 ( .A(n1158), .B(n9040), .Z(n9038) );
  XOR U12119 ( .A(n9041), .B(n9042), .Z(n9040) );
  XOR U12120 ( .A(DB[1555]), .B(DB[1548]), .Z(n9042) );
  AND U12121 ( .A(n1162), .B(n9043), .Z(n9041) );
  XOR U12122 ( .A(n9044), .B(n9045), .Z(n9043) );
  XOR U12123 ( .A(DB[1548]), .B(DB[1541]), .Z(n9045) );
  AND U12124 ( .A(n1166), .B(n9046), .Z(n9044) );
  XOR U12125 ( .A(n9047), .B(n9048), .Z(n9046) );
  XOR U12126 ( .A(DB[1541]), .B(DB[1534]), .Z(n9048) );
  AND U12127 ( .A(n1170), .B(n9049), .Z(n9047) );
  XOR U12128 ( .A(n9050), .B(n9051), .Z(n9049) );
  XOR U12129 ( .A(DB[1534]), .B(DB[1527]), .Z(n9051) );
  AND U12130 ( .A(n1174), .B(n9052), .Z(n9050) );
  XOR U12131 ( .A(n9053), .B(n9054), .Z(n9052) );
  XOR U12132 ( .A(DB[1527]), .B(DB[1520]), .Z(n9054) );
  AND U12133 ( .A(n1178), .B(n9055), .Z(n9053) );
  XOR U12134 ( .A(n9056), .B(n9057), .Z(n9055) );
  XOR U12135 ( .A(DB[1520]), .B(DB[1513]), .Z(n9057) );
  AND U12136 ( .A(n1182), .B(n9058), .Z(n9056) );
  XOR U12137 ( .A(n9059), .B(n9060), .Z(n9058) );
  XOR U12138 ( .A(DB[1513]), .B(DB[1506]), .Z(n9060) );
  AND U12139 ( .A(n1186), .B(n9061), .Z(n9059) );
  XOR U12140 ( .A(n9062), .B(n9063), .Z(n9061) );
  XOR U12141 ( .A(DB[1506]), .B(DB[1499]), .Z(n9063) );
  AND U12142 ( .A(n1190), .B(n9064), .Z(n9062) );
  XOR U12143 ( .A(n9065), .B(n9066), .Z(n9064) );
  XOR U12144 ( .A(DB[1499]), .B(DB[1492]), .Z(n9066) );
  AND U12145 ( .A(n1194), .B(n9067), .Z(n9065) );
  XOR U12146 ( .A(n9068), .B(n9069), .Z(n9067) );
  XOR U12147 ( .A(DB[1492]), .B(DB[1485]), .Z(n9069) );
  AND U12148 ( .A(n1198), .B(n9070), .Z(n9068) );
  XOR U12149 ( .A(n9071), .B(n9072), .Z(n9070) );
  XOR U12150 ( .A(DB[1485]), .B(DB[1478]), .Z(n9072) );
  AND U12151 ( .A(n1202), .B(n9073), .Z(n9071) );
  XOR U12152 ( .A(n9074), .B(n9075), .Z(n9073) );
  XOR U12153 ( .A(DB[1478]), .B(DB[1471]), .Z(n9075) );
  AND U12154 ( .A(n1206), .B(n9076), .Z(n9074) );
  XOR U12155 ( .A(n9077), .B(n9078), .Z(n9076) );
  XOR U12156 ( .A(DB[1471]), .B(DB[1464]), .Z(n9078) );
  AND U12157 ( .A(n1210), .B(n9079), .Z(n9077) );
  XOR U12158 ( .A(n9080), .B(n9081), .Z(n9079) );
  XOR U12159 ( .A(DB[1464]), .B(DB[1457]), .Z(n9081) );
  AND U12160 ( .A(n1214), .B(n9082), .Z(n9080) );
  XOR U12161 ( .A(n9083), .B(n9084), .Z(n9082) );
  XOR U12162 ( .A(DB[1457]), .B(DB[1450]), .Z(n9084) );
  AND U12163 ( .A(n1218), .B(n9085), .Z(n9083) );
  XOR U12164 ( .A(n9086), .B(n9087), .Z(n9085) );
  XOR U12165 ( .A(DB[1450]), .B(DB[1443]), .Z(n9087) );
  AND U12166 ( .A(n1222), .B(n9088), .Z(n9086) );
  XOR U12167 ( .A(n9089), .B(n9090), .Z(n9088) );
  XOR U12168 ( .A(DB[1443]), .B(DB[1436]), .Z(n9090) );
  AND U12169 ( .A(n1226), .B(n9091), .Z(n9089) );
  XOR U12170 ( .A(n9092), .B(n9093), .Z(n9091) );
  XOR U12171 ( .A(DB[1436]), .B(DB[1429]), .Z(n9093) );
  AND U12172 ( .A(n1230), .B(n9094), .Z(n9092) );
  XOR U12173 ( .A(n9095), .B(n9096), .Z(n9094) );
  XOR U12174 ( .A(DB[1429]), .B(DB[1422]), .Z(n9096) );
  AND U12175 ( .A(n1234), .B(n9097), .Z(n9095) );
  XOR U12176 ( .A(n9098), .B(n9099), .Z(n9097) );
  XOR U12177 ( .A(DB[1422]), .B(DB[1415]), .Z(n9099) );
  AND U12178 ( .A(n1238), .B(n9100), .Z(n9098) );
  XOR U12179 ( .A(n9101), .B(n9102), .Z(n9100) );
  XOR U12180 ( .A(DB[1415]), .B(DB[1408]), .Z(n9102) );
  AND U12181 ( .A(n1242), .B(n9103), .Z(n9101) );
  XOR U12182 ( .A(n9104), .B(n9105), .Z(n9103) );
  XOR U12183 ( .A(DB[1408]), .B(DB[1401]), .Z(n9105) );
  AND U12184 ( .A(n1246), .B(n9106), .Z(n9104) );
  XOR U12185 ( .A(n9107), .B(n9108), .Z(n9106) );
  XOR U12186 ( .A(DB[1401]), .B(DB[1394]), .Z(n9108) );
  AND U12187 ( .A(n1250), .B(n9109), .Z(n9107) );
  XOR U12188 ( .A(n9110), .B(n9111), .Z(n9109) );
  XOR U12189 ( .A(DB[1394]), .B(DB[1387]), .Z(n9111) );
  AND U12190 ( .A(n1254), .B(n9112), .Z(n9110) );
  XOR U12191 ( .A(n9113), .B(n9114), .Z(n9112) );
  XOR U12192 ( .A(DB[1387]), .B(DB[1380]), .Z(n9114) );
  AND U12193 ( .A(n1258), .B(n9115), .Z(n9113) );
  XOR U12194 ( .A(n9116), .B(n9117), .Z(n9115) );
  XOR U12195 ( .A(DB[1380]), .B(DB[1373]), .Z(n9117) );
  AND U12196 ( .A(n1262), .B(n9118), .Z(n9116) );
  XOR U12197 ( .A(n9119), .B(n9120), .Z(n9118) );
  XOR U12198 ( .A(DB[1373]), .B(DB[1366]), .Z(n9120) );
  AND U12199 ( .A(n1266), .B(n9121), .Z(n9119) );
  XOR U12200 ( .A(n9122), .B(n9123), .Z(n9121) );
  XOR U12201 ( .A(DB[1366]), .B(DB[1359]), .Z(n9123) );
  AND U12202 ( .A(n1270), .B(n9124), .Z(n9122) );
  XOR U12203 ( .A(n9125), .B(n9126), .Z(n9124) );
  XOR U12204 ( .A(DB[1359]), .B(DB[1352]), .Z(n9126) );
  AND U12205 ( .A(n1274), .B(n9127), .Z(n9125) );
  XOR U12206 ( .A(n9128), .B(n9129), .Z(n9127) );
  XOR U12207 ( .A(DB[1352]), .B(DB[1345]), .Z(n9129) );
  AND U12208 ( .A(n1278), .B(n9130), .Z(n9128) );
  XOR U12209 ( .A(n9131), .B(n9132), .Z(n9130) );
  XOR U12210 ( .A(DB[1345]), .B(DB[1338]), .Z(n9132) );
  AND U12211 ( .A(n1282), .B(n9133), .Z(n9131) );
  XOR U12212 ( .A(n9134), .B(n9135), .Z(n9133) );
  XOR U12213 ( .A(DB[1338]), .B(DB[1331]), .Z(n9135) );
  AND U12214 ( .A(n1286), .B(n9136), .Z(n9134) );
  XOR U12215 ( .A(n9137), .B(n9138), .Z(n9136) );
  XOR U12216 ( .A(DB[1331]), .B(DB[1324]), .Z(n9138) );
  AND U12217 ( .A(n1290), .B(n9139), .Z(n9137) );
  XOR U12218 ( .A(n9140), .B(n9141), .Z(n9139) );
  XOR U12219 ( .A(DB[1324]), .B(DB[1317]), .Z(n9141) );
  AND U12220 ( .A(n1294), .B(n9142), .Z(n9140) );
  XOR U12221 ( .A(n9143), .B(n9144), .Z(n9142) );
  XOR U12222 ( .A(DB[1317]), .B(DB[1310]), .Z(n9144) );
  AND U12223 ( .A(n1298), .B(n9145), .Z(n9143) );
  XOR U12224 ( .A(n9146), .B(n9147), .Z(n9145) );
  XOR U12225 ( .A(DB[1310]), .B(DB[1303]), .Z(n9147) );
  AND U12226 ( .A(n1302), .B(n9148), .Z(n9146) );
  XOR U12227 ( .A(n9149), .B(n9150), .Z(n9148) );
  XOR U12228 ( .A(DB[1303]), .B(DB[1296]), .Z(n9150) );
  AND U12229 ( .A(n1306), .B(n9151), .Z(n9149) );
  XOR U12230 ( .A(n9152), .B(n9153), .Z(n9151) );
  XOR U12231 ( .A(DB[1296]), .B(DB[1289]), .Z(n9153) );
  AND U12232 ( .A(n1310), .B(n9154), .Z(n9152) );
  XOR U12233 ( .A(n9155), .B(n9156), .Z(n9154) );
  XOR U12234 ( .A(DB[1289]), .B(DB[1282]), .Z(n9156) );
  AND U12235 ( .A(n1314), .B(n9157), .Z(n9155) );
  XOR U12236 ( .A(n9158), .B(n9159), .Z(n9157) );
  XOR U12237 ( .A(DB[1282]), .B(DB[1275]), .Z(n9159) );
  AND U12238 ( .A(n1318), .B(n9160), .Z(n9158) );
  XOR U12239 ( .A(n9161), .B(n9162), .Z(n9160) );
  XOR U12240 ( .A(DB[1275]), .B(DB[1268]), .Z(n9162) );
  AND U12241 ( .A(n1322), .B(n9163), .Z(n9161) );
  XOR U12242 ( .A(n9164), .B(n9165), .Z(n9163) );
  XOR U12243 ( .A(DB[1268]), .B(DB[1261]), .Z(n9165) );
  AND U12244 ( .A(n1326), .B(n9166), .Z(n9164) );
  XOR U12245 ( .A(n9167), .B(n9168), .Z(n9166) );
  XOR U12246 ( .A(DB[1261]), .B(DB[1254]), .Z(n9168) );
  AND U12247 ( .A(n1330), .B(n9169), .Z(n9167) );
  XOR U12248 ( .A(n9170), .B(n9171), .Z(n9169) );
  XOR U12249 ( .A(DB[1254]), .B(DB[1247]), .Z(n9171) );
  AND U12250 ( .A(n1334), .B(n9172), .Z(n9170) );
  XOR U12251 ( .A(n9173), .B(n9174), .Z(n9172) );
  XOR U12252 ( .A(DB[1247]), .B(DB[1240]), .Z(n9174) );
  AND U12253 ( .A(n1338), .B(n9175), .Z(n9173) );
  XOR U12254 ( .A(n9176), .B(n9177), .Z(n9175) );
  XOR U12255 ( .A(DB[1240]), .B(DB[1233]), .Z(n9177) );
  AND U12256 ( .A(n1342), .B(n9178), .Z(n9176) );
  XOR U12257 ( .A(n9179), .B(n9180), .Z(n9178) );
  XOR U12258 ( .A(DB[1233]), .B(DB[1226]), .Z(n9180) );
  AND U12259 ( .A(n1346), .B(n9181), .Z(n9179) );
  XOR U12260 ( .A(n9182), .B(n9183), .Z(n9181) );
  XOR U12261 ( .A(DB[1226]), .B(DB[1219]), .Z(n9183) );
  AND U12262 ( .A(n1350), .B(n9184), .Z(n9182) );
  XOR U12263 ( .A(n9185), .B(n9186), .Z(n9184) );
  XOR U12264 ( .A(DB[1219]), .B(DB[1212]), .Z(n9186) );
  AND U12265 ( .A(n1354), .B(n9187), .Z(n9185) );
  XOR U12266 ( .A(n9188), .B(n9189), .Z(n9187) );
  XOR U12267 ( .A(DB[1212]), .B(DB[1205]), .Z(n9189) );
  AND U12268 ( .A(n1358), .B(n9190), .Z(n9188) );
  XOR U12269 ( .A(n9191), .B(n9192), .Z(n9190) );
  XOR U12270 ( .A(DB[1205]), .B(DB[1198]), .Z(n9192) );
  AND U12271 ( .A(n1362), .B(n9193), .Z(n9191) );
  XOR U12272 ( .A(n9194), .B(n9195), .Z(n9193) );
  XOR U12273 ( .A(DB[1198]), .B(DB[1191]), .Z(n9195) );
  AND U12274 ( .A(n1366), .B(n9196), .Z(n9194) );
  XOR U12275 ( .A(n9197), .B(n9198), .Z(n9196) );
  XOR U12276 ( .A(DB[1191]), .B(DB[1184]), .Z(n9198) );
  AND U12277 ( .A(n1370), .B(n9199), .Z(n9197) );
  XOR U12278 ( .A(n9200), .B(n9201), .Z(n9199) );
  XOR U12279 ( .A(DB[1184]), .B(DB[1177]), .Z(n9201) );
  AND U12280 ( .A(n1374), .B(n9202), .Z(n9200) );
  XOR U12281 ( .A(n9203), .B(n9204), .Z(n9202) );
  XOR U12282 ( .A(DB[1177]), .B(DB[1170]), .Z(n9204) );
  AND U12283 ( .A(n1378), .B(n9205), .Z(n9203) );
  XOR U12284 ( .A(n9206), .B(n9207), .Z(n9205) );
  XOR U12285 ( .A(DB[1170]), .B(DB[1163]), .Z(n9207) );
  AND U12286 ( .A(n1382), .B(n9208), .Z(n9206) );
  XOR U12287 ( .A(n9209), .B(n9210), .Z(n9208) );
  XOR U12288 ( .A(DB[1163]), .B(DB[1156]), .Z(n9210) );
  AND U12289 ( .A(n1386), .B(n9211), .Z(n9209) );
  XOR U12290 ( .A(n9212), .B(n9213), .Z(n9211) );
  XOR U12291 ( .A(DB[1156]), .B(DB[1149]), .Z(n9213) );
  AND U12292 ( .A(n1390), .B(n9214), .Z(n9212) );
  XOR U12293 ( .A(n9215), .B(n9216), .Z(n9214) );
  XOR U12294 ( .A(DB[1149]), .B(DB[1142]), .Z(n9216) );
  AND U12295 ( .A(n1394), .B(n9217), .Z(n9215) );
  XOR U12296 ( .A(n9218), .B(n9219), .Z(n9217) );
  XOR U12297 ( .A(DB[1142]), .B(DB[1135]), .Z(n9219) );
  AND U12298 ( .A(n1398), .B(n9220), .Z(n9218) );
  XOR U12299 ( .A(n9221), .B(n9222), .Z(n9220) );
  XOR U12300 ( .A(DB[1135]), .B(DB[1128]), .Z(n9222) );
  AND U12301 ( .A(n1402), .B(n9223), .Z(n9221) );
  XOR U12302 ( .A(n9224), .B(n9225), .Z(n9223) );
  XOR U12303 ( .A(DB[1128]), .B(DB[1121]), .Z(n9225) );
  AND U12304 ( .A(n1406), .B(n9226), .Z(n9224) );
  XOR U12305 ( .A(n9227), .B(n9228), .Z(n9226) );
  XOR U12306 ( .A(DB[1121]), .B(DB[1114]), .Z(n9228) );
  AND U12307 ( .A(n1410), .B(n9229), .Z(n9227) );
  XOR U12308 ( .A(n9230), .B(n9231), .Z(n9229) );
  XOR U12309 ( .A(DB[1114]), .B(DB[1107]), .Z(n9231) );
  AND U12310 ( .A(n1414), .B(n9232), .Z(n9230) );
  XOR U12311 ( .A(n9233), .B(n9234), .Z(n9232) );
  XOR U12312 ( .A(DB[1107]), .B(DB[1100]), .Z(n9234) );
  AND U12313 ( .A(n1418), .B(n9235), .Z(n9233) );
  XOR U12314 ( .A(n9236), .B(n9237), .Z(n9235) );
  XOR U12315 ( .A(DB[1100]), .B(DB[1093]), .Z(n9237) );
  AND U12316 ( .A(n1422), .B(n9238), .Z(n9236) );
  XOR U12317 ( .A(n9239), .B(n9240), .Z(n9238) );
  XOR U12318 ( .A(DB[1093]), .B(DB[1086]), .Z(n9240) );
  AND U12319 ( .A(n1426), .B(n9241), .Z(n9239) );
  XOR U12320 ( .A(n9242), .B(n9243), .Z(n9241) );
  XOR U12321 ( .A(DB[1086]), .B(DB[1079]), .Z(n9243) );
  AND U12322 ( .A(n1430), .B(n9244), .Z(n9242) );
  XOR U12323 ( .A(n9245), .B(n9246), .Z(n9244) );
  XOR U12324 ( .A(DB[1079]), .B(DB[1072]), .Z(n9246) );
  AND U12325 ( .A(n1434), .B(n9247), .Z(n9245) );
  XOR U12326 ( .A(n9248), .B(n9249), .Z(n9247) );
  XOR U12327 ( .A(DB[1072]), .B(DB[1065]), .Z(n9249) );
  AND U12328 ( .A(n1438), .B(n9250), .Z(n9248) );
  XOR U12329 ( .A(n9251), .B(n9252), .Z(n9250) );
  XOR U12330 ( .A(DB[1065]), .B(DB[1058]), .Z(n9252) );
  AND U12331 ( .A(n1442), .B(n9253), .Z(n9251) );
  XOR U12332 ( .A(n9254), .B(n9255), .Z(n9253) );
  XOR U12333 ( .A(DB[1058]), .B(DB[1051]), .Z(n9255) );
  AND U12334 ( .A(n1446), .B(n9256), .Z(n9254) );
  XOR U12335 ( .A(n9257), .B(n9258), .Z(n9256) );
  XOR U12336 ( .A(DB[1051]), .B(DB[1044]), .Z(n9258) );
  AND U12337 ( .A(n1450), .B(n9259), .Z(n9257) );
  XOR U12338 ( .A(n9260), .B(n9261), .Z(n9259) );
  XOR U12339 ( .A(DB[1044]), .B(DB[1037]), .Z(n9261) );
  AND U12340 ( .A(n1454), .B(n9262), .Z(n9260) );
  XOR U12341 ( .A(n9263), .B(n9264), .Z(n9262) );
  XOR U12342 ( .A(DB[1037]), .B(DB[1030]), .Z(n9264) );
  AND U12343 ( .A(n1458), .B(n9265), .Z(n9263) );
  XOR U12344 ( .A(n9266), .B(n9267), .Z(n9265) );
  XOR U12345 ( .A(DB[1030]), .B(DB[1023]), .Z(n9267) );
  AND U12346 ( .A(n1462), .B(n9268), .Z(n9266) );
  XOR U12347 ( .A(n9269), .B(n9270), .Z(n9268) );
  XOR U12348 ( .A(DB[1023]), .B(DB[1016]), .Z(n9270) );
  AND U12349 ( .A(n1466), .B(n9271), .Z(n9269) );
  XOR U12350 ( .A(n9272), .B(n9273), .Z(n9271) );
  XOR U12351 ( .A(DB[1016]), .B(DB[1009]), .Z(n9273) );
  AND U12352 ( .A(n1470), .B(n9274), .Z(n9272) );
  XOR U12353 ( .A(n9275), .B(n9276), .Z(n9274) );
  XOR U12354 ( .A(DB[1009]), .B(DB[1002]), .Z(n9276) );
  AND U12355 ( .A(n1474), .B(n9277), .Z(n9275) );
  XOR U12356 ( .A(n9278), .B(n9279), .Z(n9277) );
  XOR U12357 ( .A(DB[995]), .B(DB[1002]), .Z(n9279) );
  AND U12358 ( .A(n1478), .B(n9280), .Z(n9278) );
  XOR U12359 ( .A(n9281), .B(n9282), .Z(n9280) );
  XOR U12360 ( .A(DB[995]), .B(DB[988]), .Z(n9282) );
  AND U12361 ( .A(n1482), .B(n9283), .Z(n9281) );
  XOR U12362 ( .A(n9284), .B(n9285), .Z(n9283) );
  XOR U12363 ( .A(DB[988]), .B(DB[981]), .Z(n9285) );
  AND U12364 ( .A(n1486), .B(n9286), .Z(n9284) );
  XOR U12365 ( .A(n9287), .B(n9288), .Z(n9286) );
  XOR U12366 ( .A(DB[981]), .B(DB[974]), .Z(n9288) );
  AND U12367 ( .A(n1490), .B(n9289), .Z(n9287) );
  XOR U12368 ( .A(n9290), .B(n9291), .Z(n9289) );
  XOR U12369 ( .A(DB[974]), .B(DB[967]), .Z(n9291) );
  AND U12370 ( .A(n1494), .B(n9292), .Z(n9290) );
  XOR U12371 ( .A(n9293), .B(n9294), .Z(n9292) );
  XOR U12372 ( .A(DB[967]), .B(DB[960]), .Z(n9294) );
  AND U12373 ( .A(n1498), .B(n9295), .Z(n9293) );
  XOR U12374 ( .A(n9296), .B(n9297), .Z(n9295) );
  XOR U12375 ( .A(DB[960]), .B(DB[953]), .Z(n9297) );
  AND U12376 ( .A(n1502), .B(n9298), .Z(n9296) );
  XOR U12377 ( .A(n9299), .B(n9300), .Z(n9298) );
  XOR U12378 ( .A(DB[953]), .B(DB[946]), .Z(n9300) );
  AND U12379 ( .A(n1506), .B(n9301), .Z(n9299) );
  XOR U12380 ( .A(n9302), .B(n9303), .Z(n9301) );
  XOR U12381 ( .A(DB[946]), .B(DB[939]), .Z(n9303) );
  AND U12382 ( .A(n1510), .B(n9304), .Z(n9302) );
  XOR U12383 ( .A(n9305), .B(n9306), .Z(n9304) );
  XOR U12384 ( .A(DB[939]), .B(DB[932]), .Z(n9306) );
  AND U12385 ( .A(n1514), .B(n9307), .Z(n9305) );
  XOR U12386 ( .A(n9308), .B(n9309), .Z(n9307) );
  XOR U12387 ( .A(DB[932]), .B(DB[925]), .Z(n9309) );
  AND U12388 ( .A(n1518), .B(n9310), .Z(n9308) );
  XOR U12389 ( .A(n9311), .B(n9312), .Z(n9310) );
  XOR U12390 ( .A(DB[925]), .B(DB[918]), .Z(n9312) );
  AND U12391 ( .A(n1522), .B(n9313), .Z(n9311) );
  XOR U12392 ( .A(n9314), .B(n9315), .Z(n9313) );
  XOR U12393 ( .A(DB[918]), .B(DB[911]), .Z(n9315) );
  AND U12394 ( .A(n1526), .B(n9316), .Z(n9314) );
  XOR U12395 ( .A(n9317), .B(n9318), .Z(n9316) );
  XOR U12396 ( .A(DB[911]), .B(DB[904]), .Z(n9318) );
  AND U12397 ( .A(n1530), .B(n9319), .Z(n9317) );
  XOR U12398 ( .A(n9320), .B(n9321), .Z(n9319) );
  XOR U12399 ( .A(DB[904]), .B(DB[897]), .Z(n9321) );
  AND U12400 ( .A(n1534), .B(n9322), .Z(n9320) );
  XOR U12401 ( .A(n9323), .B(n9324), .Z(n9322) );
  XOR U12402 ( .A(DB[897]), .B(DB[890]), .Z(n9324) );
  AND U12403 ( .A(n1538), .B(n9325), .Z(n9323) );
  XOR U12404 ( .A(n9326), .B(n9327), .Z(n9325) );
  XOR U12405 ( .A(DB[890]), .B(DB[883]), .Z(n9327) );
  AND U12406 ( .A(n1542), .B(n9328), .Z(n9326) );
  XOR U12407 ( .A(n9329), .B(n9330), .Z(n9328) );
  XOR U12408 ( .A(DB[883]), .B(DB[876]), .Z(n9330) );
  AND U12409 ( .A(n1546), .B(n9331), .Z(n9329) );
  XOR U12410 ( .A(n9332), .B(n9333), .Z(n9331) );
  XOR U12411 ( .A(DB[876]), .B(DB[869]), .Z(n9333) );
  AND U12412 ( .A(n1550), .B(n9334), .Z(n9332) );
  XOR U12413 ( .A(n9335), .B(n9336), .Z(n9334) );
  XOR U12414 ( .A(DB[869]), .B(DB[862]), .Z(n9336) );
  AND U12415 ( .A(n1554), .B(n9337), .Z(n9335) );
  XOR U12416 ( .A(n9338), .B(n9339), .Z(n9337) );
  XOR U12417 ( .A(DB[862]), .B(DB[855]), .Z(n9339) );
  AND U12418 ( .A(n1558), .B(n9340), .Z(n9338) );
  XOR U12419 ( .A(n9341), .B(n9342), .Z(n9340) );
  XOR U12420 ( .A(DB[855]), .B(DB[848]), .Z(n9342) );
  AND U12421 ( .A(n1562), .B(n9343), .Z(n9341) );
  XOR U12422 ( .A(n9344), .B(n9345), .Z(n9343) );
  XOR U12423 ( .A(DB[848]), .B(DB[841]), .Z(n9345) );
  AND U12424 ( .A(n1566), .B(n9346), .Z(n9344) );
  XOR U12425 ( .A(n9347), .B(n9348), .Z(n9346) );
  XOR U12426 ( .A(DB[841]), .B(DB[834]), .Z(n9348) );
  AND U12427 ( .A(n1570), .B(n9349), .Z(n9347) );
  XOR U12428 ( .A(n9350), .B(n9351), .Z(n9349) );
  XOR U12429 ( .A(DB[834]), .B(DB[827]), .Z(n9351) );
  AND U12430 ( .A(n1574), .B(n9352), .Z(n9350) );
  XOR U12431 ( .A(n9353), .B(n9354), .Z(n9352) );
  XOR U12432 ( .A(DB[827]), .B(DB[820]), .Z(n9354) );
  AND U12433 ( .A(n1578), .B(n9355), .Z(n9353) );
  XOR U12434 ( .A(n9356), .B(n9357), .Z(n9355) );
  XOR U12435 ( .A(DB[820]), .B(DB[813]), .Z(n9357) );
  AND U12436 ( .A(n1582), .B(n9358), .Z(n9356) );
  XOR U12437 ( .A(n9359), .B(n9360), .Z(n9358) );
  XOR U12438 ( .A(DB[813]), .B(DB[806]), .Z(n9360) );
  AND U12439 ( .A(n1586), .B(n9361), .Z(n9359) );
  XOR U12440 ( .A(n9362), .B(n9363), .Z(n9361) );
  XOR U12441 ( .A(DB[806]), .B(DB[799]), .Z(n9363) );
  AND U12442 ( .A(n1590), .B(n9364), .Z(n9362) );
  XOR U12443 ( .A(n9365), .B(n9366), .Z(n9364) );
  XOR U12444 ( .A(DB[799]), .B(DB[792]), .Z(n9366) );
  AND U12445 ( .A(n1594), .B(n9367), .Z(n9365) );
  XOR U12446 ( .A(n9368), .B(n9369), .Z(n9367) );
  XOR U12447 ( .A(DB[792]), .B(DB[785]), .Z(n9369) );
  AND U12448 ( .A(n1598), .B(n9370), .Z(n9368) );
  XOR U12449 ( .A(n9371), .B(n9372), .Z(n9370) );
  XOR U12450 ( .A(DB[785]), .B(DB[778]), .Z(n9372) );
  AND U12451 ( .A(n1602), .B(n9373), .Z(n9371) );
  XOR U12452 ( .A(n9374), .B(n9375), .Z(n9373) );
  XOR U12453 ( .A(DB[778]), .B(DB[771]), .Z(n9375) );
  AND U12454 ( .A(n1606), .B(n9376), .Z(n9374) );
  XOR U12455 ( .A(n9377), .B(n9378), .Z(n9376) );
  XOR U12456 ( .A(DB[771]), .B(DB[764]), .Z(n9378) );
  AND U12457 ( .A(n1610), .B(n9379), .Z(n9377) );
  XOR U12458 ( .A(n9380), .B(n9381), .Z(n9379) );
  XOR U12459 ( .A(DB[764]), .B(DB[757]), .Z(n9381) );
  AND U12460 ( .A(n1614), .B(n9382), .Z(n9380) );
  XOR U12461 ( .A(n9383), .B(n9384), .Z(n9382) );
  XOR U12462 ( .A(DB[757]), .B(DB[750]), .Z(n9384) );
  AND U12463 ( .A(n1618), .B(n9385), .Z(n9383) );
  XOR U12464 ( .A(n9386), .B(n9387), .Z(n9385) );
  XOR U12465 ( .A(DB[750]), .B(DB[743]), .Z(n9387) );
  AND U12466 ( .A(n1622), .B(n9388), .Z(n9386) );
  XOR U12467 ( .A(n9389), .B(n9390), .Z(n9388) );
  XOR U12468 ( .A(DB[743]), .B(DB[736]), .Z(n9390) );
  AND U12469 ( .A(n1626), .B(n9391), .Z(n9389) );
  XOR U12470 ( .A(n9392), .B(n9393), .Z(n9391) );
  XOR U12471 ( .A(DB[736]), .B(DB[729]), .Z(n9393) );
  AND U12472 ( .A(n1630), .B(n9394), .Z(n9392) );
  XOR U12473 ( .A(n9395), .B(n9396), .Z(n9394) );
  XOR U12474 ( .A(DB[729]), .B(DB[722]), .Z(n9396) );
  AND U12475 ( .A(n1634), .B(n9397), .Z(n9395) );
  XOR U12476 ( .A(n9398), .B(n9399), .Z(n9397) );
  XOR U12477 ( .A(DB[722]), .B(DB[715]), .Z(n9399) );
  AND U12478 ( .A(n1638), .B(n9400), .Z(n9398) );
  XOR U12479 ( .A(n9401), .B(n9402), .Z(n9400) );
  XOR U12480 ( .A(DB[715]), .B(DB[708]), .Z(n9402) );
  AND U12481 ( .A(n1642), .B(n9403), .Z(n9401) );
  XOR U12482 ( .A(n9404), .B(n9405), .Z(n9403) );
  XOR U12483 ( .A(DB[708]), .B(DB[701]), .Z(n9405) );
  AND U12484 ( .A(n1646), .B(n9406), .Z(n9404) );
  XOR U12485 ( .A(n9407), .B(n9408), .Z(n9406) );
  XOR U12486 ( .A(DB[701]), .B(DB[694]), .Z(n9408) );
  AND U12487 ( .A(n1650), .B(n9409), .Z(n9407) );
  XOR U12488 ( .A(n9410), .B(n9411), .Z(n9409) );
  XOR U12489 ( .A(DB[694]), .B(DB[687]), .Z(n9411) );
  AND U12490 ( .A(n1654), .B(n9412), .Z(n9410) );
  XOR U12491 ( .A(n9413), .B(n9414), .Z(n9412) );
  XOR U12492 ( .A(DB[687]), .B(DB[680]), .Z(n9414) );
  AND U12493 ( .A(n1658), .B(n9415), .Z(n9413) );
  XOR U12494 ( .A(n9416), .B(n9417), .Z(n9415) );
  XOR U12495 ( .A(DB[680]), .B(DB[673]), .Z(n9417) );
  AND U12496 ( .A(n1662), .B(n9418), .Z(n9416) );
  XOR U12497 ( .A(n9419), .B(n9420), .Z(n9418) );
  XOR U12498 ( .A(DB[673]), .B(DB[666]), .Z(n9420) );
  AND U12499 ( .A(n1666), .B(n9421), .Z(n9419) );
  XOR U12500 ( .A(n9422), .B(n9423), .Z(n9421) );
  XOR U12501 ( .A(DB[666]), .B(DB[659]), .Z(n9423) );
  AND U12502 ( .A(n1670), .B(n9424), .Z(n9422) );
  XOR U12503 ( .A(n9425), .B(n9426), .Z(n9424) );
  XOR U12504 ( .A(DB[659]), .B(DB[652]), .Z(n9426) );
  AND U12505 ( .A(n1674), .B(n9427), .Z(n9425) );
  XOR U12506 ( .A(n9428), .B(n9429), .Z(n9427) );
  XOR U12507 ( .A(DB[652]), .B(DB[645]), .Z(n9429) );
  AND U12508 ( .A(n1678), .B(n9430), .Z(n9428) );
  XOR U12509 ( .A(n9431), .B(n9432), .Z(n9430) );
  XOR U12510 ( .A(DB[645]), .B(DB[638]), .Z(n9432) );
  AND U12511 ( .A(n1682), .B(n9433), .Z(n9431) );
  XOR U12512 ( .A(n9434), .B(n9435), .Z(n9433) );
  XOR U12513 ( .A(DB[638]), .B(DB[631]), .Z(n9435) );
  AND U12514 ( .A(n1686), .B(n9436), .Z(n9434) );
  XOR U12515 ( .A(n9437), .B(n9438), .Z(n9436) );
  XOR U12516 ( .A(DB[631]), .B(DB[624]), .Z(n9438) );
  AND U12517 ( .A(n1690), .B(n9439), .Z(n9437) );
  XOR U12518 ( .A(n9440), .B(n9441), .Z(n9439) );
  XOR U12519 ( .A(DB[624]), .B(DB[617]), .Z(n9441) );
  AND U12520 ( .A(n1694), .B(n9442), .Z(n9440) );
  XOR U12521 ( .A(n9443), .B(n9444), .Z(n9442) );
  XOR U12522 ( .A(DB[617]), .B(DB[610]), .Z(n9444) );
  AND U12523 ( .A(n1698), .B(n9445), .Z(n9443) );
  XOR U12524 ( .A(n9446), .B(n9447), .Z(n9445) );
  XOR U12525 ( .A(DB[610]), .B(DB[603]), .Z(n9447) );
  AND U12526 ( .A(n1702), .B(n9448), .Z(n9446) );
  XOR U12527 ( .A(n9449), .B(n9450), .Z(n9448) );
  XOR U12528 ( .A(DB[603]), .B(DB[596]), .Z(n9450) );
  AND U12529 ( .A(n1706), .B(n9451), .Z(n9449) );
  XOR U12530 ( .A(n9452), .B(n9453), .Z(n9451) );
  XOR U12531 ( .A(DB[596]), .B(DB[589]), .Z(n9453) );
  AND U12532 ( .A(n1710), .B(n9454), .Z(n9452) );
  XOR U12533 ( .A(n9455), .B(n9456), .Z(n9454) );
  XOR U12534 ( .A(DB[589]), .B(DB[582]), .Z(n9456) );
  AND U12535 ( .A(n1714), .B(n9457), .Z(n9455) );
  XOR U12536 ( .A(n9458), .B(n9459), .Z(n9457) );
  XOR U12537 ( .A(DB[582]), .B(DB[575]), .Z(n9459) );
  AND U12538 ( .A(n1718), .B(n9460), .Z(n9458) );
  XOR U12539 ( .A(n9461), .B(n9462), .Z(n9460) );
  XOR U12540 ( .A(DB[575]), .B(DB[568]), .Z(n9462) );
  AND U12541 ( .A(n1722), .B(n9463), .Z(n9461) );
  XOR U12542 ( .A(n9464), .B(n9465), .Z(n9463) );
  XOR U12543 ( .A(DB[568]), .B(DB[561]), .Z(n9465) );
  AND U12544 ( .A(n1726), .B(n9466), .Z(n9464) );
  XOR U12545 ( .A(n9467), .B(n9468), .Z(n9466) );
  XOR U12546 ( .A(DB[561]), .B(DB[554]), .Z(n9468) );
  AND U12547 ( .A(n1730), .B(n9469), .Z(n9467) );
  XOR U12548 ( .A(n9470), .B(n9471), .Z(n9469) );
  XOR U12549 ( .A(DB[554]), .B(DB[547]), .Z(n9471) );
  AND U12550 ( .A(n1734), .B(n9472), .Z(n9470) );
  XOR U12551 ( .A(n9473), .B(n9474), .Z(n9472) );
  XOR U12552 ( .A(DB[547]), .B(DB[540]), .Z(n9474) );
  AND U12553 ( .A(n1738), .B(n9475), .Z(n9473) );
  XOR U12554 ( .A(n9476), .B(n9477), .Z(n9475) );
  XOR U12555 ( .A(DB[540]), .B(DB[533]), .Z(n9477) );
  AND U12556 ( .A(n1742), .B(n9478), .Z(n9476) );
  XOR U12557 ( .A(n9479), .B(n9480), .Z(n9478) );
  XOR U12558 ( .A(DB[533]), .B(DB[526]), .Z(n9480) );
  AND U12559 ( .A(n1746), .B(n9481), .Z(n9479) );
  XOR U12560 ( .A(n9482), .B(n9483), .Z(n9481) );
  XOR U12561 ( .A(DB[526]), .B(DB[519]), .Z(n9483) );
  AND U12562 ( .A(n1750), .B(n9484), .Z(n9482) );
  XOR U12563 ( .A(n9485), .B(n9486), .Z(n9484) );
  XOR U12564 ( .A(DB[519]), .B(DB[512]), .Z(n9486) );
  AND U12565 ( .A(n1754), .B(n9487), .Z(n9485) );
  XOR U12566 ( .A(n9488), .B(n9489), .Z(n9487) );
  XOR U12567 ( .A(DB[512]), .B(DB[505]), .Z(n9489) );
  AND U12568 ( .A(n1758), .B(n9490), .Z(n9488) );
  XOR U12569 ( .A(n9491), .B(n9492), .Z(n9490) );
  XOR U12570 ( .A(DB[505]), .B(DB[498]), .Z(n9492) );
  AND U12571 ( .A(n1762), .B(n9493), .Z(n9491) );
  XOR U12572 ( .A(n9494), .B(n9495), .Z(n9493) );
  XOR U12573 ( .A(DB[498]), .B(DB[491]), .Z(n9495) );
  AND U12574 ( .A(n1766), .B(n9496), .Z(n9494) );
  XOR U12575 ( .A(n9497), .B(n9498), .Z(n9496) );
  XOR U12576 ( .A(DB[491]), .B(DB[484]), .Z(n9498) );
  AND U12577 ( .A(n1770), .B(n9499), .Z(n9497) );
  XOR U12578 ( .A(n9500), .B(n9501), .Z(n9499) );
  XOR U12579 ( .A(DB[484]), .B(DB[477]), .Z(n9501) );
  AND U12580 ( .A(n1774), .B(n9502), .Z(n9500) );
  XOR U12581 ( .A(n9503), .B(n9504), .Z(n9502) );
  XOR U12582 ( .A(DB[477]), .B(DB[470]), .Z(n9504) );
  AND U12583 ( .A(n1778), .B(n9505), .Z(n9503) );
  XOR U12584 ( .A(n9506), .B(n9507), .Z(n9505) );
  XOR U12585 ( .A(DB[470]), .B(DB[463]), .Z(n9507) );
  AND U12586 ( .A(n1782), .B(n9508), .Z(n9506) );
  XOR U12587 ( .A(n9509), .B(n9510), .Z(n9508) );
  XOR U12588 ( .A(DB[463]), .B(DB[456]), .Z(n9510) );
  AND U12589 ( .A(n1786), .B(n9511), .Z(n9509) );
  XOR U12590 ( .A(n9512), .B(n9513), .Z(n9511) );
  XOR U12591 ( .A(DB[456]), .B(DB[449]), .Z(n9513) );
  AND U12592 ( .A(n1790), .B(n9514), .Z(n9512) );
  XOR U12593 ( .A(n9515), .B(n9516), .Z(n9514) );
  XOR U12594 ( .A(DB[449]), .B(DB[442]), .Z(n9516) );
  AND U12595 ( .A(n1794), .B(n9517), .Z(n9515) );
  XOR U12596 ( .A(n9518), .B(n9519), .Z(n9517) );
  XOR U12597 ( .A(DB[442]), .B(DB[435]), .Z(n9519) );
  AND U12598 ( .A(n1798), .B(n9520), .Z(n9518) );
  XOR U12599 ( .A(n9521), .B(n9522), .Z(n9520) );
  XOR U12600 ( .A(DB[435]), .B(DB[428]), .Z(n9522) );
  AND U12601 ( .A(n1802), .B(n9523), .Z(n9521) );
  XOR U12602 ( .A(n9524), .B(n9525), .Z(n9523) );
  XOR U12603 ( .A(DB[428]), .B(DB[421]), .Z(n9525) );
  AND U12604 ( .A(n1806), .B(n9526), .Z(n9524) );
  XOR U12605 ( .A(n9527), .B(n9528), .Z(n9526) );
  XOR U12606 ( .A(DB[421]), .B(DB[414]), .Z(n9528) );
  AND U12607 ( .A(n1810), .B(n9529), .Z(n9527) );
  XOR U12608 ( .A(n9530), .B(n9531), .Z(n9529) );
  XOR U12609 ( .A(DB[414]), .B(DB[407]), .Z(n9531) );
  AND U12610 ( .A(n1814), .B(n9532), .Z(n9530) );
  XOR U12611 ( .A(n9533), .B(n9534), .Z(n9532) );
  XOR U12612 ( .A(DB[407]), .B(DB[400]), .Z(n9534) );
  AND U12613 ( .A(n1818), .B(n9535), .Z(n9533) );
  XOR U12614 ( .A(n9536), .B(n9537), .Z(n9535) );
  XOR U12615 ( .A(DB[400]), .B(DB[393]), .Z(n9537) );
  AND U12616 ( .A(n1822), .B(n9538), .Z(n9536) );
  XOR U12617 ( .A(n9539), .B(n9540), .Z(n9538) );
  XOR U12618 ( .A(DB[393]), .B(DB[386]), .Z(n9540) );
  AND U12619 ( .A(n1826), .B(n9541), .Z(n9539) );
  XOR U12620 ( .A(n9542), .B(n9543), .Z(n9541) );
  XOR U12621 ( .A(DB[386]), .B(DB[379]), .Z(n9543) );
  AND U12622 ( .A(n1830), .B(n9544), .Z(n9542) );
  XOR U12623 ( .A(n9545), .B(n9546), .Z(n9544) );
  XOR U12624 ( .A(DB[379]), .B(DB[372]), .Z(n9546) );
  AND U12625 ( .A(n1834), .B(n9547), .Z(n9545) );
  XOR U12626 ( .A(n9548), .B(n9549), .Z(n9547) );
  XOR U12627 ( .A(DB[372]), .B(DB[365]), .Z(n9549) );
  AND U12628 ( .A(n1838), .B(n9550), .Z(n9548) );
  XOR U12629 ( .A(n9551), .B(n9552), .Z(n9550) );
  XOR U12630 ( .A(DB[365]), .B(DB[358]), .Z(n9552) );
  AND U12631 ( .A(n1842), .B(n9553), .Z(n9551) );
  XOR U12632 ( .A(n9554), .B(n9555), .Z(n9553) );
  XOR U12633 ( .A(DB[358]), .B(DB[351]), .Z(n9555) );
  AND U12634 ( .A(n1846), .B(n9556), .Z(n9554) );
  XOR U12635 ( .A(n9557), .B(n9558), .Z(n9556) );
  XOR U12636 ( .A(DB[351]), .B(DB[344]), .Z(n9558) );
  AND U12637 ( .A(n1850), .B(n9559), .Z(n9557) );
  XOR U12638 ( .A(n9560), .B(n9561), .Z(n9559) );
  XOR U12639 ( .A(DB[344]), .B(DB[337]), .Z(n9561) );
  AND U12640 ( .A(n1854), .B(n9562), .Z(n9560) );
  XOR U12641 ( .A(n9563), .B(n9564), .Z(n9562) );
  XOR U12642 ( .A(DB[337]), .B(DB[330]), .Z(n9564) );
  AND U12643 ( .A(n1858), .B(n9565), .Z(n9563) );
  XOR U12644 ( .A(n9566), .B(n9567), .Z(n9565) );
  XOR U12645 ( .A(DB[330]), .B(DB[323]), .Z(n9567) );
  AND U12646 ( .A(n1862), .B(n9568), .Z(n9566) );
  XOR U12647 ( .A(n9569), .B(n9570), .Z(n9568) );
  XOR U12648 ( .A(DB[323]), .B(DB[316]), .Z(n9570) );
  AND U12649 ( .A(n1866), .B(n9571), .Z(n9569) );
  XOR U12650 ( .A(n9572), .B(n9573), .Z(n9571) );
  XOR U12651 ( .A(DB[316]), .B(DB[309]), .Z(n9573) );
  AND U12652 ( .A(n1870), .B(n9574), .Z(n9572) );
  XOR U12653 ( .A(n9575), .B(n9576), .Z(n9574) );
  XOR U12654 ( .A(DB[309]), .B(DB[302]), .Z(n9576) );
  AND U12655 ( .A(n1874), .B(n9577), .Z(n9575) );
  XOR U12656 ( .A(n9578), .B(n9579), .Z(n9577) );
  XOR U12657 ( .A(DB[302]), .B(DB[295]), .Z(n9579) );
  AND U12658 ( .A(n1878), .B(n9580), .Z(n9578) );
  XOR U12659 ( .A(n9581), .B(n9582), .Z(n9580) );
  XOR U12660 ( .A(DB[295]), .B(DB[288]), .Z(n9582) );
  AND U12661 ( .A(n1882), .B(n9583), .Z(n9581) );
  XOR U12662 ( .A(n9584), .B(n9585), .Z(n9583) );
  XOR U12663 ( .A(DB[288]), .B(DB[281]), .Z(n9585) );
  AND U12664 ( .A(n1886), .B(n9586), .Z(n9584) );
  XOR U12665 ( .A(n9587), .B(n9588), .Z(n9586) );
  XOR U12666 ( .A(DB[281]), .B(DB[274]), .Z(n9588) );
  AND U12667 ( .A(n1890), .B(n9589), .Z(n9587) );
  XOR U12668 ( .A(n9590), .B(n9591), .Z(n9589) );
  XOR U12669 ( .A(DB[274]), .B(DB[267]), .Z(n9591) );
  AND U12670 ( .A(n1894), .B(n9592), .Z(n9590) );
  XOR U12671 ( .A(n9593), .B(n9594), .Z(n9592) );
  XOR U12672 ( .A(DB[267]), .B(DB[260]), .Z(n9594) );
  AND U12673 ( .A(n1898), .B(n9595), .Z(n9593) );
  XOR U12674 ( .A(n9596), .B(n9597), .Z(n9595) );
  XOR U12675 ( .A(DB[260]), .B(DB[253]), .Z(n9597) );
  AND U12676 ( .A(n1902), .B(n9598), .Z(n9596) );
  XOR U12677 ( .A(n9599), .B(n9600), .Z(n9598) );
  XOR U12678 ( .A(DB[253]), .B(DB[246]), .Z(n9600) );
  AND U12679 ( .A(n1906), .B(n9601), .Z(n9599) );
  XOR U12680 ( .A(n9602), .B(n9603), .Z(n9601) );
  XOR U12681 ( .A(DB[246]), .B(DB[239]), .Z(n9603) );
  AND U12682 ( .A(n1910), .B(n9604), .Z(n9602) );
  XOR U12683 ( .A(n9605), .B(n9606), .Z(n9604) );
  XOR U12684 ( .A(DB[239]), .B(DB[232]), .Z(n9606) );
  AND U12685 ( .A(n1914), .B(n9607), .Z(n9605) );
  XOR U12686 ( .A(n9608), .B(n9609), .Z(n9607) );
  XOR U12687 ( .A(DB[232]), .B(DB[225]), .Z(n9609) );
  AND U12688 ( .A(n1918), .B(n9610), .Z(n9608) );
  XOR U12689 ( .A(n9611), .B(n9612), .Z(n9610) );
  XOR U12690 ( .A(DB[225]), .B(DB[218]), .Z(n9612) );
  AND U12691 ( .A(n1922), .B(n9613), .Z(n9611) );
  XOR U12692 ( .A(n9614), .B(n9615), .Z(n9613) );
  XOR U12693 ( .A(DB[218]), .B(DB[211]), .Z(n9615) );
  AND U12694 ( .A(n1926), .B(n9616), .Z(n9614) );
  XOR U12695 ( .A(n9617), .B(n9618), .Z(n9616) );
  XOR U12696 ( .A(DB[211]), .B(DB[204]), .Z(n9618) );
  AND U12697 ( .A(n1930), .B(n9619), .Z(n9617) );
  XOR U12698 ( .A(n9620), .B(n9621), .Z(n9619) );
  XOR U12699 ( .A(DB[204]), .B(DB[197]), .Z(n9621) );
  AND U12700 ( .A(n1934), .B(n9622), .Z(n9620) );
  XOR U12701 ( .A(n9623), .B(n9624), .Z(n9622) );
  XOR U12702 ( .A(DB[197]), .B(DB[190]), .Z(n9624) );
  AND U12703 ( .A(n1938), .B(n9625), .Z(n9623) );
  XOR U12704 ( .A(n9626), .B(n9627), .Z(n9625) );
  XOR U12705 ( .A(DB[190]), .B(DB[183]), .Z(n9627) );
  AND U12706 ( .A(n1942), .B(n9628), .Z(n9626) );
  XOR U12707 ( .A(n9629), .B(n9630), .Z(n9628) );
  XOR U12708 ( .A(DB[183]), .B(DB[176]), .Z(n9630) );
  AND U12709 ( .A(n1946), .B(n9631), .Z(n9629) );
  XOR U12710 ( .A(n9632), .B(n9633), .Z(n9631) );
  XOR U12711 ( .A(DB[176]), .B(DB[169]), .Z(n9633) );
  AND U12712 ( .A(n1950), .B(n9634), .Z(n9632) );
  XOR U12713 ( .A(n9635), .B(n9636), .Z(n9634) );
  XOR U12714 ( .A(DB[169]), .B(DB[162]), .Z(n9636) );
  AND U12715 ( .A(n1954), .B(n9637), .Z(n9635) );
  XOR U12716 ( .A(n9638), .B(n9639), .Z(n9637) );
  XOR U12717 ( .A(DB[162]), .B(DB[155]), .Z(n9639) );
  AND U12718 ( .A(n1958), .B(n9640), .Z(n9638) );
  XOR U12719 ( .A(n9641), .B(n9642), .Z(n9640) );
  XOR U12720 ( .A(DB[155]), .B(DB[148]), .Z(n9642) );
  AND U12721 ( .A(n1962), .B(n9643), .Z(n9641) );
  XOR U12722 ( .A(n9644), .B(n9645), .Z(n9643) );
  XOR U12723 ( .A(DB[148]), .B(DB[141]), .Z(n9645) );
  AND U12724 ( .A(n1966), .B(n9646), .Z(n9644) );
  XOR U12725 ( .A(n9647), .B(n9648), .Z(n9646) );
  XOR U12726 ( .A(DB[141]), .B(DB[134]), .Z(n9648) );
  AND U12727 ( .A(n1970), .B(n9649), .Z(n9647) );
  XOR U12728 ( .A(n9650), .B(n9651), .Z(n9649) );
  XOR U12729 ( .A(DB[134]), .B(DB[127]), .Z(n9651) );
  AND U12730 ( .A(n1974), .B(n9652), .Z(n9650) );
  XOR U12731 ( .A(n9653), .B(n9654), .Z(n9652) );
  XOR U12732 ( .A(DB[127]), .B(DB[120]), .Z(n9654) );
  AND U12733 ( .A(n1978), .B(n9655), .Z(n9653) );
  XOR U12734 ( .A(n9656), .B(n9657), .Z(n9655) );
  XOR U12735 ( .A(DB[120]), .B(DB[113]), .Z(n9657) );
  AND U12736 ( .A(n1982), .B(n9658), .Z(n9656) );
  XOR U12737 ( .A(n9659), .B(n9660), .Z(n9658) );
  XOR U12738 ( .A(DB[113]), .B(DB[106]), .Z(n9660) );
  AND U12739 ( .A(n1986), .B(n9661), .Z(n9659) );
  XOR U12740 ( .A(n9662), .B(n9663), .Z(n9661) );
  XOR U12741 ( .A(DB[99]), .B(DB[106]), .Z(n9663) );
  AND U12742 ( .A(n1990), .B(n9664), .Z(n9662) );
  XOR U12743 ( .A(n9665), .B(n9666), .Z(n9664) );
  XOR U12744 ( .A(DB[99]), .B(DB[92]), .Z(n9666) );
  AND U12745 ( .A(n1994), .B(n9667), .Z(n9665) );
  XOR U12746 ( .A(n9668), .B(n9669), .Z(n9667) );
  XOR U12747 ( .A(DB[92]), .B(DB[85]), .Z(n9669) );
  AND U12748 ( .A(n1998), .B(n9670), .Z(n9668) );
  XOR U12749 ( .A(n9671), .B(n9672), .Z(n9670) );
  XOR U12750 ( .A(DB[85]), .B(DB[78]), .Z(n9672) );
  AND U12751 ( .A(n2002), .B(n9673), .Z(n9671) );
  XOR U12752 ( .A(n9674), .B(n9675), .Z(n9673) );
  XOR U12753 ( .A(DB[78]), .B(DB[71]), .Z(n9675) );
  AND U12754 ( .A(n2006), .B(n9676), .Z(n9674) );
  XOR U12755 ( .A(n9677), .B(n9678), .Z(n9676) );
  XOR U12756 ( .A(DB[71]), .B(DB[64]), .Z(n9678) );
  AND U12757 ( .A(n2010), .B(n9679), .Z(n9677) );
  XOR U12758 ( .A(n9680), .B(n9681), .Z(n9679) );
  XOR U12759 ( .A(DB[64]), .B(DB[57]), .Z(n9681) );
  AND U12760 ( .A(n2014), .B(n9682), .Z(n9680) );
  XOR U12761 ( .A(n9683), .B(n9684), .Z(n9682) );
  XOR U12762 ( .A(DB[57]), .B(DB[50]), .Z(n9684) );
  AND U12763 ( .A(n2018), .B(n9685), .Z(n9683) );
  XOR U12764 ( .A(n9686), .B(n9687), .Z(n9685) );
  XOR U12765 ( .A(DB[50]), .B(DB[43]), .Z(n9687) );
  AND U12766 ( .A(n2022), .B(n9688), .Z(n9686) );
  XOR U12767 ( .A(n9689), .B(n9690), .Z(n9688) );
  XOR U12768 ( .A(DB[43]), .B(DB[36]), .Z(n9690) );
  AND U12769 ( .A(n2026), .B(n9691), .Z(n9689) );
  XOR U12770 ( .A(n9692), .B(n9693), .Z(n9691) );
  XOR U12771 ( .A(DB[36]), .B(DB[29]), .Z(n9693) );
  AND U12772 ( .A(n2030), .B(n9694), .Z(n9692) );
  XOR U12773 ( .A(n9695), .B(n9696), .Z(n9694) );
  XOR U12774 ( .A(DB[29]), .B(DB[22]), .Z(n9696) );
  AND U12775 ( .A(n2034), .B(n9697), .Z(n9695) );
  XOR U12776 ( .A(n9698), .B(n9699), .Z(n9697) );
  XOR U12777 ( .A(DB[22]), .B(DB[15]), .Z(n9699) );
  AND U12778 ( .A(n2038), .B(n9700), .Z(n9698) );
  XOR U12779 ( .A(n9701), .B(n9702), .Z(n9700) );
  XOR U12780 ( .A(DB[8]), .B(DB[15]), .Z(n9702) );
  AND U12781 ( .A(n2042), .B(n9703), .Z(n9701) );
  XOR U12782 ( .A(DB[8]), .B(DB[1]), .Z(n9703) );
  XOR U12783 ( .A(DB[3577]), .B(n9704), .Z(min_val_out[0]) );
  AND U12784 ( .A(n2), .B(n9705), .Z(n9704) );
  XOR U12785 ( .A(n9706), .B(n9707), .Z(n9705) );
  XOR U12786 ( .A(DB[3577]), .B(DB[3570]), .Z(n9707) );
  AND U12787 ( .A(n6), .B(n9708), .Z(n9706) );
  XOR U12788 ( .A(n9709), .B(n9710), .Z(n9708) );
  XOR U12789 ( .A(DB[3570]), .B(DB[3563]), .Z(n9710) );
  AND U12790 ( .A(n10), .B(n9711), .Z(n9709) );
  XOR U12791 ( .A(n9712), .B(n9713), .Z(n9711) );
  XOR U12792 ( .A(DB[3563]), .B(DB[3556]), .Z(n9713) );
  AND U12793 ( .A(n14), .B(n9714), .Z(n9712) );
  XOR U12794 ( .A(n9715), .B(n9716), .Z(n9714) );
  XOR U12795 ( .A(DB[3556]), .B(DB[3549]), .Z(n9716) );
  AND U12796 ( .A(n18), .B(n9717), .Z(n9715) );
  XOR U12797 ( .A(n9718), .B(n9719), .Z(n9717) );
  XOR U12798 ( .A(DB[3549]), .B(DB[3542]), .Z(n9719) );
  AND U12799 ( .A(n22), .B(n9720), .Z(n9718) );
  XOR U12800 ( .A(n9721), .B(n9722), .Z(n9720) );
  XOR U12801 ( .A(DB[3542]), .B(DB[3535]), .Z(n9722) );
  AND U12802 ( .A(n26), .B(n9723), .Z(n9721) );
  XOR U12803 ( .A(n9724), .B(n9725), .Z(n9723) );
  XOR U12804 ( .A(DB[3535]), .B(DB[3528]), .Z(n9725) );
  AND U12805 ( .A(n30), .B(n9726), .Z(n9724) );
  XOR U12806 ( .A(n9727), .B(n9728), .Z(n9726) );
  XOR U12807 ( .A(DB[3528]), .B(DB[3521]), .Z(n9728) );
  AND U12808 ( .A(n34), .B(n9729), .Z(n9727) );
  XOR U12809 ( .A(n9730), .B(n9731), .Z(n9729) );
  XOR U12810 ( .A(DB[3521]), .B(DB[3514]), .Z(n9731) );
  AND U12811 ( .A(n38), .B(n9732), .Z(n9730) );
  XOR U12812 ( .A(n9733), .B(n9734), .Z(n9732) );
  XOR U12813 ( .A(DB[3514]), .B(DB[3507]), .Z(n9734) );
  AND U12814 ( .A(n42), .B(n9735), .Z(n9733) );
  XOR U12815 ( .A(n9736), .B(n9737), .Z(n9735) );
  XOR U12816 ( .A(DB[3507]), .B(DB[3500]), .Z(n9737) );
  AND U12817 ( .A(n46), .B(n9738), .Z(n9736) );
  XOR U12818 ( .A(n9739), .B(n9740), .Z(n9738) );
  XOR U12819 ( .A(DB[3500]), .B(DB[3493]), .Z(n9740) );
  AND U12820 ( .A(n50), .B(n9741), .Z(n9739) );
  XOR U12821 ( .A(n9742), .B(n9743), .Z(n9741) );
  XOR U12822 ( .A(DB[3493]), .B(DB[3486]), .Z(n9743) );
  AND U12823 ( .A(n54), .B(n9744), .Z(n9742) );
  XOR U12824 ( .A(n9745), .B(n9746), .Z(n9744) );
  XOR U12825 ( .A(DB[3486]), .B(DB[3479]), .Z(n9746) );
  AND U12826 ( .A(n58), .B(n9747), .Z(n9745) );
  XOR U12827 ( .A(n9748), .B(n9749), .Z(n9747) );
  XOR U12828 ( .A(DB[3479]), .B(DB[3472]), .Z(n9749) );
  AND U12829 ( .A(n62), .B(n9750), .Z(n9748) );
  XOR U12830 ( .A(n9751), .B(n9752), .Z(n9750) );
  XOR U12831 ( .A(DB[3472]), .B(DB[3465]), .Z(n9752) );
  AND U12832 ( .A(n66), .B(n9753), .Z(n9751) );
  XOR U12833 ( .A(n9754), .B(n9755), .Z(n9753) );
  XOR U12834 ( .A(DB[3465]), .B(DB[3458]), .Z(n9755) );
  AND U12835 ( .A(n70), .B(n9756), .Z(n9754) );
  XOR U12836 ( .A(n9757), .B(n9758), .Z(n9756) );
  XOR U12837 ( .A(DB[3458]), .B(DB[3451]), .Z(n9758) );
  AND U12838 ( .A(n74), .B(n9759), .Z(n9757) );
  XOR U12839 ( .A(n9760), .B(n9761), .Z(n9759) );
  XOR U12840 ( .A(DB[3451]), .B(DB[3444]), .Z(n9761) );
  AND U12841 ( .A(n78), .B(n9762), .Z(n9760) );
  XOR U12842 ( .A(n9763), .B(n9764), .Z(n9762) );
  XOR U12843 ( .A(DB[3444]), .B(DB[3437]), .Z(n9764) );
  AND U12844 ( .A(n82), .B(n9765), .Z(n9763) );
  XOR U12845 ( .A(n9766), .B(n9767), .Z(n9765) );
  XOR U12846 ( .A(DB[3437]), .B(DB[3430]), .Z(n9767) );
  AND U12847 ( .A(n86), .B(n9768), .Z(n9766) );
  XOR U12848 ( .A(n9769), .B(n9770), .Z(n9768) );
  XOR U12849 ( .A(DB[3430]), .B(DB[3423]), .Z(n9770) );
  AND U12850 ( .A(n90), .B(n9771), .Z(n9769) );
  XOR U12851 ( .A(n9772), .B(n9773), .Z(n9771) );
  XOR U12852 ( .A(DB[3423]), .B(DB[3416]), .Z(n9773) );
  AND U12853 ( .A(n94), .B(n9774), .Z(n9772) );
  XOR U12854 ( .A(n9775), .B(n9776), .Z(n9774) );
  XOR U12855 ( .A(DB[3416]), .B(DB[3409]), .Z(n9776) );
  AND U12856 ( .A(n98), .B(n9777), .Z(n9775) );
  XOR U12857 ( .A(n9778), .B(n9779), .Z(n9777) );
  XOR U12858 ( .A(DB[3409]), .B(DB[3402]), .Z(n9779) );
  AND U12859 ( .A(n102), .B(n9780), .Z(n9778) );
  XOR U12860 ( .A(n9781), .B(n9782), .Z(n9780) );
  XOR U12861 ( .A(DB[3402]), .B(DB[3395]), .Z(n9782) );
  AND U12862 ( .A(n106), .B(n9783), .Z(n9781) );
  XOR U12863 ( .A(n9784), .B(n9785), .Z(n9783) );
  XOR U12864 ( .A(DB[3395]), .B(DB[3388]), .Z(n9785) );
  AND U12865 ( .A(n110), .B(n9786), .Z(n9784) );
  XOR U12866 ( .A(n9787), .B(n9788), .Z(n9786) );
  XOR U12867 ( .A(DB[3388]), .B(DB[3381]), .Z(n9788) );
  AND U12868 ( .A(n114), .B(n9789), .Z(n9787) );
  XOR U12869 ( .A(n9790), .B(n9791), .Z(n9789) );
  XOR U12870 ( .A(DB[3381]), .B(DB[3374]), .Z(n9791) );
  AND U12871 ( .A(n118), .B(n9792), .Z(n9790) );
  XOR U12872 ( .A(n9793), .B(n9794), .Z(n9792) );
  XOR U12873 ( .A(DB[3374]), .B(DB[3367]), .Z(n9794) );
  AND U12874 ( .A(n122), .B(n9795), .Z(n9793) );
  XOR U12875 ( .A(n9796), .B(n9797), .Z(n9795) );
  XOR U12876 ( .A(DB[3367]), .B(DB[3360]), .Z(n9797) );
  AND U12877 ( .A(n126), .B(n9798), .Z(n9796) );
  XOR U12878 ( .A(n9799), .B(n9800), .Z(n9798) );
  XOR U12879 ( .A(DB[3360]), .B(DB[3353]), .Z(n9800) );
  AND U12880 ( .A(n130), .B(n9801), .Z(n9799) );
  XOR U12881 ( .A(n9802), .B(n9803), .Z(n9801) );
  XOR U12882 ( .A(DB[3353]), .B(DB[3346]), .Z(n9803) );
  AND U12883 ( .A(n134), .B(n9804), .Z(n9802) );
  XOR U12884 ( .A(n9805), .B(n9806), .Z(n9804) );
  XOR U12885 ( .A(DB[3346]), .B(DB[3339]), .Z(n9806) );
  AND U12886 ( .A(n138), .B(n9807), .Z(n9805) );
  XOR U12887 ( .A(n9808), .B(n9809), .Z(n9807) );
  XOR U12888 ( .A(DB[3339]), .B(DB[3332]), .Z(n9809) );
  AND U12889 ( .A(n142), .B(n9810), .Z(n9808) );
  XOR U12890 ( .A(n9811), .B(n9812), .Z(n9810) );
  XOR U12891 ( .A(DB[3332]), .B(DB[3325]), .Z(n9812) );
  AND U12892 ( .A(n146), .B(n9813), .Z(n9811) );
  XOR U12893 ( .A(n9814), .B(n9815), .Z(n9813) );
  XOR U12894 ( .A(DB[3325]), .B(DB[3318]), .Z(n9815) );
  AND U12895 ( .A(n150), .B(n9816), .Z(n9814) );
  XOR U12896 ( .A(n9817), .B(n9818), .Z(n9816) );
  XOR U12897 ( .A(DB[3318]), .B(DB[3311]), .Z(n9818) );
  AND U12898 ( .A(n154), .B(n9819), .Z(n9817) );
  XOR U12899 ( .A(n9820), .B(n9821), .Z(n9819) );
  XOR U12900 ( .A(DB[3311]), .B(DB[3304]), .Z(n9821) );
  AND U12901 ( .A(n158), .B(n9822), .Z(n9820) );
  XOR U12902 ( .A(n9823), .B(n9824), .Z(n9822) );
  XOR U12903 ( .A(DB[3304]), .B(DB[3297]), .Z(n9824) );
  AND U12904 ( .A(n162), .B(n9825), .Z(n9823) );
  XOR U12905 ( .A(n9826), .B(n9827), .Z(n9825) );
  XOR U12906 ( .A(DB[3297]), .B(DB[3290]), .Z(n9827) );
  AND U12907 ( .A(n166), .B(n9828), .Z(n9826) );
  XOR U12908 ( .A(n9829), .B(n9830), .Z(n9828) );
  XOR U12909 ( .A(DB[3290]), .B(DB[3283]), .Z(n9830) );
  AND U12910 ( .A(n170), .B(n9831), .Z(n9829) );
  XOR U12911 ( .A(n9832), .B(n9833), .Z(n9831) );
  XOR U12912 ( .A(DB[3283]), .B(DB[3276]), .Z(n9833) );
  AND U12913 ( .A(n174), .B(n9834), .Z(n9832) );
  XOR U12914 ( .A(n9835), .B(n9836), .Z(n9834) );
  XOR U12915 ( .A(DB[3276]), .B(DB[3269]), .Z(n9836) );
  AND U12916 ( .A(n178), .B(n9837), .Z(n9835) );
  XOR U12917 ( .A(n9838), .B(n9839), .Z(n9837) );
  XOR U12918 ( .A(DB[3269]), .B(DB[3262]), .Z(n9839) );
  AND U12919 ( .A(n182), .B(n9840), .Z(n9838) );
  XOR U12920 ( .A(n9841), .B(n9842), .Z(n9840) );
  XOR U12921 ( .A(DB[3262]), .B(DB[3255]), .Z(n9842) );
  AND U12922 ( .A(n186), .B(n9843), .Z(n9841) );
  XOR U12923 ( .A(n9844), .B(n9845), .Z(n9843) );
  XOR U12924 ( .A(DB[3255]), .B(DB[3248]), .Z(n9845) );
  AND U12925 ( .A(n190), .B(n9846), .Z(n9844) );
  XOR U12926 ( .A(n9847), .B(n9848), .Z(n9846) );
  XOR U12927 ( .A(DB[3248]), .B(DB[3241]), .Z(n9848) );
  AND U12928 ( .A(n194), .B(n9849), .Z(n9847) );
  XOR U12929 ( .A(n9850), .B(n9851), .Z(n9849) );
  XOR U12930 ( .A(DB[3241]), .B(DB[3234]), .Z(n9851) );
  AND U12931 ( .A(n198), .B(n9852), .Z(n9850) );
  XOR U12932 ( .A(n9853), .B(n9854), .Z(n9852) );
  XOR U12933 ( .A(DB[3234]), .B(DB[3227]), .Z(n9854) );
  AND U12934 ( .A(n202), .B(n9855), .Z(n9853) );
  XOR U12935 ( .A(n9856), .B(n9857), .Z(n9855) );
  XOR U12936 ( .A(DB[3227]), .B(DB[3220]), .Z(n9857) );
  AND U12937 ( .A(n206), .B(n9858), .Z(n9856) );
  XOR U12938 ( .A(n9859), .B(n9860), .Z(n9858) );
  XOR U12939 ( .A(DB[3220]), .B(DB[3213]), .Z(n9860) );
  AND U12940 ( .A(n210), .B(n9861), .Z(n9859) );
  XOR U12941 ( .A(n9862), .B(n9863), .Z(n9861) );
  XOR U12942 ( .A(DB[3213]), .B(DB[3206]), .Z(n9863) );
  AND U12943 ( .A(n214), .B(n9864), .Z(n9862) );
  XOR U12944 ( .A(n9865), .B(n9866), .Z(n9864) );
  XOR U12945 ( .A(DB[3206]), .B(DB[3199]), .Z(n9866) );
  AND U12946 ( .A(n218), .B(n9867), .Z(n9865) );
  XOR U12947 ( .A(n9868), .B(n9869), .Z(n9867) );
  XOR U12948 ( .A(DB[3199]), .B(DB[3192]), .Z(n9869) );
  AND U12949 ( .A(n222), .B(n9870), .Z(n9868) );
  XOR U12950 ( .A(n9871), .B(n9872), .Z(n9870) );
  XOR U12951 ( .A(DB[3192]), .B(DB[3185]), .Z(n9872) );
  AND U12952 ( .A(n226), .B(n9873), .Z(n9871) );
  XOR U12953 ( .A(n9874), .B(n9875), .Z(n9873) );
  XOR U12954 ( .A(DB[3185]), .B(DB[3178]), .Z(n9875) );
  AND U12955 ( .A(n230), .B(n9876), .Z(n9874) );
  XOR U12956 ( .A(n9877), .B(n9878), .Z(n9876) );
  XOR U12957 ( .A(DB[3178]), .B(DB[3171]), .Z(n9878) );
  AND U12958 ( .A(n234), .B(n9879), .Z(n9877) );
  XOR U12959 ( .A(n9880), .B(n9881), .Z(n9879) );
  XOR U12960 ( .A(DB[3171]), .B(DB[3164]), .Z(n9881) );
  AND U12961 ( .A(n238), .B(n9882), .Z(n9880) );
  XOR U12962 ( .A(n9883), .B(n9884), .Z(n9882) );
  XOR U12963 ( .A(DB[3164]), .B(DB[3157]), .Z(n9884) );
  AND U12964 ( .A(n242), .B(n9885), .Z(n9883) );
  XOR U12965 ( .A(n9886), .B(n9887), .Z(n9885) );
  XOR U12966 ( .A(DB[3157]), .B(DB[3150]), .Z(n9887) );
  AND U12967 ( .A(n246), .B(n9888), .Z(n9886) );
  XOR U12968 ( .A(n9889), .B(n9890), .Z(n9888) );
  XOR U12969 ( .A(DB[3150]), .B(DB[3143]), .Z(n9890) );
  AND U12970 ( .A(n250), .B(n9891), .Z(n9889) );
  XOR U12971 ( .A(n9892), .B(n9893), .Z(n9891) );
  XOR U12972 ( .A(DB[3143]), .B(DB[3136]), .Z(n9893) );
  AND U12973 ( .A(n254), .B(n9894), .Z(n9892) );
  XOR U12974 ( .A(n9895), .B(n9896), .Z(n9894) );
  XOR U12975 ( .A(DB[3136]), .B(DB[3129]), .Z(n9896) );
  AND U12976 ( .A(n258), .B(n9897), .Z(n9895) );
  XOR U12977 ( .A(n9898), .B(n9899), .Z(n9897) );
  XOR U12978 ( .A(DB[3129]), .B(DB[3122]), .Z(n9899) );
  AND U12979 ( .A(n262), .B(n9900), .Z(n9898) );
  XOR U12980 ( .A(n9901), .B(n9902), .Z(n9900) );
  XOR U12981 ( .A(DB[3122]), .B(DB[3115]), .Z(n9902) );
  AND U12982 ( .A(n266), .B(n9903), .Z(n9901) );
  XOR U12983 ( .A(n9904), .B(n9905), .Z(n9903) );
  XOR U12984 ( .A(DB[3115]), .B(DB[3108]), .Z(n9905) );
  AND U12985 ( .A(n270), .B(n9906), .Z(n9904) );
  XOR U12986 ( .A(n9907), .B(n9908), .Z(n9906) );
  XOR U12987 ( .A(DB[3108]), .B(DB[3101]), .Z(n9908) );
  AND U12988 ( .A(n274), .B(n9909), .Z(n9907) );
  XOR U12989 ( .A(n9910), .B(n9911), .Z(n9909) );
  XOR U12990 ( .A(DB[3101]), .B(DB[3094]), .Z(n9911) );
  AND U12991 ( .A(n278), .B(n9912), .Z(n9910) );
  XOR U12992 ( .A(n9913), .B(n9914), .Z(n9912) );
  XOR U12993 ( .A(DB[3094]), .B(DB[3087]), .Z(n9914) );
  AND U12994 ( .A(n282), .B(n9915), .Z(n9913) );
  XOR U12995 ( .A(n9916), .B(n9917), .Z(n9915) );
  XOR U12996 ( .A(DB[3087]), .B(DB[3080]), .Z(n9917) );
  AND U12997 ( .A(n286), .B(n9918), .Z(n9916) );
  XOR U12998 ( .A(n9919), .B(n9920), .Z(n9918) );
  XOR U12999 ( .A(DB[3080]), .B(DB[3073]), .Z(n9920) );
  AND U13000 ( .A(n290), .B(n9921), .Z(n9919) );
  XOR U13001 ( .A(n9922), .B(n9923), .Z(n9921) );
  XOR U13002 ( .A(DB[3073]), .B(DB[3066]), .Z(n9923) );
  AND U13003 ( .A(n294), .B(n9924), .Z(n9922) );
  XOR U13004 ( .A(n9925), .B(n9926), .Z(n9924) );
  XOR U13005 ( .A(DB[3066]), .B(DB[3059]), .Z(n9926) );
  AND U13006 ( .A(n298), .B(n9927), .Z(n9925) );
  XOR U13007 ( .A(n9928), .B(n9929), .Z(n9927) );
  XOR U13008 ( .A(DB[3059]), .B(DB[3052]), .Z(n9929) );
  AND U13009 ( .A(n302), .B(n9930), .Z(n9928) );
  XOR U13010 ( .A(n9931), .B(n9932), .Z(n9930) );
  XOR U13011 ( .A(DB[3052]), .B(DB[3045]), .Z(n9932) );
  AND U13012 ( .A(n306), .B(n9933), .Z(n9931) );
  XOR U13013 ( .A(n9934), .B(n9935), .Z(n9933) );
  XOR U13014 ( .A(DB[3045]), .B(DB[3038]), .Z(n9935) );
  AND U13015 ( .A(n310), .B(n9936), .Z(n9934) );
  XOR U13016 ( .A(n9937), .B(n9938), .Z(n9936) );
  XOR U13017 ( .A(DB[3038]), .B(DB[3031]), .Z(n9938) );
  AND U13018 ( .A(n314), .B(n9939), .Z(n9937) );
  XOR U13019 ( .A(n9940), .B(n9941), .Z(n9939) );
  XOR U13020 ( .A(DB[3031]), .B(DB[3024]), .Z(n9941) );
  AND U13021 ( .A(n318), .B(n9942), .Z(n9940) );
  XOR U13022 ( .A(n9943), .B(n9944), .Z(n9942) );
  XOR U13023 ( .A(DB[3024]), .B(DB[3017]), .Z(n9944) );
  AND U13024 ( .A(n322), .B(n9945), .Z(n9943) );
  XOR U13025 ( .A(n9946), .B(n9947), .Z(n9945) );
  XOR U13026 ( .A(DB[3017]), .B(DB[3010]), .Z(n9947) );
  AND U13027 ( .A(n326), .B(n9948), .Z(n9946) );
  XOR U13028 ( .A(n9949), .B(n9950), .Z(n9948) );
  XOR U13029 ( .A(DB[3010]), .B(DB[3003]), .Z(n9950) );
  AND U13030 ( .A(n330), .B(n9951), .Z(n9949) );
  XOR U13031 ( .A(n9952), .B(n9953), .Z(n9951) );
  XOR U13032 ( .A(DB[3003]), .B(DB[2996]), .Z(n9953) );
  AND U13033 ( .A(n334), .B(n9954), .Z(n9952) );
  XOR U13034 ( .A(n9955), .B(n9956), .Z(n9954) );
  XOR U13035 ( .A(DB[2996]), .B(DB[2989]), .Z(n9956) );
  AND U13036 ( .A(n338), .B(n9957), .Z(n9955) );
  XOR U13037 ( .A(n9958), .B(n9959), .Z(n9957) );
  XOR U13038 ( .A(DB[2989]), .B(DB[2982]), .Z(n9959) );
  AND U13039 ( .A(n342), .B(n9960), .Z(n9958) );
  XOR U13040 ( .A(n9961), .B(n9962), .Z(n9960) );
  XOR U13041 ( .A(DB[2982]), .B(DB[2975]), .Z(n9962) );
  AND U13042 ( .A(n346), .B(n9963), .Z(n9961) );
  XOR U13043 ( .A(n9964), .B(n9965), .Z(n9963) );
  XOR U13044 ( .A(DB[2975]), .B(DB[2968]), .Z(n9965) );
  AND U13045 ( .A(n350), .B(n9966), .Z(n9964) );
  XOR U13046 ( .A(n9967), .B(n9968), .Z(n9966) );
  XOR U13047 ( .A(DB[2968]), .B(DB[2961]), .Z(n9968) );
  AND U13048 ( .A(n354), .B(n9969), .Z(n9967) );
  XOR U13049 ( .A(n9970), .B(n9971), .Z(n9969) );
  XOR U13050 ( .A(DB[2961]), .B(DB[2954]), .Z(n9971) );
  AND U13051 ( .A(n358), .B(n9972), .Z(n9970) );
  XOR U13052 ( .A(n9973), .B(n9974), .Z(n9972) );
  XOR U13053 ( .A(DB[2954]), .B(DB[2947]), .Z(n9974) );
  AND U13054 ( .A(n362), .B(n9975), .Z(n9973) );
  XOR U13055 ( .A(n9976), .B(n9977), .Z(n9975) );
  XOR U13056 ( .A(DB[2947]), .B(DB[2940]), .Z(n9977) );
  AND U13057 ( .A(n366), .B(n9978), .Z(n9976) );
  XOR U13058 ( .A(n9979), .B(n9980), .Z(n9978) );
  XOR U13059 ( .A(DB[2940]), .B(DB[2933]), .Z(n9980) );
  AND U13060 ( .A(n370), .B(n9981), .Z(n9979) );
  XOR U13061 ( .A(n9982), .B(n9983), .Z(n9981) );
  XOR U13062 ( .A(DB[2933]), .B(DB[2926]), .Z(n9983) );
  AND U13063 ( .A(n374), .B(n9984), .Z(n9982) );
  XOR U13064 ( .A(n9985), .B(n9986), .Z(n9984) );
  XOR U13065 ( .A(DB[2926]), .B(DB[2919]), .Z(n9986) );
  AND U13066 ( .A(n378), .B(n9987), .Z(n9985) );
  XOR U13067 ( .A(n9988), .B(n9989), .Z(n9987) );
  XOR U13068 ( .A(DB[2919]), .B(DB[2912]), .Z(n9989) );
  AND U13069 ( .A(n382), .B(n9990), .Z(n9988) );
  XOR U13070 ( .A(n9991), .B(n9992), .Z(n9990) );
  XOR U13071 ( .A(DB[2912]), .B(DB[2905]), .Z(n9992) );
  AND U13072 ( .A(n386), .B(n9993), .Z(n9991) );
  XOR U13073 ( .A(n9994), .B(n9995), .Z(n9993) );
  XOR U13074 ( .A(DB[2905]), .B(DB[2898]), .Z(n9995) );
  AND U13075 ( .A(n390), .B(n9996), .Z(n9994) );
  XOR U13076 ( .A(n9997), .B(n9998), .Z(n9996) );
  XOR U13077 ( .A(DB[2898]), .B(DB[2891]), .Z(n9998) );
  AND U13078 ( .A(n394), .B(n9999), .Z(n9997) );
  XOR U13079 ( .A(n10000), .B(n10001), .Z(n9999) );
  XOR U13080 ( .A(DB[2891]), .B(DB[2884]), .Z(n10001) );
  AND U13081 ( .A(n398), .B(n10002), .Z(n10000) );
  XOR U13082 ( .A(n10003), .B(n10004), .Z(n10002) );
  XOR U13083 ( .A(DB[2884]), .B(DB[2877]), .Z(n10004) );
  AND U13084 ( .A(n402), .B(n10005), .Z(n10003) );
  XOR U13085 ( .A(n10006), .B(n10007), .Z(n10005) );
  XOR U13086 ( .A(DB[2877]), .B(DB[2870]), .Z(n10007) );
  AND U13087 ( .A(n406), .B(n10008), .Z(n10006) );
  XOR U13088 ( .A(n10009), .B(n10010), .Z(n10008) );
  XOR U13089 ( .A(DB[2870]), .B(DB[2863]), .Z(n10010) );
  AND U13090 ( .A(n410), .B(n10011), .Z(n10009) );
  XOR U13091 ( .A(n10012), .B(n10013), .Z(n10011) );
  XOR U13092 ( .A(DB[2863]), .B(DB[2856]), .Z(n10013) );
  AND U13093 ( .A(n414), .B(n10014), .Z(n10012) );
  XOR U13094 ( .A(n10015), .B(n10016), .Z(n10014) );
  XOR U13095 ( .A(DB[2856]), .B(DB[2849]), .Z(n10016) );
  AND U13096 ( .A(n418), .B(n10017), .Z(n10015) );
  XOR U13097 ( .A(n10018), .B(n10019), .Z(n10017) );
  XOR U13098 ( .A(DB[2849]), .B(DB[2842]), .Z(n10019) );
  AND U13099 ( .A(n422), .B(n10020), .Z(n10018) );
  XOR U13100 ( .A(n10021), .B(n10022), .Z(n10020) );
  XOR U13101 ( .A(DB[2842]), .B(DB[2835]), .Z(n10022) );
  AND U13102 ( .A(n426), .B(n10023), .Z(n10021) );
  XOR U13103 ( .A(n10024), .B(n10025), .Z(n10023) );
  XOR U13104 ( .A(DB[2835]), .B(DB[2828]), .Z(n10025) );
  AND U13105 ( .A(n430), .B(n10026), .Z(n10024) );
  XOR U13106 ( .A(n10027), .B(n10028), .Z(n10026) );
  XOR U13107 ( .A(DB[2828]), .B(DB[2821]), .Z(n10028) );
  AND U13108 ( .A(n434), .B(n10029), .Z(n10027) );
  XOR U13109 ( .A(n10030), .B(n10031), .Z(n10029) );
  XOR U13110 ( .A(DB[2821]), .B(DB[2814]), .Z(n10031) );
  AND U13111 ( .A(n438), .B(n10032), .Z(n10030) );
  XOR U13112 ( .A(n10033), .B(n10034), .Z(n10032) );
  XOR U13113 ( .A(DB[2814]), .B(DB[2807]), .Z(n10034) );
  AND U13114 ( .A(n442), .B(n10035), .Z(n10033) );
  XOR U13115 ( .A(n10036), .B(n10037), .Z(n10035) );
  XOR U13116 ( .A(DB[2807]), .B(DB[2800]), .Z(n10037) );
  AND U13117 ( .A(n446), .B(n10038), .Z(n10036) );
  XOR U13118 ( .A(n10039), .B(n10040), .Z(n10038) );
  XOR U13119 ( .A(DB[2800]), .B(DB[2793]), .Z(n10040) );
  AND U13120 ( .A(n450), .B(n10041), .Z(n10039) );
  XOR U13121 ( .A(n10042), .B(n10043), .Z(n10041) );
  XOR U13122 ( .A(DB[2793]), .B(DB[2786]), .Z(n10043) );
  AND U13123 ( .A(n454), .B(n10044), .Z(n10042) );
  XOR U13124 ( .A(n10045), .B(n10046), .Z(n10044) );
  XOR U13125 ( .A(DB[2786]), .B(DB[2779]), .Z(n10046) );
  AND U13126 ( .A(n458), .B(n10047), .Z(n10045) );
  XOR U13127 ( .A(n10048), .B(n10049), .Z(n10047) );
  XOR U13128 ( .A(DB[2779]), .B(DB[2772]), .Z(n10049) );
  AND U13129 ( .A(n462), .B(n10050), .Z(n10048) );
  XOR U13130 ( .A(n10051), .B(n10052), .Z(n10050) );
  XOR U13131 ( .A(DB[2772]), .B(DB[2765]), .Z(n10052) );
  AND U13132 ( .A(n466), .B(n10053), .Z(n10051) );
  XOR U13133 ( .A(n10054), .B(n10055), .Z(n10053) );
  XOR U13134 ( .A(DB[2765]), .B(DB[2758]), .Z(n10055) );
  AND U13135 ( .A(n470), .B(n10056), .Z(n10054) );
  XOR U13136 ( .A(n10057), .B(n10058), .Z(n10056) );
  XOR U13137 ( .A(DB[2758]), .B(DB[2751]), .Z(n10058) );
  AND U13138 ( .A(n474), .B(n10059), .Z(n10057) );
  XOR U13139 ( .A(n10060), .B(n10061), .Z(n10059) );
  XOR U13140 ( .A(DB[2751]), .B(DB[2744]), .Z(n10061) );
  AND U13141 ( .A(n478), .B(n10062), .Z(n10060) );
  XOR U13142 ( .A(n10063), .B(n10064), .Z(n10062) );
  XOR U13143 ( .A(DB[2744]), .B(DB[2737]), .Z(n10064) );
  AND U13144 ( .A(n482), .B(n10065), .Z(n10063) );
  XOR U13145 ( .A(n10066), .B(n10067), .Z(n10065) );
  XOR U13146 ( .A(DB[2737]), .B(DB[2730]), .Z(n10067) );
  AND U13147 ( .A(n486), .B(n10068), .Z(n10066) );
  XOR U13148 ( .A(n10069), .B(n10070), .Z(n10068) );
  XOR U13149 ( .A(DB[2730]), .B(DB[2723]), .Z(n10070) );
  AND U13150 ( .A(n490), .B(n10071), .Z(n10069) );
  XOR U13151 ( .A(n10072), .B(n10073), .Z(n10071) );
  XOR U13152 ( .A(DB[2723]), .B(DB[2716]), .Z(n10073) );
  AND U13153 ( .A(n494), .B(n10074), .Z(n10072) );
  XOR U13154 ( .A(n10075), .B(n10076), .Z(n10074) );
  XOR U13155 ( .A(DB[2716]), .B(DB[2709]), .Z(n10076) );
  AND U13156 ( .A(n498), .B(n10077), .Z(n10075) );
  XOR U13157 ( .A(n10078), .B(n10079), .Z(n10077) );
  XOR U13158 ( .A(DB[2709]), .B(DB[2702]), .Z(n10079) );
  AND U13159 ( .A(n502), .B(n10080), .Z(n10078) );
  XOR U13160 ( .A(n10081), .B(n10082), .Z(n10080) );
  XOR U13161 ( .A(DB[2702]), .B(DB[2695]), .Z(n10082) );
  AND U13162 ( .A(n506), .B(n10083), .Z(n10081) );
  XOR U13163 ( .A(n10084), .B(n10085), .Z(n10083) );
  XOR U13164 ( .A(DB[2695]), .B(DB[2688]), .Z(n10085) );
  AND U13165 ( .A(n510), .B(n10086), .Z(n10084) );
  XOR U13166 ( .A(n10087), .B(n10088), .Z(n10086) );
  XOR U13167 ( .A(DB[2688]), .B(DB[2681]), .Z(n10088) );
  AND U13168 ( .A(n514), .B(n10089), .Z(n10087) );
  XOR U13169 ( .A(n10090), .B(n10091), .Z(n10089) );
  XOR U13170 ( .A(DB[2681]), .B(DB[2674]), .Z(n10091) );
  AND U13171 ( .A(n518), .B(n10092), .Z(n10090) );
  XOR U13172 ( .A(n10093), .B(n10094), .Z(n10092) );
  XOR U13173 ( .A(DB[2674]), .B(DB[2667]), .Z(n10094) );
  AND U13174 ( .A(n522), .B(n10095), .Z(n10093) );
  XOR U13175 ( .A(n10096), .B(n10097), .Z(n10095) );
  XOR U13176 ( .A(DB[2667]), .B(DB[2660]), .Z(n10097) );
  AND U13177 ( .A(n526), .B(n10098), .Z(n10096) );
  XOR U13178 ( .A(n10099), .B(n10100), .Z(n10098) );
  XOR U13179 ( .A(DB[2660]), .B(DB[2653]), .Z(n10100) );
  AND U13180 ( .A(n530), .B(n10101), .Z(n10099) );
  XOR U13181 ( .A(n10102), .B(n10103), .Z(n10101) );
  XOR U13182 ( .A(DB[2653]), .B(DB[2646]), .Z(n10103) );
  AND U13183 ( .A(n534), .B(n10104), .Z(n10102) );
  XOR U13184 ( .A(n10105), .B(n10106), .Z(n10104) );
  XOR U13185 ( .A(DB[2646]), .B(DB[2639]), .Z(n10106) );
  AND U13186 ( .A(n538), .B(n10107), .Z(n10105) );
  XOR U13187 ( .A(n10108), .B(n10109), .Z(n10107) );
  XOR U13188 ( .A(DB[2639]), .B(DB[2632]), .Z(n10109) );
  AND U13189 ( .A(n542), .B(n10110), .Z(n10108) );
  XOR U13190 ( .A(n10111), .B(n10112), .Z(n10110) );
  XOR U13191 ( .A(DB[2632]), .B(DB[2625]), .Z(n10112) );
  AND U13192 ( .A(n546), .B(n10113), .Z(n10111) );
  XOR U13193 ( .A(n10114), .B(n10115), .Z(n10113) );
  XOR U13194 ( .A(DB[2625]), .B(DB[2618]), .Z(n10115) );
  AND U13195 ( .A(n550), .B(n10116), .Z(n10114) );
  XOR U13196 ( .A(n10117), .B(n10118), .Z(n10116) );
  XOR U13197 ( .A(DB[2618]), .B(DB[2611]), .Z(n10118) );
  AND U13198 ( .A(n554), .B(n10119), .Z(n10117) );
  XOR U13199 ( .A(n10120), .B(n10121), .Z(n10119) );
  XOR U13200 ( .A(DB[2611]), .B(DB[2604]), .Z(n10121) );
  AND U13201 ( .A(n558), .B(n10122), .Z(n10120) );
  XOR U13202 ( .A(n10123), .B(n10124), .Z(n10122) );
  XOR U13203 ( .A(DB[2604]), .B(DB[2597]), .Z(n10124) );
  AND U13204 ( .A(n562), .B(n10125), .Z(n10123) );
  XOR U13205 ( .A(n10126), .B(n10127), .Z(n10125) );
  XOR U13206 ( .A(DB[2597]), .B(DB[2590]), .Z(n10127) );
  AND U13207 ( .A(n566), .B(n10128), .Z(n10126) );
  XOR U13208 ( .A(n10129), .B(n10130), .Z(n10128) );
  XOR U13209 ( .A(DB[2590]), .B(DB[2583]), .Z(n10130) );
  AND U13210 ( .A(n570), .B(n10131), .Z(n10129) );
  XOR U13211 ( .A(n10132), .B(n10133), .Z(n10131) );
  XOR U13212 ( .A(DB[2583]), .B(DB[2576]), .Z(n10133) );
  AND U13213 ( .A(n574), .B(n10134), .Z(n10132) );
  XOR U13214 ( .A(n10135), .B(n10136), .Z(n10134) );
  XOR U13215 ( .A(DB[2576]), .B(DB[2569]), .Z(n10136) );
  AND U13216 ( .A(n578), .B(n10137), .Z(n10135) );
  XOR U13217 ( .A(n10138), .B(n10139), .Z(n10137) );
  XOR U13218 ( .A(DB[2569]), .B(DB[2562]), .Z(n10139) );
  AND U13219 ( .A(n582), .B(n10140), .Z(n10138) );
  XOR U13220 ( .A(n10141), .B(n10142), .Z(n10140) );
  XOR U13221 ( .A(DB[2562]), .B(DB[2555]), .Z(n10142) );
  AND U13222 ( .A(n586), .B(n10143), .Z(n10141) );
  XOR U13223 ( .A(n10144), .B(n10145), .Z(n10143) );
  XOR U13224 ( .A(DB[2555]), .B(DB[2548]), .Z(n10145) );
  AND U13225 ( .A(n590), .B(n10146), .Z(n10144) );
  XOR U13226 ( .A(n10147), .B(n10148), .Z(n10146) );
  XOR U13227 ( .A(DB[2548]), .B(DB[2541]), .Z(n10148) );
  AND U13228 ( .A(n594), .B(n10149), .Z(n10147) );
  XOR U13229 ( .A(n10150), .B(n10151), .Z(n10149) );
  XOR U13230 ( .A(DB[2541]), .B(DB[2534]), .Z(n10151) );
  AND U13231 ( .A(n598), .B(n10152), .Z(n10150) );
  XOR U13232 ( .A(n10153), .B(n10154), .Z(n10152) );
  XOR U13233 ( .A(DB[2534]), .B(DB[2527]), .Z(n10154) );
  AND U13234 ( .A(n602), .B(n10155), .Z(n10153) );
  XOR U13235 ( .A(n10156), .B(n10157), .Z(n10155) );
  XOR U13236 ( .A(DB[2527]), .B(DB[2520]), .Z(n10157) );
  AND U13237 ( .A(n606), .B(n10158), .Z(n10156) );
  XOR U13238 ( .A(n10159), .B(n10160), .Z(n10158) );
  XOR U13239 ( .A(DB[2520]), .B(DB[2513]), .Z(n10160) );
  AND U13240 ( .A(n610), .B(n10161), .Z(n10159) );
  XOR U13241 ( .A(n10162), .B(n10163), .Z(n10161) );
  XOR U13242 ( .A(DB[2513]), .B(DB[2506]), .Z(n10163) );
  AND U13243 ( .A(n614), .B(n10164), .Z(n10162) );
  XOR U13244 ( .A(n10165), .B(n10166), .Z(n10164) );
  XOR U13245 ( .A(DB[2506]), .B(DB[2499]), .Z(n10166) );
  AND U13246 ( .A(n618), .B(n10167), .Z(n10165) );
  XOR U13247 ( .A(n10168), .B(n10169), .Z(n10167) );
  XOR U13248 ( .A(DB[2499]), .B(DB[2492]), .Z(n10169) );
  AND U13249 ( .A(n622), .B(n10170), .Z(n10168) );
  XOR U13250 ( .A(n10171), .B(n10172), .Z(n10170) );
  XOR U13251 ( .A(DB[2492]), .B(DB[2485]), .Z(n10172) );
  AND U13252 ( .A(n626), .B(n10173), .Z(n10171) );
  XOR U13253 ( .A(n10174), .B(n10175), .Z(n10173) );
  XOR U13254 ( .A(DB[2485]), .B(DB[2478]), .Z(n10175) );
  AND U13255 ( .A(n630), .B(n10176), .Z(n10174) );
  XOR U13256 ( .A(n10177), .B(n10178), .Z(n10176) );
  XOR U13257 ( .A(DB[2478]), .B(DB[2471]), .Z(n10178) );
  AND U13258 ( .A(n634), .B(n10179), .Z(n10177) );
  XOR U13259 ( .A(n10180), .B(n10181), .Z(n10179) );
  XOR U13260 ( .A(DB[2471]), .B(DB[2464]), .Z(n10181) );
  AND U13261 ( .A(n638), .B(n10182), .Z(n10180) );
  XOR U13262 ( .A(n10183), .B(n10184), .Z(n10182) );
  XOR U13263 ( .A(DB[2464]), .B(DB[2457]), .Z(n10184) );
  AND U13264 ( .A(n642), .B(n10185), .Z(n10183) );
  XOR U13265 ( .A(n10186), .B(n10187), .Z(n10185) );
  XOR U13266 ( .A(DB[2457]), .B(DB[2450]), .Z(n10187) );
  AND U13267 ( .A(n646), .B(n10188), .Z(n10186) );
  XOR U13268 ( .A(n10189), .B(n10190), .Z(n10188) );
  XOR U13269 ( .A(DB[2450]), .B(DB[2443]), .Z(n10190) );
  AND U13270 ( .A(n650), .B(n10191), .Z(n10189) );
  XOR U13271 ( .A(n10192), .B(n10193), .Z(n10191) );
  XOR U13272 ( .A(DB[2443]), .B(DB[2436]), .Z(n10193) );
  AND U13273 ( .A(n654), .B(n10194), .Z(n10192) );
  XOR U13274 ( .A(n10195), .B(n10196), .Z(n10194) );
  XOR U13275 ( .A(DB[2436]), .B(DB[2429]), .Z(n10196) );
  AND U13276 ( .A(n658), .B(n10197), .Z(n10195) );
  XOR U13277 ( .A(n10198), .B(n10199), .Z(n10197) );
  XOR U13278 ( .A(DB[2429]), .B(DB[2422]), .Z(n10199) );
  AND U13279 ( .A(n662), .B(n10200), .Z(n10198) );
  XOR U13280 ( .A(n10201), .B(n10202), .Z(n10200) );
  XOR U13281 ( .A(DB[2422]), .B(DB[2415]), .Z(n10202) );
  AND U13282 ( .A(n666), .B(n10203), .Z(n10201) );
  XOR U13283 ( .A(n10204), .B(n10205), .Z(n10203) );
  XOR U13284 ( .A(DB[2415]), .B(DB[2408]), .Z(n10205) );
  AND U13285 ( .A(n670), .B(n10206), .Z(n10204) );
  XOR U13286 ( .A(n10207), .B(n10208), .Z(n10206) );
  XOR U13287 ( .A(DB[2408]), .B(DB[2401]), .Z(n10208) );
  AND U13288 ( .A(n674), .B(n10209), .Z(n10207) );
  XOR U13289 ( .A(n10210), .B(n10211), .Z(n10209) );
  XOR U13290 ( .A(DB[2401]), .B(DB[2394]), .Z(n10211) );
  AND U13291 ( .A(n678), .B(n10212), .Z(n10210) );
  XOR U13292 ( .A(n10213), .B(n10214), .Z(n10212) );
  XOR U13293 ( .A(DB[2394]), .B(DB[2387]), .Z(n10214) );
  AND U13294 ( .A(n682), .B(n10215), .Z(n10213) );
  XOR U13295 ( .A(n10216), .B(n10217), .Z(n10215) );
  XOR U13296 ( .A(DB[2387]), .B(DB[2380]), .Z(n10217) );
  AND U13297 ( .A(n686), .B(n10218), .Z(n10216) );
  XOR U13298 ( .A(n10219), .B(n10220), .Z(n10218) );
  XOR U13299 ( .A(DB[2380]), .B(DB[2373]), .Z(n10220) );
  AND U13300 ( .A(n690), .B(n10221), .Z(n10219) );
  XOR U13301 ( .A(n10222), .B(n10223), .Z(n10221) );
  XOR U13302 ( .A(DB[2373]), .B(DB[2366]), .Z(n10223) );
  AND U13303 ( .A(n694), .B(n10224), .Z(n10222) );
  XOR U13304 ( .A(n10225), .B(n10226), .Z(n10224) );
  XOR U13305 ( .A(DB[2366]), .B(DB[2359]), .Z(n10226) );
  AND U13306 ( .A(n698), .B(n10227), .Z(n10225) );
  XOR U13307 ( .A(n10228), .B(n10229), .Z(n10227) );
  XOR U13308 ( .A(DB[2359]), .B(DB[2352]), .Z(n10229) );
  AND U13309 ( .A(n702), .B(n10230), .Z(n10228) );
  XOR U13310 ( .A(n10231), .B(n10232), .Z(n10230) );
  XOR U13311 ( .A(DB[2352]), .B(DB[2345]), .Z(n10232) );
  AND U13312 ( .A(n706), .B(n10233), .Z(n10231) );
  XOR U13313 ( .A(n10234), .B(n10235), .Z(n10233) );
  XOR U13314 ( .A(DB[2345]), .B(DB[2338]), .Z(n10235) );
  AND U13315 ( .A(n710), .B(n10236), .Z(n10234) );
  XOR U13316 ( .A(n10237), .B(n10238), .Z(n10236) );
  XOR U13317 ( .A(DB[2338]), .B(DB[2331]), .Z(n10238) );
  AND U13318 ( .A(n714), .B(n10239), .Z(n10237) );
  XOR U13319 ( .A(n10240), .B(n10241), .Z(n10239) );
  XOR U13320 ( .A(DB[2331]), .B(DB[2324]), .Z(n10241) );
  AND U13321 ( .A(n718), .B(n10242), .Z(n10240) );
  XOR U13322 ( .A(n10243), .B(n10244), .Z(n10242) );
  XOR U13323 ( .A(DB[2324]), .B(DB[2317]), .Z(n10244) );
  AND U13324 ( .A(n722), .B(n10245), .Z(n10243) );
  XOR U13325 ( .A(n10246), .B(n10247), .Z(n10245) );
  XOR U13326 ( .A(DB[2317]), .B(DB[2310]), .Z(n10247) );
  AND U13327 ( .A(n726), .B(n10248), .Z(n10246) );
  XOR U13328 ( .A(n10249), .B(n10250), .Z(n10248) );
  XOR U13329 ( .A(DB[2310]), .B(DB[2303]), .Z(n10250) );
  AND U13330 ( .A(n730), .B(n10251), .Z(n10249) );
  XOR U13331 ( .A(n10252), .B(n10253), .Z(n10251) );
  XOR U13332 ( .A(DB[2303]), .B(DB[2296]), .Z(n10253) );
  AND U13333 ( .A(n734), .B(n10254), .Z(n10252) );
  XOR U13334 ( .A(n10255), .B(n10256), .Z(n10254) );
  XOR U13335 ( .A(DB[2296]), .B(DB[2289]), .Z(n10256) );
  AND U13336 ( .A(n738), .B(n10257), .Z(n10255) );
  XOR U13337 ( .A(n10258), .B(n10259), .Z(n10257) );
  XOR U13338 ( .A(DB[2289]), .B(DB[2282]), .Z(n10259) );
  AND U13339 ( .A(n742), .B(n10260), .Z(n10258) );
  XOR U13340 ( .A(n10261), .B(n10262), .Z(n10260) );
  XOR U13341 ( .A(DB[2282]), .B(DB[2275]), .Z(n10262) );
  AND U13342 ( .A(n746), .B(n10263), .Z(n10261) );
  XOR U13343 ( .A(n10264), .B(n10265), .Z(n10263) );
  XOR U13344 ( .A(DB[2275]), .B(DB[2268]), .Z(n10265) );
  AND U13345 ( .A(n750), .B(n10266), .Z(n10264) );
  XOR U13346 ( .A(n10267), .B(n10268), .Z(n10266) );
  XOR U13347 ( .A(DB[2268]), .B(DB[2261]), .Z(n10268) );
  AND U13348 ( .A(n754), .B(n10269), .Z(n10267) );
  XOR U13349 ( .A(n10270), .B(n10271), .Z(n10269) );
  XOR U13350 ( .A(DB[2261]), .B(DB[2254]), .Z(n10271) );
  AND U13351 ( .A(n758), .B(n10272), .Z(n10270) );
  XOR U13352 ( .A(n10273), .B(n10274), .Z(n10272) );
  XOR U13353 ( .A(DB[2254]), .B(DB[2247]), .Z(n10274) );
  AND U13354 ( .A(n762), .B(n10275), .Z(n10273) );
  XOR U13355 ( .A(n10276), .B(n10277), .Z(n10275) );
  XOR U13356 ( .A(DB[2247]), .B(DB[2240]), .Z(n10277) );
  AND U13357 ( .A(n766), .B(n10278), .Z(n10276) );
  XOR U13358 ( .A(n10279), .B(n10280), .Z(n10278) );
  XOR U13359 ( .A(DB[2240]), .B(DB[2233]), .Z(n10280) );
  AND U13360 ( .A(n770), .B(n10281), .Z(n10279) );
  XOR U13361 ( .A(n10282), .B(n10283), .Z(n10281) );
  XOR U13362 ( .A(DB[2233]), .B(DB[2226]), .Z(n10283) );
  AND U13363 ( .A(n774), .B(n10284), .Z(n10282) );
  XOR U13364 ( .A(n10285), .B(n10286), .Z(n10284) );
  XOR U13365 ( .A(DB[2226]), .B(DB[2219]), .Z(n10286) );
  AND U13366 ( .A(n778), .B(n10287), .Z(n10285) );
  XOR U13367 ( .A(n10288), .B(n10289), .Z(n10287) );
  XOR U13368 ( .A(DB[2219]), .B(DB[2212]), .Z(n10289) );
  AND U13369 ( .A(n782), .B(n10290), .Z(n10288) );
  XOR U13370 ( .A(n10291), .B(n10292), .Z(n10290) );
  XOR U13371 ( .A(DB[2212]), .B(DB[2205]), .Z(n10292) );
  AND U13372 ( .A(n786), .B(n10293), .Z(n10291) );
  XOR U13373 ( .A(n10294), .B(n10295), .Z(n10293) );
  XOR U13374 ( .A(DB[2205]), .B(DB[2198]), .Z(n10295) );
  AND U13375 ( .A(n790), .B(n10296), .Z(n10294) );
  XOR U13376 ( .A(n10297), .B(n10298), .Z(n10296) );
  XOR U13377 ( .A(DB[2198]), .B(DB[2191]), .Z(n10298) );
  AND U13378 ( .A(n794), .B(n10299), .Z(n10297) );
  XOR U13379 ( .A(n10300), .B(n10301), .Z(n10299) );
  XOR U13380 ( .A(DB[2191]), .B(DB[2184]), .Z(n10301) );
  AND U13381 ( .A(n798), .B(n10302), .Z(n10300) );
  XOR U13382 ( .A(n10303), .B(n10304), .Z(n10302) );
  XOR U13383 ( .A(DB[2184]), .B(DB[2177]), .Z(n10304) );
  AND U13384 ( .A(n802), .B(n10305), .Z(n10303) );
  XOR U13385 ( .A(n10306), .B(n10307), .Z(n10305) );
  XOR U13386 ( .A(DB[2177]), .B(DB[2170]), .Z(n10307) );
  AND U13387 ( .A(n806), .B(n10308), .Z(n10306) );
  XOR U13388 ( .A(n10309), .B(n10310), .Z(n10308) );
  XOR U13389 ( .A(DB[2170]), .B(DB[2163]), .Z(n10310) );
  AND U13390 ( .A(n810), .B(n10311), .Z(n10309) );
  XOR U13391 ( .A(n10312), .B(n10313), .Z(n10311) );
  XOR U13392 ( .A(DB[2163]), .B(DB[2156]), .Z(n10313) );
  AND U13393 ( .A(n814), .B(n10314), .Z(n10312) );
  XOR U13394 ( .A(n10315), .B(n10316), .Z(n10314) );
  XOR U13395 ( .A(DB[2156]), .B(DB[2149]), .Z(n10316) );
  AND U13396 ( .A(n818), .B(n10317), .Z(n10315) );
  XOR U13397 ( .A(n10318), .B(n10319), .Z(n10317) );
  XOR U13398 ( .A(DB[2149]), .B(DB[2142]), .Z(n10319) );
  AND U13399 ( .A(n822), .B(n10320), .Z(n10318) );
  XOR U13400 ( .A(n10321), .B(n10322), .Z(n10320) );
  XOR U13401 ( .A(DB[2142]), .B(DB[2135]), .Z(n10322) );
  AND U13402 ( .A(n826), .B(n10323), .Z(n10321) );
  XOR U13403 ( .A(n10324), .B(n10325), .Z(n10323) );
  XOR U13404 ( .A(DB[2135]), .B(DB[2128]), .Z(n10325) );
  AND U13405 ( .A(n830), .B(n10326), .Z(n10324) );
  XOR U13406 ( .A(n10327), .B(n10328), .Z(n10326) );
  XOR U13407 ( .A(DB[2128]), .B(DB[2121]), .Z(n10328) );
  AND U13408 ( .A(n834), .B(n10329), .Z(n10327) );
  XOR U13409 ( .A(n10330), .B(n10331), .Z(n10329) );
  XOR U13410 ( .A(DB[2121]), .B(DB[2114]), .Z(n10331) );
  AND U13411 ( .A(n838), .B(n10332), .Z(n10330) );
  XOR U13412 ( .A(n10333), .B(n10334), .Z(n10332) );
  XOR U13413 ( .A(DB[2114]), .B(DB[2107]), .Z(n10334) );
  AND U13414 ( .A(n842), .B(n10335), .Z(n10333) );
  XOR U13415 ( .A(n10336), .B(n10337), .Z(n10335) );
  XOR U13416 ( .A(DB[2107]), .B(DB[2100]), .Z(n10337) );
  AND U13417 ( .A(n846), .B(n10338), .Z(n10336) );
  XOR U13418 ( .A(n10339), .B(n10340), .Z(n10338) );
  XOR U13419 ( .A(DB[2100]), .B(DB[2093]), .Z(n10340) );
  AND U13420 ( .A(n850), .B(n10341), .Z(n10339) );
  XOR U13421 ( .A(n10342), .B(n10343), .Z(n10341) );
  XOR U13422 ( .A(DB[2093]), .B(DB[2086]), .Z(n10343) );
  AND U13423 ( .A(n854), .B(n10344), .Z(n10342) );
  XOR U13424 ( .A(n10345), .B(n10346), .Z(n10344) );
  XOR U13425 ( .A(DB[2086]), .B(DB[2079]), .Z(n10346) );
  AND U13426 ( .A(n858), .B(n10347), .Z(n10345) );
  XOR U13427 ( .A(n10348), .B(n10349), .Z(n10347) );
  XOR U13428 ( .A(DB[2079]), .B(DB[2072]), .Z(n10349) );
  AND U13429 ( .A(n862), .B(n10350), .Z(n10348) );
  XOR U13430 ( .A(n10351), .B(n10352), .Z(n10350) );
  XOR U13431 ( .A(DB[2072]), .B(DB[2065]), .Z(n10352) );
  AND U13432 ( .A(n866), .B(n10353), .Z(n10351) );
  XOR U13433 ( .A(n10354), .B(n10355), .Z(n10353) );
  XOR U13434 ( .A(DB[2065]), .B(DB[2058]), .Z(n10355) );
  AND U13435 ( .A(n870), .B(n10356), .Z(n10354) );
  XOR U13436 ( .A(n10357), .B(n10358), .Z(n10356) );
  XOR U13437 ( .A(DB[2058]), .B(DB[2051]), .Z(n10358) );
  AND U13438 ( .A(n874), .B(n10359), .Z(n10357) );
  XOR U13439 ( .A(n10360), .B(n10361), .Z(n10359) );
  XOR U13440 ( .A(DB[2051]), .B(DB[2044]), .Z(n10361) );
  AND U13441 ( .A(n878), .B(n10362), .Z(n10360) );
  XOR U13442 ( .A(n10363), .B(n10364), .Z(n10362) );
  XOR U13443 ( .A(DB[2044]), .B(DB[2037]), .Z(n10364) );
  AND U13444 ( .A(n882), .B(n10365), .Z(n10363) );
  XOR U13445 ( .A(n10366), .B(n10367), .Z(n10365) );
  XOR U13446 ( .A(DB[2037]), .B(DB[2030]), .Z(n10367) );
  AND U13447 ( .A(n886), .B(n10368), .Z(n10366) );
  XOR U13448 ( .A(n10369), .B(n10370), .Z(n10368) );
  XOR U13449 ( .A(DB[2030]), .B(DB[2023]), .Z(n10370) );
  AND U13450 ( .A(n890), .B(n10371), .Z(n10369) );
  XOR U13451 ( .A(n10372), .B(n10373), .Z(n10371) );
  XOR U13452 ( .A(DB[2023]), .B(DB[2016]), .Z(n10373) );
  AND U13453 ( .A(n894), .B(n10374), .Z(n10372) );
  XOR U13454 ( .A(n10375), .B(n10376), .Z(n10374) );
  XOR U13455 ( .A(DB[2016]), .B(DB[2009]), .Z(n10376) );
  AND U13456 ( .A(n898), .B(n10377), .Z(n10375) );
  XOR U13457 ( .A(n10378), .B(n10379), .Z(n10377) );
  XOR U13458 ( .A(DB[2009]), .B(DB[2002]), .Z(n10379) );
  AND U13459 ( .A(n902), .B(n10380), .Z(n10378) );
  XOR U13460 ( .A(n10381), .B(n10382), .Z(n10380) );
  XOR U13461 ( .A(DB[2002]), .B(DB[1995]), .Z(n10382) );
  AND U13462 ( .A(n906), .B(n10383), .Z(n10381) );
  XOR U13463 ( .A(n10384), .B(n10385), .Z(n10383) );
  XOR U13464 ( .A(DB[1995]), .B(DB[1988]), .Z(n10385) );
  AND U13465 ( .A(n910), .B(n10386), .Z(n10384) );
  XOR U13466 ( .A(n10387), .B(n10388), .Z(n10386) );
  XOR U13467 ( .A(DB[1988]), .B(DB[1981]), .Z(n10388) );
  AND U13468 ( .A(n914), .B(n10389), .Z(n10387) );
  XOR U13469 ( .A(n10390), .B(n10391), .Z(n10389) );
  XOR U13470 ( .A(DB[1981]), .B(DB[1974]), .Z(n10391) );
  AND U13471 ( .A(n918), .B(n10392), .Z(n10390) );
  XOR U13472 ( .A(n10393), .B(n10394), .Z(n10392) );
  XOR U13473 ( .A(DB[1974]), .B(DB[1967]), .Z(n10394) );
  AND U13474 ( .A(n922), .B(n10395), .Z(n10393) );
  XOR U13475 ( .A(n10396), .B(n10397), .Z(n10395) );
  XOR U13476 ( .A(DB[1967]), .B(DB[1960]), .Z(n10397) );
  AND U13477 ( .A(n926), .B(n10398), .Z(n10396) );
  XOR U13478 ( .A(n10399), .B(n10400), .Z(n10398) );
  XOR U13479 ( .A(DB[1960]), .B(DB[1953]), .Z(n10400) );
  AND U13480 ( .A(n930), .B(n10401), .Z(n10399) );
  XOR U13481 ( .A(n10402), .B(n10403), .Z(n10401) );
  XOR U13482 ( .A(DB[1953]), .B(DB[1946]), .Z(n10403) );
  AND U13483 ( .A(n934), .B(n10404), .Z(n10402) );
  XOR U13484 ( .A(n10405), .B(n10406), .Z(n10404) );
  XOR U13485 ( .A(DB[1946]), .B(DB[1939]), .Z(n10406) );
  AND U13486 ( .A(n938), .B(n10407), .Z(n10405) );
  XOR U13487 ( .A(n10408), .B(n10409), .Z(n10407) );
  XOR U13488 ( .A(DB[1939]), .B(DB[1932]), .Z(n10409) );
  AND U13489 ( .A(n942), .B(n10410), .Z(n10408) );
  XOR U13490 ( .A(n10411), .B(n10412), .Z(n10410) );
  XOR U13491 ( .A(DB[1932]), .B(DB[1925]), .Z(n10412) );
  AND U13492 ( .A(n946), .B(n10413), .Z(n10411) );
  XOR U13493 ( .A(n10414), .B(n10415), .Z(n10413) );
  XOR U13494 ( .A(DB[1925]), .B(DB[1918]), .Z(n10415) );
  AND U13495 ( .A(n950), .B(n10416), .Z(n10414) );
  XOR U13496 ( .A(n10417), .B(n10418), .Z(n10416) );
  XOR U13497 ( .A(DB[1918]), .B(DB[1911]), .Z(n10418) );
  AND U13498 ( .A(n954), .B(n10419), .Z(n10417) );
  XOR U13499 ( .A(n10420), .B(n10421), .Z(n10419) );
  XOR U13500 ( .A(DB[1911]), .B(DB[1904]), .Z(n10421) );
  AND U13501 ( .A(n958), .B(n10422), .Z(n10420) );
  XOR U13502 ( .A(n10423), .B(n10424), .Z(n10422) );
  XOR U13503 ( .A(DB[1904]), .B(DB[1897]), .Z(n10424) );
  AND U13504 ( .A(n962), .B(n10425), .Z(n10423) );
  XOR U13505 ( .A(n10426), .B(n10427), .Z(n10425) );
  XOR U13506 ( .A(DB[1897]), .B(DB[1890]), .Z(n10427) );
  AND U13507 ( .A(n966), .B(n10428), .Z(n10426) );
  XOR U13508 ( .A(n10429), .B(n10430), .Z(n10428) );
  XOR U13509 ( .A(DB[1890]), .B(DB[1883]), .Z(n10430) );
  AND U13510 ( .A(n970), .B(n10431), .Z(n10429) );
  XOR U13511 ( .A(n10432), .B(n10433), .Z(n10431) );
  XOR U13512 ( .A(DB[1883]), .B(DB[1876]), .Z(n10433) );
  AND U13513 ( .A(n974), .B(n10434), .Z(n10432) );
  XOR U13514 ( .A(n10435), .B(n10436), .Z(n10434) );
  XOR U13515 ( .A(DB[1876]), .B(DB[1869]), .Z(n10436) );
  AND U13516 ( .A(n978), .B(n10437), .Z(n10435) );
  XOR U13517 ( .A(n10438), .B(n10439), .Z(n10437) );
  XOR U13518 ( .A(DB[1869]), .B(DB[1862]), .Z(n10439) );
  AND U13519 ( .A(n982), .B(n10440), .Z(n10438) );
  XOR U13520 ( .A(n10441), .B(n10442), .Z(n10440) );
  XOR U13521 ( .A(DB[1862]), .B(DB[1855]), .Z(n10442) );
  AND U13522 ( .A(n986), .B(n10443), .Z(n10441) );
  XOR U13523 ( .A(n10444), .B(n10445), .Z(n10443) );
  XOR U13524 ( .A(DB[1855]), .B(DB[1848]), .Z(n10445) );
  AND U13525 ( .A(n990), .B(n10446), .Z(n10444) );
  XOR U13526 ( .A(n10447), .B(n10448), .Z(n10446) );
  XOR U13527 ( .A(DB[1848]), .B(DB[1841]), .Z(n10448) );
  AND U13528 ( .A(n994), .B(n10449), .Z(n10447) );
  XOR U13529 ( .A(n10450), .B(n10451), .Z(n10449) );
  XOR U13530 ( .A(DB[1841]), .B(DB[1834]), .Z(n10451) );
  AND U13531 ( .A(n998), .B(n10452), .Z(n10450) );
  XOR U13532 ( .A(n10453), .B(n10454), .Z(n10452) );
  XOR U13533 ( .A(DB[1834]), .B(DB[1827]), .Z(n10454) );
  AND U13534 ( .A(n1002), .B(n10455), .Z(n10453) );
  XOR U13535 ( .A(n10456), .B(n10457), .Z(n10455) );
  XOR U13536 ( .A(DB[1827]), .B(DB[1820]), .Z(n10457) );
  AND U13537 ( .A(n1006), .B(n10458), .Z(n10456) );
  XOR U13538 ( .A(n10459), .B(n10460), .Z(n10458) );
  XOR U13539 ( .A(DB[1820]), .B(DB[1813]), .Z(n10460) );
  AND U13540 ( .A(n1010), .B(n10461), .Z(n10459) );
  XOR U13541 ( .A(n10462), .B(n10463), .Z(n10461) );
  XOR U13542 ( .A(DB[1813]), .B(DB[1806]), .Z(n10463) );
  AND U13543 ( .A(n1014), .B(n10464), .Z(n10462) );
  XOR U13544 ( .A(n10465), .B(n10466), .Z(n10464) );
  XOR U13545 ( .A(DB[1806]), .B(DB[1799]), .Z(n10466) );
  AND U13546 ( .A(n1018), .B(n10467), .Z(n10465) );
  XOR U13547 ( .A(n10468), .B(n10469), .Z(n10467) );
  XOR U13548 ( .A(DB[1799]), .B(DB[1792]), .Z(n10469) );
  AND U13549 ( .A(n1022), .B(n10470), .Z(n10468) );
  XOR U13550 ( .A(n10471), .B(n10472), .Z(n10470) );
  XOR U13551 ( .A(DB[1792]), .B(DB[1785]), .Z(n10472) );
  AND U13552 ( .A(n1026), .B(n10473), .Z(n10471) );
  XOR U13553 ( .A(n10474), .B(n10475), .Z(n10473) );
  XOR U13554 ( .A(DB[1785]), .B(DB[1778]), .Z(n10475) );
  AND U13555 ( .A(n1030), .B(n10476), .Z(n10474) );
  XOR U13556 ( .A(n10477), .B(n10478), .Z(n10476) );
  XOR U13557 ( .A(DB[1778]), .B(DB[1771]), .Z(n10478) );
  AND U13558 ( .A(n1034), .B(n10479), .Z(n10477) );
  XOR U13559 ( .A(n10480), .B(n10481), .Z(n10479) );
  XOR U13560 ( .A(DB[1771]), .B(DB[1764]), .Z(n10481) );
  AND U13561 ( .A(n1038), .B(n10482), .Z(n10480) );
  XOR U13562 ( .A(n10483), .B(n10484), .Z(n10482) );
  XOR U13563 ( .A(DB[1764]), .B(DB[1757]), .Z(n10484) );
  AND U13564 ( .A(n1042), .B(n10485), .Z(n10483) );
  XOR U13565 ( .A(n10486), .B(n10487), .Z(n10485) );
  XOR U13566 ( .A(DB[1757]), .B(DB[1750]), .Z(n10487) );
  AND U13567 ( .A(n1046), .B(n10488), .Z(n10486) );
  XOR U13568 ( .A(n10489), .B(n10490), .Z(n10488) );
  XOR U13569 ( .A(DB[1750]), .B(DB[1743]), .Z(n10490) );
  AND U13570 ( .A(n1050), .B(n10491), .Z(n10489) );
  XOR U13571 ( .A(n10492), .B(n10493), .Z(n10491) );
  XOR U13572 ( .A(DB[1743]), .B(DB[1736]), .Z(n10493) );
  AND U13573 ( .A(n1054), .B(n10494), .Z(n10492) );
  XOR U13574 ( .A(n10495), .B(n10496), .Z(n10494) );
  XOR U13575 ( .A(DB[1736]), .B(DB[1729]), .Z(n10496) );
  AND U13576 ( .A(n1058), .B(n10497), .Z(n10495) );
  XOR U13577 ( .A(n10498), .B(n10499), .Z(n10497) );
  XOR U13578 ( .A(DB[1729]), .B(DB[1722]), .Z(n10499) );
  AND U13579 ( .A(n1062), .B(n10500), .Z(n10498) );
  XOR U13580 ( .A(n10501), .B(n10502), .Z(n10500) );
  XOR U13581 ( .A(DB[1722]), .B(DB[1715]), .Z(n10502) );
  AND U13582 ( .A(n1066), .B(n10503), .Z(n10501) );
  XOR U13583 ( .A(n10504), .B(n10505), .Z(n10503) );
  XOR U13584 ( .A(DB[1715]), .B(DB[1708]), .Z(n10505) );
  AND U13585 ( .A(n1070), .B(n10506), .Z(n10504) );
  XOR U13586 ( .A(n10507), .B(n10508), .Z(n10506) );
  XOR U13587 ( .A(DB[1708]), .B(DB[1701]), .Z(n10508) );
  AND U13588 ( .A(n1074), .B(n10509), .Z(n10507) );
  XOR U13589 ( .A(n10510), .B(n10511), .Z(n10509) );
  XOR U13590 ( .A(DB[1701]), .B(DB[1694]), .Z(n10511) );
  AND U13591 ( .A(n1078), .B(n10512), .Z(n10510) );
  XOR U13592 ( .A(n10513), .B(n10514), .Z(n10512) );
  XOR U13593 ( .A(DB[1694]), .B(DB[1687]), .Z(n10514) );
  AND U13594 ( .A(n1082), .B(n10515), .Z(n10513) );
  XOR U13595 ( .A(n10516), .B(n10517), .Z(n10515) );
  XOR U13596 ( .A(DB[1687]), .B(DB[1680]), .Z(n10517) );
  AND U13597 ( .A(n1086), .B(n10518), .Z(n10516) );
  XOR U13598 ( .A(n10519), .B(n10520), .Z(n10518) );
  XOR U13599 ( .A(DB[1680]), .B(DB[1673]), .Z(n10520) );
  AND U13600 ( .A(n1090), .B(n10521), .Z(n10519) );
  XOR U13601 ( .A(n10522), .B(n10523), .Z(n10521) );
  XOR U13602 ( .A(DB[1673]), .B(DB[1666]), .Z(n10523) );
  AND U13603 ( .A(n1094), .B(n10524), .Z(n10522) );
  XOR U13604 ( .A(n10525), .B(n10526), .Z(n10524) );
  XOR U13605 ( .A(DB[1666]), .B(DB[1659]), .Z(n10526) );
  AND U13606 ( .A(n1098), .B(n10527), .Z(n10525) );
  XOR U13607 ( .A(n10528), .B(n10529), .Z(n10527) );
  XOR U13608 ( .A(DB[1659]), .B(DB[1652]), .Z(n10529) );
  AND U13609 ( .A(n1102), .B(n10530), .Z(n10528) );
  XOR U13610 ( .A(n10531), .B(n10532), .Z(n10530) );
  XOR U13611 ( .A(DB[1652]), .B(DB[1645]), .Z(n10532) );
  AND U13612 ( .A(n1106), .B(n10533), .Z(n10531) );
  XOR U13613 ( .A(n10534), .B(n10535), .Z(n10533) );
  XOR U13614 ( .A(DB[1645]), .B(DB[1638]), .Z(n10535) );
  AND U13615 ( .A(n1110), .B(n10536), .Z(n10534) );
  XOR U13616 ( .A(n10537), .B(n10538), .Z(n10536) );
  XOR U13617 ( .A(DB[1638]), .B(DB[1631]), .Z(n10538) );
  AND U13618 ( .A(n1114), .B(n10539), .Z(n10537) );
  XOR U13619 ( .A(n10540), .B(n10541), .Z(n10539) );
  XOR U13620 ( .A(DB[1631]), .B(DB[1624]), .Z(n10541) );
  AND U13621 ( .A(n1118), .B(n10542), .Z(n10540) );
  XOR U13622 ( .A(n10543), .B(n10544), .Z(n10542) );
  XOR U13623 ( .A(DB[1624]), .B(DB[1617]), .Z(n10544) );
  AND U13624 ( .A(n1122), .B(n10545), .Z(n10543) );
  XOR U13625 ( .A(n10546), .B(n10547), .Z(n10545) );
  XOR U13626 ( .A(DB[1617]), .B(DB[1610]), .Z(n10547) );
  AND U13627 ( .A(n1126), .B(n10548), .Z(n10546) );
  XOR U13628 ( .A(n10549), .B(n10550), .Z(n10548) );
  XOR U13629 ( .A(DB[1610]), .B(DB[1603]), .Z(n10550) );
  AND U13630 ( .A(n1130), .B(n10551), .Z(n10549) );
  XOR U13631 ( .A(n10552), .B(n10553), .Z(n10551) );
  XOR U13632 ( .A(DB[1603]), .B(DB[1596]), .Z(n10553) );
  AND U13633 ( .A(n1134), .B(n10554), .Z(n10552) );
  XOR U13634 ( .A(n10555), .B(n10556), .Z(n10554) );
  XOR U13635 ( .A(DB[1596]), .B(DB[1589]), .Z(n10556) );
  AND U13636 ( .A(n1138), .B(n10557), .Z(n10555) );
  XOR U13637 ( .A(n10558), .B(n10559), .Z(n10557) );
  XOR U13638 ( .A(DB[1589]), .B(DB[1582]), .Z(n10559) );
  AND U13639 ( .A(n1142), .B(n10560), .Z(n10558) );
  XOR U13640 ( .A(n10561), .B(n10562), .Z(n10560) );
  XOR U13641 ( .A(DB[1582]), .B(DB[1575]), .Z(n10562) );
  AND U13642 ( .A(n1146), .B(n10563), .Z(n10561) );
  XOR U13643 ( .A(n10564), .B(n10565), .Z(n10563) );
  XOR U13644 ( .A(DB[1575]), .B(DB[1568]), .Z(n10565) );
  AND U13645 ( .A(n1150), .B(n10566), .Z(n10564) );
  XOR U13646 ( .A(n10567), .B(n10568), .Z(n10566) );
  XOR U13647 ( .A(DB[1568]), .B(DB[1561]), .Z(n10568) );
  AND U13648 ( .A(n1154), .B(n10569), .Z(n10567) );
  XOR U13649 ( .A(n10570), .B(n10571), .Z(n10569) );
  XOR U13650 ( .A(DB[1561]), .B(DB[1554]), .Z(n10571) );
  AND U13651 ( .A(n1158), .B(n10572), .Z(n10570) );
  XOR U13652 ( .A(n10573), .B(n10574), .Z(n10572) );
  XOR U13653 ( .A(DB[1554]), .B(DB[1547]), .Z(n10574) );
  AND U13654 ( .A(n1162), .B(n10575), .Z(n10573) );
  XOR U13655 ( .A(n10576), .B(n10577), .Z(n10575) );
  XOR U13656 ( .A(DB[1547]), .B(DB[1540]), .Z(n10577) );
  AND U13657 ( .A(n1166), .B(n10578), .Z(n10576) );
  XOR U13658 ( .A(n10579), .B(n10580), .Z(n10578) );
  XOR U13659 ( .A(DB[1540]), .B(DB[1533]), .Z(n10580) );
  AND U13660 ( .A(n1170), .B(n10581), .Z(n10579) );
  XOR U13661 ( .A(n10582), .B(n10583), .Z(n10581) );
  XOR U13662 ( .A(DB[1533]), .B(DB[1526]), .Z(n10583) );
  AND U13663 ( .A(n1174), .B(n10584), .Z(n10582) );
  XOR U13664 ( .A(n10585), .B(n10586), .Z(n10584) );
  XOR U13665 ( .A(DB[1526]), .B(DB[1519]), .Z(n10586) );
  AND U13666 ( .A(n1178), .B(n10587), .Z(n10585) );
  XOR U13667 ( .A(n10588), .B(n10589), .Z(n10587) );
  XOR U13668 ( .A(DB[1519]), .B(DB[1512]), .Z(n10589) );
  AND U13669 ( .A(n1182), .B(n10590), .Z(n10588) );
  XOR U13670 ( .A(n10591), .B(n10592), .Z(n10590) );
  XOR U13671 ( .A(DB[1512]), .B(DB[1505]), .Z(n10592) );
  AND U13672 ( .A(n1186), .B(n10593), .Z(n10591) );
  XOR U13673 ( .A(n10594), .B(n10595), .Z(n10593) );
  XOR U13674 ( .A(DB[1505]), .B(DB[1498]), .Z(n10595) );
  AND U13675 ( .A(n1190), .B(n10596), .Z(n10594) );
  XOR U13676 ( .A(n10597), .B(n10598), .Z(n10596) );
  XOR U13677 ( .A(DB[1498]), .B(DB[1491]), .Z(n10598) );
  AND U13678 ( .A(n1194), .B(n10599), .Z(n10597) );
  XOR U13679 ( .A(n10600), .B(n10601), .Z(n10599) );
  XOR U13680 ( .A(DB[1491]), .B(DB[1484]), .Z(n10601) );
  AND U13681 ( .A(n1198), .B(n10602), .Z(n10600) );
  XOR U13682 ( .A(n10603), .B(n10604), .Z(n10602) );
  XOR U13683 ( .A(DB[1484]), .B(DB[1477]), .Z(n10604) );
  AND U13684 ( .A(n1202), .B(n10605), .Z(n10603) );
  XOR U13685 ( .A(n10606), .B(n10607), .Z(n10605) );
  XOR U13686 ( .A(DB[1477]), .B(DB[1470]), .Z(n10607) );
  AND U13687 ( .A(n1206), .B(n10608), .Z(n10606) );
  XOR U13688 ( .A(n10609), .B(n10610), .Z(n10608) );
  XOR U13689 ( .A(DB[1470]), .B(DB[1463]), .Z(n10610) );
  AND U13690 ( .A(n1210), .B(n10611), .Z(n10609) );
  XOR U13691 ( .A(n10612), .B(n10613), .Z(n10611) );
  XOR U13692 ( .A(DB[1463]), .B(DB[1456]), .Z(n10613) );
  AND U13693 ( .A(n1214), .B(n10614), .Z(n10612) );
  XOR U13694 ( .A(n10615), .B(n10616), .Z(n10614) );
  XOR U13695 ( .A(DB[1456]), .B(DB[1449]), .Z(n10616) );
  AND U13696 ( .A(n1218), .B(n10617), .Z(n10615) );
  XOR U13697 ( .A(n10618), .B(n10619), .Z(n10617) );
  XOR U13698 ( .A(DB[1449]), .B(DB[1442]), .Z(n10619) );
  AND U13699 ( .A(n1222), .B(n10620), .Z(n10618) );
  XOR U13700 ( .A(n10621), .B(n10622), .Z(n10620) );
  XOR U13701 ( .A(DB[1442]), .B(DB[1435]), .Z(n10622) );
  AND U13702 ( .A(n1226), .B(n10623), .Z(n10621) );
  XOR U13703 ( .A(n10624), .B(n10625), .Z(n10623) );
  XOR U13704 ( .A(DB[1435]), .B(DB[1428]), .Z(n10625) );
  AND U13705 ( .A(n1230), .B(n10626), .Z(n10624) );
  XOR U13706 ( .A(n10627), .B(n10628), .Z(n10626) );
  XOR U13707 ( .A(DB[1428]), .B(DB[1421]), .Z(n10628) );
  AND U13708 ( .A(n1234), .B(n10629), .Z(n10627) );
  XOR U13709 ( .A(n10630), .B(n10631), .Z(n10629) );
  XOR U13710 ( .A(DB[1421]), .B(DB[1414]), .Z(n10631) );
  AND U13711 ( .A(n1238), .B(n10632), .Z(n10630) );
  XOR U13712 ( .A(n10633), .B(n10634), .Z(n10632) );
  XOR U13713 ( .A(DB[1414]), .B(DB[1407]), .Z(n10634) );
  AND U13714 ( .A(n1242), .B(n10635), .Z(n10633) );
  XOR U13715 ( .A(n10636), .B(n10637), .Z(n10635) );
  XOR U13716 ( .A(DB[1407]), .B(DB[1400]), .Z(n10637) );
  AND U13717 ( .A(n1246), .B(n10638), .Z(n10636) );
  XOR U13718 ( .A(n10639), .B(n10640), .Z(n10638) );
  XOR U13719 ( .A(DB[1400]), .B(DB[1393]), .Z(n10640) );
  AND U13720 ( .A(n1250), .B(n10641), .Z(n10639) );
  XOR U13721 ( .A(n10642), .B(n10643), .Z(n10641) );
  XOR U13722 ( .A(DB[1393]), .B(DB[1386]), .Z(n10643) );
  AND U13723 ( .A(n1254), .B(n10644), .Z(n10642) );
  XOR U13724 ( .A(n10645), .B(n10646), .Z(n10644) );
  XOR U13725 ( .A(DB[1386]), .B(DB[1379]), .Z(n10646) );
  AND U13726 ( .A(n1258), .B(n10647), .Z(n10645) );
  XOR U13727 ( .A(n10648), .B(n10649), .Z(n10647) );
  XOR U13728 ( .A(DB[1379]), .B(DB[1372]), .Z(n10649) );
  AND U13729 ( .A(n1262), .B(n10650), .Z(n10648) );
  XOR U13730 ( .A(n10651), .B(n10652), .Z(n10650) );
  XOR U13731 ( .A(DB[1372]), .B(DB[1365]), .Z(n10652) );
  AND U13732 ( .A(n1266), .B(n10653), .Z(n10651) );
  XOR U13733 ( .A(n10654), .B(n10655), .Z(n10653) );
  XOR U13734 ( .A(DB[1365]), .B(DB[1358]), .Z(n10655) );
  AND U13735 ( .A(n1270), .B(n10656), .Z(n10654) );
  XOR U13736 ( .A(n10657), .B(n10658), .Z(n10656) );
  XOR U13737 ( .A(DB[1358]), .B(DB[1351]), .Z(n10658) );
  AND U13738 ( .A(n1274), .B(n10659), .Z(n10657) );
  XOR U13739 ( .A(n10660), .B(n10661), .Z(n10659) );
  XOR U13740 ( .A(DB[1351]), .B(DB[1344]), .Z(n10661) );
  AND U13741 ( .A(n1278), .B(n10662), .Z(n10660) );
  XOR U13742 ( .A(n10663), .B(n10664), .Z(n10662) );
  XOR U13743 ( .A(DB[1344]), .B(DB[1337]), .Z(n10664) );
  AND U13744 ( .A(n1282), .B(n10665), .Z(n10663) );
  XOR U13745 ( .A(n10666), .B(n10667), .Z(n10665) );
  XOR U13746 ( .A(DB[1337]), .B(DB[1330]), .Z(n10667) );
  AND U13747 ( .A(n1286), .B(n10668), .Z(n10666) );
  XOR U13748 ( .A(n10669), .B(n10670), .Z(n10668) );
  XOR U13749 ( .A(DB[1330]), .B(DB[1323]), .Z(n10670) );
  AND U13750 ( .A(n1290), .B(n10671), .Z(n10669) );
  XOR U13751 ( .A(n10672), .B(n10673), .Z(n10671) );
  XOR U13752 ( .A(DB[1323]), .B(DB[1316]), .Z(n10673) );
  AND U13753 ( .A(n1294), .B(n10674), .Z(n10672) );
  XOR U13754 ( .A(n10675), .B(n10676), .Z(n10674) );
  XOR U13755 ( .A(DB[1316]), .B(DB[1309]), .Z(n10676) );
  AND U13756 ( .A(n1298), .B(n10677), .Z(n10675) );
  XOR U13757 ( .A(n10678), .B(n10679), .Z(n10677) );
  XOR U13758 ( .A(DB[1309]), .B(DB[1302]), .Z(n10679) );
  AND U13759 ( .A(n1302), .B(n10680), .Z(n10678) );
  XOR U13760 ( .A(n10681), .B(n10682), .Z(n10680) );
  XOR U13761 ( .A(DB[1302]), .B(DB[1295]), .Z(n10682) );
  AND U13762 ( .A(n1306), .B(n10683), .Z(n10681) );
  XOR U13763 ( .A(n10684), .B(n10685), .Z(n10683) );
  XOR U13764 ( .A(DB[1295]), .B(DB[1288]), .Z(n10685) );
  AND U13765 ( .A(n1310), .B(n10686), .Z(n10684) );
  XOR U13766 ( .A(n10687), .B(n10688), .Z(n10686) );
  XOR U13767 ( .A(DB[1288]), .B(DB[1281]), .Z(n10688) );
  AND U13768 ( .A(n1314), .B(n10689), .Z(n10687) );
  XOR U13769 ( .A(n10690), .B(n10691), .Z(n10689) );
  XOR U13770 ( .A(DB[1281]), .B(DB[1274]), .Z(n10691) );
  AND U13771 ( .A(n1318), .B(n10692), .Z(n10690) );
  XOR U13772 ( .A(n10693), .B(n10694), .Z(n10692) );
  XOR U13773 ( .A(DB[1274]), .B(DB[1267]), .Z(n10694) );
  AND U13774 ( .A(n1322), .B(n10695), .Z(n10693) );
  XOR U13775 ( .A(n10696), .B(n10697), .Z(n10695) );
  XOR U13776 ( .A(DB[1267]), .B(DB[1260]), .Z(n10697) );
  AND U13777 ( .A(n1326), .B(n10698), .Z(n10696) );
  XOR U13778 ( .A(n10699), .B(n10700), .Z(n10698) );
  XOR U13779 ( .A(DB[1260]), .B(DB[1253]), .Z(n10700) );
  AND U13780 ( .A(n1330), .B(n10701), .Z(n10699) );
  XOR U13781 ( .A(n10702), .B(n10703), .Z(n10701) );
  XOR U13782 ( .A(DB[1253]), .B(DB[1246]), .Z(n10703) );
  AND U13783 ( .A(n1334), .B(n10704), .Z(n10702) );
  XOR U13784 ( .A(n10705), .B(n10706), .Z(n10704) );
  XOR U13785 ( .A(DB[1246]), .B(DB[1239]), .Z(n10706) );
  AND U13786 ( .A(n1338), .B(n10707), .Z(n10705) );
  XOR U13787 ( .A(n10708), .B(n10709), .Z(n10707) );
  XOR U13788 ( .A(DB[1239]), .B(DB[1232]), .Z(n10709) );
  AND U13789 ( .A(n1342), .B(n10710), .Z(n10708) );
  XOR U13790 ( .A(n10711), .B(n10712), .Z(n10710) );
  XOR U13791 ( .A(DB[1232]), .B(DB[1225]), .Z(n10712) );
  AND U13792 ( .A(n1346), .B(n10713), .Z(n10711) );
  XOR U13793 ( .A(n10714), .B(n10715), .Z(n10713) );
  XOR U13794 ( .A(DB[1225]), .B(DB[1218]), .Z(n10715) );
  AND U13795 ( .A(n1350), .B(n10716), .Z(n10714) );
  XOR U13796 ( .A(n10717), .B(n10718), .Z(n10716) );
  XOR U13797 ( .A(DB[1218]), .B(DB[1211]), .Z(n10718) );
  AND U13798 ( .A(n1354), .B(n10719), .Z(n10717) );
  XOR U13799 ( .A(n10720), .B(n10721), .Z(n10719) );
  XOR U13800 ( .A(DB[1211]), .B(DB[1204]), .Z(n10721) );
  AND U13801 ( .A(n1358), .B(n10722), .Z(n10720) );
  XOR U13802 ( .A(n10723), .B(n10724), .Z(n10722) );
  XOR U13803 ( .A(DB[1204]), .B(DB[1197]), .Z(n10724) );
  AND U13804 ( .A(n1362), .B(n10725), .Z(n10723) );
  XOR U13805 ( .A(n10726), .B(n10727), .Z(n10725) );
  XOR U13806 ( .A(DB[1197]), .B(DB[1190]), .Z(n10727) );
  AND U13807 ( .A(n1366), .B(n10728), .Z(n10726) );
  XOR U13808 ( .A(n10729), .B(n10730), .Z(n10728) );
  XOR U13809 ( .A(DB[1190]), .B(DB[1183]), .Z(n10730) );
  AND U13810 ( .A(n1370), .B(n10731), .Z(n10729) );
  XOR U13811 ( .A(n10732), .B(n10733), .Z(n10731) );
  XOR U13812 ( .A(DB[1183]), .B(DB[1176]), .Z(n10733) );
  AND U13813 ( .A(n1374), .B(n10734), .Z(n10732) );
  XOR U13814 ( .A(n10735), .B(n10736), .Z(n10734) );
  XOR U13815 ( .A(DB[1176]), .B(DB[1169]), .Z(n10736) );
  AND U13816 ( .A(n1378), .B(n10737), .Z(n10735) );
  XOR U13817 ( .A(n10738), .B(n10739), .Z(n10737) );
  XOR U13818 ( .A(DB[1169]), .B(DB[1162]), .Z(n10739) );
  AND U13819 ( .A(n1382), .B(n10740), .Z(n10738) );
  XOR U13820 ( .A(n10741), .B(n10742), .Z(n10740) );
  XOR U13821 ( .A(DB[1162]), .B(DB[1155]), .Z(n10742) );
  AND U13822 ( .A(n1386), .B(n10743), .Z(n10741) );
  XOR U13823 ( .A(n10744), .B(n10745), .Z(n10743) );
  XOR U13824 ( .A(DB[1155]), .B(DB[1148]), .Z(n10745) );
  AND U13825 ( .A(n1390), .B(n10746), .Z(n10744) );
  XOR U13826 ( .A(n10747), .B(n10748), .Z(n10746) );
  XOR U13827 ( .A(DB[1148]), .B(DB[1141]), .Z(n10748) );
  AND U13828 ( .A(n1394), .B(n10749), .Z(n10747) );
  XOR U13829 ( .A(n10750), .B(n10751), .Z(n10749) );
  XOR U13830 ( .A(DB[1141]), .B(DB[1134]), .Z(n10751) );
  AND U13831 ( .A(n1398), .B(n10752), .Z(n10750) );
  XOR U13832 ( .A(n10753), .B(n10754), .Z(n10752) );
  XOR U13833 ( .A(DB[1134]), .B(DB[1127]), .Z(n10754) );
  AND U13834 ( .A(n1402), .B(n10755), .Z(n10753) );
  XOR U13835 ( .A(n10756), .B(n10757), .Z(n10755) );
  XOR U13836 ( .A(DB[1127]), .B(DB[1120]), .Z(n10757) );
  AND U13837 ( .A(n1406), .B(n10758), .Z(n10756) );
  XOR U13838 ( .A(n10759), .B(n10760), .Z(n10758) );
  XOR U13839 ( .A(DB[1120]), .B(DB[1113]), .Z(n10760) );
  AND U13840 ( .A(n1410), .B(n10761), .Z(n10759) );
  XOR U13841 ( .A(n10762), .B(n10763), .Z(n10761) );
  XOR U13842 ( .A(DB[1113]), .B(DB[1106]), .Z(n10763) );
  AND U13843 ( .A(n1414), .B(n10764), .Z(n10762) );
  XOR U13844 ( .A(n10765), .B(n10766), .Z(n10764) );
  XOR U13845 ( .A(DB[1106]), .B(DB[1099]), .Z(n10766) );
  AND U13846 ( .A(n1418), .B(n10767), .Z(n10765) );
  XOR U13847 ( .A(n10768), .B(n10769), .Z(n10767) );
  XOR U13848 ( .A(DB[1099]), .B(DB[1092]), .Z(n10769) );
  AND U13849 ( .A(n1422), .B(n10770), .Z(n10768) );
  XOR U13850 ( .A(n10771), .B(n10772), .Z(n10770) );
  XOR U13851 ( .A(DB[1092]), .B(DB[1085]), .Z(n10772) );
  AND U13852 ( .A(n1426), .B(n10773), .Z(n10771) );
  XOR U13853 ( .A(n10774), .B(n10775), .Z(n10773) );
  XOR U13854 ( .A(DB[1085]), .B(DB[1078]), .Z(n10775) );
  AND U13855 ( .A(n1430), .B(n10776), .Z(n10774) );
  XOR U13856 ( .A(n10777), .B(n10778), .Z(n10776) );
  XOR U13857 ( .A(DB[1078]), .B(DB[1071]), .Z(n10778) );
  AND U13858 ( .A(n1434), .B(n10779), .Z(n10777) );
  XOR U13859 ( .A(n10780), .B(n10781), .Z(n10779) );
  XOR U13860 ( .A(DB[1071]), .B(DB[1064]), .Z(n10781) );
  AND U13861 ( .A(n1438), .B(n10782), .Z(n10780) );
  XOR U13862 ( .A(n10783), .B(n10784), .Z(n10782) );
  XOR U13863 ( .A(DB[1064]), .B(DB[1057]), .Z(n10784) );
  AND U13864 ( .A(n1442), .B(n10785), .Z(n10783) );
  XOR U13865 ( .A(n10786), .B(n10787), .Z(n10785) );
  XOR U13866 ( .A(DB[1057]), .B(DB[1050]), .Z(n10787) );
  AND U13867 ( .A(n1446), .B(n10788), .Z(n10786) );
  XOR U13868 ( .A(n10789), .B(n10790), .Z(n10788) );
  XOR U13869 ( .A(DB[1050]), .B(DB[1043]), .Z(n10790) );
  AND U13870 ( .A(n1450), .B(n10791), .Z(n10789) );
  XOR U13871 ( .A(n10792), .B(n10793), .Z(n10791) );
  XOR U13872 ( .A(DB[1043]), .B(DB[1036]), .Z(n10793) );
  AND U13873 ( .A(n1454), .B(n10794), .Z(n10792) );
  XOR U13874 ( .A(n10795), .B(n10796), .Z(n10794) );
  XOR U13875 ( .A(DB[1036]), .B(DB[1029]), .Z(n10796) );
  AND U13876 ( .A(n1458), .B(n10797), .Z(n10795) );
  XOR U13877 ( .A(n10798), .B(n10799), .Z(n10797) );
  XOR U13878 ( .A(DB[1029]), .B(DB[1022]), .Z(n10799) );
  AND U13879 ( .A(n1462), .B(n10800), .Z(n10798) );
  XOR U13880 ( .A(n10801), .B(n10802), .Z(n10800) );
  XOR U13881 ( .A(DB[1022]), .B(DB[1015]), .Z(n10802) );
  AND U13882 ( .A(n1466), .B(n10803), .Z(n10801) );
  XOR U13883 ( .A(n10804), .B(n10805), .Z(n10803) );
  XOR U13884 ( .A(DB[1015]), .B(DB[1008]), .Z(n10805) );
  AND U13885 ( .A(n1470), .B(n10806), .Z(n10804) );
  XOR U13886 ( .A(n10807), .B(n10808), .Z(n10806) );
  XOR U13887 ( .A(DB[1008]), .B(DB[1001]), .Z(n10808) );
  AND U13888 ( .A(n1474), .B(n10809), .Z(n10807) );
  XOR U13889 ( .A(n10810), .B(n10811), .Z(n10809) );
  XOR U13890 ( .A(DB[994]), .B(DB[1001]), .Z(n10811) );
  AND U13891 ( .A(n1478), .B(n10812), .Z(n10810) );
  XOR U13892 ( .A(n10813), .B(n10814), .Z(n10812) );
  XOR U13893 ( .A(DB[994]), .B(DB[987]), .Z(n10814) );
  AND U13894 ( .A(n1482), .B(n10815), .Z(n10813) );
  XOR U13895 ( .A(n10816), .B(n10817), .Z(n10815) );
  XOR U13896 ( .A(DB[987]), .B(DB[980]), .Z(n10817) );
  AND U13897 ( .A(n1486), .B(n10818), .Z(n10816) );
  XOR U13898 ( .A(n10819), .B(n10820), .Z(n10818) );
  XOR U13899 ( .A(DB[980]), .B(DB[973]), .Z(n10820) );
  AND U13900 ( .A(n1490), .B(n10821), .Z(n10819) );
  XOR U13901 ( .A(n10822), .B(n10823), .Z(n10821) );
  XOR U13902 ( .A(DB[973]), .B(DB[966]), .Z(n10823) );
  AND U13903 ( .A(n1494), .B(n10824), .Z(n10822) );
  XOR U13904 ( .A(n10825), .B(n10826), .Z(n10824) );
  XOR U13905 ( .A(DB[966]), .B(DB[959]), .Z(n10826) );
  AND U13906 ( .A(n1498), .B(n10827), .Z(n10825) );
  XOR U13907 ( .A(n10828), .B(n10829), .Z(n10827) );
  XOR U13908 ( .A(DB[959]), .B(DB[952]), .Z(n10829) );
  AND U13909 ( .A(n1502), .B(n10830), .Z(n10828) );
  XOR U13910 ( .A(n10831), .B(n10832), .Z(n10830) );
  XOR U13911 ( .A(DB[952]), .B(DB[945]), .Z(n10832) );
  AND U13912 ( .A(n1506), .B(n10833), .Z(n10831) );
  XOR U13913 ( .A(n10834), .B(n10835), .Z(n10833) );
  XOR U13914 ( .A(DB[945]), .B(DB[938]), .Z(n10835) );
  AND U13915 ( .A(n1510), .B(n10836), .Z(n10834) );
  XOR U13916 ( .A(n10837), .B(n10838), .Z(n10836) );
  XOR U13917 ( .A(DB[938]), .B(DB[931]), .Z(n10838) );
  AND U13918 ( .A(n1514), .B(n10839), .Z(n10837) );
  XOR U13919 ( .A(n10840), .B(n10841), .Z(n10839) );
  XOR U13920 ( .A(DB[931]), .B(DB[924]), .Z(n10841) );
  AND U13921 ( .A(n1518), .B(n10842), .Z(n10840) );
  XOR U13922 ( .A(n10843), .B(n10844), .Z(n10842) );
  XOR U13923 ( .A(DB[924]), .B(DB[917]), .Z(n10844) );
  AND U13924 ( .A(n1522), .B(n10845), .Z(n10843) );
  XOR U13925 ( .A(n10846), .B(n10847), .Z(n10845) );
  XOR U13926 ( .A(DB[917]), .B(DB[910]), .Z(n10847) );
  AND U13927 ( .A(n1526), .B(n10848), .Z(n10846) );
  XOR U13928 ( .A(n10849), .B(n10850), .Z(n10848) );
  XOR U13929 ( .A(DB[910]), .B(DB[903]), .Z(n10850) );
  AND U13930 ( .A(n1530), .B(n10851), .Z(n10849) );
  XOR U13931 ( .A(n10852), .B(n10853), .Z(n10851) );
  XOR U13932 ( .A(DB[903]), .B(DB[896]), .Z(n10853) );
  AND U13933 ( .A(n1534), .B(n10854), .Z(n10852) );
  XOR U13934 ( .A(n10855), .B(n10856), .Z(n10854) );
  XOR U13935 ( .A(DB[896]), .B(DB[889]), .Z(n10856) );
  AND U13936 ( .A(n1538), .B(n10857), .Z(n10855) );
  XOR U13937 ( .A(n10858), .B(n10859), .Z(n10857) );
  XOR U13938 ( .A(DB[889]), .B(DB[882]), .Z(n10859) );
  AND U13939 ( .A(n1542), .B(n10860), .Z(n10858) );
  XOR U13940 ( .A(n10861), .B(n10862), .Z(n10860) );
  XOR U13941 ( .A(DB[882]), .B(DB[875]), .Z(n10862) );
  AND U13942 ( .A(n1546), .B(n10863), .Z(n10861) );
  XOR U13943 ( .A(n10864), .B(n10865), .Z(n10863) );
  XOR U13944 ( .A(DB[875]), .B(DB[868]), .Z(n10865) );
  AND U13945 ( .A(n1550), .B(n10866), .Z(n10864) );
  XOR U13946 ( .A(n10867), .B(n10868), .Z(n10866) );
  XOR U13947 ( .A(DB[868]), .B(DB[861]), .Z(n10868) );
  AND U13948 ( .A(n1554), .B(n10869), .Z(n10867) );
  XOR U13949 ( .A(n10870), .B(n10871), .Z(n10869) );
  XOR U13950 ( .A(DB[861]), .B(DB[854]), .Z(n10871) );
  AND U13951 ( .A(n1558), .B(n10872), .Z(n10870) );
  XOR U13952 ( .A(n10873), .B(n10874), .Z(n10872) );
  XOR U13953 ( .A(DB[854]), .B(DB[847]), .Z(n10874) );
  AND U13954 ( .A(n1562), .B(n10875), .Z(n10873) );
  XOR U13955 ( .A(n10876), .B(n10877), .Z(n10875) );
  XOR U13956 ( .A(DB[847]), .B(DB[840]), .Z(n10877) );
  AND U13957 ( .A(n1566), .B(n10878), .Z(n10876) );
  XOR U13958 ( .A(n10879), .B(n10880), .Z(n10878) );
  XOR U13959 ( .A(DB[840]), .B(DB[833]), .Z(n10880) );
  AND U13960 ( .A(n1570), .B(n10881), .Z(n10879) );
  XOR U13961 ( .A(n10882), .B(n10883), .Z(n10881) );
  XOR U13962 ( .A(DB[833]), .B(DB[826]), .Z(n10883) );
  AND U13963 ( .A(n1574), .B(n10884), .Z(n10882) );
  XOR U13964 ( .A(n10885), .B(n10886), .Z(n10884) );
  XOR U13965 ( .A(DB[826]), .B(DB[819]), .Z(n10886) );
  AND U13966 ( .A(n1578), .B(n10887), .Z(n10885) );
  XOR U13967 ( .A(n10888), .B(n10889), .Z(n10887) );
  XOR U13968 ( .A(DB[819]), .B(DB[812]), .Z(n10889) );
  AND U13969 ( .A(n1582), .B(n10890), .Z(n10888) );
  XOR U13970 ( .A(n10891), .B(n10892), .Z(n10890) );
  XOR U13971 ( .A(DB[812]), .B(DB[805]), .Z(n10892) );
  AND U13972 ( .A(n1586), .B(n10893), .Z(n10891) );
  XOR U13973 ( .A(n10894), .B(n10895), .Z(n10893) );
  XOR U13974 ( .A(DB[805]), .B(DB[798]), .Z(n10895) );
  AND U13975 ( .A(n1590), .B(n10896), .Z(n10894) );
  XOR U13976 ( .A(n10897), .B(n10898), .Z(n10896) );
  XOR U13977 ( .A(DB[798]), .B(DB[791]), .Z(n10898) );
  AND U13978 ( .A(n1594), .B(n10899), .Z(n10897) );
  XOR U13979 ( .A(n10900), .B(n10901), .Z(n10899) );
  XOR U13980 ( .A(DB[791]), .B(DB[784]), .Z(n10901) );
  AND U13981 ( .A(n1598), .B(n10902), .Z(n10900) );
  XOR U13982 ( .A(n10903), .B(n10904), .Z(n10902) );
  XOR U13983 ( .A(DB[784]), .B(DB[777]), .Z(n10904) );
  AND U13984 ( .A(n1602), .B(n10905), .Z(n10903) );
  XOR U13985 ( .A(n10906), .B(n10907), .Z(n10905) );
  XOR U13986 ( .A(DB[777]), .B(DB[770]), .Z(n10907) );
  AND U13987 ( .A(n1606), .B(n10908), .Z(n10906) );
  XOR U13988 ( .A(n10909), .B(n10910), .Z(n10908) );
  XOR U13989 ( .A(DB[770]), .B(DB[763]), .Z(n10910) );
  AND U13990 ( .A(n1610), .B(n10911), .Z(n10909) );
  XOR U13991 ( .A(n10912), .B(n10913), .Z(n10911) );
  XOR U13992 ( .A(DB[763]), .B(DB[756]), .Z(n10913) );
  AND U13993 ( .A(n1614), .B(n10914), .Z(n10912) );
  XOR U13994 ( .A(n10915), .B(n10916), .Z(n10914) );
  XOR U13995 ( .A(DB[756]), .B(DB[749]), .Z(n10916) );
  AND U13996 ( .A(n1618), .B(n10917), .Z(n10915) );
  XOR U13997 ( .A(n10918), .B(n10919), .Z(n10917) );
  XOR U13998 ( .A(DB[749]), .B(DB[742]), .Z(n10919) );
  AND U13999 ( .A(n1622), .B(n10920), .Z(n10918) );
  XOR U14000 ( .A(n10921), .B(n10922), .Z(n10920) );
  XOR U14001 ( .A(DB[742]), .B(DB[735]), .Z(n10922) );
  AND U14002 ( .A(n1626), .B(n10923), .Z(n10921) );
  XOR U14003 ( .A(n10924), .B(n10925), .Z(n10923) );
  XOR U14004 ( .A(DB[735]), .B(DB[728]), .Z(n10925) );
  AND U14005 ( .A(n1630), .B(n10926), .Z(n10924) );
  XOR U14006 ( .A(n10927), .B(n10928), .Z(n10926) );
  XOR U14007 ( .A(DB[728]), .B(DB[721]), .Z(n10928) );
  AND U14008 ( .A(n1634), .B(n10929), .Z(n10927) );
  XOR U14009 ( .A(n10930), .B(n10931), .Z(n10929) );
  XOR U14010 ( .A(DB[721]), .B(DB[714]), .Z(n10931) );
  AND U14011 ( .A(n1638), .B(n10932), .Z(n10930) );
  XOR U14012 ( .A(n10933), .B(n10934), .Z(n10932) );
  XOR U14013 ( .A(DB[714]), .B(DB[707]), .Z(n10934) );
  AND U14014 ( .A(n1642), .B(n10935), .Z(n10933) );
  XOR U14015 ( .A(n10936), .B(n10937), .Z(n10935) );
  XOR U14016 ( .A(DB[707]), .B(DB[700]), .Z(n10937) );
  AND U14017 ( .A(n1646), .B(n10938), .Z(n10936) );
  XOR U14018 ( .A(n10939), .B(n10940), .Z(n10938) );
  XOR U14019 ( .A(DB[700]), .B(DB[693]), .Z(n10940) );
  AND U14020 ( .A(n1650), .B(n10941), .Z(n10939) );
  XOR U14021 ( .A(n10942), .B(n10943), .Z(n10941) );
  XOR U14022 ( .A(DB[693]), .B(DB[686]), .Z(n10943) );
  AND U14023 ( .A(n1654), .B(n10944), .Z(n10942) );
  XOR U14024 ( .A(n10945), .B(n10946), .Z(n10944) );
  XOR U14025 ( .A(DB[686]), .B(DB[679]), .Z(n10946) );
  AND U14026 ( .A(n1658), .B(n10947), .Z(n10945) );
  XOR U14027 ( .A(n10948), .B(n10949), .Z(n10947) );
  XOR U14028 ( .A(DB[679]), .B(DB[672]), .Z(n10949) );
  AND U14029 ( .A(n1662), .B(n10950), .Z(n10948) );
  XOR U14030 ( .A(n10951), .B(n10952), .Z(n10950) );
  XOR U14031 ( .A(DB[672]), .B(DB[665]), .Z(n10952) );
  AND U14032 ( .A(n1666), .B(n10953), .Z(n10951) );
  XOR U14033 ( .A(n10954), .B(n10955), .Z(n10953) );
  XOR U14034 ( .A(DB[665]), .B(DB[658]), .Z(n10955) );
  AND U14035 ( .A(n1670), .B(n10956), .Z(n10954) );
  XOR U14036 ( .A(n10957), .B(n10958), .Z(n10956) );
  XOR U14037 ( .A(DB[658]), .B(DB[651]), .Z(n10958) );
  AND U14038 ( .A(n1674), .B(n10959), .Z(n10957) );
  XOR U14039 ( .A(n10960), .B(n10961), .Z(n10959) );
  XOR U14040 ( .A(DB[651]), .B(DB[644]), .Z(n10961) );
  AND U14041 ( .A(n1678), .B(n10962), .Z(n10960) );
  XOR U14042 ( .A(n10963), .B(n10964), .Z(n10962) );
  XOR U14043 ( .A(DB[644]), .B(DB[637]), .Z(n10964) );
  AND U14044 ( .A(n1682), .B(n10965), .Z(n10963) );
  XOR U14045 ( .A(n10966), .B(n10967), .Z(n10965) );
  XOR U14046 ( .A(DB[637]), .B(DB[630]), .Z(n10967) );
  AND U14047 ( .A(n1686), .B(n10968), .Z(n10966) );
  XOR U14048 ( .A(n10969), .B(n10970), .Z(n10968) );
  XOR U14049 ( .A(DB[630]), .B(DB[623]), .Z(n10970) );
  AND U14050 ( .A(n1690), .B(n10971), .Z(n10969) );
  XOR U14051 ( .A(n10972), .B(n10973), .Z(n10971) );
  XOR U14052 ( .A(DB[623]), .B(DB[616]), .Z(n10973) );
  AND U14053 ( .A(n1694), .B(n10974), .Z(n10972) );
  XOR U14054 ( .A(n10975), .B(n10976), .Z(n10974) );
  XOR U14055 ( .A(DB[616]), .B(DB[609]), .Z(n10976) );
  AND U14056 ( .A(n1698), .B(n10977), .Z(n10975) );
  XOR U14057 ( .A(n10978), .B(n10979), .Z(n10977) );
  XOR U14058 ( .A(DB[609]), .B(DB[602]), .Z(n10979) );
  AND U14059 ( .A(n1702), .B(n10980), .Z(n10978) );
  XOR U14060 ( .A(n10981), .B(n10982), .Z(n10980) );
  XOR U14061 ( .A(DB[602]), .B(DB[595]), .Z(n10982) );
  AND U14062 ( .A(n1706), .B(n10983), .Z(n10981) );
  XOR U14063 ( .A(n10984), .B(n10985), .Z(n10983) );
  XOR U14064 ( .A(DB[595]), .B(DB[588]), .Z(n10985) );
  AND U14065 ( .A(n1710), .B(n10986), .Z(n10984) );
  XOR U14066 ( .A(n10987), .B(n10988), .Z(n10986) );
  XOR U14067 ( .A(DB[588]), .B(DB[581]), .Z(n10988) );
  AND U14068 ( .A(n1714), .B(n10989), .Z(n10987) );
  XOR U14069 ( .A(n10990), .B(n10991), .Z(n10989) );
  XOR U14070 ( .A(DB[581]), .B(DB[574]), .Z(n10991) );
  AND U14071 ( .A(n1718), .B(n10992), .Z(n10990) );
  XOR U14072 ( .A(n10993), .B(n10994), .Z(n10992) );
  XOR U14073 ( .A(DB[574]), .B(DB[567]), .Z(n10994) );
  AND U14074 ( .A(n1722), .B(n10995), .Z(n10993) );
  XOR U14075 ( .A(n10996), .B(n10997), .Z(n10995) );
  XOR U14076 ( .A(DB[567]), .B(DB[560]), .Z(n10997) );
  AND U14077 ( .A(n1726), .B(n10998), .Z(n10996) );
  XOR U14078 ( .A(n10999), .B(n11000), .Z(n10998) );
  XOR U14079 ( .A(DB[560]), .B(DB[553]), .Z(n11000) );
  AND U14080 ( .A(n1730), .B(n11001), .Z(n10999) );
  XOR U14081 ( .A(n11002), .B(n11003), .Z(n11001) );
  XOR U14082 ( .A(DB[553]), .B(DB[546]), .Z(n11003) );
  AND U14083 ( .A(n1734), .B(n11004), .Z(n11002) );
  XOR U14084 ( .A(n11005), .B(n11006), .Z(n11004) );
  XOR U14085 ( .A(DB[546]), .B(DB[539]), .Z(n11006) );
  AND U14086 ( .A(n1738), .B(n11007), .Z(n11005) );
  XOR U14087 ( .A(n11008), .B(n11009), .Z(n11007) );
  XOR U14088 ( .A(DB[539]), .B(DB[532]), .Z(n11009) );
  AND U14089 ( .A(n1742), .B(n11010), .Z(n11008) );
  XOR U14090 ( .A(n11011), .B(n11012), .Z(n11010) );
  XOR U14091 ( .A(DB[532]), .B(DB[525]), .Z(n11012) );
  AND U14092 ( .A(n1746), .B(n11013), .Z(n11011) );
  XOR U14093 ( .A(n11014), .B(n11015), .Z(n11013) );
  XOR U14094 ( .A(DB[525]), .B(DB[518]), .Z(n11015) );
  AND U14095 ( .A(n1750), .B(n11016), .Z(n11014) );
  XOR U14096 ( .A(n11017), .B(n11018), .Z(n11016) );
  XOR U14097 ( .A(DB[518]), .B(DB[511]), .Z(n11018) );
  AND U14098 ( .A(n1754), .B(n11019), .Z(n11017) );
  XOR U14099 ( .A(n11020), .B(n11021), .Z(n11019) );
  XOR U14100 ( .A(DB[511]), .B(DB[504]), .Z(n11021) );
  AND U14101 ( .A(n1758), .B(n11022), .Z(n11020) );
  XOR U14102 ( .A(n11023), .B(n11024), .Z(n11022) );
  XOR U14103 ( .A(DB[504]), .B(DB[497]), .Z(n11024) );
  AND U14104 ( .A(n1762), .B(n11025), .Z(n11023) );
  XOR U14105 ( .A(n11026), .B(n11027), .Z(n11025) );
  XOR U14106 ( .A(DB[497]), .B(DB[490]), .Z(n11027) );
  AND U14107 ( .A(n1766), .B(n11028), .Z(n11026) );
  XOR U14108 ( .A(n11029), .B(n11030), .Z(n11028) );
  XOR U14109 ( .A(DB[490]), .B(DB[483]), .Z(n11030) );
  AND U14110 ( .A(n1770), .B(n11031), .Z(n11029) );
  XOR U14111 ( .A(n11032), .B(n11033), .Z(n11031) );
  XOR U14112 ( .A(DB[483]), .B(DB[476]), .Z(n11033) );
  AND U14113 ( .A(n1774), .B(n11034), .Z(n11032) );
  XOR U14114 ( .A(n11035), .B(n11036), .Z(n11034) );
  XOR U14115 ( .A(DB[476]), .B(DB[469]), .Z(n11036) );
  AND U14116 ( .A(n1778), .B(n11037), .Z(n11035) );
  XOR U14117 ( .A(n11038), .B(n11039), .Z(n11037) );
  XOR U14118 ( .A(DB[469]), .B(DB[462]), .Z(n11039) );
  AND U14119 ( .A(n1782), .B(n11040), .Z(n11038) );
  XOR U14120 ( .A(n11041), .B(n11042), .Z(n11040) );
  XOR U14121 ( .A(DB[462]), .B(DB[455]), .Z(n11042) );
  AND U14122 ( .A(n1786), .B(n11043), .Z(n11041) );
  XOR U14123 ( .A(n11044), .B(n11045), .Z(n11043) );
  XOR U14124 ( .A(DB[455]), .B(DB[448]), .Z(n11045) );
  AND U14125 ( .A(n1790), .B(n11046), .Z(n11044) );
  XOR U14126 ( .A(n11047), .B(n11048), .Z(n11046) );
  XOR U14127 ( .A(DB[448]), .B(DB[441]), .Z(n11048) );
  AND U14128 ( .A(n1794), .B(n11049), .Z(n11047) );
  XOR U14129 ( .A(n11050), .B(n11051), .Z(n11049) );
  XOR U14130 ( .A(DB[441]), .B(DB[434]), .Z(n11051) );
  AND U14131 ( .A(n1798), .B(n11052), .Z(n11050) );
  XOR U14132 ( .A(n11053), .B(n11054), .Z(n11052) );
  XOR U14133 ( .A(DB[434]), .B(DB[427]), .Z(n11054) );
  AND U14134 ( .A(n1802), .B(n11055), .Z(n11053) );
  XOR U14135 ( .A(n11056), .B(n11057), .Z(n11055) );
  XOR U14136 ( .A(DB[427]), .B(DB[420]), .Z(n11057) );
  AND U14137 ( .A(n1806), .B(n11058), .Z(n11056) );
  XOR U14138 ( .A(n11059), .B(n11060), .Z(n11058) );
  XOR U14139 ( .A(DB[420]), .B(DB[413]), .Z(n11060) );
  AND U14140 ( .A(n1810), .B(n11061), .Z(n11059) );
  XOR U14141 ( .A(n11062), .B(n11063), .Z(n11061) );
  XOR U14142 ( .A(DB[413]), .B(DB[406]), .Z(n11063) );
  AND U14143 ( .A(n1814), .B(n11064), .Z(n11062) );
  XOR U14144 ( .A(n11065), .B(n11066), .Z(n11064) );
  XOR U14145 ( .A(DB[406]), .B(DB[399]), .Z(n11066) );
  AND U14146 ( .A(n1818), .B(n11067), .Z(n11065) );
  XOR U14147 ( .A(n11068), .B(n11069), .Z(n11067) );
  XOR U14148 ( .A(DB[399]), .B(DB[392]), .Z(n11069) );
  AND U14149 ( .A(n1822), .B(n11070), .Z(n11068) );
  XOR U14150 ( .A(n11071), .B(n11072), .Z(n11070) );
  XOR U14151 ( .A(DB[392]), .B(DB[385]), .Z(n11072) );
  AND U14152 ( .A(n1826), .B(n11073), .Z(n11071) );
  XOR U14153 ( .A(n11074), .B(n11075), .Z(n11073) );
  XOR U14154 ( .A(DB[385]), .B(DB[378]), .Z(n11075) );
  AND U14155 ( .A(n1830), .B(n11076), .Z(n11074) );
  XOR U14156 ( .A(n11077), .B(n11078), .Z(n11076) );
  XOR U14157 ( .A(DB[378]), .B(DB[371]), .Z(n11078) );
  AND U14158 ( .A(n1834), .B(n11079), .Z(n11077) );
  XOR U14159 ( .A(n11080), .B(n11081), .Z(n11079) );
  XOR U14160 ( .A(DB[371]), .B(DB[364]), .Z(n11081) );
  AND U14161 ( .A(n1838), .B(n11082), .Z(n11080) );
  XOR U14162 ( .A(n11083), .B(n11084), .Z(n11082) );
  XOR U14163 ( .A(DB[364]), .B(DB[357]), .Z(n11084) );
  AND U14164 ( .A(n1842), .B(n11085), .Z(n11083) );
  XOR U14165 ( .A(n11086), .B(n11087), .Z(n11085) );
  XOR U14166 ( .A(DB[357]), .B(DB[350]), .Z(n11087) );
  AND U14167 ( .A(n1846), .B(n11088), .Z(n11086) );
  XOR U14168 ( .A(n11089), .B(n11090), .Z(n11088) );
  XOR U14169 ( .A(DB[350]), .B(DB[343]), .Z(n11090) );
  AND U14170 ( .A(n1850), .B(n11091), .Z(n11089) );
  XOR U14171 ( .A(n11092), .B(n11093), .Z(n11091) );
  XOR U14172 ( .A(DB[343]), .B(DB[336]), .Z(n11093) );
  AND U14173 ( .A(n1854), .B(n11094), .Z(n11092) );
  XOR U14174 ( .A(n11095), .B(n11096), .Z(n11094) );
  XOR U14175 ( .A(DB[336]), .B(DB[329]), .Z(n11096) );
  AND U14176 ( .A(n1858), .B(n11097), .Z(n11095) );
  XOR U14177 ( .A(n11098), .B(n11099), .Z(n11097) );
  XOR U14178 ( .A(DB[329]), .B(DB[322]), .Z(n11099) );
  AND U14179 ( .A(n1862), .B(n11100), .Z(n11098) );
  XOR U14180 ( .A(n11101), .B(n11102), .Z(n11100) );
  XOR U14181 ( .A(DB[322]), .B(DB[315]), .Z(n11102) );
  AND U14182 ( .A(n1866), .B(n11103), .Z(n11101) );
  XOR U14183 ( .A(n11104), .B(n11105), .Z(n11103) );
  XOR U14184 ( .A(DB[315]), .B(DB[308]), .Z(n11105) );
  AND U14185 ( .A(n1870), .B(n11106), .Z(n11104) );
  XOR U14186 ( .A(n11107), .B(n11108), .Z(n11106) );
  XOR U14187 ( .A(DB[308]), .B(DB[301]), .Z(n11108) );
  AND U14188 ( .A(n1874), .B(n11109), .Z(n11107) );
  XOR U14189 ( .A(n11110), .B(n11111), .Z(n11109) );
  XOR U14190 ( .A(DB[301]), .B(DB[294]), .Z(n11111) );
  AND U14191 ( .A(n1878), .B(n11112), .Z(n11110) );
  XOR U14192 ( .A(n11113), .B(n11114), .Z(n11112) );
  XOR U14193 ( .A(DB[294]), .B(DB[287]), .Z(n11114) );
  AND U14194 ( .A(n1882), .B(n11115), .Z(n11113) );
  XOR U14195 ( .A(n11116), .B(n11117), .Z(n11115) );
  XOR U14196 ( .A(DB[287]), .B(DB[280]), .Z(n11117) );
  AND U14197 ( .A(n1886), .B(n11118), .Z(n11116) );
  XOR U14198 ( .A(n11119), .B(n11120), .Z(n11118) );
  XOR U14199 ( .A(DB[280]), .B(DB[273]), .Z(n11120) );
  AND U14200 ( .A(n1890), .B(n11121), .Z(n11119) );
  XOR U14201 ( .A(n11122), .B(n11123), .Z(n11121) );
  XOR U14202 ( .A(DB[273]), .B(DB[266]), .Z(n11123) );
  AND U14203 ( .A(n1894), .B(n11124), .Z(n11122) );
  XOR U14204 ( .A(n11125), .B(n11126), .Z(n11124) );
  XOR U14205 ( .A(DB[266]), .B(DB[259]), .Z(n11126) );
  AND U14206 ( .A(n1898), .B(n11127), .Z(n11125) );
  XOR U14207 ( .A(n11128), .B(n11129), .Z(n11127) );
  XOR U14208 ( .A(DB[259]), .B(DB[252]), .Z(n11129) );
  AND U14209 ( .A(n1902), .B(n11130), .Z(n11128) );
  XOR U14210 ( .A(n11131), .B(n11132), .Z(n11130) );
  XOR U14211 ( .A(DB[252]), .B(DB[245]), .Z(n11132) );
  AND U14212 ( .A(n1906), .B(n11133), .Z(n11131) );
  XOR U14213 ( .A(n11134), .B(n11135), .Z(n11133) );
  XOR U14214 ( .A(DB[245]), .B(DB[238]), .Z(n11135) );
  AND U14215 ( .A(n1910), .B(n11136), .Z(n11134) );
  XOR U14216 ( .A(n11137), .B(n11138), .Z(n11136) );
  XOR U14217 ( .A(DB[238]), .B(DB[231]), .Z(n11138) );
  AND U14218 ( .A(n1914), .B(n11139), .Z(n11137) );
  XOR U14219 ( .A(n11140), .B(n11141), .Z(n11139) );
  XOR U14220 ( .A(DB[231]), .B(DB[224]), .Z(n11141) );
  AND U14221 ( .A(n1918), .B(n11142), .Z(n11140) );
  XOR U14222 ( .A(n11143), .B(n11144), .Z(n11142) );
  XOR U14223 ( .A(DB[224]), .B(DB[217]), .Z(n11144) );
  AND U14224 ( .A(n1922), .B(n11145), .Z(n11143) );
  XOR U14225 ( .A(n11146), .B(n11147), .Z(n11145) );
  XOR U14226 ( .A(DB[217]), .B(DB[210]), .Z(n11147) );
  AND U14227 ( .A(n1926), .B(n11148), .Z(n11146) );
  XOR U14228 ( .A(n11149), .B(n11150), .Z(n11148) );
  XOR U14229 ( .A(DB[210]), .B(DB[203]), .Z(n11150) );
  AND U14230 ( .A(n1930), .B(n11151), .Z(n11149) );
  XOR U14231 ( .A(n11152), .B(n11153), .Z(n11151) );
  XOR U14232 ( .A(DB[203]), .B(DB[196]), .Z(n11153) );
  AND U14233 ( .A(n1934), .B(n11154), .Z(n11152) );
  XOR U14234 ( .A(n11155), .B(n11156), .Z(n11154) );
  XOR U14235 ( .A(DB[196]), .B(DB[189]), .Z(n11156) );
  AND U14236 ( .A(n1938), .B(n11157), .Z(n11155) );
  XOR U14237 ( .A(n11158), .B(n11159), .Z(n11157) );
  XOR U14238 ( .A(DB[189]), .B(DB[182]), .Z(n11159) );
  AND U14239 ( .A(n1942), .B(n11160), .Z(n11158) );
  XOR U14240 ( .A(n11161), .B(n11162), .Z(n11160) );
  XOR U14241 ( .A(DB[182]), .B(DB[175]), .Z(n11162) );
  AND U14242 ( .A(n1946), .B(n11163), .Z(n11161) );
  XOR U14243 ( .A(n11164), .B(n11165), .Z(n11163) );
  XOR U14244 ( .A(DB[175]), .B(DB[168]), .Z(n11165) );
  AND U14245 ( .A(n1950), .B(n11166), .Z(n11164) );
  XOR U14246 ( .A(n11167), .B(n11168), .Z(n11166) );
  XOR U14247 ( .A(DB[168]), .B(DB[161]), .Z(n11168) );
  AND U14248 ( .A(n1954), .B(n11169), .Z(n11167) );
  XOR U14249 ( .A(n11170), .B(n11171), .Z(n11169) );
  XOR U14250 ( .A(DB[161]), .B(DB[154]), .Z(n11171) );
  AND U14251 ( .A(n1958), .B(n11172), .Z(n11170) );
  XOR U14252 ( .A(n11173), .B(n11174), .Z(n11172) );
  XOR U14253 ( .A(DB[154]), .B(DB[147]), .Z(n11174) );
  AND U14254 ( .A(n1962), .B(n11175), .Z(n11173) );
  XOR U14255 ( .A(n11176), .B(n11177), .Z(n11175) );
  XOR U14256 ( .A(DB[147]), .B(DB[140]), .Z(n11177) );
  AND U14257 ( .A(n1966), .B(n11178), .Z(n11176) );
  XOR U14258 ( .A(n11179), .B(n11180), .Z(n11178) );
  XOR U14259 ( .A(DB[140]), .B(DB[133]), .Z(n11180) );
  AND U14260 ( .A(n1970), .B(n11181), .Z(n11179) );
  XOR U14261 ( .A(n11182), .B(n11183), .Z(n11181) );
  XOR U14262 ( .A(DB[133]), .B(DB[126]), .Z(n11183) );
  AND U14263 ( .A(n1974), .B(n11184), .Z(n11182) );
  XOR U14264 ( .A(n11185), .B(n11186), .Z(n11184) );
  XOR U14265 ( .A(DB[126]), .B(DB[119]), .Z(n11186) );
  AND U14266 ( .A(n1978), .B(n11187), .Z(n11185) );
  XOR U14267 ( .A(n11188), .B(n11189), .Z(n11187) );
  XOR U14268 ( .A(DB[119]), .B(DB[112]), .Z(n11189) );
  AND U14269 ( .A(n1982), .B(n11190), .Z(n11188) );
  XOR U14270 ( .A(n11191), .B(n11192), .Z(n11190) );
  XOR U14271 ( .A(DB[112]), .B(DB[105]), .Z(n11192) );
  AND U14272 ( .A(n1986), .B(n11193), .Z(n11191) );
  XOR U14273 ( .A(n11194), .B(n11195), .Z(n11193) );
  XOR U14274 ( .A(DB[98]), .B(DB[105]), .Z(n11195) );
  AND U14275 ( .A(n1990), .B(n11196), .Z(n11194) );
  XOR U14276 ( .A(n11197), .B(n11198), .Z(n11196) );
  XOR U14277 ( .A(DB[98]), .B(DB[91]), .Z(n11198) );
  AND U14278 ( .A(n1994), .B(n11199), .Z(n11197) );
  XOR U14279 ( .A(n11200), .B(n11201), .Z(n11199) );
  XOR U14280 ( .A(DB[91]), .B(DB[84]), .Z(n11201) );
  AND U14281 ( .A(n1998), .B(n11202), .Z(n11200) );
  XOR U14282 ( .A(n11203), .B(n11204), .Z(n11202) );
  XOR U14283 ( .A(DB[84]), .B(DB[77]), .Z(n11204) );
  AND U14284 ( .A(n2002), .B(n11205), .Z(n11203) );
  XOR U14285 ( .A(n11206), .B(n11207), .Z(n11205) );
  XOR U14286 ( .A(DB[77]), .B(DB[70]), .Z(n11207) );
  AND U14287 ( .A(n2006), .B(n11208), .Z(n11206) );
  XOR U14288 ( .A(n11209), .B(n11210), .Z(n11208) );
  XOR U14289 ( .A(DB[70]), .B(DB[63]), .Z(n11210) );
  AND U14290 ( .A(n2010), .B(n11211), .Z(n11209) );
  XOR U14291 ( .A(n11212), .B(n11213), .Z(n11211) );
  XOR U14292 ( .A(DB[63]), .B(DB[56]), .Z(n11213) );
  AND U14293 ( .A(n2014), .B(n11214), .Z(n11212) );
  XOR U14294 ( .A(n11215), .B(n11216), .Z(n11214) );
  XOR U14295 ( .A(DB[56]), .B(DB[49]), .Z(n11216) );
  AND U14296 ( .A(n2018), .B(n11217), .Z(n11215) );
  XOR U14297 ( .A(n11218), .B(n11219), .Z(n11217) );
  XOR U14298 ( .A(DB[49]), .B(DB[42]), .Z(n11219) );
  AND U14299 ( .A(n2022), .B(n11220), .Z(n11218) );
  XOR U14300 ( .A(n11221), .B(n11222), .Z(n11220) );
  XOR U14301 ( .A(DB[42]), .B(DB[35]), .Z(n11222) );
  AND U14302 ( .A(n2026), .B(n11223), .Z(n11221) );
  XOR U14303 ( .A(n11224), .B(n11225), .Z(n11223) );
  XOR U14304 ( .A(DB[35]), .B(DB[28]), .Z(n11225) );
  AND U14305 ( .A(n2030), .B(n11226), .Z(n11224) );
  XOR U14306 ( .A(n11227), .B(n11228), .Z(n11226) );
  XOR U14307 ( .A(DB[28]), .B(DB[21]), .Z(n11228) );
  AND U14308 ( .A(n2034), .B(n11229), .Z(n11227) );
  XOR U14309 ( .A(n11230), .B(n11231), .Z(n11229) );
  XOR U14310 ( .A(DB[21]), .B(DB[14]), .Z(n11231) );
  AND U14311 ( .A(n2038), .B(n11232), .Z(n11230) );
  XOR U14312 ( .A(n11233), .B(n11234), .Z(n11232) );
  XOR U14313 ( .A(DB[7]), .B(DB[14]), .Z(n11234) );
  AND U14314 ( .A(n2042), .B(n11235), .Z(n11233) );
  XOR U14315 ( .A(DB[7]), .B(DB[0]), .Z(n11235) );
  XOR U14316 ( .A(n11236), .B(n11237), .Z(n2) );
  AND U14317 ( .A(n11238), .B(n11239), .Z(n11236) );
  XNOR U14318 ( .A(n11237), .B(n11240), .Z(n11239) );
  XOR U14319 ( .A(n11241), .B(n11242), .Z(n11240) );
  AND U14320 ( .A(n11243), .B(n11244), .Z(n11241) );
  XNOR U14321 ( .A(n11245), .B(n11246), .Z(n11244) );
  XNOR U14322 ( .A(n11237), .B(n11247), .Z(n11238) );
  XNOR U14323 ( .A(n11248), .B(n11249), .Z(n11247) );
  AND U14324 ( .A(n6), .B(n11250), .Z(n11248) );
  XOR U14325 ( .A(n11251), .B(n11249), .Z(n11250) );
  XNOR U14326 ( .A(n11252), .B(n11253), .Z(n11237) );
  NAND U14327 ( .A(n11254), .B(n11255), .Z(n11253) );
  XOR U14328 ( .A(n11243), .B(n11256), .Z(n11255) );
  XNOR U14329 ( .A(n11252), .B(n11245), .Z(n11256) );
  XOR U14330 ( .A(n11257), .B(n11258), .Z(n11245) );
  ANDN U14331 ( .B(n11259), .A(n11260), .Z(n11257) );
  XNOR U14332 ( .A(n11258), .B(n11261), .Z(n11259) );
  XNOR U14333 ( .A(n11242), .B(n11262), .Z(n11243) );
  XNOR U14334 ( .A(n11263), .B(n11264), .Z(n11262) );
  ANDN U14335 ( .B(n11265), .A(n11266), .Z(n11263) );
  XNOR U14336 ( .A(n11267), .B(n11268), .Z(n11265) );
  IV U14337 ( .A(n11264), .Z(n11268) );
  IV U14338 ( .A(n11246), .Z(n11242) );
  XNOR U14339 ( .A(n11269), .B(n11270), .Z(n11246) );
  AND U14340 ( .A(n11271), .B(n11272), .Z(n11269) );
  XNOR U14341 ( .A(n11270), .B(n11273), .Z(n11272) );
  XOR U14342 ( .A(n11274), .B(n11275), .Z(n11254) );
  XNOR U14343 ( .A(n11252), .B(n11276), .Z(n11275) );
  NAND U14344 ( .A(n11277), .B(n6), .Z(n11276) );
  XOR U14345 ( .A(n11278), .B(n11274), .Z(n11277) );
  NAND U14346 ( .A(n11279), .B(n11280), .Z(n11252) );
  XNOR U14347 ( .A(n11271), .B(n11273), .Z(n11280) );
  XOR U14348 ( .A(n11281), .B(n11261), .Z(n11273) );
  XNOR U14349 ( .A(q[6]), .B(DB[3583]), .Z(n11261) );
  IV U14350 ( .A(n11260), .Z(n11281) );
  XOR U14351 ( .A(n11258), .B(n11282), .Z(n11260) );
  XNOR U14352 ( .A(q[5]), .B(DB[3582]), .Z(n11282) );
  XOR U14353 ( .A(q[4]), .B(DB[3581]), .Z(n11258) );
  XNOR U14354 ( .A(n11283), .B(n11284), .Z(n11271) );
  XNOR U14355 ( .A(n11267), .B(n11270), .Z(n11284) );
  XOR U14356 ( .A(q[0]), .B(DB[3577]), .Z(n11270) );
  XOR U14357 ( .A(q[3]), .B(DB[3580]), .Z(n11267) );
  IV U14358 ( .A(n11266), .Z(n11283) );
  XOR U14359 ( .A(n11264), .B(n11285), .Z(n11266) );
  XNOR U14360 ( .A(q[2]), .B(DB[3579]), .Z(n11285) );
  XOR U14361 ( .A(q[1]), .B(DB[3578]), .Z(n11264) );
  XOR U14362 ( .A(n11286), .B(n11287), .Z(n11279) );
  AND U14363 ( .A(n6), .B(n11288), .Z(n11286) );
  XOR U14364 ( .A(n11287), .B(n11289), .Z(n11288) );
  XOR U14365 ( .A(n11290), .B(n11291), .Z(n6) );
  AND U14366 ( .A(n11292), .B(n11293), .Z(n11290) );
  XNOR U14367 ( .A(n11291), .B(n11249), .Z(n11293) );
  XNOR U14368 ( .A(n11294), .B(n11295), .Z(n11249) );
  ANDN U14369 ( .B(n11296), .A(n11297), .Z(n11294) );
  XOR U14370 ( .A(n11295), .B(n11298), .Z(n11296) );
  XOR U14371 ( .A(n11291), .B(n11251), .Z(n11292) );
  XOR U14372 ( .A(n11299), .B(n11300), .Z(n11251) );
  AND U14373 ( .A(n10), .B(n11301), .Z(n11299) );
  XOR U14374 ( .A(n11302), .B(n11300), .Z(n11301) );
  XNOR U14375 ( .A(n11303), .B(n11304), .Z(n11291) );
  NAND U14376 ( .A(n11305), .B(n11306), .Z(n11304) );
  XOR U14377 ( .A(n11307), .B(n11274), .Z(n11306) );
  XNOR U14378 ( .A(n11308), .B(n11298), .Z(n11274) );
  XOR U14379 ( .A(n11309), .B(n11310), .Z(n11298) );
  ANDN U14380 ( .B(n11311), .A(n11312), .Z(n11309) );
  XOR U14381 ( .A(n11310), .B(n11313), .Z(n11311) );
  IV U14382 ( .A(n11297), .Z(n11308) );
  XOR U14383 ( .A(n11314), .B(n11315), .Z(n11297) );
  XOR U14384 ( .A(n11316), .B(n11317), .Z(n11315) );
  ANDN U14385 ( .B(n11318), .A(n11319), .Z(n11316) );
  XOR U14386 ( .A(n11320), .B(n11317), .Z(n11318) );
  IV U14387 ( .A(n11295), .Z(n11314) );
  XOR U14388 ( .A(n11321), .B(n11322), .Z(n11295) );
  ANDN U14389 ( .B(n11323), .A(n11324), .Z(n11321) );
  XOR U14390 ( .A(n11322), .B(n11325), .Z(n11323) );
  IV U14391 ( .A(n11303), .Z(n11307) );
  XOR U14392 ( .A(n11303), .B(n11278), .Z(n11305) );
  XOR U14393 ( .A(n11326), .B(n11327), .Z(n11278) );
  AND U14394 ( .A(n10), .B(n11328), .Z(n11326) );
  XOR U14395 ( .A(n11329), .B(n11327), .Z(n11328) );
  NANDN U14396 ( .A(n11287), .B(n11289), .Z(n11303) );
  XOR U14397 ( .A(n11330), .B(n11331), .Z(n11289) );
  AND U14398 ( .A(n10), .B(n11332), .Z(n11330) );
  XOR U14399 ( .A(n11331), .B(n11333), .Z(n11332) );
  XOR U14400 ( .A(n11334), .B(n11335), .Z(n10) );
  AND U14401 ( .A(n11336), .B(n11337), .Z(n11334) );
  XNOR U14402 ( .A(n11335), .B(n11300), .Z(n11337) );
  XNOR U14403 ( .A(n11338), .B(n11339), .Z(n11300) );
  ANDN U14404 ( .B(n11340), .A(n11341), .Z(n11338) );
  XOR U14405 ( .A(n11339), .B(n11342), .Z(n11340) );
  XOR U14406 ( .A(n11335), .B(n11302), .Z(n11336) );
  XOR U14407 ( .A(n11343), .B(n11344), .Z(n11302) );
  AND U14408 ( .A(n14), .B(n11345), .Z(n11343) );
  XOR U14409 ( .A(n11346), .B(n11344), .Z(n11345) );
  XNOR U14410 ( .A(n11347), .B(n11348), .Z(n11335) );
  NAND U14411 ( .A(n11349), .B(n11350), .Z(n11348) );
  XOR U14412 ( .A(n11351), .B(n11327), .Z(n11350) );
  XOR U14413 ( .A(n11341), .B(n11342), .Z(n11327) );
  XOR U14414 ( .A(n11352), .B(n11353), .Z(n11342) );
  ANDN U14415 ( .B(n11354), .A(n11355), .Z(n11352) );
  XOR U14416 ( .A(n11353), .B(n11356), .Z(n11354) );
  XOR U14417 ( .A(n11357), .B(n11358), .Z(n11341) );
  XOR U14418 ( .A(n11359), .B(n11360), .Z(n11358) );
  ANDN U14419 ( .B(n11361), .A(n11362), .Z(n11359) );
  XOR U14420 ( .A(n11363), .B(n11360), .Z(n11361) );
  IV U14421 ( .A(n11339), .Z(n11357) );
  XOR U14422 ( .A(n11364), .B(n11365), .Z(n11339) );
  ANDN U14423 ( .B(n11366), .A(n11367), .Z(n11364) );
  XOR U14424 ( .A(n11365), .B(n11368), .Z(n11366) );
  IV U14425 ( .A(n11347), .Z(n11351) );
  XOR U14426 ( .A(n11347), .B(n11329), .Z(n11349) );
  XOR U14427 ( .A(n11369), .B(n11370), .Z(n11329) );
  AND U14428 ( .A(n14), .B(n11371), .Z(n11369) );
  XOR U14429 ( .A(n11372), .B(n11370), .Z(n11371) );
  NANDN U14430 ( .A(n11331), .B(n11333), .Z(n11347) );
  XOR U14431 ( .A(n11373), .B(n11374), .Z(n11333) );
  AND U14432 ( .A(n14), .B(n11375), .Z(n11373) );
  XOR U14433 ( .A(n11374), .B(n11376), .Z(n11375) );
  XOR U14434 ( .A(n11377), .B(n11378), .Z(n14) );
  AND U14435 ( .A(n11379), .B(n11380), .Z(n11377) );
  XNOR U14436 ( .A(n11378), .B(n11344), .Z(n11380) );
  XNOR U14437 ( .A(n11381), .B(n11382), .Z(n11344) );
  ANDN U14438 ( .B(n11383), .A(n11384), .Z(n11381) );
  XOR U14439 ( .A(n11382), .B(n11385), .Z(n11383) );
  XOR U14440 ( .A(n11378), .B(n11346), .Z(n11379) );
  XOR U14441 ( .A(n11386), .B(n11387), .Z(n11346) );
  AND U14442 ( .A(n18), .B(n11388), .Z(n11386) );
  XOR U14443 ( .A(n11389), .B(n11387), .Z(n11388) );
  XNOR U14444 ( .A(n11390), .B(n11391), .Z(n11378) );
  NAND U14445 ( .A(n11392), .B(n11393), .Z(n11391) );
  XOR U14446 ( .A(n11394), .B(n11370), .Z(n11393) );
  XOR U14447 ( .A(n11384), .B(n11385), .Z(n11370) );
  XOR U14448 ( .A(n11395), .B(n11396), .Z(n11385) );
  ANDN U14449 ( .B(n11397), .A(n11398), .Z(n11395) );
  XOR U14450 ( .A(n11396), .B(n11399), .Z(n11397) );
  XOR U14451 ( .A(n11400), .B(n11401), .Z(n11384) );
  XOR U14452 ( .A(n11402), .B(n11403), .Z(n11401) );
  ANDN U14453 ( .B(n11404), .A(n11405), .Z(n11402) );
  XOR U14454 ( .A(n11406), .B(n11403), .Z(n11404) );
  IV U14455 ( .A(n11382), .Z(n11400) );
  XOR U14456 ( .A(n11407), .B(n11408), .Z(n11382) );
  ANDN U14457 ( .B(n11409), .A(n11410), .Z(n11407) );
  XOR U14458 ( .A(n11408), .B(n11411), .Z(n11409) );
  IV U14459 ( .A(n11390), .Z(n11394) );
  XOR U14460 ( .A(n11390), .B(n11372), .Z(n11392) );
  XOR U14461 ( .A(n11412), .B(n11413), .Z(n11372) );
  AND U14462 ( .A(n18), .B(n11414), .Z(n11412) );
  XOR U14463 ( .A(n11415), .B(n11413), .Z(n11414) );
  NANDN U14464 ( .A(n11374), .B(n11376), .Z(n11390) );
  XOR U14465 ( .A(n11416), .B(n11417), .Z(n11376) );
  AND U14466 ( .A(n18), .B(n11418), .Z(n11416) );
  XOR U14467 ( .A(n11417), .B(n11419), .Z(n11418) );
  XOR U14468 ( .A(n11420), .B(n11421), .Z(n18) );
  AND U14469 ( .A(n11422), .B(n11423), .Z(n11420) );
  XNOR U14470 ( .A(n11421), .B(n11387), .Z(n11423) );
  XNOR U14471 ( .A(n11424), .B(n11425), .Z(n11387) );
  ANDN U14472 ( .B(n11426), .A(n11427), .Z(n11424) );
  XOR U14473 ( .A(n11425), .B(n11428), .Z(n11426) );
  XOR U14474 ( .A(n11421), .B(n11389), .Z(n11422) );
  XOR U14475 ( .A(n11429), .B(n11430), .Z(n11389) );
  AND U14476 ( .A(n22), .B(n11431), .Z(n11429) );
  XOR U14477 ( .A(n11432), .B(n11430), .Z(n11431) );
  XNOR U14478 ( .A(n11433), .B(n11434), .Z(n11421) );
  NAND U14479 ( .A(n11435), .B(n11436), .Z(n11434) );
  XOR U14480 ( .A(n11437), .B(n11413), .Z(n11436) );
  XOR U14481 ( .A(n11427), .B(n11428), .Z(n11413) );
  XOR U14482 ( .A(n11438), .B(n11439), .Z(n11428) );
  ANDN U14483 ( .B(n11440), .A(n11441), .Z(n11438) );
  XOR U14484 ( .A(n11439), .B(n11442), .Z(n11440) );
  XOR U14485 ( .A(n11443), .B(n11444), .Z(n11427) );
  XOR U14486 ( .A(n11445), .B(n11446), .Z(n11444) );
  ANDN U14487 ( .B(n11447), .A(n11448), .Z(n11445) );
  XOR U14488 ( .A(n11449), .B(n11446), .Z(n11447) );
  IV U14489 ( .A(n11425), .Z(n11443) );
  XOR U14490 ( .A(n11450), .B(n11451), .Z(n11425) );
  ANDN U14491 ( .B(n11452), .A(n11453), .Z(n11450) );
  XOR U14492 ( .A(n11451), .B(n11454), .Z(n11452) );
  IV U14493 ( .A(n11433), .Z(n11437) );
  XOR U14494 ( .A(n11433), .B(n11415), .Z(n11435) );
  XOR U14495 ( .A(n11455), .B(n11456), .Z(n11415) );
  AND U14496 ( .A(n22), .B(n11457), .Z(n11455) );
  XOR U14497 ( .A(n11458), .B(n11456), .Z(n11457) );
  NANDN U14498 ( .A(n11417), .B(n11419), .Z(n11433) );
  XOR U14499 ( .A(n11459), .B(n11460), .Z(n11419) );
  AND U14500 ( .A(n22), .B(n11461), .Z(n11459) );
  XOR U14501 ( .A(n11460), .B(n11462), .Z(n11461) );
  XOR U14502 ( .A(n11463), .B(n11464), .Z(n22) );
  AND U14503 ( .A(n11465), .B(n11466), .Z(n11463) );
  XNOR U14504 ( .A(n11464), .B(n11430), .Z(n11466) );
  XNOR U14505 ( .A(n11467), .B(n11468), .Z(n11430) );
  ANDN U14506 ( .B(n11469), .A(n11470), .Z(n11467) );
  XOR U14507 ( .A(n11468), .B(n11471), .Z(n11469) );
  XOR U14508 ( .A(n11464), .B(n11432), .Z(n11465) );
  XOR U14509 ( .A(n11472), .B(n11473), .Z(n11432) );
  AND U14510 ( .A(n26), .B(n11474), .Z(n11472) );
  XOR U14511 ( .A(n11475), .B(n11473), .Z(n11474) );
  XNOR U14512 ( .A(n11476), .B(n11477), .Z(n11464) );
  NAND U14513 ( .A(n11478), .B(n11479), .Z(n11477) );
  XOR U14514 ( .A(n11480), .B(n11456), .Z(n11479) );
  XOR U14515 ( .A(n11470), .B(n11471), .Z(n11456) );
  XOR U14516 ( .A(n11481), .B(n11482), .Z(n11471) );
  ANDN U14517 ( .B(n11483), .A(n11484), .Z(n11481) );
  XOR U14518 ( .A(n11482), .B(n11485), .Z(n11483) );
  XOR U14519 ( .A(n11486), .B(n11487), .Z(n11470) );
  XOR U14520 ( .A(n11488), .B(n11489), .Z(n11487) );
  ANDN U14521 ( .B(n11490), .A(n11491), .Z(n11488) );
  XOR U14522 ( .A(n11492), .B(n11489), .Z(n11490) );
  IV U14523 ( .A(n11468), .Z(n11486) );
  XOR U14524 ( .A(n11493), .B(n11494), .Z(n11468) );
  ANDN U14525 ( .B(n11495), .A(n11496), .Z(n11493) );
  XOR U14526 ( .A(n11494), .B(n11497), .Z(n11495) );
  IV U14527 ( .A(n11476), .Z(n11480) );
  XOR U14528 ( .A(n11476), .B(n11458), .Z(n11478) );
  XOR U14529 ( .A(n11498), .B(n11499), .Z(n11458) );
  AND U14530 ( .A(n26), .B(n11500), .Z(n11498) );
  XOR U14531 ( .A(n11501), .B(n11499), .Z(n11500) );
  NANDN U14532 ( .A(n11460), .B(n11462), .Z(n11476) );
  XOR U14533 ( .A(n11502), .B(n11503), .Z(n11462) );
  AND U14534 ( .A(n26), .B(n11504), .Z(n11502) );
  XOR U14535 ( .A(n11503), .B(n11505), .Z(n11504) );
  XOR U14536 ( .A(n11506), .B(n11507), .Z(n26) );
  AND U14537 ( .A(n11508), .B(n11509), .Z(n11506) );
  XNOR U14538 ( .A(n11507), .B(n11473), .Z(n11509) );
  XNOR U14539 ( .A(n11510), .B(n11511), .Z(n11473) );
  ANDN U14540 ( .B(n11512), .A(n11513), .Z(n11510) );
  XOR U14541 ( .A(n11511), .B(n11514), .Z(n11512) );
  XOR U14542 ( .A(n11507), .B(n11475), .Z(n11508) );
  XOR U14543 ( .A(n11515), .B(n11516), .Z(n11475) );
  AND U14544 ( .A(n30), .B(n11517), .Z(n11515) );
  XOR U14545 ( .A(n11518), .B(n11516), .Z(n11517) );
  XNOR U14546 ( .A(n11519), .B(n11520), .Z(n11507) );
  NAND U14547 ( .A(n11521), .B(n11522), .Z(n11520) );
  XOR U14548 ( .A(n11523), .B(n11499), .Z(n11522) );
  XOR U14549 ( .A(n11513), .B(n11514), .Z(n11499) );
  XOR U14550 ( .A(n11524), .B(n11525), .Z(n11514) );
  ANDN U14551 ( .B(n11526), .A(n11527), .Z(n11524) );
  XOR U14552 ( .A(n11525), .B(n11528), .Z(n11526) );
  XOR U14553 ( .A(n11529), .B(n11530), .Z(n11513) );
  XOR U14554 ( .A(n11531), .B(n11532), .Z(n11530) );
  ANDN U14555 ( .B(n11533), .A(n11534), .Z(n11531) );
  XOR U14556 ( .A(n11535), .B(n11532), .Z(n11533) );
  IV U14557 ( .A(n11511), .Z(n11529) );
  XOR U14558 ( .A(n11536), .B(n11537), .Z(n11511) );
  ANDN U14559 ( .B(n11538), .A(n11539), .Z(n11536) );
  XOR U14560 ( .A(n11537), .B(n11540), .Z(n11538) );
  IV U14561 ( .A(n11519), .Z(n11523) );
  XOR U14562 ( .A(n11519), .B(n11501), .Z(n11521) );
  XOR U14563 ( .A(n11541), .B(n11542), .Z(n11501) );
  AND U14564 ( .A(n30), .B(n11543), .Z(n11541) );
  XOR U14565 ( .A(n11544), .B(n11542), .Z(n11543) );
  NANDN U14566 ( .A(n11503), .B(n11505), .Z(n11519) );
  XOR U14567 ( .A(n11545), .B(n11546), .Z(n11505) );
  AND U14568 ( .A(n30), .B(n11547), .Z(n11545) );
  XOR U14569 ( .A(n11546), .B(n11548), .Z(n11547) );
  XOR U14570 ( .A(n11549), .B(n11550), .Z(n30) );
  AND U14571 ( .A(n11551), .B(n11552), .Z(n11549) );
  XNOR U14572 ( .A(n11550), .B(n11516), .Z(n11552) );
  XNOR U14573 ( .A(n11553), .B(n11554), .Z(n11516) );
  ANDN U14574 ( .B(n11555), .A(n11556), .Z(n11553) );
  XOR U14575 ( .A(n11554), .B(n11557), .Z(n11555) );
  XOR U14576 ( .A(n11550), .B(n11518), .Z(n11551) );
  XOR U14577 ( .A(n11558), .B(n11559), .Z(n11518) );
  AND U14578 ( .A(n34), .B(n11560), .Z(n11558) );
  XOR U14579 ( .A(n11561), .B(n11559), .Z(n11560) );
  XNOR U14580 ( .A(n11562), .B(n11563), .Z(n11550) );
  NAND U14581 ( .A(n11564), .B(n11565), .Z(n11563) );
  XOR U14582 ( .A(n11566), .B(n11542), .Z(n11565) );
  XOR U14583 ( .A(n11556), .B(n11557), .Z(n11542) );
  XOR U14584 ( .A(n11567), .B(n11568), .Z(n11557) );
  ANDN U14585 ( .B(n11569), .A(n11570), .Z(n11567) );
  XOR U14586 ( .A(n11568), .B(n11571), .Z(n11569) );
  XOR U14587 ( .A(n11572), .B(n11573), .Z(n11556) );
  XOR U14588 ( .A(n11574), .B(n11575), .Z(n11573) );
  ANDN U14589 ( .B(n11576), .A(n11577), .Z(n11574) );
  XOR U14590 ( .A(n11578), .B(n11575), .Z(n11576) );
  IV U14591 ( .A(n11554), .Z(n11572) );
  XOR U14592 ( .A(n11579), .B(n11580), .Z(n11554) );
  ANDN U14593 ( .B(n11581), .A(n11582), .Z(n11579) );
  XOR U14594 ( .A(n11580), .B(n11583), .Z(n11581) );
  IV U14595 ( .A(n11562), .Z(n11566) );
  XOR U14596 ( .A(n11562), .B(n11544), .Z(n11564) );
  XOR U14597 ( .A(n11584), .B(n11585), .Z(n11544) );
  AND U14598 ( .A(n34), .B(n11586), .Z(n11584) );
  XOR U14599 ( .A(n11587), .B(n11585), .Z(n11586) );
  NANDN U14600 ( .A(n11546), .B(n11548), .Z(n11562) );
  XOR U14601 ( .A(n11588), .B(n11589), .Z(n11548) );
  AND U14602 ( .A(n34), .B(n11590), .Z(n11588) );
  XOR U14603 ( .A(n11589), .B(n11591), .Z(n11590) );
  XOR U14604 ( .A(n11592), .B(n11593), .Z(n34) );
  AND U14605 ( .A(n11594), .B(n11595), .Z(n11592) );
  XNOR U14606 ( .A(n11593), .B(n11559), .Z(n11595) );
  XNOR U14607 ( .A(n11596), .B(n11597), .Z(n11559) );
  ANDN U14608 ( .B(n11598), .A(n11599), .Z(n11596) );
  XOR U14609 ( .A(n11597), .B(n11600), .Z(n11598) );
  XOR U14610 ( .A(n11593), .B(n11561), .Z(n11594) );
  XOR U14611 ( .A(n11601), .B(n11602), .Z(n11561) );
  AND U14612 ( .A(n38), .B(n11603), .Z(n11601) );
  XOR U14613 ( .A(n11604), .B(n11602), .Z(n11603) );
  XNOR U14614 ( .A(n11605), .B(n11606), .Z(n11593) );
  NAND U14615 ( .A(n11607), .B(n11608), .Z(n11606) );
  XOR U14616 ( .A(n11609), .B(n11585), .Z(n11608) );
  XOR U14617 ( .A(n11599), .B(n11600), .Z(n11585) );
  XOR U14618 ( .A(n11610), .B(n11611), .Z(n11600) );
  ANDN U14619 ( .B(n11612), .A(n11613), .Z(n11610) );
  XOR U14620 ( .A(n11611), .B(n11614), .Z(n11612) );
  XOR U14621 ( .A(n11615), .B(n11616), .Z(n11599) );
  XOR U14622 ( .A(n11617), .B(n11618), .Z(n11616) );
  ANDN U14623 ( .B(n11619), .A(n11620), .Z(n11617) );
  XOR U14624 ( .A(n11621), .B(n11618), .Z(n11619) );
  IV U14625 ( .A(n11597), .Z(n11615) );
  XOR U14626 ( .A(n11622), .B(n11623), .Z(n11597) );
  ANDN U14627 ( .B(n11624), .A(n11625), .Z(n11622) );
  XOR U14628 ( .A(n11623), .B(n11626), .Z(n11624) );
  IV U14629 ( .A(n11605), .Z(n11609) );
  XOR U14630 ( .A(n11605), .B(n11587), .Z(n11607) );
  XOR U14631 ( .A(n11627), .B(n11628), .Z(n11587) );
  AND U14632 ( .A(n38), .B(n11629), .Z(n11627) );
  XOR U14633 ( .A(n11630), .B(n11628), .Z(n11629) );
  NANDN U14634 ( .A(n11589), .B(n11591), .Z(n11605) );
  XOR U14635 ( .A(n11631), .B(n11632), .Z(n11591) );
  AND U14636 ( .A(n38), .B(n11633), .Z(n11631) );
  XOR U14637 ( .A(n11632), .B(n11634), .Z(n11633) );
  XOR U14638 ( .A(n11635), .B(n11636), .Z(n38) );
  AND U14639 ( .A(n11637), .B(n11638), .Z(n11635) );
  XNOR U14640 ( .A(n11636), .B(n11602), .Z(n11638) );
  XNOR U14641 ( .A(n11639), .B(n11640), .Z(n11602) );
  ANDN U14642 ( .B(n11641), .A(n11642), .Z(n11639) );
  XOR U14643 ( .A(n11640), .B(n11643), .Z(n11641) );
  XOR U14644 ( .A(n11636), .B(n11604), .Z(n11637) );
  XOR U14645 ( .A(n11644), .B(n11645), .Z(n11604) );
  AND U14646 ( .A(n42), .B(n11646), .Z(n11644) );
  XOR U14647 ( .A(n11647), .B(n11645), .Z(n11646) );
  XNOR U14648 ( .A(n11648), .B(n11649), .Z(n11636) );
  NAND U14649 ( .A(n11650), .B(n11651), .Z(n11649) );
  XOR U14650 ( .A(n11652), .B(n11628), .Z(n11651) );
  XOR U14651 ( .A(n11642), .B(n11643), .Z(n11628) );
  XOR U14652 ( .A(n11653), .B(n11654), .Z(n11643) );
  ANDN U14653 ( .B(n11655), .A(n11656), .Z(n11653) );
  XOR U14654 ( .A(n11654), .B(n11657), .Z(n11655) );
  XOR U14655 ( .A(n11658), .B(n11659), .Z(n11642) );
  XOR U14656 ( .A(n11660), .B(n11661), .Z(n11659) );
  ANDN U14657 ( .B(n11662), .A(n11663), .Z(n11660) );
  XOR U14658 ( .A(n11664), .B(n11661), .Z(n11662) );
  IV U14659 ( .A(n11640), .Z(n11658) );
  XOR U14660 ( .A(n11665), .B(n11666), .Z(n11640) );
  ANDN U14661 ( .B(n11667), .A(n11668), .Z(n11665) );
  XOR U14662 ( .A(n11666), .B(n11669), .Z(n11667) );
  IV U14663 ( .A(n11648), .Z(n11652) );
  XOR U14664 ( .A(n11648), .B(n11630), .Z(n11650) );
  XOR U14665 ( .A(n11670), .B(n11671), .Z(n11630) );
  AND U14666 ( .A(n42), .B(n11672), .Z(n11670) );
  XOR U14667 ( .A(n11673), .B(n11671), .Z(n11672) );
  NANDN U14668 ( .A(n11632), .B(n11634), .Z(n11648) );
  XOR U14669 ( .A(n11674), .B(n11675), .Z(n11634) );
  AND U14670 ( .A(n42), .B(n11676), .Z(n11674) );
  XOR U14671 ( .A(n11675), .B(n11677), .Z(n11676) );
  XOR U14672 ( .A(n11678), .B(n11679), .Z(n42) );
  AND U14673 ( .A(n11680), .B(n11681), .Z(n11678) );
  XNOR U14674 ( .A(n11679), .B(n11645), .Z(n11681) );
  XNOR U14675 ( .A(n11682), .B(n11683), .Z(n11645) );
  ANDN U14676 ( .B(n11684), .A(n11685), .Z(n11682) );
  XOR U14677 ( .A(n11683), .B(n11686), .Z(n11684) );
  XOR U14678 ( .A(n11679), .B(n11647), .Z(n11680) );
  XOR U14679 ( .A(n11687), .B(n11688), .Z(n11647) );
  AND U14680 ( .A(n46), .B(n11689), .Z(n11687) );
  XOR U14681 ( .A(n11690), .B(n11688), .Z(n11689) );
  XNOR U14682 ( .A(n11691), .B(n11692), .Z(n11679) );
  NAND U14683 ( .A(n11693), .B(n11694), .Z(n11692) );
  XOR U14684 ( .A(n11695), .B(n11671), .Z(n11694) );
  XOR U14685 ( .A(n11685), .B(n11686), .Z(n11671) );
  XOR U14686 ( .A(n11696), .B(n11697), .Z(n11686) );
  ANDN U14687 ( .B(n11698), .A(n11699), .Z(n11696) );
  XOR U14688 ( .A(n11697), .B(n11700), .Z(n11698) );
  XOR U14689 ( .A(n11701), .B(n11702), .Z(n11685) );
  XOR U14690 ( .A(n11703), .B(n11704), .Z(n11702) );
  ANDN U14691 ( .B(n11705), .A(n11706), .Z(n11703) );
  XOR U14692 ( .A(n11707), .B(n11704), .Z(n11705) );
  IV U14693 ( .A(n11683), .Z(n11701) );
  XOR U14694 ( .A(n11708), .B(n11709), .Z(n11683) );
  ANDN U14695 ( .B(n11710), .A(n11711), .Z(n11708) );
  XOR U14696 ( .A(n11709), .B(n11712), .Z(n11710) );
  IV U14697 ( .A(n11691), .Z(n11695) );
  XOR U14698 ( .A(n11691), .B(n11673), .Z(n11693) );
  XOR U14699 ( .A(n11713), .B(n11714), .Z(n11673) );
  AND U14700 ( .A(n46), .B(n11715), .Z(n11713) );
  XOR U14701 ( .A(n11716), .B(n11714), .Z(n11715) );
  NANDN U14702 ( .A(n11675), .B(n11677), .Z(n11691) );
  XOR U14703 ( .A(n11717), .B(n11718), .Z(n11677) );
  AND U14704 ( .A(n46), .B(n11719), .Z(n11717) );
  XOR U14705 ( .A(n11718), .B(n11720), .Z(n11719) );
  XOR U14706 ( .A(n11721), .B(n11722), .Z(n46) );
  AND U14707 ( .A(n11723), .B(n11724), .Z(n11721) );
  XNOR U14708 ( .A(n11722), .B(n11688), .Z(n11724) );
  XNOR U14709 ( .A(n11725), .B(n11726), .Z(n11688) );
  ANDN U14710 ( .B(n11727), .A(n11728), .Z(n11725) );
  XOR U14711 ( .A(n11726), .B(n11729), .Z(n11727) );
  XOR U14712 ( .A(n11722), .B(n11690), .Z(n11723) );
  XOR U14713 ( .A(n11730), .B(n11731), .Z(n11690) );
  AND U14714 ( .A(n50), .B(n11732), .Z(n11730) );
  XOR U14715 ( .A(n11733), .B(n11731), .Z(n11732) );
  XNOR U14716 ( .A(n11734), .B(n11735), .Z(n11722) );
  NAND U14717 ( .A(n11736), .B(n11737), .Z(n11735) );
  XOR U14718 ( .A(n11738), .B(n11714), .Z(n11737) );
  XOR U14719 ( .A(n11728), .B(n11729), .Z(n11714) );
  XOR U14720 ( .A(n11739), .B(n11740), .Z(n11729) );
  ANDN U14721 ( .B(n11741), .A(n11742), .Z(n11739) );
  XOR U14722 ( .A(n11740), .B(n11743), .Z(n11741) );
  XOR U14723 ( .A(n11744), .B(n11745), .Z(n11728) );
  XOR U14724 ( .A(n11746), .B(n11747), .Z(n11745) );
  ANDN U14725 ( .B(n11748), .A(n11749), .Z(n11746) );
  XOR U14726 ( .A(n11750), .B(n11747), .Z(n11748) );
  IV U14727 ( .A(n11726), .Z(n11744) );
  XOR U14728 ( .A(n11751), .B(n11752), .Z(n11726) );
  ANDN U14729 ( .B(n11753), .A(n11754), .Z(n11751) );
  XOR U14730 ( .A(n11752), .B(n11755), .Z(n11753) );
  IV U14731 ( .A(n11734), .Z(n11738) );
  XOR U14732 ( .A(n11734), .B(n11716), .Z(n11736) );
  XOR U14733 ( .A(n11756), .B(n11757), .Z(n11716) );
  AND U14734 ( .A(n50), .B(n11758), .Z(n11756) );
  XOR U14735 ( .A(n11759), .B(n11757), .Z(n11758) );
  NANDN U14736 ( .A(n11718), .B(n11720), .Z(n11734) );
  XOR U14737 ( .A(n11760), .B(n11761), .Z(n11720) );
  AND U14738 ( .A(n50), .B(n11762), .Z(n11760) );
  XOR U14739 ( .A(n11761), .B(n11763), .Z(n11762) );
  XOR U14740 ( .A(n11764), .B(n11765), .Z(n50) );
  AND U14741 ( .A(n11766), .B(n11767), .Z(n11764) );
  XNOR U14742 ( .A(n11765), .B(n11731), .Z(n11767) );
  XNOR U14743 ( .A(n11768), .B(n11769), .Z(n11731) );
  ANDN U14744 ( .B(n11770), .A(n11771), .Z(n11768) );
  XOR U14745 ( .A(n11769), .B(n11772), .Z(n11770) );
  XOR U14746 ( .A(n11765), .B(n11733), .Z(n11766) );
  XOR U14747 ( .A(n11773), .B(n11774), .Z(n11733) );
  AND U14748 ( .A(n54), .B(n11775), .Z(n11773) );
  XOR U14749 ( .A(n11776), .B(n11774), .Z(n11775) );
  XNOR U14750 ( .A(n11777), .B(n11778), .Z(n11765) );
  NAND U14751 ( .A(n11779), .B(n11780), .Z(n11778) );
  XOR U14752 ( .A(n11781), .B(n11757), .Z(n11780) );
  XOR U14753 ( .A(n11771), .B(n11772), .Z(n11757) );
  XOR U14754 ( .A(n11782), .B(n11783), .Z(n11772) );
  ANDN U14755 ( .B(n11784), .A(n11785), .Z(n11782) );
  XOR U14756 ( .A(n11783), .B(n11786), .Z(n11784) );
  XOR U14757 ( .A(n11787), .B(n11788), .Z(n11771) );
  XOR U14758 ( .A(n11789), .B(n11790), .Z(n11788) );
  ANDN U14759 ( .B(n11791), .A(n11792), .Z(n11789) );
  XOR U14760 ( .A(n11793), .B(n11790), .Z(n11791) );
  IV U14761 ( .A(n11769), .Z(n11787) );
  XOR U14762 ( .A(n11794), .B(n11795), .Z(n11769) );
  ANDN U14763 ( .B(n11796), .A(n11797), .Z(n11794) );
  XOR U14764 ( .A(n11795), .B(n11798), .Z(n11796) );
  IV U14765 ( .A(n11777), .Z(n11781) );
  XOR U14766 ( .A(n11777), .B(n11759), .Z(n11779) );
  XOR U14767 ( .A(n11799), .B(n11800), .Z(n11759) );
  AND U14768 ( .A(n54), .B(n11801), .Z(n11799) );
  XOR U14769 ( .A(n11802), .B(n11800), .Z(n11801) );
  NANDN U14770 ( .A(n11761), .B(n11763), .Z(n11777) );
  XOR U14771 ( .A(n11803), .B(n11804), .Z(n11763) );
  AND U14772 ( .A(n54), .B(n11805), .Z(n11803) );
  XOR U14773 ( .A(n11804), .B(n11806), .Z(n11805) );
  XOR U14774 ( .A(n11807), .B(n11808), .Z(n54) );
  AND U14775 ( .A(n11809), .B(n11810), .Z(n11807) );
  XNOR U14776 ( .A(n11808), .B(n11774), .Z(n11810) );
  XNOR U14777 ( .A(n11811), .B(n11812), .Z(n11774) );
  ANDN U14778 ( .B(n11813), .A(n11814), .Z(n11811) );
  XOR U14779 ( .A(n11812), .B(n11815), .Z(n11813) );
  XOR U14780 ( .A(n11808), .B(n11776), .Z(n11809) );
  XOR U14781 ( .A(n11816), .B(n11817), .Z(n11776) );
  AND U14782 ( .A(n58), .B(n11818), .Z(n11816) );
  XOR U14783 ( .A(n11819), .B(n11817), .Z(n11818) );
  XNOR U14784 ( .A(n11820), .B(n11821), .Z(n11808) );
  NAND U14785 ( .A(n11822), .B(n11823), .Z(n11821) );
  XOR U14786 ( .A(n11824), .B(n11800), .Z(n11823) );
  XOR U14787 ( .A(n11814), .B(n11815), .Z(n11800) );
  XOR U14788 ( .A(n11825), .B(n11826), .Z(n11815) );
  ANDN U14789 ( .B(n11827), .A(n11828), .Z(n11825) );
  XOR U14790 ( .A(n11826), .B(n11829), .Z(n11827) );
  XOR U14791 ( .A(n11830), .B(n11831), .Z(n11814) );
  XOR U14792 ( .A(n11832), .B(n11833), .Z(n11831) );
  ANDN U14793 ( .B(n11834), .A(n11835), .Z(n11832) );
  XOR U14794 ( .A(n11836), .B(n11833), .Z(n11834) );
  IV U14795 ( .A(n11812), .Z(n11830) );
  XOR U14796 ( .A(n11837), .B(n11838), .Z(n11812) );
  ANDN U14797 ( .B(n11839), .A(n11840), .Z(n11837) );
  XOR U14798 ( .A(n11838), .B(n11841), .Z(n11839) );
  IV U14799 ( .A(n11820), .Z(n11824) );
  XOR U14800 ( .A(n11820), .B(n11802), .Z(n11822) );
  XOR U14801 ( .A(n11842), .B(n11843), .Z(n11802) );
  AND U14802 ( .A(n58), .B(n11844), .Z(n11842) );
  XOR U14803 ( .A(n11845), .B(n11843), .Z(n11844) );
  NANDN U14804 ( .A(n11804), .B(n11806), .Z(n11820) );
  XOR U14805 ( .A(n11846), .B(n11847), .Z(n11806) );
  AND U14806 ( .A(n58), .B(n11848), .Z(n11846) );
  XOR U14807 ( .A(n11847), .B(n11849), .Z(n11848) );
  XOR U14808 ( .A(n11850), .B(n11851), .Z(n58) );
  AND U14809 ( .A(n11852), .B(n11853), .Z(n11850) );
  XNOR U14810 ( .A(n11851), .B(n11817), .Z(n11853) );
  XNOR U14811 ( .A(n11854), .B(n11855), .Z(n11817) );
  ANDN U14812 ( .B(n11856), .A(n11857), .Z(n11854) );
  XOR U14813 ( .A(n11855), .B(n11858), .Z(n11856) );
  XOR U14814 ( .A(n11851), .B(n11819), .Z(n11852) );
  XOR U14815 ( .A(n11859), .B(n11860), .Z(n11819) );
  AND U14816 ( .A(n62), .B(n11861), .Z(n11859) );
  XOR U14817 ( .A(n11862), .B(n11860), .Z(n11861) );
  XNOR U14818 ( .A(n11863), .B(n11864), .Z(n11851) );
  NAND U14819 ( .A(n11865), .B(n11866), .Z(n11864) );
  XOR U14820 ( .A(n11867), .B(n11843), .Z(n11866) );
  XOR U14821 ( .A(n11857), .B(n11858), .Z(n11843) );
  XOR U14822 ( .A(n11868), .B(n11869), .Z(n11858) );
  ANDN U14823 ( .B(n11870), .A(n11871), .Z(n11868) );
  XOR U14824 ( .A(n11869), .B(n11872), .Z(n11870) );
  XOR U14825 ( .A(n11873), .B(n11874), .Z(n11857) );
  XOR U14826 ( .A(n11875), .B(n11876), .Z(n11874) );
  ANDN U14827 ( .B(n11877), .A(n11878), .Z(n11875) );
  XOR U14828 ( .A(n11879), .B(n11876), .Z(n11877) );
  IV U14829 ( .A(n11855), .Z(n11873) );
  XOR U14830 ( .A(n11880), .B(n11881), .Z(n11855) );
  ANDN U14831 ( .B(n11882), .A(n11883), .Z(n11880) );
  XOR U14832 ( .A(n11881), .B(n11884), .Z(n11882) );
  IV U14833 ( .A(n11863), .Z(n11867) );
  XOR U14834 ( .A(n11863), .B(n11845), .Z(n11865) );
  XOR U14835 ( .A(n11885), .B(n11886), .Z(n11845) );
  AND U14836 ( .A(n62), .B(n11887), .Z(n11885) );
  XOR U14837 ( .A(n11888), .B(n11886), .Z(n11887) );
  NANDN U14838 ( .A(n11847), .B(n11849), .Z(n11863) );
  XOR U14839 ( .A(n11889), .B(n11890), .Z(n11849) );
  AND U14840 ( .A(n62), .B(n11891), .Z(n11889) );
  XOR U14841 ( .A(n11890), .B(n11892), .Z(n11891) );
  XOR U14842 ( .A(n11893), .B(n11894), .Z(n62) );
  AND U14843 ( .A(n11895), .B(n11896), .Z(n11893) );
  XNOR U14844 ( .A(n11894), .B(n11860), .Z(n11896) );
  XNOR U14845 ( .A(n11897), .B(n11898), .Z(n11860) );
  ANDN U14846 ( .B(n11899), .A(n11900), .Z(n11897) );
  XOR U14847 ( .A(n11898), .B(n11901), .Z(n11899) );
  XOR U14848 ( .A(n11894), .B(n11862), .Z(n11895) );
  XOR U14849 ( .A(n11902), .B(n11903), .Z(n11862) );
  AND U14850 ( .A(n66), .B(n11904), .Z(n11902) );
  XOR U14851 ( .A(n11905), .B(n11903), .Z(n11904) );
  XNOR U14852 ( .A(n11906), .B(n11907), .Z(n11894) );
  NAND U14853 ( .A(n11908), .B(n11909), .Z(n11907) );
  XOR U14854 ( .A(n11910), .B(n11886), .Z(n11909) );
  XOR U14855 ( .A(n11900), .B(n11901), .Z(n11886) );
  XOR U14856 ( .A(n11911), .B(n11912), .Z(n11901) );
  ANDN U14857 ( .B(n11913), .A(n11914), .Z(n11911) );
  XOR U14858 ( .A(n11912), .B(n11915), .Z(n11913) );
  XOR U14859 ( .A(n11916), .B(n11917), .Z(n11900) );
  XOR U14860 ( .A(n11918), .B(n11919), .Z(n11917) );
  ANDN U14861 ( .B(n11920), .A(n11921), .Z(n11918) );
  XOR U14862 ( .A(n11922), .B(n11919), .Z(n11920) );
  IV U14863 ( .A(n11898), .Z(n11916) );
  XOR U14864 ( .A(n11923), .B(n11924), .Z(n11898) );
  ANDN U14865 ( .B(n11925), .A(n11926), .Z(n11923) );
  XOR U14866 ( .A(n11924), .B(n11927), .Z(n11925) );
  IV U14867 ( .A(n11906), .Z(n11910) );
  XOR U14868 ( .A(n11906), .B(n11888), .Z(n11908) );
  XOR U14869 ( .A(n11928), .B(n11929), .Z(n11888) );
  AND U14870 ( .A(n66), .B(n11930), .Z(n11928) );
  XOR U14871 ( .A(n11931), .B(n11929), .Z(n11930) );
  NANDN U14872 ( .A(n11890), .B(n11892), .Z(n11906) );
  XOR U14873 ( .A(n11932), .B(n11933), .Z(n11892) );
  AND U14874 ( .A(n66), .B(n11934), .Z(n11932) );
  XOR U14875 ( .A(n11933), .B(n11935), .Z(n11934) );
  XOR U14876 ( .A(n11936), .B(n11937), .Z(n66) );
  AND U14877 ( .A(n11938), .B(n11939), .Z(n11936) );
  XNOR U14878 ( .A(n11937), .B(n11903), .Z(n11939) );
  XNOR U14879 ( .A(n11940), .B(n11941), .Z(n11903) );
  ANDN U14880 ( .B(n11942), .A(n11943), .Z(n11940) );
  XOR U14881 ( .A(n11941), .B(n11944), .Z(n11942) );
  XOR U14882 ( .A(n11937), .B(n11905), .Z(n11938) );
  XOR U14883 ( .A(n11945), .B(n11946), .Z(n11905) );
  AND U14884 ( .A(n70), .B(n11947), .Z(n11945) );
  XOR U14885 ( .A(n11948), .B(n11946), .Z(n11947) );
  XNOR U14886 ( .A(n11949), .B(n11950), .Z(n11937) );
  NAND U14887 ( .A(n11951), .B(n11952), .Z(n11950) );
  XOR U14888 ( .A(n11953), .B(n11929), .Z(n11952) );
  XOR U14889 ( .A(n11943), .B(n11944), .Z(n11929) );
  XOR U14890 ( .A(n11954), .B(n11955), .Z(n11944) );
  ANDN U14891 ( .B(n11956), .A(n11957), .Z(n11954) );
  XOR U14892 ( .A(n11955), .B(n11958), .Z(n11956) );
  XOR U14893 ( .A(n11959), .B(n11960), .Z(n11943) );
  XOR U14894 ( .A(n11961), .B(n11962), .Z(n11960) );
  ANDN U14895 ( .B(n11963), .A(n11964), .Z(n11961) );
  XOR U14896 ( .A(n11965), .B(n11962), .Z(n11963) );
  IV U14897 ( .A(n11941), .Z(n11959) );
  XOR U14898 ( .A(n11966), .B(n11967), .Z(n11941) );
  ANDN U14899 ( .B(n11968), .A(n11969), .Z(n11966) );
  XOR U14900 ( .A(n11967), .B(n11970), .Z(n11968) );
  IV U14901 ( .A(n11949), .Z(n11953) );
  XOR U14902 ( .A(n11949), .B(n11931), .Z(n11951) );
  XOR U14903 ( .A(n11971), .B(n11972), .Z(n11931) );
  AND U14904 ( .A(n70), .B(n11973), .Z(n11971) );
  XOR U14905 ( .A(n11974), .B(n11972), .Z(n11973) );
  NANDN U14906 ( .A(n11933), .B(n11935), .Z(n11949) );
  XOR U14907 ( .A(n11975), .B(n11976), .Z(n11935) );
  AND U14908 ( .A(n70), .B(n11977), .Z(n11975) );
  XOR U14909 ( .A(n11976), .B(n11978), .Z(n11977) );
  XOR U14910 ( .A(n11979), .B(n11980), .Z(n70) );
  AND U14911 ( .A(n11981), .B(n11982), .Z(n11979) );
  XNOR U14912 ( .A(n11980), .B(n11946), .Z(n11982) );
  XNOR U14913 ( .A(n11983), .B(n11984), .Z(n11946) );
  ANDN U14914 ( .B(n11985), .A(n11986), .Z(n11983) );
  XOR U14915 ( .A(n11984), .B(n11987), .Z(n11985) );
  XOR U14916 ( .A(n11980), .B(n11948), .Z(n11981) );
  XOR U14917 ( .A(n11988), .B(n11989), .Z(n11948) );
  AND U14918 ( .A(n74), .B(n11990), .Z(n11988) );
  XOR U14919 ( .A(n11991), .B(n11989), .Z(n11990) );
  XNOR U14920 ( .A(n11992), .B(n11993), .Z(n11980) );
  NAND U14921 ( .A(n11994), .B(n11995), .Z(n11993) );
  XOR U14922 ( .A(n11996), .B(n11972), .Z(n11995) );
  XOR U14923 ( .A(n11986), .B(n11987), .Z(n11972) );
  XOR U14924 ( .A(n11997), .B(n11998), .Z(n11987) );
  ANDN U14925 ( .B(n11999), .A(n12000), .Z(n11997) );
  XOR U14926 ( .A(n11998), .B(n12001), .Z(n11999) );
  XOR U14927 ( .A(n12002), .B(n12003), .Z(n11986) );
  XOR U14928 ( .A(n12004), .B(n12005), .Z(n12003) );
  ANDN U14929 ( .B(n12006), .A(n12007), .Z(n12004) );
  XOR U14930 ( .A(n12008), .B(n12005), .Z(n12006) );
  IV U14931 ( .A(n11984), .Z(n12002) );
  XOR U14932 ( .A(n12009), .B(n12010), .Z(n11984) );
  ANDN U14933 ( .B(n12011), .A(n12012), .Z(n12009) );
  XOR U14934 ( .A(n12010), .B(n12013), .Z(n12011) );
  IV U14935 ( .A(n11992), .Z(n11996) );
  XOR U14936 ( .A(n11992), .B(n11974), .Z(n11994) );
  XOR U14937 ( .A(n12014), .B(n12015), .Z(n11974) );
  AND U14938 ( .A(n74), .B(n12016), .Z(n12014) );
  XOR U14939 ( .A(n12017), .B(n12015), .Z(n12016) );
  NANDN U14940 ( .A(n11976), .B(n11978), .Z(n11992) );
  XOR U14941 ( .A(n12018), .B(n12019), .Z(n11978) );
  AND U14942 ( .A(n74), .B(n12020), .Z(n12018) );
  XOR U14943 ( .A(n12019), .B(n12021), .Z(n12020) );
  XOR U14944 ( .A(n12022), .B(n12023), .Z(n74) );
  AND U14945 ( .A(n12024), .B(n12025), .Z(n12022) );
  XNOR U14946 ( .A(n12023), .B(n11989), .Z(n12025) );
  XNOR U14947 ( .A(n12026), .B(n12027), .Z(n11989) );
  ANDN U14948 ( .B(n12028), .A(n12029), .Z(n12026) );
  XOR U14949 ( .A(n12027), .B(n12030), .Z(n12028) );
  XOR U14950 ( .A(n12023), .B(n11991), .Z(n12024) );
  XOR U14951 ( .A(n12031), .B(n12032), .Z(n11991) );
  AND U14952 ( .A(n78), .B(n12033), .Z(n12031) );
  XOR U14953 ( .A(n12034), .B(n12032), .Z(n12033) );
  XNOR U14954 ( .A(n12035), .B(n12036), .Z(n12023) );
  NAND U14955 ( .A(n12037), .B(n12038), .Z(n12036) );
  XOR U14956 ( .A(n12039), .B(n12015), .Z(n12038) );
  XOR U14957 ( .A(n12029), .B(n12030), .Z(n12015) );
  XOR U14958 ( .A(n12040), .B(n12041), .Z(n12030) );
  ANDN U14959 ( .B(n12042), .A(n12043), .Z(n12040) );
  XOR U14960 ( .A(n12041), .B(n12044), .Z(n12042) );
  XOR U14961 ( .A(n12045), .B(n12046), .Z(n12029) );
  XOR U14962 ( .A(n12047), .B(n12048), .Z(n12046) );
  ANDN U14963 ( .B(n12049), .A(n12050), .Z(n12047) );
  XOR U14964 ( .A(n12051), .B(n12048), .Z(n12049) );
  IV U14965 ( .A(n12027), .Z(n12045) );
  XOR U14966 ( .A(n12052), .B(n12053), .Z(n12027) );
  ANDN U14967 ( .B(n12054), .A(n12055), .Z(n12052) );
  XOR U14968 ( .A(n12053), .B(n12056), .Z(n12054) );
  IV U14969 ( .A(n12035), .Z(n12039) );
  XOR U14970 ( .A(n12035), .B(n12017), .Z(n12037) );
  XOR U14971 ( .A(n12057), .B(n12058), .Z(n12017) );
  AND U14972 ( .A(n78), .B(n12059), .Z(n12057) );
  XOR U14973 ( .A(n12060), .B(n12058), .Z(n12059) );
  NANDN U14974 ( .A(n12019), .B(n12021), .Z(n12035) );
  XOR U14975 ( .A(n12061), .B(n12062), .Z(n12021) );
  AND U14976 ( .A(n78), .B(n12063), .Z(n12061) );
  XOR U14977 ( .A(n12062), .B(n12064), .Z(n12063) );
  XOR U14978 ( .A(n12065), .B(n12066), .Z(n78) );
  AND U14979 ( .A(n12067), .B(n12068), .Z(n12065) );
  XNOR U14980 ( .A(n12066), .B(n12032), .Z(n12068) );
  XNOR U14981 ( .A(n12069), .B(n12070), .Z(n12032) );
  ANDN U14982 ( .B(n12071), .A(n12072), .Z(n12069) );
  XOR U14983 ( .A(n12070), .B(n12073), .Z(n12071) );
  XOR U14984 ( .A(n12066), .B(n12034), .Z(n12067) );
  XOR U14985 ( .A(n12074), .B(n12075), .Z(n12034) );
  AND U14986 ( .A(n82), .B(n12076), .Z(n12074) );
  XOR U14987 ( .A(n12077), .B(n12075), .Z(n12076) );
  XNOR U14988 ( .A(n12078), .B(n12079), .Z(n12066) );
  NAND U14989 ( .A(n12080), .B(n12081), .Z(n12079) );
  XOR U14990 ( .A(n12082), .B(n12058), .Z(n12081) );
  XOR U14991 ( .A(n12072), .B(n12073), .Z(n12058) );
  XOR U14992 ( .A(n12083), .B(n12084), .Z(n12073) );
  ANDN U14993 ( .B(n12085), .A(n12086), .Z(n12083) );
  XOR U14994 ( .A(n12084), .B(n12087), .Z(n12085) );
  XOR U14995 ( .A(n12088), .B(n12089), .Z(n12072) );
  XOR U14996 ( .A(n12090), .B(n12091), .Z(n12089) );
  ANDN U14997 ( .B(n12092), .A(n12093), .Z(n12090) );
  XOR U14998 ( .A(n12094), .B(n12091), .Z(n12092) );
  IV U14999 ( .A(n12070), .Z(n12088) );
  XOR U15000 ( .A(n12095), .B(n12096), .Z(n12070) );
  ANDN U15001 ( .B(n12097), .A(n12098), .Z(n12095) );
  XOR U15002 ( .A(n12096), .B(n12099), .Z(n12097) );
  IV U15003 ( .A(n12078), .Z(n12082) );
  XOR U15004 ( .A(n12078), .B(n12060), .Z(n12080) );
  XOR U15005 ( .A(n12100), .B(n12101), .Z(n12060) );
  AND U15006 ( .A(n82), .B(n12102), .Z(n12100) );
  XOR U15007 ( .A(n12103), .B(n12101), .Z(n12102) );
  NANDN U15008 ( .A(n12062), .B(n12064), .Z(n12078) );
  XOR U15009 ( .A(n12104), .B(n12105), .Z(n12064) );
  AND U15010 ( .A(n82), .B(n12106), .Z(n12104) );
  XOR U15011 ( .A(n12105), .B(n12107), .Z(n12106) );
  XOR U15012 ( .A(n12108), .B(n12109), .Z(n82) );
  AND U15013 ( .A(n12110), .B(n12111), .Z(n12108) );
  XNOR U15014 ( .A(n12109), .B(n12075), .Z(n12111) );
  XNOR U15015 ( .A(n12112), .B(n12113), .Z(n12075) );
  ANDN U15016 ( .B(n12114), .A(n12115), .Z(n12112) );
  XOR U15017 ( .A(n12113), .B(n12116), .Z(n12114) );
  XOR U15018 ( .A(n12109), .B(n12077), .Z(n12110) );
  XOR U15019 ( .A(n12117), .B(n12118), .Z(n12077) );
  AND U15020 ( .A(n86), .B(n12119), .Z(n12117) );
  XOR U15021 ( .A(n12120), .B(n12118), .Z(n12119) );
  XNOR U15022 ( .A(n12121), .B(n12122), .Z(n12109) );
  NAND U15023 ( .A(n12123), .B(n12124), .Z(n12122) );
  XOR U15024 ( .A(n12125), .B(n12101), .Z(n12124) );
  XOR U15025 ( .A(n12115), .B(n12116), .Z(n12101) );
  XOR U15026 ( .A(n12126), .B(n12127), .Z(n12116) );
  ANDN U15027 ( .B(n12128), .A(n12129), .Z(n12126) );
  XOR U15028 ( .A(n12127), .B(n12130), .Z(n12128) );
  XOR U15029 ( .A(n12131), .B(n12132), .Z(n12115) );
  XOR U15030 ( .A(n12133), .B(n12134), .Z(n12132) );
  ANDN U15031 ( .B(n12135), .A(n12136), .Z(n12133) );
  XOR U15032 ( .A(n12137), .B(n12134), .Z(n12135) );
  IV U15033 ( .A(n12113), .Z(n12131) );
  XOR U15034 ( .A(n12138), .B(n12139), .Z(n12113) );
  ANDN U15035 ( .B(n12140), .A(n12141), .Z(n12138) );
  XOR U15036 ( .A(n12139), .B(n12142), .Z(n12140) );
  IV U15037 ( .A(n12121), .Z(n12125) );
  XOR U15038 ( .A(n12121), .B(n12103), .Z(n12123) );
  XOR U15039 ( .A(n12143), .B(n12144), .Z(n12103) );
  AND U15040 ( .A(n86), .B(n12145), .Z(n12143) );
  XOR U15041 ( .A(n12146), .B(n12144), .Z(n12145) );
  NANDN U15042 ( .A(n12105), .B(n12107), .Z(n12121) );
  XOR U15043 ( .A(n12147), .B(n12148), .Z(n12107) );
  AND U15044 ( .A(n86), .B(n12149), .Z(n12147) );
  XOR U15045 ( .A(n12148), .B(n12150), .Z(n12149) );
  XOR U15046 ( .A(n12151), .B(n12152), .Z(n86) );
  AND U15047 ( .A(n12153), .B(n12154), .Z(n12151) );
  XNOR U15048 ( .A(n12152), .B(n12118), .Z(n12154) );
  XNOR U15049 ( .A(n12155), .B(n12156), .Z(n12118) );
  ANDN U15050 ( .B(n12157), .A(n12158), .Z(n12155) );
  XOR U15051 ( .A(n12156), .B(n12159), .Z(n12157) );
  XOR U15052 ( .A(n12152), .B(n12120), .Z(n12153) );
  XOR U15053 ( .A(n12160), .B(n12161), .Z(n12120) );
  AND U15054 ( .A(n90), .B(n12162), .Z(n12160) );
  XOR U15055 ( .A(n12163), .B(n12161), .Z(n12162) );
  XNOR U15056 ( .A(n12164), .B(n12165), .Z(n12152) );
  NAND U15057 ( .A(n12166), .B(n12167), .Z(n12165) );
  XOR U15058 ( .A(n12168), .B(n12144), .Z(n12167) );
  XOR U15059 ( .A(n12158), .B(n12159), .Z(n12144) );
  XOR U15060 ( .A(n12169), .B(n12170), .Z(n12159) );
  ANDN U15061 ( .B(n12171), .A(n12172), .Z(n12169) );
  XOR U15062 ( .A(n12170), .B(n12173), .Z(n12171) );
  XOR U15063 ( .A(n12174), .B(n12175), .Z(n12158) );
  XOR U15064 ( .A(n12176), .B(n12177), .Z(n12175) );
  ANDN U15065 ( .B(n12178), .A(n12179), .Z(n12176) );
  XOR U15066 ( .A(n12180), .B(n12177), .Z(n12178) );
  IV U15067 ( .A(n12156), .Z(n12174) );
  XOR U15068 ( .A(n12181), .B(n12182), .Z(n12156) );
  ANDN U15069 ( .B(n12183), .A(n12184), .Z(n12181) );
  XOR U15070 ( .A(n12182), .B(n12185), .Z(n12183) );
  IV U15071 ( .A(n12164), .Z(n12168) );
  XOR U15072 ( .A(n12164), .B(n12146), .Z(n12166) );
  XOR U15073 ( .A(n12186), .B(n12187), .Z(n12146) );
  AND U15074 ( .A(n90), .B(n12188), .Z(n12186) );
  XOR U15075 ( .A(n12189), .B(n12187), .Z(n12188) );
  NANDN U15076 ( .A(n12148), .B(n12150), .Z(n12164) );
  XOR U15077 ( .A(n12190), .B(n12191), .Z(n12150) );
  AND U15078 ( .A(n90), .B(n12192), .Z(n12190) );
  XOR U15079 ( .A(n12191), .B(n12193), .Z(n12192) );
  XOR U15080 ( .A(n12194), .B(n12195), .Z(n90) );
  AND U15081 ( .A(n12196), .B(n12197), .Z(n12194) );
  XNOR U15082 ( .A(n12195), .B(n12161), .Z(n12197) );
  XNOR U15083 ( .A(n12198), .B(n12199), .Z(n12161) );
  ANDN U15084 ( .B(n12200), .A(n12201), .Z(n12198) );
  XOR U15085 ( .A(n12199), .B(n12202), .Z(n12200) );
  XOR U15086 ( .A(n12195), .B(n12163), .Z(n12196) );
  XOR U15087 ( .A(n12203), .B(n12204), .Z(n12163) );
  AND U15088 ( .A(n94), .B(n12205), .Z(n12203) );
  XOR U15089 ( .A(n12206), .B(n12204), .Z(n12205) );
  XNOR U15090 ( .A(n12207), .B(n12208), .Z(n12195) );
  NAND U15091 ( .A(n12209), .B(n12210), .Z(n12208) );
  XOR U15092 ( .A(n12211), .B(n12187), .Z(n12210) );
  XOR U15093 ( .A(n12201), .B(n12202), .Z(n12187) );
  XOR U15094 ( .A(n12212), .B(n12213), .Z(n12202) );
  ANDN U15095 ( .B(n12214), .A(n12215), .Z(n12212) );
  XOR U15096 ( .A(n12213), .B(n12216), .Z(n12214) );
  XOR U15097 ( .A(n12217), .B(n12218), .Z(n12201) );
  XOR U15098 ( .A(n12219), .B(n12220), .Z(n12218) );
  ANDN U15099 ( .B(n12221), .A(n12222), .Z(n12219) );
  XOR U15100 ( .A(n12223), .B(n12220), .Z(n12221) );
  IV U15101 ( .A(n12199), .Z(n12217) );
  XOR U15102 ( .A(n12224), .B(n12225), .Z(n12199) );
  ANDN U15103 ( .B(n12226), .A(n12227), .Z(n12224) );
  XOR U15104 ( .A(n12225), .B(n12228), .Z(n12226) );
  IV U15105 ( .A(n12207), .Z(n12211) );
  XOR U15106 ( .A(n12207), .B(n12189), .Z(n12209) );
  XOR U15107 ( .A(n12229), .B(n12230), .Z(n12189) );
  AND U15108 ( .A(n94), .B(n12231), .Z(n12229) );
  XOR U15109 ( .A(n12232), .B(n12230), .Z(n12231) );
  NANDN U15110 ( .A(n12191), .B(n12193), .Z(n12207) );
  XOR U15111 ( .A(n12233), .B(n12234), .Z(n12193) );
  AND U15112 ( .A(n94), .B(n12235), .Z(n12233) );
  XOR U15113 ( .A(n12234), .B(n12236), .Z(n12235) );
  XOR U15114 ( .A(n12237), .B(n12238), .Z(n94) );
  AND U15115 ( .A(n12239), .B(n12240), .Z(n12237) );
  XNOR U15116 ( .A(n12238), .B(n12204), .Z(n12240) );
  XNOR U15117 ( .A(n12241), .B(n12242), .Z(n12204) );
  ANDN U15118 ( .B(n12243), .A(n12244), .Z(n12241) );
  XOR U15119 ( .A(n12242), .B(n12245), .Z(n12243) );
  XOR U15120 ( .A(n12238), .B(n12206), .Z(n12239) );
  XOR U15121 ( .A(n12246), .B(n12247), .Z(n12206) );
  AND U15122 ( .A(n98), .B(n12248), .Z(n12246) );
  XOR U15123 ( .A(n12249), .B(n12247), .Z(n12248) );
  XNOR U15124 ( .A(n12250), .B(n12251), .Z(n12238) );
  NAND U15125 ( .A(n12252), .B(n12253), .Z(n12251) );
  XOR U15126 ( .A(n12254), .B(n12230), .Z(n12253) );
  XOR U15127 ( .A(n12244), .B(n12245), .Z(n12230) );
  XOR U15128 ( .A(n12255), .B(n12256), .Z(n12245) );
  ANDN U15129 ( .B(n12257), .A(n12258), .Z(n12255) );
  XOR U15130 ( .A(n12256), .B(n12259), .Z(n12257) );
  XOR U15131 ( .A(n12260), .B(n12261), .Z(n12244) );
  XOR U15132 ( .A(n12262), .B(n12263), .Z(n12261) );
  ANDN U15133 ( .B(n12264), .A(n12265), .Z(n12262) );
  XOR U15134 ( .A(n12266), .B(n12263), .Z(n12264) );
  IV U15135 ( .A(n12242), .Z(n12260) );
  XOR U15136 ( .A(n12267), .B(n12268), .Z(n12242) );
  ANDN U15137 ( .B(n12269), .A(n12270), .Z(n12267) );
  XOR U15138 ( .A(n12268), .B(n12271), .Z(n12269) );
  IV U15139 ( .A(n12250), .Z(n12254) );
  XOR U15140 ( .A(n12250), .B(n12232), .Z(n12252) );
  XOR U15141 ( .A(n12272), .B(n12273), .Z(n12232) );
  AND U15142 ( .A(n98), .B(n12274), .Z(n12272) );
  XOR U15143 ( .A(n12275), .B(n12273), .Z(n12274) );
  NANDN U15144 ( .A(n12234), .B(n12236), .Z(n12250) );
  XOR U15145 ( .A(n12276), .B(n12277), .Z(n12236) );
  AND U15146 ( .A(n98), .B(n12278), .Z(n12276) );
  XOR U15147 ( .A(n12277), .B(n12279), .Z(n12278) );
  XOR U15148 ( .A(n12280), .B(n12281), .Z(n98) );
  AND U15149 ( .A(n12282), .B(n12283), .Z(n12280) );
  XNOR U15150 ( .A(n12281), .B(n12247), .Z(n12283) );
  XNOR U15151 ( .A(n12284), .B(n12285), .Z(n12247) );
  ANDN U15152 ( .B(n12286), .A(n12287), .Z(n12284) );
  XOR U15153 ( .A(n12285), .B(n12288), .Z(n12286) );
  XOR U15154 ( .A(n12281), .B(n12249), .Z(n12282) );
  XOR U15155 ( .A(n12289), .B(n12290), .Z(n12249) );
  AND U15156 ( .A(n102), .B(n12291), .Z(n12289) );
  XOR U15157 ( .A(n12292), .B(n12290), .Z(n12291) );
  XNOR U15158 ( .A(n12293), .B(n12294), .Z(n12281) );
  NAND U15159 ( .A(n12295), .B(n12296), .Z(n12294) );
  XOR U15160 ( .A(n12297), .B(n12273), .Z(n12296) );
  XOR U15161 ( .A(n12287), .B(n12288), .Z(n12273) );
  XOR U15162 ( .A(n12298), .B(n12299), .Z(n12288) );
  ANDN U15163 ( .B(n12300), .A(n12301), .Z(n12298) );
  XOR U15164 ( .A(n12299), .B(n12302), .Z(n12300) );
  XOR U15165 ( .A(n12303), .B(n12304), .Z(n12287) );
  XOR U15166 ( .A(n12305), .B(n12306), .Z(n12304) );
  ANDN U15167 ( .B(n12307), .A(n12308), .Z(n12305) );
  XOR U15168 ( .A(n12309), .B(n12306), .Z(n12307) );
  IV U15169 ( .A(n12285), .Z(n12303) );
  XOR U15170 ( .A(n12310), .B(n12311), .Z(n12285) );
  ANDN U15171 ( .B(n12312), .A(n12313), .Z(n12310) );
  XOR U15172 ( .A(n12311), .B(n12314), .Z(n12312) );
  IV U15173 ( .A(n12293), .Z(n12297) );
  XOR U15174 ( .A(n12293), .B(n12275), .Z(n12295) );
  XOR U15175 ( .A(n12315), .B(n12316), .Z(n12275) );
  AND U15176 ( .A(n102), .B(n12317), .Z(n12315) );
  XOR U15177 ( .A(n12318), .B(n12316), .Z(n12317) );
  NANDN U15178 ( .A(n12277), .B(n12279), .Z(n12293) );
  XOR U15179 ( .A(n12319), .B(n12320), .Z(n12279) );
  AND U15180 ( .A(n102), .B(n12321), .Z(n12319) );
  XOR U15181 ( .A(n12320), .B(n12322), .Z(n12321) );
  XOR U15182 ( .A(n12323), .B(n12324), .Z(n102) );
  AND U15183 ( .A(n12325), .B(n12326), .Z(n12323) );
  XNOR U15184 ( .A(n12324), .B(n12290), .Z(n12326) );
  XNOR U15185 ( .A(n12327), .B(n12328), .Z(n12290) );
  ANDN U15186 ( .B(n12329), .A(n12330), .Z(n12327) );
  XOR U15187 ( .A(n12328), .B(n12331), .Z(n12329) );
  XOR U15188 ( .A(n12324), .B(n12292), .Z(n12325) );
  XOR U15189 ( .A(n12332), .B(n12333), .Z(n12292) );
  AND U15190 ( .A(n106), .B(n12334), .Z(n12332) );
  XOR U15191 ( .A(n12335), .B(n12333), .Z(n12334) );
  XNOR U15192 ( .A(n12336), .B(n12337), .Z(n12324) );
  NAND U15193 ( .A(n12338), .B(n12339), .Z(n12337) );
  XOR U15194 ( .A(n12340), .B(n12316), .Z(n12339) );
  XOR U15195 ( .A(n12330), .B(n12331), .Z(n12316) );
  XOR U15196 ( .A(n12341), .B(n12342), .Z(n12331) );
  ANDN U15197 ( .B(n12343), .A(n12344), .Z(n12341) );
  XOR U15198 ( .A(n12342), .B(n12345), .Z(n12343) );
  XOR U15199 ( .A(n12346), .B(n12347), .Z(n12330) );
  XOR U15200 ( .A(n12348), .B(n12349), .Z(n12347) );
  ANDN U15201 ( .B(n12350), .A(n12351), .Z(n12348) );
  XOR U15202 ( .A(n12352), .B(n12349), .Z(n12350) );
  IV U15203 ( .A(n12328), .Z(n12346) );
  XOR U15204 ( .A(n12353), .B(n12354), .Z(n12328) );
  ANDN U15205 ( .B(n12355), .A(n12356), .Z(n12353) );
  XOR U15206 ( .A(n12354), .B(n12357), .Z(n12355) );
  IV U15207 ( .A(n12336), .Z(n12340) );
  XOR U15208 ( .A(n12336), .B(n12318), .Z(n12338) );
  XOR U15209 ( .A(n12358), .B(n12359), .Z(n12318) );
  AND U15210 ( .A(n106), .B(n12360), .Z(n12358) );
  XOR U15211 ( .A(n12361), .B(n12359), .Z(n12360) );
  NANDN U15212 ( .A(n12320), .B(n12322), .Z(n12336) );
  XOR U15213 ( .A(n12362), .B(n12363), .Z(n12322) );
  AND U15214 ( .A(n106), .B(n12364), .Z(n12362) );
  XOR U15215 ( .A(n12363), .B(n12365), .Z(n12364) );
  XOR U15216 ( .A(n12366), .B(n12367), .Z(n106) );
  AND U15217 ( .A(n12368), .B(n12369), .Z(n12366) );
  XNOR U15218 ( .A(n12367), .B(n12333), .Z(n12369) );
  XNOR U15219 ( .A(n12370), .B(n12371), .Z(n12333) );
  ANDN U15220 ( .B(n12372), .A(n12373), .Z(n12370) );
  XOR U15221 ( .A(n12371), .B(n12374), .Z(n12372) );
  XOR U15222 ( .A(n12367), .B(n12335), .Z(n12368) );
  XOR U15223 ( .A(n12375), .B(n12376), .Z(n12335) );
  AND U15224 ( .A(n110), .B(n12377), .Z(n12375) );
  XOR U15225 ( .A(n12378), .B(n12376), .Z(n12377) );
  XNOR U15226 ( .A(n12379), .B(n12380), .Z(n12367) );
  NAND U15227 ( .A(n12381), .B(n12382), .Z(n12380) );
  XOR U15228 ( .A(n12383), .B(n12359), .Z(n12382) );
  XOR U15229 ( .A(n12373), .B(n12374), .Z(n12359) );
  XOR U15230 ( .A(n12384), .B(n12385), .Z(n12374) );
  ANDN U15231 ( .B(n12386), .A(n12387), .Z(n12384) );
  XOR U15232 ( .A(n12385), .B(n12388), .Z(n12386) );
  XOR U15233 ( .A(n12389), .B(n12390), .Z(n12373) );
  XOR U15234 ( .A(n12391), .B(n12392), .Z(n12390) );
  ANDN U15235 ( .B(n12393), .A(n12394), .Z(n12391) );
  XOR U15236 ( .A(n12395), .B(n12392), .Z(n12393) );
  IV U15237 ( .A(n12371), .Z(n12389) );
  XOR U15238 ( .A(n12396), .B(n12397), .Z(n12371) );
  ANDN U15239 ( .B(n12398), .A(n12399), .Z(n12396) );
  XOR U15240 ( .A(n12397), .B(n12400), .Z(n12398) );
  IV U15241 ( .A(n12379), .Z(n12383) );
  XOR U15242 ( .A(n12379), .B(n12361), .Z(n12381) );
  XOR U15243 ( .A(n12401), .B(n12402), .Z(n12361) );
  AND U15244 ( .A(n110), .B(n12403), .Z(n12401) );
  XOR U15245 ( .A(n12404), .B(n12402), .Z(n12403) );
  NANDN U15246 ( .A(n12363), .B(n12365), .Z(n12379) );
  XOR U15247 ( .A(n12405), .B(n12406), .Z(n12365) );
  AND U15248 ( .A(n110), .B(n12407), .Z(n12405) );
  XOR U15249 ( .A(n12406), .B(n12408), .Z(n12407) );
  XOR U15250 ( .A(n12409), .B(n12410), .Z(n110) );
  AND U15251 ( .A(n12411), .B(n12412), .Z(n12409) );
  XNOR U15252 ( .A(n12410), .B(n12376), .Z(n12412) );
  XNOR U15253 ( .A(n12413), .B(n12414), .Z(n12376) );
  ANDN U15254 ( .B(n12415), .A(n12416), .Z(n12413) );
  XOR U15255 ( .A(n12414), .B(n12417), .Z(n12415) );
  XOR U15256 ( .A(n12410), .B(n12378), .Z(n12411) );
  XOR U15257 ( .A(n12418), .B(n12419), .Z(n12378) );
  AND U15258 ( .A(n114), .B(n12420), .Z(n12418) );
  XOR U15259 ( .A(n12421), .B(n12419), .Z(n12420) );
  XNOR U15260 ( .A(n12422), .B(n12423), .Z(n12410) );
  NAND U15261 ( .A(n12424), .B(n12425), .Z(n12423) );
  XOR U15262 ( .A(n12426), .B(n12402), .Z(n12425) );
  XOR U15263 ( .A(n12416), .B(n12417), .Z(n12402) );
  XOR U15264 ( .A(n12427), .B(n12428), .Z(n12417) );
  ANDN U15265 ( .B(n12429), .A(n12430), .Z(n12427) );
  XOR U15266 ( .A(n12428), .B(n12431), .Z(n12429) );
  XOR U15267 ( .A(n12432), .B(n12433), .Z(n12416) );
  XOR U15268 ( .A(n12434), .B(n12435), .Z(n12433) );
  ANDN U15269 ( .B(n12436), .A(n12437), .Z(n12434) );
  XOR U15270 ( .A(n12438), .B(n12435), .Z(n12436) );
  IV U15271 ( .A(n12414), .Z(n12432) );
  XOR U15272 ( .A(n12439), .B(n12440), .Z(n12414) );
  ANDN U15273 ( .B(n12441), .A(n12442), .Z(n12439) );
  XOR U15274 ( .A(n12440), .B(n12443), .Z(n12441) );
  IV U15275 ( .A(n12422), .Z(n12426) );
  XOR U15276 ( .A(n12422), .B(n12404), .Z(n12424) );
  XOR U15277 ( .A(n12444), .B(n12445), .Z(n12404) );
  AND U15278 ( .A(n114), .B(n12446), .Z(n12444) );
  XOR U15279 ( .A(n12447), .B(n12445), .Z(n12446) );
  NANDN U15280 ( .A(n12406), .B(n12408), .Z(n12422) );
  XOR U15281 ( .A(n12448), .B(n12449), .Z(n12408) );
  AND U15282 ( .A(n114), .B(n12450), .Z(n12448) );
  XOR U15283 ( .A(n12449), .B(n12451), .Z(n12450) );
  XOR U15284 ( .A(n12452), .B(n12453), .Z(n114) );
  AND U15285 ( .A(n12454), .B(n12455), .Z(n12452) );
  XNOR U15286 ( .A(n12453), .B(n12419), .Z(n12455) );
  XNOR U15287 ( .A(n12456), .B(n12457), .Z(n12419) );
  ANDN U15288 ( .B(n12458), .A(n12459), .Z(n12456) );
  XOR U15289 ( .A(n12457), .B(n12460), .Z(n12458) );
  XOR U15290 ( .A(n12453), .B(n12421), .Z(n12454) );
  XOR U15291 ( .A(n12461), .B(n12462), .Z(n12421) );
  AND U15292 ( .A(n118), .B(n12463), .Z(n12461) );
  XOR U15293 ( .A(n12464), .B(n12462), .Z(n12463) );
  XNOR U15294 ( .A(n12465), .B(n12466), .Z(n12453) );
  NAND U15295 ( .A(n12467), .B(n12468), .Z(n12466) );
  XOR U15296 ( .A(n12469), .B(n12445), .Z(n12468) );
  XOR U15297 ( .A(n12459), .B(n12460), .Z(n12445) );
  XOR U15298 ( .A(n12470), .B(n12471), .Z(n12460) );
  ANDN U15299 ( .B(n12472), .A(n12473), .Z(n12470) );
  XOR U15300 ( .A(n12471), .B(n12474), .Z(n12472) );
  XOR U15301 ( .A(n12475), .B(n12476), .Z(n12459) );
  XOR U15302 ( .A(n12477), .B(n12478), .Z(n12476) );
  ANDN U15303 ( .B(n12479), .A(n12480), .Z(n12477) );
  XOR U15304 ( .A(n12481), .B(n12478), .Z(n12479) );
  IV U15305 ( .A(n12457), .Z(n12475) );
  XOR U15306 ( .A(n12482), .B(n12483), .Z(n12457) );
  ANDN U15307 ( .B(n12484), .A(n12485), .Z(n12482) );
  XOR U15308 ( .A(n12483), .B(n12486), .Z(n12484) );
  IV U15309 ( .A(n12465), .Z(n12469) );
  XOR U15310 ( .A(n12465), .B(n12447), .Z(n12467) );
  XOR U15311 ( .A(n12487), .B(n12488), .Z(n12447) );
  AND U15312 ( .A(n118), .B(n12489), .Z(n12487) );
  XOR U15313 ( .A(n12490), .B(n12488), .Z(n12489) );
  NANDN U15314 ( .A(n12449), .B(n12451), .Z(n12465) );
  XOR U15315 ( .A(n12491), .B(n12492), .Z(n12451) );
  AND U15316 ( .A(n118), .B(n12493), .Z(n12491) );
  XOR U15317 ( .A(n12492), .B(n12494), .Z(n12493) );
  XOR U15318 ( .A(n12495), .B(n12496), .Z(n118) );
  AND U15319 ( .A(n12497), .B(n12498), .Z(n12495) );
  XNOR U15320 ( .A(n12496), .B(n12462), .Z(n12498) );
  XNOR U15321 ( .A(n12499), .B(n12500), .Z(n12462) );
  ANDN U15322 ( .B(n12501), .A(n12502), .Z(n12499) );
  XOR U15323 ( .A(n12500), .B(n12503), .Z(n12501) );
  XOR U15324 ( .A(n12496), .B(n12464), .Z(n12497) );
  XOR U15325 ( .A(n12504), .B(n12505), .Z(n12464) );
  AND U15326 ( .A(n122), .B(n12506), .Z(n12504) );
  XOR U15327 ( .A(n12507), .B(n12505), .Z(n12506) );
  XNOR U15328 ( .A(n12508), .B(n12509), .Z(n12496) );
  NAND U15329 ( .A(n12510), .B(n12511), .Z(n12509) );
  XOR U15330 ( .A(n12512), .B(n12488), .Z(n12511) );
  XOR U15331 ( .A(n12502), .B(n12503), .Z(n12488) );
  XOR U15332 ( .A(n12513), .B(n12514), .Z(n12503) );
  ANDN U15333 ( .B(n12515), .A(n12516), .Z(n12513) );
  XOR U15334 ( .A(n12514), .B(n12517), .Z(n12515) );
  XOR U15335 ( .A(n12518), .B(n12519), .Z(n12502) );
  XOR U15336 ( .A(n12520), .B(n12521), .Z(n12519) );
  ANDN U15337 ( .B(n12522), .A(n12523), .Z(n12520) );
  XOR U15338 ( .A(n12524), .B(n12521), .Z(n12522) );
  IV U15339 ( .A(n12500), .Z(n12518) );
  XOR U15340 ( .A(n12525), .B(n12526), .Z(n12500) );
  ANDN U15341 ( .B(n12527), .A(n12528), .Z(n12525) );
  XOR U15342 ( .A(n12526), .B(n12529), .Z(n12527) );
  IV U15343 ( .A(n12508), .Z(n12512) );
  XOR U15344 ( .A(n12508), .B(n12490), .Z(n12510) );
  XOR U15345 ( .A(n12530), .B(n12531), .Z(n12490) );
  AND U15346 ( .A(n122), .B(n12532), .Z(n12530) );
  XOR U15347 ( .A(n12533), .B(n12531), .Z(n12532) );
  NANDN U15348 ( .A(n12492), .B(n12494), .Z(n12508) );
  XOR U15349 ( .A(n12534), .B(n12535), .Z(n12494) );
  AND U15350 ( .A(n122), .B(n12536), .Z(n12534) );
  XOR U15351 ( .A(n12535), .B(n12537), .Z(n12536) );
  XOR U15352 ( .A(n12538), .B(n12539), .Z(n122) );
  AND U15353 ( .A(n12540), .B(n12541), .Z(n12538) );
  XNOR U15354 ( .A(n12539), .B(n12505), .Z(n12541) );
  XNOR U15355 ( .A(n12542), .B(n12543), .Z(n12505) );
  ANDN U15356 ( .B(n12544), .A(n12545), .Z(n12542) );
  XOR U15357 ( .A(n12543), .B(n12546), .Z(n12544) );
  XOR U15358 ( .A(n12539), .B(n12507), .Z(n12540) );
  XOR U15359 ( .A(n12547), .B(n12548), .Z(n12507) );
  AND U15360 ( .A(n126), .B(n12549), .Z(n12547) );
  XOR U15361 ( .A(n12550), .B(n12548), .Z(n12549) );
  XNOR U15362 ( .A(n12551), .B(n12552), .Z(n12539) );
  NAND U15363 ( .A(n12553), .B(n12554), .Z(n12552) );
  XOR U15364 ( .A(n12555), .B(n12531), .Z(n12554) );
  XOR U15365 ( .A(n12545), .B(n12546), .Z(n12531) );
  XOR U15366 ( .A(n12556), .B(n12557), .Z(n12546) );
  ANDN U15367 ( .B(n12558), .A(n12559), .Z(n12556) );
  XOR U15368 ( .A(n12557), .B(n12560), .Z(n12558) );
  XOR U15369 ( .A(n12561), .B(n12562), .Z(n12545) );
  XOR U15370 ( .A(n12563), .B(n12564), .Z(n12562) );
  ANDN U15371 ( .B(n12565), .A(n12566), .Z(n12563) );
  XOR U15372 ( .A(n12567), .B(n12564), .Z(n12565) );
  IV U15373 ( .A(n12543), .Z(n12561) );
  XOR U15374 ( .A(n12568), .B(n12569), .Z(n12543) );
  ANDN U15375 ( .B(n12570), .A(n12571), .Z(n12568) );
  XOR U15376 ( .A(n12569), .B(n12572), .Z(n12570) );
  IV U15377 ( .A(n12551), .Z(n12555) );
  XOR U15378 ( .A(n12551), .B(n12533), .Z(n12553) );
  XOR U15379 ( .A(n12573), .B(n12574), .Z(n12533) );
  AND U15380 ( .A(n126), .B(n12575), .Z(n12573) );
  XOR U15381 ( .A(n12576), .B(n12574), .Z(n12575) );
  NANDN U15382 ( .A(n12535), .B(n12537), .Z(n12551) );
  XOR U15383 ( .A(n12577), .B(n12578), .Z(n12537) );
  AND U15384 ( .A(n126), .B(n12579), .Z(n12577) );
  XOR U15385 ( .A(n12578), .B(n12580), .Z(n12579) );
  XOR U15386 ( .A(n12581), .B(n12582), .Z(n126) );
  AND U15387 ( .A(n12583), .B(n12584), .Z(n12581) );
  XNOR U15388 ( .A(n12582), .B(n12548), .Z(n12584) );
  XNOR U15389 ( .A(n12585), .B(n12586), .Z(n12548) );
  ANDN U15390 ( .B(n12587), .A(n12588), .Z(n12585) );
  XOR U15391 ( .A(n12586), .B(n12589), .Z(n12587) );
  XOR U15392 ( .A(n12582), .B(n12550), .Z(n12583) );
  XOR U15393 ( .A(n12590), .B(n12591), .Z(n12550) );
  AND U15394 ( .A(n130), .B(n12592), .Z(n12590) );
  XOR U15395 ( .A(n12593), .B(n12591), .Z(n12592) );
  XNOR U15396 ( .A(n12594), .B(n12595), .Z(n12582) );
  NAND U15397 ( .A(n12596), .B(n12597), .Z(n12595) );
  XOR U15398 ( .A(n12598), .B(n12574), .Z(n12597) );
  XOR U15399 ( .A(n12588), .B(n12589), .Z(n12574) );
  XOR U15400 ( .A(n12599), .B(n12600), .Z(n12589) );
  ANDN U15401 ( .B(n12601), .A(n12602), .Z(n12599) );
  XOR U15402 ( .A(n12600), .B(n12603), .Z(n12601) );
  XOR U15403 ( .A(n12604), .B(n12605), .Z(n12588) );
  XOR U15404 ( .A(n12606), .B(n12607), .Z(n12605) );
  ANDN U15405 ( .B(n12608), .A(n12609), .Z(n12606) );
  XOR U15406 ( .A(n12610), .B(n12607), .Z(n12608) );
  IV U15407 ( .A(n12586), .Z(n12604) );
  XOR U15408 ( .A(n12611), .B(n12612), .Z(n12586) );
  ANDN U15409 ( .B(n12613), .A(n12614), .Z(n12611) );
  XOR U15410 ( .A(n12612), .B(n12615), .Z(n12613) );
  IV U15411 ( .A(n12594), .Z(n12598) );
  XOR U15412 ( .A(n12594), .B(n12576), .Z(n12596) );
  XOR U15413 ( .A(n12616), .B(n12617), .Z(n12576) );
  AND U15414 ( .A(n130), .B(n12618), .Z(n12616) );
  XOR U15415 ( .A(n12619), .B(n12617), .Z(n12618) );
  NANDN U15416 ( .A(n12578), .B(n12580), .Z(n12594) );
  XOR U15417 ( .A(n12620), .B(n12621), .Z(n12580) );
  AND U15418 ( .A(n130), .B(n12622), .Z(n12620) );
  XOR U15419 ( .A(n12621), .B(n12623), .Z(n12622) );
  XOR U15420 ( .A(n12624), .B(n12625), .Z(n130) );
  AND U15421 ( .A(n12626), .B(n12627), .Z(n12624) );
  XNOR U15422 ( .A(n12625), .B(n12591), .Z(n12627) );
  XNOR U15423 ( .A(n12628), .B(n12629), .Z(n12591) );
  ANDN U15424 ( .B(n12630), .A(n12631), .Z(n12628) );
  XOR U15425 ( .A(n12629), .B(n12632), .Z(n12630) );
  XOR U15426 ( .A(n12625), .B(n12593), .Z(n12626) );
  XOR U15427 ( .A(n12633), .B(n12634), .Z(n12593) );
  AND U15428 ( .A(n134), .B(n12635), .Z(n12633) );
  XOR U15429 ( .A(n12636), .B(n12634), .Z(n12635) );
  XNOR U15430 ( .A(n12637), .B(n12638), .Z(n12625) );
  NAND U15431 ( .A(n12639), .B(n12640), .Z(n12638) );
  XOR U15432 ( .A(n12641), .B(n12617), .Z(n12640) );
  XOR U15433 ( .A(n12631), .B(n12632), .Z(n12617) );
  XOR U15434 ( .A(n12642), .B(n12643), .Z(n12632) );
  ANDN U15435 ( .B(n12644), .A(n12645), .Z(n12642) );
  XOR U15436 ( .A(n12643), .B(n12646), .Z(n12644) );
  XOR U15437 ( .A(n12647), .B(n12648), .Z(n12631) );
  XOR U15438 ( .A(n12649), .B(n12650), .Z(n12648) );
  ANDN U15439 ( .B(n12651), .A(n12652), .Z(n12649) );
  XOR U15440 ( .A(n12653), .B(n12650), .Z(n12651) );
  IV U15441 ( .A(n12629), .Z(n12647) );
  XOR U15442 ( .A(n12654), .B(n12655), .Z(n12629) );
  ANDN U15443 ( .B(n12656), .A(n12657), .Z(n12654) );
  XOR U15444 ( .A(n12655), .B(n12658), .Z(n12656) );
  IV U15445 ( .A(n12637), .Z(n12641) );
  XOR U15446 ( .A(n12637), .B(n12619), .Z(n12639) );
  XOR U15447 ( .A(n12659), .B(n12660), .Z(n12619) );
  AND U15448 ( .A(n134), .B(n12661), .Z(n12659) );
  XOR U15449 ( .A(n12662), .B(n12660), .Z(n12661) );
  NANDN U15450 ( .A(n12621), .B(n12623), .Z(n12637) );
  XOR U15451 ( .A(n12663), .B(n12664), .Z(n12623) );
  AND U15452 ( .A(n134), .B(n12665), .Z(n12663) );
  XOR U15453 ( .A(n12664), .B(n12666), .Z(n12665) );
  XOR U15454 ( .A(n12667), .B(n12668), .Z(n134) );
  AND U15455 ( .A(n12669), .B(n12670), .Z(n12667) );
  XNOR U15456 ( .A(n12668), .B(n12634), .Z(n12670) );
  XNOR U15457 ( .A(n12671), .B(n12672), .Z(n12634) );
  ANDN U15458 ( .B(n12673), .A(n12674), .Z(n12671) );
  XOR U15459 ( .A(n12672), .B(n12675), .Z(n12673) );
  XOR U15460 ( .A(n12668), .B(n12636), .Z(n12669) );
  XOR U15461 ( .A(n12676), .B(n12677), .Z(n12636) );
  AND U15462 ( .A(n138), .B(n12678), .Z(n12676) );
  XOR U15463 ( .A(n12679), .B(n12677), .Z(n12678) );
  XNOR U15464 ( .A(n12680), .B(n12681), .Z(n12668) );
  NAND U15465 ( .A(n12682), .B(n12683), .Z(n12681) );
  XOR U15466 ( .A(n12684), .B(n12660), .Z(n12683) );
  XOR U15467 ( .A(n12674), .B(n12675), .Z(n12660) );
  XOR U15468 ( .A(n12685), .B(n12686), .Z(n12675) );
  ANDN U15469 ( .B(n12687), .A(n12688), .Z(n12685) );
  XOR U15470 ( .A(n12686), .B(n12689), .Z(n12687) );
  XOR U15471 ( .A(n12690), .B(n12691), .Z(n12674) );
  XOR U15472 ( .A(n12692), .B(n12693), .Z(n12691) );
  ANDN U15473 ( .B(n12694), .A(n12695), .Z(n12692) );
  XOR U15474 ( .A(n12696), .B(n12693), .Z(n12694) );
  IV U15475 ( .A(n12672), .Z(n12690) );
  XOR U15476 ( .A(n12697), .B(n12698), .Z(n12672) );
  ANDN U15477 ( .B(n12699), .A(n12700), .Z(n12697) );
  XOR U15478 ( .A(n12698), .B(n12701), .Z(n12699) );
  IV U15479 ( .A(n12680), .Z(n12684) );
  XOR U15480 ( .A(n12680), .B(n12662), .Z(n12682) );
  XOR U15481 ( .A(n12702), .B(n12703), .Z(n12662) );
  AND U15482 ( .A(n138), .B(n12704), .Z(n12702) );
  XOR U15483 ( .A(n12705), .B(n12703), .Z(n12704) );
  NANDN U15484 ( .A(n12664), .B(n12666), .Z(n12680) );
  XOR U15485 ( .A(n12706), .B(n12707), .Z(n12666) );
  AND U15486 ( .A(n138), .B(n12708), .Z(n12706) );
  XOR U15487 ( .A(n12707), .B(n12709), .Z(n12708) );
  XOR U15488 ( .A(n12710), .B(n12711), .Z(n138) );
  AND U15489 ( .A(n12712), .B(n12713), .Z(n12710) );
  XNOR U15490 ( .A(n12711), .B(n12677), .Z(n12713) );
  XNOR U15491 ( .A(n12714), .B(n12715), .Z(n12677) );
  ANDN U15492 ( .B(n12716), .A(n12717), .Z(n12714) );
  XOR U15493 ( .A(n12715), .B(n12718), .Z(n12716) );
  XOR U15494 ( .A(n12711), .B(n12679), .Z(n12712) );
  XOR U15495 ( .A(n12719), .B(n12720), .Z(n12679) );
  AND U15496 ( .A(n142), .B(n12721), .Z(n12719) );
  XOR U15497 ( .A(n12722), .B(n12720), .Z(n12721) );
  XNOR U15498 ( .A(n12723), .B(n12724), .Z(n12711) );
  NAND U15499 ( .A(n12725), .B(n12726), .Z(n12724) );
  XOR U15500 ( .A(n12727), .B(n12703), .Z(n12726) );
  XOR U15501 ( .A(n12717), .B(n12718), .Z(n12703) );
  XOR U15502 ( .A(n12728), .B(n12729), .Z(n12718) );
  ANDN U15503 ( .B(n12730), .A(n12731), .Z(n12728) );
  XOR U15504 ( .A(n12729), .B(n12732), .Z(n12730) );
  XOR U15505 ( .A(n12733), .B(n12734), .Z(n12717) );
  XOR U15506 ( .A(n12735), .B(n12736), .Z(n12734) );
  ANDN U15507 ( .B(n12737), .A(n12738), .Z(n12735) );
  XOR U15508 ( .A(n12739), .B(n12736), .Z(n12737) );
  IV U15509 ( .A(n12715), .Z(n12733) );
  XOR U15510 ( .A(n12740), .B(n12741), .Z(n12715) );
  ANDN U15511 ( .B(n12742), .A(n12743), .Z(n12740) );
  XOR U15512 ( .A(n12741), .B(n12744), .Z(n12742) );
  IV U15513 ( .A(n12723), .Z(n12727) );
  XOR U15514 ( .A(n12723), .B(n12705), .Z(n12725) );
  XOR U15515 ( .A(n12745), .B(n12746), .Z(n12705) );
  AND U15516 ( .A(n142), .B(n12747), .Z(n12745) );
  XOR U15517 ( .A(n12748), .B(n12746), .Z(n12747) );
  NANDN U15518 ( .A(n12707), .B(n12709), .Z(n12723) );
  XOR U15519 ( .A(n12749), .B(n12750), .Z(n12709) );
  AND U15520 ( .A(n142), .B(n12751), .Z(n12749) );
  XOR U15521 ( .A(n12750), .B(n12752), .Z(n12751) );
  XOR U15522 ( .A(n12753), .B(n12754), .Z(n142) );
  AND U15523 ( .A(n12755), .B(n12756), .Z(n12753) );
  XNOR U15524 ( .A(n12754), .B(n12720), .Z(n12756) );
  XNOR U15525 ( .A(n12757), .B(n12758), .Z(n12720) );
  ANDN U15526 ( .B(n12759), .A(n12760), .Z(n12757) );
  XOR U15527 ( .A(n12758), .B(n12761), .Z(n12759) );
  XOR U15528 ( .A(n12754), .B(n12722), .Z(n12755) );
  XOR U15529 ( .A(n12762), .B(n12763), .Z(n12722) );
  AND U15530 ( .A(n146), .B(n12764), .Z(n12762) );
  XOR U15531 ( .A(n12765), .B(n12763), .Z(n12764) );
  XNOR U15532 ( .A(n12766), .B(n12767), .Z(n12754) );
  NAND U15533 ( .A(n12768), .B(n12769), .Z(n12767) );
  XOR U15534 ( .A(n12770), .B(n12746), .Z(n12769) );
  XOR U15535 ( .A(n12760), .B(n12761), .Z(n12746) );
  XOR U15536 ( .A(n12771), .B(n12772), .Z(n12761) );
  ANDN U15537 ( .B(n12773), .A(n12774), .Z(n12771) );
  XOR U15538 ( .A(n12772), .B(n12775), .Z(n12773) );
  XOR U15539 ( .A(n12776), .B(n12777), .Z(n12760) );
  XOR U15540 ( .A(n12778), .B(n12779), .Z(n12777) );
  ANDN U15541 ( .B(n12780), .A(n12781), .Z(n12778) );
  XOR U15542 ( .A(n12782), .B(n12779), .Z(n12780) );
  IV U15543 ( .A(n12758), .Z(n12776) );
  XOR U15544 ( .A(n12783), .B(n12784), .Z(n12758) );
  ANDN U15545 ( .B(n12785), .A(n12786), .Z(n12783) );
  XOR U15546 ( .A(n12784), .B(n12787), .Z(n12785) );
  IV U15547 ( .A(n12766), .Z(n12770) );
  XOR U15548 ( .A(n12766), .B(n12748), .Z(n12768) );
  XOR U15549 ( .A(n12788), .B(n12789), .Z(n12748) );
  AND U15550 ( .A(n146), .B(n12790), .Z(n12788) );
  XOR U15551 ( .A(n12791), .B(n12789), .Z(n12790) );
  NANDN U15552 ( .A(n12750), .B(n12752), .Z(n12766) );
  XOR U15553 ( .A(n12792), .B(n12793), .Z(n12752) );
  AND U15554 ( .A(n146), .B(n12794), .Z(n12792) );
  XOR U15555 ( .A(n12793), .B(n12795), .Z(n12794) );
  XOR U15556 ( .A(n12796), .B(n12797), .Z(n146) );
  AND U15557 ( .A(n12798), .B(n12799), .Z(n12796) );
  XNOR U15558 ( .A(n12797), .B(n12763), .Z(n12799) );
  XNOR U15559 ( .A(n12800), .B(n12801), .Z(n12763) );
  ANDN U15560 ( .B(n12802), .A(n12803), .Z(n12800) );
  XOR U15561 ( .A(n12801), .B(n12804), .Z(n12802) );
  XOR U15562 ( .A(n12797), .B(n12765), .Z(n12798) );
  XOR U15563 ( .A(n12805), .B(n12806), .Z(n12765) );
  AND U15564 ( .A(n150), .B(n12807), .Z(n12805) );
  XOR U15565 ( .A(n12808), .B(n12806), .Z(n12807) );
  XNOR U15566 ( .A(n12809), .B(n12810), .Z(n12797) );
  NAND U15567 ( .A(n12811), .B(n12812), .Z(n12810) );
  XOR U15568 ( .A(n12813), .B(n12789), .Z(n12812) );
  XOR U15569 ( .A(n12803), .B(n12804), .Z(n12789) );
  XOR U15570 ( .A(n12814), .B(n12815), .Z(n12804) );
  ANDN U15571 ( .B(n12816), .A(n12817), .Z(n12814) );
  XOR U15572 ( .A(n12815), .B(n12818), .Z(n12816) );
  XOR U15573 ( .A(n12819), .B(n12820), .Z(n12803) );
  XOR U15574 ( .A(n12821), .B(n12822), .Z(n12820) );
  ANDN U15575 ( .B(n12823), .A(n12824), .Z(n12821) );
  XOR U15576 ( .A(n12825), .B(n12822), .Z(n12823) );
  IV U15577 ( .A(n12801), .Z(n12819) );
  XOR U15578 ( .A(n12826), .B(n12827), .Z(n12801) );
  ANDN U15579 ( .B(n12828), .A(n12829), .Z(n12826) );
  XOR U15580 ( .A(n12827), .B(n12830), .Z(n12828) );
  IV U15581 ( .A(n12809), .Z(n12813) );
  XOR U15582 ( .A(n12809), .B(n12791), .Z(n12811) );
  XOR U15583 ( .A(n12831), .B(n12832), .Z(n12791) );
  AND U15584 ( .A(n150), .B(n12833), .Z(n12831) );
  XOR U15585 ( .A(n12834), .B(n12832), .Z(n12833) );
  NANDN U15586 ( .A(n12793), .B(n12795), .Z(n12809) );
  XOR U15587 ( .A(n12835), .B(n12836), .Z(n12795) );
  AND U15588 ( .A(n150), .B(n12837), .Z(n12835) );
  XOR U15589 ( .A(n12836), .B(n12838), .Z(n12837) );
  XOR U15590 ( .A(n12839), .B(n12840), .Z(n150) );
  AND U15591 ( .A(n12841), .B(n12842), .Z(n12839) );
  XNOR U15592 ( .A(n12840), .B(n12806), .Z(n12842) );
  XNOR U15593 ( .A(n12843), .B(n12844), .Z(n12806) );
  ANDN U15594 ( .B(n12845), .A(n12846), .Z(n12843) );
  XOR U15595 ( .A(n12844), .B(n12847), .Z(n12845) );
  XOR U15596 ( .A(n12840), .B(n12808), .Z(n12841) );
  XOR U15597 ( .A(n12848), .B(n12849), .Z(n12808) );
  AND U15598 ( .A(n154), .B(n12850), .Z(n12848) );
  XOR U15599 ( .A(n12851), .B(n12849), .Z(n12850) );
  XNOR U15600 ( .A(n12852), .B(n12853), .Z(n12840) );
  NAND U15601 ( .A(n12854), .B(n12855), .Z(n12853) );
  XOR U15602 ( .A(n12856), .B(n12832), .Z(n12855) );
  XOR U15603 ( .A(n12846), .B(n12847), .Z(n12832) );
  XOR U15604 ( .A(n12857), .B(n12858), .Z(n12847) );
  ANDN U15605 ( .B(n12859), .A(n12860), .Z(n12857) );
  XOR U15606 ( .A(n12858), .B(n12861), .Z(n12859) );
  XOR U15607 ( .A(n12862), .B(n12863), .Z(n12846) );
  XOR U15608 ( .A(n12864), .B(n12865), .Z(n12863) );
  ANDN U15609 ( .B(n12866), .A(n12867), .Z(n12864) );
  XOR U15610 ( .A(n12868), .B(n12865), .Z(n12866) );
  IV U15611 ( .A(n12844), .Z(n12862) );
  XOR U15612 ( .A(n12869), .B(n12870), .Z(n12844) );
  ANDN U15613 ( .B(n12871), .A(n12872), .Z(n12869) );
  XOR U15614 ( .A(n12870), .B(n12873), .Z(n12871) );
  IV U15615 ( .A(n12852), .Z(n12856) );
  XOR U15616 ( .A(n12852), .B(n12834), .Z(n12854) );
  XOR U15617 ( .A(n12874), .B(n12875), .Z(n12834) );
  AND U15618 ( .A(n154), .B(n12876), .Z(n12874) );
  XOR U15619 ( .A(n12877), .B(n12875), .Z(n12876) );
  NANDN U15620 ( .A(n12836), .B(n12838), .Z(n12852) );
  XOR U15621 ( .A(n12878), .B(n12879), .Z(n12838) );
  AND U15622 ( .A(n154), .B(n12880), .Z(n12878) );
  XOR U15623 ( .A(n12879), .B(n12881), .Z(n12880) );
  XOR U15624 ( .A(n12882), .B(n12883), .Z(n154) );
  AND U15625 ( .A(n12884), .B(n12885), .Z(n12882) );
  XNOR U15626 ( .A(n12883), .B(n12849), .Z(n12885) );
  XNOR U15627 ( .A(n12886), .B(n12887), .Z(n12849) );
  ANDN U15628 ( .B(n12888), .A(n12889), .Z(n12886) );
  XOR U15629 ( .A(n12887), .B(n12890), .Z(n12888) );
  XOR U15630 ( .A(n12883), .B(n12851), .Z(n12884) );
  XOR U15631 ( .A(n12891), .B(n12892), .Z(n12851) );
  AND U15632 ( .A(n158), .B(n12893), .Z(n12891) );
  XOR U15633 ( .A(n12894), .B(n12892), .Z(n12893) );
  XNOR U15634 ( .A(n12895), .B(n12896), .Z(n12883) );
  NAND U15635 ( .A(n12897), .B(n12898), .Z(n12896) );
  XOR U15636 ( .A(n12899), .B(n12875), .Z(n12898) );
  XOR U15637 ( .A(n12889), .B(n12890), .Z(n12875) );
  XOR U15638 ( .A(n12900), .B(n12901), .Z(n12890) );
  ANDN U15639 ( .B(n12902), .A(n12903), .Z(n12900) );
  XOR U15640 ( .A(n12901), .B(n12904), .Z(n12902) );
  XOR U15641 ( .A(n12905), .B(n12906), .Z(n12889) );
  XOR U15642 ( .A(n12907), .B(n12908), .Z(n12906) );
  ANDN U15643 ( .B(n12909), .A(n12910), .Z(n12907) );
  XOR U15644 ( .A(n12911), .B(n12908), .Z(n12909) );
  IV U15645 ( .A(n12887), .Z(n12905) );
  XOR U15646 ( .A(n12912), .B(n12913), .Z(n12887) );
  ANDN U15647 ( .B(n12914), .A(n12915), .Z(n12912) );
  XOR U15648 ( .A(n12913), .B(n12916), .Z(n12914) );
  IV U15649 ( .A(n12895), .Z(n12899) );
  XOR U15650 ( .A(n12895), .B(n12877), .Z(n12897) );
  XOR U15651 ( .A(n12917), .B(n12918), .Z(n12877) );
  AND U15652 ( .A(n158), .B(n12919), .Z(n12917) );
  XOR U15653 ( .A(n12920), .B(n12918), .Z(n12919) );
  NANDN U15654 ( .A(n12879), .B(n12881), .Z(n12895) );
  XOR U15655 ( .A(n12921), .B(n12922), .Z(n12881) );
  AND U15656 ( .A(n158), .B(n12923), .Z(n12921) );
  XOR U15657 ( .A(n12922), .B(n12924), .Z(n12923) );
  XOR U15658 ( .A(n12925), .B(n12926), .Z(n158) );
  AND U15659 ( .A(n12927), .B(n12928), .Z(n12925) );
  XNOR U15660 ( .A(n12926), .B(n12892), .Z(n12928) );
  XNOR U15661 ( .A(n12929), .B(n12930), .Z(n12892) );
  ANDN U15662 ( .B(n12931), .A(n12932), .Z(n12929) );
  XOR U15663 ( .A(n12930), .B(n12933), .Z(n12931) );
  XOR U15664 ( .A(n12926), .B(n12894), .Z(n12927) );
  XOR U15665 ( .A(n12934), .B(n12935), .Z(n12894) );
  AND U15666 ( .A(n162), .B(n12936), .Z(n12934) );
  XOR U15667 ( .A(n12937), .B(n12935), .Z(n12936) );
  XNOR U15668 ( .A(n12938), .B(n12939), .Z(n12926) );
  NAND U15669 ( .A(n12940), .B(n12941), .Z(n12939) );
  XOR U15670 ( .A(n12942), .B(n12918), .Z(n12941) );
  XOR U15671 ( .A(n12932), .B(n12933), .Z(n12918) );
  XOR U15672 ( .A(n12943), .B(n12944), .Z(n12933) );
  ANDN U15673 ( .B(n12945), .A(n12946), .Z(n12943) );
  XOR U15674 ( .A(n12944), .B(n12947), .Z(n12945) );
  XOR U15675 ( .A(n12948), .B(n12949), .Z(n12932) );
  XOR U15676 ( .A(n12950), .B(n12951), .Z(n12949) );
  ANDN U15677 ( .B(n12952), .A(n12953), .Z(n12950) );
  XOR U15678 ( .A(n12954), .B(n12951), .Z(n12952) );
  IV U15679 ( .A(n12930), .Z(n12948) );
  XOR U15680 ( .A(n12955), .B(n12956), .Z(n12930) );
  ANDN U15681 ( .B(n12957), .A(n12958), .Z(n12955) );
  XOR U15682 ( .A(n12956), .B(n12959), .Z(n12957) );
  IV U15683 ( .A(n12938), .Z(n12942) );
  XOR U15684 ( .A(n12938), .B(n12920), .Z(n12940) );
  XOR U15685 ( .A(n12960), .B(n12961), .Z(n12920) );
  AND U15686 ( .A(n162), .B(n12962), .Z(n12960) );
  XOR U15687 ( .A(n12963), .B(n12961), .Z(n12962) );
  NANDN U15688 ( .A(n12922), .B(n12924), .Z(n12938) );
  XOR U15689 ( .A(n12964), .B(n12965), .Z(n12924) );
  AND U15690 ( .A(n162), .B(n12966), .Z(n12964) );
  XOR U15691 ( .A(n12965), .B(n12967), .Z(n12966) );
  XOR U15692 ( .A(n12968), .B(n12969), .Z(n162) );
  AND U15693 ( .A(n12970), .B(n12971), .Z(n12968) );
  XNOR U15694 ( .A(n12969), .B(n12935), .Z(n12971) );
  XNOR U15695 ( .A(n12972), .B(n12973), .Z(n12935) );
  ANDN U15696 ( .B(n12974), .A(n12975), .Z(n12972) );
  XOR U15697 ( .A(n12973), .B(n12976), .Z(n12974) );
  XOR U15698 ( .A(n12969), .B(n12937), .Z(n12970) );
  XOR U15699 ( .A(n12977), .B(n12978), .Z(n12937) );
  AND U15700 ( .A(n166), .B(n12979), .Z(n12977) );
  XOR U15701 ( .A(n12980), .B(n12978), .Z(n12979) );
  XNOR U15702 ( .A(n12981), .B(n12982), .Z(n12969) );
  NAND U15703 ( .A(n12983), .B(n12984), .Z(n12982) );
  XOR U15704 ( .A(n12985), .B(n12961), .Z(n12984) );
  XOR U15705 ( .A(n12975), .B(n12976), .Z(n12961) );
  XOR U15706 ( .A(n12986), .B(n12987), .Z(n12976) );
  ANDN U15707 ( .B(n12988), .A(n12989), .Z(n12986) );
  XOR U15708 ( .A(n12987), .B(n12990), .Z(n12988) );
  XOR U15709 ( .A(n12991), .B(n12992), .Z(n12975) );
  XOR U15710 ( .A(n12993), .B(n12994), .Z(n12992) );
  ANDN U15711 ( .B(n12995), .A(n12996), .Z(n12993) );
  XOR U15712 ( .A(n12997), .B(n12994), .Z(n12995) );
  IV U15713 ( .A(n12973), .Z(n12991) );
  XOR U15714 ( .A(n12998), .B(n12999), .Z(n12973) );
  ANDN U15715 ( .B(n13000), .A(n13001), .Z(n12998) );
  XOR U15716 ( .A(n12999), .B(n13002), .Z(n13000) );
  IV U15717 ( .A(n12981), .Z(n12985) );
  XOR U15718 ( .A(n12981), .B(n12963), .Z(n12983) );
  XOR U15719 ( .A(n13003), .B(n13004), .Z(n12963) );
  AND U15720 ( .A(n166), .B(n13005), .Z(n13003) );
  XOR U15721 ( .A(n13006), .B(n13004), .Z(n13005) );
  NANDN U15722 ( .A(n12965), .B(n12967), .Z(n12981) );
  XOR U15723 ( .A(n13007), .B(n13008), .Z(n12967) );
  AND U15724 ( .A(n166), .B(n13009), .Z(n13007) );
  XOR U15725 ( .A(n13008), .B(n13010), .Z(n13009) );
  XOR U15726 ( .A(n13011), .B(n13012), .Z(n166) );
  AND U15727 ( .A(n13013), .B(n13014), .Z(n13011) );
  XNOR U15728 ( .A(n13012), .B(n12978), .Z(n13014) );
  XNOR U15729 ( .A(n13015), .B(n13016), .Z(n12978) );
  ANDN U15730 ( .B(n13017), .A(n13018), .Z(n13015) );
  XOR U15731 ( .A(n13016), .B(n13019), .Z(n13017) );
  XOR U15732 ( .A(n13012), .B(n12980), .Z(n13013) );
  XOR U15733 ( .A(n13020), .B(n13021), .Z(n12980) );
  AND U15734 ( .A(n170), .B(n13022), .Z(n13020) );
  XOR U15735 ( .A(n13023), .B(n13021), .Z(n13022) );
  XNOR U15736 ( .A(n13024), .B(n13025), .Z(n13012) );
  NAND U15737 ( .A(n13026), .B(n13027), .Z(n13025) );
  XOR U15738 ( .A(n13028), .B(n13004), .Z(n13027) );
  XOR U15739 ( .A(n13018), .B(n13019), .Z(n13004) );
  XOR U15740 ( .A(n13029), .B(n13030), .Z(n13019) );
  ANDN U15741 ( .B(n13031), .A(n13032), .Z(n13029) );
  XOR U15742 ( .A(n13030), .B(n13033), .Z(n13031) );
  XOR U15743 ( .A(n13034), .B(n13035), .Z(n13018) );
  XOR U15744 ( .A(n13036), .B(n13037), .Z(n13035) );
  ANDN U15745 ( .B(n13038), .A(n13039), .Z(n13036) );
  XOR U15746 ( .A(n13040), .B(n13037), .Z(n13038) );
  IV U15747 ( .A(n13016), .Z(n13034) );
  XOR U15748 ( .A(n13041), .B(n13042), .Z(n13016) );
  ANDN U15749 ( .B(n13043), .A(n13044), .Z(n13041) );
  XOR U15750 ( .A(n13042), .B(n13045), .Z(n13043) );
  IV U15751 ( .A(n13024), .Z(n13028) );
  XOR U15752 ( .A(n13024), .B(n13006), .Z(n13026) );
  XOR U15753 ( .A(n13046), .B(n13047), .Z(n13006) );
  AND U15754 ( .A(n170), .B(n13048), .Z(n13046) );
  XOR U15755 ( .A(n13049), .B(n13047), .Z(n13048) );
  NANDN U15756 ( .A(n13008), .B(n13010), .Z(n13024) );
  XOR U15757 ( .A(n13050), .B(n13051), .Z(n13010) );
  AND U15758 ( .A(n170), .B(n13052), .Z(n13050) );
  XOR U15759 ( .A(n13051), .B(n13053), .Z(n13052) );
  XOR U15760 ( .A(n13054), .B(n13055), .Z(n170) );
  AND U15761 ( .A(n13056), .B(n13057), .Z(n13054) );
  XNOR U15762 ( .A(n13055), .B(n13021), .Z(n13057) );
  XNOR U15763 ( .A(n13058), .B(n13059), .Z(n13021) );
  ANDN U15764 ( .B(n13060), .A(n13061), .Z(n13058) );
  XOR U15765 ( .A(n13059), .B(n13062), .Z(n13060) );
  XOR U15766 ( .A(n13055), .B(n13023), .Z(n13056) );
  XOR U15767 ( .A(n13063), .B(n13064), .Z(n13023) );
  AND U15768 ( .A(n174), .B(n13065), .Z(n13063) );
  XOR U15769 ( .A(n13066), .B(n13064), .Z(n13065) );
  XNOR U15770 ( .A(n13067), .B(n13068), .Z(n13055) );
  NAND U15771 ( .A(n13069), .B(n13070), .Z(n13068) );
  XOR U15772 ( .A(n13071), .B(n13047), .Z(n13070) );
  XOR U15773 ( .A(n13061), .B(n13062), .Z(n13047) );
  XOR U15774 ( .A(n13072), .B(n13073), .Z(n13062) );
  ANDN U15775 ( .B(n13074), .A(n13075), .Z(n13072) );
  XOR U15776 ( .A(n13073), .B(n13076), .Z(n13074) );
  XOR U15777 ( .A(n13077), .B(n13078), .Z(n13061) );
  XOR U15778 ( .A(n13079), .B(n13080), .Z(n13078) );
  ANDN U15779 ( .B(n13081), .A(n13082), .Z(n13079) );
  XOR U15780 ( .A(n13083), .B(n13080), .Z(n13081) );
  IV U15781 ( .A(n13059), .Z(n13077) );
  XOR U15782 ( .A(n13084), .B(n13085), .Z(n13059) );
  ANDN U15783 ( .B(n13086), .A(n13087), .Z(n13084) );
  XOR U15784 ( .A(n13085), .B(n13088), .Z(n13086) );
  IV U15785 ( .A(n13067), .Z(n13071) );
  XOR U15786 ( .A(n13067), .B(n13049), .Z(n13069) );
  XOR U15787 ( .A(n13089), .B(n13090), .Z(n13049) );
  AND U15788 ( .A(n174), .B(n13091), .Z(n13089) );
  XOR U15789 ( .A(n13092), .B(n13090), .Z(n13091) );
  NANDN U15790 ( .A(n13051), .B(n13053), .Z(n13067) );
  XOR U15791 ( .A(n13093), .B(n13094), .Z(n13053) );
  AND U15792 ( .A(n174), .B(n13095), .Z(n13093) );
  XOR U15793 ( .A(n13094), .B(n13096), .Z(n13095) );
  XOR U15794 ( .A(n13097), .B(n13098), .Z(n174) );
  AND U15795 ( .A(n13099), .B(n13100), .Z(n13097) );
  XNOR U15796 ( .A(n13098), .B(n13064), .Z(n13100) );
  XNOR U15797 ( .A(n13101), .B(n13102), .Z(n13064) );
  ANDN U15798 ( .B(n13103), .A(n13104), .Z(n13101) );
  XOR U15799 ( .A(n13102), .B(n13105), .Z(n13103) );
  XOR U15800 ( .A(n13098), .B(n13066), .Z(n13099) );
  XOR U15801 ( .A(n13106), .B(n13107), .Z(n13066) );
  AND U15802 ( .A(n178), .B(n13108), .Z(n13106) );
  XOR U15803 ( .A(n13109), .B(n13107), .Z(n13108) );
  XNOR U15804 ( .A(n13110), .B(n13111), .Z(n13098) );
  NAND U15805 ( .A(n13112), .B(n13113), .Z(n13111) );
  XOR U15806 ( .A(n13114), .B(n13090), .Z(n13113) );
  XOR U15807 ( .A(n13104), .B(n13105), .Z(n13090) );
  XOR U15808 ( .A(n13115), .B(n13116), .Z(n13105) );
  ANDN U15809 ( .B(n13117), .A(n13118), .Z(n13115) );
  XOR U15810 ( .A(n13116), .B(n13119), .Z(n13117) );
  XOR U15811 ( .A(n13120), .B(n13121), .Z(n13104) );
  XOR U15812 ( .A(n13122), .B(n13123), .Z(n13121) );
  ANDN U15813 ( .B(n13124), .A(n13125), .Z(n13122) );
  XOR U15814 ( .A(n13126), .B(n13123), .Z(n13124) );
  IV U15815 ( .A(n13102), .Z(n13120) );
  XOR U15816 ( .A(n13127), .B(n13128), .Z(n13102) );
  ANDN U15817 ( .B(n13129), .A(n13130), .Z(n13127) );
  XOR U15818 ( .A(n13128), .B(n13131), .Z(n13129) );
  IV U15819 ( .A(n13110), .Z(n13114) );
  XOR U15820 ( .A(n13110), .B(n13092), .Z(n13112) );
  XOR U15821 ( .A(n13132), .B(n13133), .Z(n13092) );
  AND U15822 ( .A(n178), .B(n13134), .Z(n13132) );
  XOR U15823 ( .A(n13135), .B(n13133), .Z(n13134) );
  NANDN U15824 ( .A(n13094), .B(n13096), .Z(n13110) );
  XOR U15825 ( .A(n13136), .B(n13137), .Z(n13096) );
  AND U15826 ( .A(n178), .B(n13138), .Z(n13136) );
  XOR U15827 ( .A(n13137), .B(n13139), .Z(n13138) );
  XOR U15828 ( .A(n13140), .B(n13141), .Z(n178) );
  AND U15829 ( .A(n13142), .B(n13143), .Z(n13140) );
  XNOR U15830 ( .A(n13141), .B(n13107), .Z(n13143) );
  XNOR U15831 ( .A(n13144), .B(n13145), .Z(n13107) );
  ANDN U15832 ( .B(n13146), .A(n13147), .Z(n13144) );
  XOR U15833 ( .A(n13145), .B(n13148), .Z(n13146) );
  XOR U15834 ( .A(n13141), .B(n13109), .Z(n13142) );
  XOR U15835 ( .A(n13149), .B(n13150), .Z(n13109) );
  AND U15836 ( .A(n182), .B(n13151), .Z(n13149) );
  XOR U15837 ( .A(n13152), .B(n13150), .Z(n13151) );
  XNOR U15838 ( .A(n13153), .B(n13154), .Z(n13141) );
  NAND U15839 ( .A(n13155), .B(n13156), .Z(n13154) );
  XOR U15840 ( .A(n13157), .B(n13133), .Z(n13156) );
  XOR U15841 ( .A(n13147), .B(n13148), .Z(n13133) );
  XOR U15842 ( .A(n13158), .B(n13159), .Z(n13148) );
  ANDN U15843 ( .B(n13160), .A(n13161), .Z(n13158) );
  XOR U15844 ( .A(n13159), .B(n13162), .Z(n13160) );
  XOR U15845 ( .A(n13163), .B(n13164), .Z(n13147) );
  XOR U15846 ( .A(n13165), .B(n13166), .Z(n13164) );
  ANDN U15847 ( .B(n13167), .A(n13168), .Z(n13165) );
  XOR U15848 ( .A(n13169), .B(n13166), .Z(n13167) );
  IV U15849 ( .A(n13145), .Z(n13163) );
  XOR U15850 ( .A(n13170), .B(n13171), .Z(n13145) );
  ANDN U15851 ( .B(n13172), .A(n13173), .Z(n13170) );
  XOR U15852 ( .A(n13171), .B(n13174), .Z(n13172) );
  IV U15853 ( .A(n13153), .Z(n13157) );
  XOR U15854 ( .A(n13153), .B(n13135), .Z(n13155) );
  XOR U15855 ( .A(n13175), .B(n13176), .Z(n13135) );
  AND U15856 ( .A(n182), .B(n13177), .Z(n13175) );
  XOR U15857 ( .A(n13178), .B(n13176), .Z(n13177) );
  NANDN U15858 ( .A(n13137), .B(n13139), .Z(n13153) );
  XOR U15859 ( .A(n13179), .B(n13180), .Z(n13139) );
  AND U15860 ( .A(n182), .B(n13181), .Z(n13179) );
  XOR U15861 ( .A(n13180), .B(n13182), .Z(n13181) );
  XOR U15862 ( .A(n13183), .B(n13184), .Z(n182) );
  AND U15863 ( .A(n13185), .B(n13186), .Z(n13183) );
  XNOR U15864 ( .A(n13184), .B(n13150), .Z(n13186) );
  XNOR U15865 ( .A(n13187), .B(n13188), .Z(n13150) );
  ANDN U15866 ( .B(n13189), .A(n13190), .Z(n13187) );
  XOR U15867 ( .A(n13188), .B(n13191), .Z(n13189) );
  XOR U15868 ( .A(n13184), .B(n13152), .Z(n13185) );
  XOR U15869 ( .A(n13192), .B(n13193), .Z(n13152) );
  AND U15870 ( .A(n186), .B(n13194), .Z(n13192) );
  XOR U15871 ( .A(n13195), .B(n13193), .Z(n13194) );
  XNOR U15872 ( .A(n13196), .B(n13197), .Z(n13184) );
  NAND U15873 ( .A(n13198), .B(n13199), .Z(n13197) );
  XOR U15874 ( .A(n13200), .B(n13176), .Z(n13199) );
  XOR U15875 ( .A(n13190), .B(n13191), .Z(n13176) );
  XOR U15876 ( .A(n13201), .B(n13202), .Z(n13191) );
  ANDN U15877 ( .B(n13203), .A(n13204), .Z(n13201) );
  XOR U15878 ( .A(n13202), .B(n13205), .Z(n13203) );
  XOR U15879 ( .A(n13206), .B(n13207), .Z(n13190) );
  XOR U15880 ( .A(n13208), .B(n13209), .Z(n13207) );
  ANDN U15881 ( .B(n13210), .A(n13211), .Z(n13208) );
  XOR U15882 ( .A(n13212), .B(n13209), .Z(n13210) );
  IV U15883 ( .A(n13188), .Z(n13206) );
  XOR U15884 ( .A(n13213), .B(n13214), .Z(n13188) );
  ANDN U15885 ( .B(n13215), .A(n13216), .Z(n13213) );
  XOR U15886 ( .A(n13214), .B(n13217), .Z(n13215) );
  IV U15887 ( .A(n13196), .Z(n13200) );
  XOR U15888 ( .A(n13196), .B(n13178), .Z(n13198) );
  XOR U15889 ( .A(n13218), .B(n13219), .Z(n13178) );
  AND U15890 ( .A(n186), .B(n13220), .Z(n13218) );
  XOR U15891 ( .A(n13221), .B(n13219), .Z(n13220) );
  NANDN U15892 ( .A(n13180), .B(n13182), .Z(n13196) );
  XOR U15893 ( .A(n13222), .B(n13223), .Z(n13182) );
  AND U15894 ( .A(n186), .B(n13224), .Z(n13222) );
  XOR U15895 ( .A(n13223), .B(n13225), .Z(n13224) );
  XOR U15896 ( .A(n13226), .B(n13227), .Z(n186) );
  AND U15897 ( .A(n13228), .B(n13229), .Z(n13226) );
  XNOR U15898 ( .A(n13227), .B(n13193), .Z(n13229) );
  XNOR U15899 ( .A(n13230), .B(n13231), .Z(n13193) );
  ANDN U15900 ( .B(n13232), .A(n13233), .Z(n13230) );
  XOR U15901 ( .A(n13231), .B(n13234), .Z(n13232) );
  XOR U15902 ( .A(n13227), .B(n13195), .Z(n13228) );
  XOR U15903 ( .A(n13235), .B(n13236), .Z(n13195) );
  AND U15904 ( .A(n190), .B(n13237), .Z(n13235) );
  XOR U15905 ( .A(n13238), .B(n13236), .Z(n13237) );
  XNOR U15906 ( .A(n13239), .B(n13240), .Z(n13227) );
  NAND U15907 ( .A(n13241), .B(n13242), .Z(n13240) );
  XOR U15908 ( .A(n13243), .B(n13219), .Z(n13242) );
  XOR U15909 ( .A(n13233), .B(n13234), .Z(n13219) );
  XOR U15910 ( .A(n13244), .B(n13245), .Z(n13234) );
  ANDN U15911 ( .B(n13246), .A(n13247), .Z(n13244) );
  XOR U15912 ( .A(n13245), .B(n13248), .Z(n13246) );
  XOR U15913 ( .A(n13249), .B(n13250), .Z(n13233) );
  XOR U15914 ( .A(n13251), .B(n13252), .Z(n13250) );
  ANDN U15915 ( .B(n13253), .A(n13254), .Z(n13251) );
  XOR U15916 ( .A(n13255), .B(n13252), .Z(n13253) );
  IV U15917 ( .A(n13231), .Z(n13249) );
  XOR U15918 ( .A(n13256), .B(n13257), .Z(n13231) );
  ANDN U15919 ( .B(n13258), .A(n13259), .Z(n13256) );
  XOR U15920 ( .A(n13257), .B(n13260), .Z(n13258) );
  IV U15921 ( .A(n13239), .Z(n13243) );
  XOR U15922 ( .A(n13239), .B(n13221), .Z(n13241) );
  XOR U15923 ( .A(n13261), .B(n13262), .Z(n13221) );
  AND U15924 ( .A(n190), .B(n13263), .Z(n13261) );
  XOR U15925 ( .A(n13264), .B(n13262), .Z(n13263) );
  NANDN U15926 ( .A(n13223), .B(n13225), .Z(n13239) );
  XOR U15927 ( .A(n13265), .B(n13266), .Z(n13225) );
  AND U15928 ( .A(n190), .B(n13267), .Z(n13265) );
  XOR U15929 ( .A(n13266), .B(n13268), .Z(n13267) );
  XOR U15930 ( .A(n13269), .B(n13270), .Z(n190) );
  AND U15931 ( .A(n13271), .B(n13272), .Z(n13269) );
  XNOR U15932 ( .A(n13270), .B(n13236), .Z(n13272) );
  XNOR U15933 ( .A(n13273), .B(n13274), .Z(n13236) );
  ANDN U15934 ( .B(n13275), .A(n13276), .Z(n13273) );
  XOR U15935 ( .A(n13274), .B(n13277), .Z(n13275) );
  XOR U15936 ( .A(n13270), .B(n13238), .Z(n13271) );
  XOR U15937 ( .A(n13278), .B(n13279), .Z(n13238) );
  AND U15938 ( .A(n194), .B(n13280), .Z(n13278) );
  XOR U15939 ( .A(n13281), .B(n13279), .Z(n13280) );
  XNOR U15940 ( .A(n13282), .B(n13283), .Z(n13270) );
  NAND U15941 ( .A(n13284), .B(n13285), .Z(n13283) );
  XOR U15942 ( .A(n13286), .B(n13262), .Z(n13285) );
  XOR U15943 ( .A(n13276), .B(n13277), .Z(n13262) );
  XOR U15944 ( .A(n13287), .B(n13288), .Z(n13277) );
  ANDN U15945 ( .B(n13289), .A(n13290), .Z(n13287) );
  XOR U15946 ( .A(n13288), .B(n13291), .Z(n13289) );
  XOR U15947 ( .A(n13292), .B(n13293), .Z(n13276) );
  XOR U15948 ( .A(n13294), .B(n13295), .Z(n13293) );
  ANDN U15949 ( .B(n13296), .A(n13297), .Z(n13294) );
  XOR U15950 ( .A(n13298), .B(n13295), .Z(n13296) );
  IV U15951 ( .A(n13274), .Z(n13292) );
  XOR U15952 ( .A(n13299), .B(n13300), .Z(n13274) );
  ANDN U15953 ( .B(n13301), .A(n13302), .Z(n13299) );
  XOR U15954 ( .A(n13300), .B(n13303), .Z(n13301) );
  IV U15955 ( .A(n13282), .Z(n13286) );
  XOR U15956 ( .A(n13282), .B(n13264), .Z(n13284) );
  XOR U15957 ( .A(n13304), .B(n13305), .Z(n13264) );
  AND U15958 ( .A(n194), .B(n13306), .Z(n13304) );
  XOR U15959 ( .A(n13307), .B(n13305), .Z(n13306) );
  NANDN U15960 ( .A(n13266), .B(n13268), .Z(n13282) );
  XOR U15961 ( .A(n13308), .B(n13309), .Z(n13268) );
  AND U15962 ( .A(n194), .B(n13310), .Z(n13308) );
  XOR U15963 ( .A(n13309), .B(n13311), .Z(n13310) );
  XOR U15964 ( .A(n13312), .B(n13313), .Z(n194) );
  AND U15965 ( .A(n13314), .B(n13315), .Z(n13312) );
  XNOR U15966 ( .A(n13313), .B(n13279), .Z(n13315) );
  XNOR U15967 ( .A(n13316), .B(n13317), .Z(n13279) );
  ANDN U15968 ( .B(n13318), .A(n13319), .Z(n13316) );
  XOR U15969 ( .A(n13317), .B(n13320), .Z(n13318) );
  XOR U15970 ( .A(n13313), .B(n13281), .Z(n13314) );
  XOR U15971 ( .A(n13321), .B(n13322), .Z(n13281) );
  AND U15972 ( .A(n198), .B(n13323), .Z(n13321) );
  XOR U15973 ( .A(n13324), .B(n13322), .Z(n13323) );
  XNOR U15974 ( .A(n13325), .B(n13326), .Z(n13313) );
  NAND U15975 ( .A(n13327), .B(n13328), .Z(n13326) );
  XOR U15976 ( .A(n13329), .B(n13305), .Z(n13328) );
  XOR U15977 ( .A(n13319), .B(n13320), .Z(n13305) );
  XOR U15978 ( .A(n13330), .B(n13331), .Z(n13320) );
  ANDN U15979 ( .B(n13332), .A(n13333), .Z(n13330) );
  XOR U15980 ( .A(n13331), .B(n13334), .Z(n13332) );
  XOR U15981 ( .A(n13335), .B(n13336), .Z(n13319) );
  XOR U15982 ( .A(n13337), .B(n13338), .Z(n13336) );
  ANDN U15983 ( .B(n13339), .A(n13340), .Z(n13337) );
  XOR U15984 ( .A(n13341), .B(n13338), .Z(n13339) );
  IV U15985 ( .A(n13317), .Z(n13335) );
  XOR U15986 ( .A(n13342), .B(n13343), .Z(n13317) );
  ANDN U15987 ( .B(n13344), .A(n13345), .Z(n13342) );
  XOR U15988 ( .A(n13343), .B(n13346), .Z(n13344) );
  IV U15989 ( .A(n13325), .Z(n13329) );
  XOR U15990 ( .A(n13325), .B(n13307), .Z(n13327) );
  XOR U15991 ( .A(n13347), .B(n13348), .Z(n13307) );
  AND U15992 ( .A(n198), .B(n13349), .Z(n13347) );
  XOR U15993 ( .A(n13350), .B(n13348), .Z(n13349) );
  NANDN U15994 ( .A(n13309), .B(n13311), .Z(n13325) );
  XOR U15995 ( .A(n13351), .B(n13352), .Z(n13311) );
  AND U15996 ( .A(n198), .B(n13353), .Z(n13351) );
  XOR U15997 ( .A(n13352), .B(n13354), .Z(n13353) );
  XOR U15998 ( .A(n13355), .B(n13356), .Z(n198) );
  AND U15999 ( .A(n13357), .B(n13358), .Z(n13355) );
  XNOR U16000 ( .A(n13356), .B(n13322), .Z(n13358) );
  XNOR U16001 ( .A(n13359), .B(n13360), .Z(n13322) );
  ANDN U16002 ( .B(n13361), .A(n13362), .Z(n13359) );
  XOR U16003 ( .A(n13360), .B(n13363), .Z(n13361) );
  XOR U16004 ( .A(n13356), .B(n13324), .Z(n13357) );
  XOR U16005 ( .A(n13364), .B(n13365), .Z(n13324) );
  AND U16006 ( .A(n202), .B(n13366), .Z(n13364) );
  XOR U16007 ( .A(n13367), .B(n13365), .Z(n13366) );
  XNOR U16008 ( .A(n13368), .B(n13369), .Z(n13356) );
  NAND U16009 ( .A(n13370), .B(n13371), .Z(n13369) );
  XOR U16010 ( .A(n13372), .B(n13348), .Z(n13371) );
  XOR U16011 ( .A(n13362), .B(n13363), .Z(n13348) );
  XOR U16012 ( .A(n13373), .B(n13374), .Z(n13363) );
  ANDN U16013 ( .B(n13375), .A(n13376), .Z(n13373) );
  XOR U16014 ( .A(n13374), .B(n13377), .Z(n13375) );
  XOR U16015 ( .A(n13378), .B(n13379), .Z(n13362) );
  XOR U16016 ( .A(n13380), .B(n13381), .Z(n13379) );
  ANDN U16017 ( .B(n13382), .A(n13383), .Z(n13380) );
  XOR U16018 ( .A(n13384), .B(n13381), .Z(n13382) );
  IV U16019 ( .A(n13360), .Z(n13378) );
  XOR U16020 ( .A(n13385), .B(n13386), .Z(n13360) );
  ANDN U16021 ( .B(n13387), .A(n13388), .Z(n13385) );
  XOR U16022 ( .A(n13386), .B(n13389), .Z(n13387) );
  IV U16023 ( .A(n13368), .Z(n13372) );
  XOR U16024 ( .A(n13368), .B(n13350), .Z(n13370) );
  XOR U16025 ( .A(n13390), .B(n13391), .Z(n13350) );
  AND U16026 ( .A(n202), .B(n13392), .Z(n13390) );
  XOR U16027 ( .A(n13393), .B(n13391), .Z(n13392) );
  NANDN U16028 ( .A(n13352), .B(n13354), .Z(n13368) );
  XOR U16029 ( .A(n13394), .B(n13395), .Z(n13354) );
  AND U16030 ( .A(n202), .B(n13396), .Z(n13394) );
  XOR U16031 ( .A(n13395), .B(n13397), .Z(n13396) );
  XOR U16032 ( .A(n13398), .B(n13399), .Z(n202) );
  AND U16033 ( .A(n13400), .B(n13401), .Z(n13398) );
  XNOR U16034 ( .A(n13399), .B(n13365), .Z(n13401) );
  XNOR U16035 ( .A(n13402), .B(n13403), .Z(n13365) );
  ANDN U16036 ( .B(n13404), .A(n13405), .Z(n13402) );
  XOR U16037 ( .A(n13403), .B(n13406), .Z(n13404) );
  XOR U16038 ( .A(n13399), .B(n13367), .Z(n13400) );
  XOR U16039 ( .A(n13407), .B(n13408), .Z(n13367) );
  AND U16040 ( .A(n206), .B(n13409), .Z(n13407) );
  XOR U16041 ( .A(n13410), .B(n13408), .Z(n13409) );
  XNOR U16042 ( .A(n13411), .B(n13412), .Z(n13399) );
  NAND U16043 ( .A(n13413), .B(n13414), .Z(n13412) );
  XOR U16044 ( .A(n13415), .B(n13391), .Z(n13414) );
  XOR U16045 ( .A(n13405), .B(n13406), .Z(n13391) );
  XOR U16046 ( .A(n13416), .B(n13417), .Z(n13406) );
  ANDN U16047 ( .B(n13418), .A(n13419), .Z(n13416) );
  XOR U16048 ( .A(n13417), .B(n13420), .Z(n13418) );
  XOR U16049 ( .A(n13421), .B(n13422), .Z(n13405) );
  XOR U16050 ( .A(n13423), .B(n13424), .Z(n13422) );
  ANDN U16051 ( .B(n13425), .A(n13426), .Z(n13423) );
  XOR U16052 ( .A(n13427), .B(n13424), .Z(n13425) );
  IV U16053 ( .A(n13403), .Z(n13421) );
  XOR U16054 ( .A(n13428), .B(n13429), .Z(n13403) );
  ANDN U16055 ( .B(n13430), .A(n13431), .Z(n13428) );
  XOR U16056 ( .A(n13429), .B(n13432), .Z(n13430) );
  IV U16057 ( .A(n13411), .Z(n13415) );
  XOR U16058 ( .A(n13411), .B(n13393), .Z(n13413) );
  XOR U16059 ( .A(n13433), .B(n13434), .Z(n13393) );
  AND U16060 ( .A(n206), .B(n13435), .Z(n13433) );
  XOR U16061 ( .A(n13436), .B(n13434), .Z(n13435) );
  NANDN U16062 ( .A(n13395), .B(n13397), .Z(n13411) );
  XOR U16063 ( .A(n13437), .B(n13438), .Z(n13397) );
  AND U16064 ( .A(n206), .B(n13439), .Z(n13437) );
  XOR U16065 ( .A(n13438), .B(n13440), .Z(n13439) );
  XOR U16066 ( .A(n13441), .B(n13442), .Z(n206) );
  AND U16067 ( .A(n13443), .B(n13444), .Z(n13441) );
  XNOR U16068 ( .A(n13442), .B(n13408), .Z(n13444) );
  XNOR U16069 ( .A(n13445), .B(n13446), .Z(n13408) );
  ANDN U16070 ( .B(n13447), .A(n13448), .Z(n13445) );
  XOR U16071 ( .A(n13446), .B(n13449), .Z(n13447) );
  XOR U16072 ( .A(n13442), .B(n13410), .Z(n13443) );
  XOR U16073 ( .A(n13450), .B(n13451), .Z(n13410) );
  AND U16074 ( .A(n210), .B(n13452), .Z(n13450) );
  XOR U16075 ( .A(n13453), .B(n13451), .Z(n13452) );
  XNOR U16076 ( .A(n13454), .B(n13455), .Z(n13442) );
  NAND U16077 ( .A(n13456), .B(n13457), .Z(n13455) );
  XOR U16078 ( .A(n13458), .B(n13434), .Z(n13457) );
  XOR U16079 ( .A(n13448), .B(n13449), .Z(n13434) );
  XOR U16080 ( .A(n13459), .B(n13460), .Z(n13449) );
  ANDN U16081 ( .B(n13461), .A(n13462), .Z(n13459) );
  XOR U16082 ( .A(n13460), .B(n13463), .Z(n13461) );
  XOR U16083 ( .A(n13464), .B(n13465), .Z(n13448) );
  XOR U16084 ( .A(n13466), .B(n13467), .Z(n13465) );
  ANDN U16085 ( .B(n13468), .A(n13469), .Z(n13466) );
  XOR U16086 ( .A(n13470), .B(n13467), .Z(n13468) );
  IV U16087 ( .A(n13446), .Z(n13464) );
  XOR U16088 ( .A(n13471), .B(n13472), .Z(n13446) );
  ANDN U16089 ( .B(n13473), .A(n13474), .Z(n13471) );
  XOR U16090 ( .A(n13472), .B(n13475), .Z(n13473) );
  IV U16091 ( .A(n13454), .Z(n13458) );
  XOR U16092 ( .A(n13454), .B(n13436), .Z(n13456) );
  XOR U16093 ( .A(n13476), .B(n13477), .Z(n13436) );
  AND U16094 ( .A(n210), .B(n13478), .Z(n13476) );
  XOR U16095 ( .A(n13479), .B(n13477), .Z(n13478) );
  NANDN U16096 ( .A(n13438), .B(n13440), .Z(n13454) );
  XOR U16097 ( .A(n13480), .B(n13481), .Z(n13440) );
  AND U16098 ( .A(n210), .B(n13482), .Z(n13480) );
  XOR U16099 ( .A(n13481), .B(n13483), .Z(n13482) );
  XOR U16100 ( .A(n13484), .B(n13485), .Z(n210) );
  AND U16101 ( .A(n13486), .B(n13487), .Z(n13484) );
  XNOR U16102 ( .A(n13485), .B(n13451), .Z(n13487) );
  XNOR U16103 ( .A(n13488), .B(n13489), .Z(n13451) );
  ANDN U16104 ( .B(n13490), .A(n13491), .Z(n13488) );
  XOR U16105 ( .A(n13489), .B(n13492), .Z(n13490) );
  XOR U16106 ( .A(n13485), .B(n13453), .Z(n13486) );
  XOR U16107 ( .A(n13493), .B(n13494), .Z(n13453) );
  AND U16108 ( .A(n214), .B(n13495), .Z(n13493) );
  XOR U16109 ( .A(n13496), .B(n13494), .Z(n13495) );
  XNOR U16110 ( .A(n13497), .B(n13498), .Z(n13485) );
  NAND U16111 ( .A(n13499), .B(n13500), .Z(n13498) );
  XOR U16112 ( .A(n13501), .B(n13477), .Z(n13500) );
  XOR U16113 ( .A(n13491), .B(n13492), .Z(n13477) );
  XOR U16114 ( .A(n13502), .B(n13503), .Z(n13492) );
  ANDN U16115 ( .B(n13504), .A(n13505), .Z(n13502) );
  XOR U16116 ( .A(n13503), .B(n13506), .Z(n13504) );
  XOR U16117 ( .A(n13507), .B(n13508), .Z(n13491) );
  XOR U16118 ( .A(n13509), .B(n13510), .Z(n13508) );
  ANDN U16119 ( .B(n13511), .A(n13512), .Z(n13509) );
  XOR U16120 ( .A(n13513), .B(n13510), .Z(n13511) );
  IV U16121 ( .A(n13489), .Z(n13507) );
  XOR U16122 ( .A(n13514), .B(n13515), .Z(n13489) );
  ANDN U16123 ( .B(n13516), .A(n13517), .Z(n13514) );
  XOR U16124 ( .A(n13515), .B(n13518), .Z(n13516) );
  IV U16125 ( .A(n13497), .Z(n13501) );
  XOR U16126 ( .A(n13497), .B(n13479), .Z(n13499) );
  XOR U16127 ( .A(n13519), .B(n13520), .Z(n13479) );
  AND U16128 ( .A(n214), .B(n13521), .Z(n13519) );
  XOR U16129 ( .A(n13522), .B(n13520), .Z(n13521) );
  NANDN U16130 ( .A(n13481), .B(n13483), .Z(n13497) );
  XOR U16131 ( .A(n13523), .B(n13524), .Z(n13483) );
  AND U16132 ( .A(n214), .B(n13525), .Z(n13523) );
  XOR U16133 ( .A(n13524), .B(n13526), .Z(n13525) );
  XOR U16134 ( .A(n13527), .B(n13528), .Z(n214) );
  AND U16135 ( .A(n13529), .B(n13530), .Z(n13527) );
  XNOR U16136 ( .A(n13528), .B(n13494), .Z(n13530) );
  XNOR U16137 ( .A(n13531), .B(n13532), .Z(n13494) );
  ANDN U16138 ( .B(n13533), .A(n13534), .Z(n13531) );
  XOR U16139 ( .A(n13532), .B(n13535), .Z(n13533) );
  XOR U16140 ( .A(n13528), .B(n13496), .Z(n13529) );
  XOR U16141 ( .A(n13536), .B(n13537), .Z(n13496) );
  AND U16142 ( .A(n218), .B(n13538), .Z(n13536) );
  XOR U16143 ( .A(n13539), .B(n13537), .Z(n13538) );
  XNOR U16144 ( .A(n13540), .B(n13541), .Z(n13528) );
  NAND U16145 ( .A(n13542), .B(n13543), .Z(n13541) );
  XOR U16146 ( .A(n13544), .B(n13520), .Z(n13543) );
  XOR U16147 ( .A(n13534), .B(n13535), .Z(n13520) );
  XOR U16148 ( .A(n13545), .B(n13546), .Z(n13535) );
  ANDN U16149 ( .B(n13547), .A(n13548), .Z(n13545) );
  XOR U16150 ( .A(n13546), .B(n13549), .Z(n13547) );
  XOR U16151 ( .A(n13550), .B(n13551), .Z(n13534) );
  XOR U16152 ( .A(n13552), .B(n13553), .Z(n13551) );
  ANDN U16153 ( .B(n13554), .A(n13555), .Z(n13552) );
  XOR U16154 ( .A(n13556), .B(n13553), .Z(n13554) );
  IV U16155 ( .A(n13532), .Z(n13550) );
  XOR U16156 ( .A(n13557), .B(n13558), .Z(n13532) );
  ANDN U16157 ( .B(n13559), .A(n13560), .Z(n13557) );
  XOR U16158 ( .A(n13558), .B(n13561), .Z(n13559) );
  IV U16159 ( .A(n13540), .Z(n13544) );
  XOR U16160 ( .A(n13540), .B(n13522), .Z(n13542) );
  XOR U16161 ( .A(n13562), .B(n13563), .Z(n13522) );
  AND U16162 ( .A(n218), .B(n13564), .Z(n13562) );
  XOR U16163 ( .A(n13565), .B(n13563), .Z(n13564) );
  NANDN U16164 ( .A(n13524), .B(n13526), .Z(n13540) );
  XOR U16165 ( .A(n13566), .B(n13567), .Z(n13526) );
  AND U16166 ( .A(n218), .B(n13568), .Z(n13566) );
  XOR U16167 ( .A(n13567), .B(n13569), .Z(n13568) );
  XOR U16168 ( .A(n13570), .B(n13571), .Z(n218) );
  AND U16169 ( .A(n13572), .B(n13573), .Z(n13570) );
  XNOR U16170 ( .A(n13571), .B(n13537), .Z(n13573) );
  XNOR U16171 ( .A(n13574), .B(n13575), .Z(n13537) );
  ANDN U16172 ( .B(n13576), .A(n13577), .Z(n13574) );
  XOR U16173 ( .A(n13575), .B(n13578), .Z(n13576) );
  XOR U16174 ( .A(n13571), .B(n13539), .Z(n13572) );
  XOR U16175 ( .A(n13579), .B(n13580), .Z(n13539) );
  AND U16176 ( .A(n222), .B(n13581), .Z(n13579) );
  XOR U16177 ( .A(n13582), .B(n13580), .Z(n13581) );
  XNOR U16178 ( .A(n13583), .B(n13584), .Z(n13571) );
  NAND U16179 ( .A(n13585), .B(n13586), .Z(n13584) );
  XOR U16180 ( .A(n13587), .B(n13563), .Z(n13586) );
  XOR U16181 ( .A(n13577), .B(n13578), .Z(n13563) );
  XOR U16182 ( .A(n13588), .B(n13589), .Z(n13578) );
  ANDN U16183 ( .B(n13590), .A(n13591), .Z(n13588) );
  XOR U16184 ( .A(n13589), .B(n13592), .Z(n13590) );
  XOR U16185 ( .A(n13593), .B(n13594), .Z(n13577) );
  XOR U16186 ( .A(n13595), .B(n13596), .Z(n13594) );
  ANDN U16187 ( .B(n13597), .A(n13598), .Z(n13595) );
  XOR U16188 ( .A(n13599), .B(n13596), .Z(n13597) );
  IV U16189 ( .A(n13575), .Z(n13593) );
  XOR U16190 ( .A(n13600), .B(n13601), .Z(n13575) );
  ANDN U16191 ( .B(n13602), .A(n13603), .Z(n13600) );
  XOR U16192 ( .A(n13601), .B(n13604), .Z(n13602) );
  IV U16193 ( .A(n13583), .Z(n13587) );
  XOR U16194 ( .A(n13583), .B(n13565), .Z(n13585) );
  XOR U16195 ( .A(n13605), .B(n13606), .Z(n13565) );
  AND U16196 ( .A(n222), .B(n13607), .Z(n13605) );
  XOR U16197 ( .A(n13608), .B(n13606), .Z(n13607) );
  NANDN U16198 ( .A(n13567), .B(n13569), .Z(n13583) );
  XOR U16199 ( .A(n13609), .B(n13610), .Z(n13569) );
  AND U16200 ( .A(n222), .B(n13611), .Z(n13609) );
  XOR U16201 ( .A(n13610), .B(n13612), .Z(n13611) );
  XOR U16202 ( .A(n13613), .B(n13614), .Z(n222) );
  AND U16203 ( .A(n13615), .B(n13616), .Z(n13613) );
  XNOR U16204 ( .A(n13614), .B(n13580), .Z(n13616) );
  XNOR U16205 ( .A(n13617), .B(n13618), .Z(n13580) );
  ANDN U16206 ( .B(n13619), .A(n13620), .Z(n13617) );
  XOR U16207 ( .A(n13618), .B(n13621), .Z(n13619) );
  XOR U16208 ( .A(n13614), .B(n13582), .Z(n13615) );
  XOR U16209 ( .A(n13622), .B(n13623), .Z(n13582) );
  AND U16210 ( .A(n226), .B(n13624), .Z(n13622) );
  XOR U16211 ( .A(n13625), .B(n13623), .Z(n13624) );
  XNOR U16212 ( .A(n13626), .B(n13627), .Z(n13614) );
  NAND U16213 ( .A(n13628), .B(n13629), .Z(n13627) );
  XOR U16214 ( .A(n13630), .B(n13606), .Z(n13629) );
  XOR U16215 ( .A(n13620), .B(n13621), .Z(n13606) );
  XOR U16216 ( .A(n13631), .B(n13632), .Z(n13621) );
  ANDN U16217 ( .B(n13633), .A(n13634), .Z(n13631) );
  XOR U16218 ( .A(n13632), .B(n13635), .Z(n13633) );
  XOR U16219 ( .A(n13636), .B(n13637), .Z(n13620) );
  XOR U16220 ( .A(n13638), .B(n13639), .Z(n13637) );
  ANDN U16221 ( .B(n13640), .A(n13641), .Z(n13638) );
  XOR U16222 ( .A(n13642), .B(n13639), .Z(n13640) );
  IV U16223 ( .A(n13618), .Z(n13636) );
  XOR U16224 ( .A(n13643), .B(n13644), .Z(n13618) );
  ANDN U16225 ( .B(n13645), .A(n13646), .Z(n13643) );
  XOR U16226 ( .A(n13644), .B(n13647), .Z(n13645) );
  IV U16227 ( .A(n13626), .Z(n13630) );
  XOR U16228 ( .A(n13626), .B(n13608), .Z(n13628) );
  XOR U16229 ( .A(n13648), .B(n13649), .Z(n13608) );
  AND U16230 ( .A(n226), .B(n13650), .Z(n13648) );
  XOR U16231 ( .A(n13651), .B(n13649), .Z(n13650) );
  NANDN U16232 ( .A(n13610), .B(n13612), .Z(n13626) );
  XOR U16233 ( .A(n13652), .B(n13653), .Z(n13612) );
  AND U16234 ( .A(n226), .B(n13654), .Z(n13652) );
  XOR U16235 ( .A(n13653), .B(n13655), .Z(n13654) );
  XOR U16236 ( .A(n13656), .B(n13657), .Z(n226) );
  AND U16237 ( .A(n13658), .B(n13659), .Z(n13656) );
  XNOR U16238 ( .A(n13657), .B(n13623), .Z(n13659) );
  XNOR U16239 ( .A(n13660), .B(n13661), .Z(n13623) );
  ANDN U16240 ( .B(n13662), .A(n13663), .Z(n13660) );
  XOR U16241 ( .A(n13661), .B(n13664), .Z(n13662) );
  XOR U16242 ( .A(n13657), .B(n13625), .Z(n13658) );
  XOR U16243 ( .A(n13665), .B(n13666), .Z(n13625) );
  AND U16244 ( .A(n230), .B(n13667), .Z(n13665) );
  XOR U16245 ( .A(n13668), .B(n13666), .Z(n13667) );
  XNOR U16246 ( .A(n13669), .B(n13670), .Z(n13657) );
  NAND U16247 ( .A(n13671), .B(n13672), .Z(n13670) );
  XOR U16248 ( .A(n13673), .B(n13649), .Z(n13672) );
  XOR U16249 ( .A(n13663), .B(n13664), .Z(n13649) );
  XOR U16250 ( .A(n13674), .B(n13675), .Z(n13664) );
  ANDN U16251 ( .B(n13676), .A(n13677), .Z(n13674) );
  XOR U16252 ( .A(n13675), .B(n13678), .Z(n13676) );
  XOR U16253 ( .A(n13679), .B(n13680), .Z(n13663) );
  XOR U16254 ( .A(n13681), .B(n13682), .Z(n13680) );
  ANDN U16255 ( .B(n13683), .A(n13684), .Z(n13681) );
  XOR U16256 ( .A(n13685), .B(n13682), .Z(n13683) );
  IV U16257 ( .A(n13661), .Z(n13679) );
  XOR U16258 ( .A(n13686), .B(n13687), .Z(n13661) );
  ANDN U16259 ( .B(n13688), .A(n13689), .Z(n13686) );
  XOR U16260 ( .A(n13687), .B(n13690), .Z(n13688) );
  IV U16261 ( .A(n13669), .Z(n13673) );
  XOR U16262 ( .A(n13669), .B(n13651), .Z(n13671) );
  XOR U16263 ( .A(n13691), .B(n13692), .Z(n13651) );
  AND U16264 ( .A(n230), .B(n13693), .Z(n13691) );
  XOR U16265 ( .A(n13694), .B(n13692), .Z(n13693) );
  NANDN U16266 ( .A(n13653), .B(n13655), .Z(n13669) );
  XOR U16267 ( .A(n13695), .B(n13696), .Z(n13655) );
  AND U16268 ( .A(n230), .B(n13697), .Z(n13695) );
  XOR U16269 ( .A(n13696), .B(n13698), .Z(n13697) );
  XOR U16270 ( .A(n13699), .B(n13700), .Z(n230) );
  AND U16271 ( .A(n13701), .B(n13702), .Z(n13699) );
  XNOR U16272 ( .A(n13700), .B(n13666), .Z(n13702) );
  XNOR U16273 ( .A(n13703), .B(n13704), .Z(n13666) );
  ANDN U16274 ( .B(n13705), .A(n13706), .Z(n13703) );
  XOR U16275 ( .A(n13704), .B(n13707), .Z(n13705) );
  XOR U16276 ( .A(n13700), .B(n13668), .Z(n13701) );
  XOR U16277 ( .A(n13708), .B(n13709), .Z(n13668) );
  AND U16278 ( .A(n234), .B(n13710), .Z(n13708) );
  XOR U16279 ( .A(n13711), .B(n13709), .Z(n13710) );
  XNOR U16280 ( .A(n13712), .B(n13713), .Z(n13700) );
  NAND U16281 ( .A(n13714), .B(n13715), .Z(n13713) );
  XOR U16282 ( .A(n13716), .B(n13692), .Z(n13715) );
  XOR U16283 ( .A(n13706), .B(n13707), .Z(n13692) );
  XOR U16284 ( .A(n13717), .B(n13718), .Z(n13707) );
  ANDN U16285 ( .B(n13719), .A(n13720), .Z(n13717) );
  XOR U16286 ( .A(n13718), .B(n13721), .Z(n13719) );
  XOR U16287 ( .A(n13722), .B(n13723), .Z(n13706) );
  XOR U16288 ( .A(n13724), .B(n13725), .Z(n13723) );
  ANDN U16289 ( .B(n13726), .A(n13727), .Z(n13724) );
  XOR U16290 ( .A(n13728), .B(n13725), .Z(n13726) );
  IV U16291 ( .A(n13704), .Z(n13722) );
  XOR U16292 ( .A(n13729), .B(n13730), .Z(n13704) );
  ANDN U16293 ( .B(n13731), .A(n13732), .Z(n13729) );
  XOR U16294 ( .A(n13730), .B(n13733), .Z(n13731) );
  IV U16295 ( .A(n13712), .Z(n13716) );
  XOR U16296 ( .A(n13712), .B(n13694), .Z(n13714) );
  XOR U16297 ( .A(n13734), .B(n13735), .Z(n13694) );
  AND U16298 ( .A(n234), .B(n13736), .Z(n13734) );
  XOR U16299 ( .A(n13737), .B(n13735), .Z(n13736) );
  NANDN U16300 ( .A(n13696), .B(n13698), .Z(n13712) );
  XOR U16301 ( .A(n13738), .B(n13739), .Z(n13698) );
  AND U16302 ( .A(n234), .B(n13740), .Z(n13738) );
  XOR U16303 ( .A(n13739), .B(n13741), .Z(n13740) );
  XOR U16304 ( .A(n13742), .B(n13743), .Z(n234) );
  AND U16305 ( .A(n13744), .B(n13745), .Z(n13742) );
  XNOR U16306 ( .A(n13743), .B(n13709), .Z(n13745) );
  XNOR U16307 ( .A(n13746), .B(n13747), .Z(n13709) );
  ANDN U16308 ( .B(n13748), .A(n13749), .Z(n13746) );
  XOR U16309 ( .A(n13747), .B(n13750), .Z(n13748) );
  XOR U16310 ( .A(n13743), .B(n13711), .Z(n13744) );
  XOR U16311 ( .A(n13751), .B(n13752), .Z(n13711) );
  AND U16312 ( .A(n238), .B(n13753), .Z(n13751) );
  XOR U16313 ( .A(n13754), .B(n13752), .Z(n13753) );
  XNOR U16314 ( .A(n13755), .B(n13756), .Z(n13743) );
  NAND U16315 ( .A(n13757), .B(n13758), .Z(n13756) );
  XOR U16316 ( .A(n13759), .B(n13735), .Z(n13758) );
  XOR U16317 ( .A(n13749), .B(n13750), .Z(n13735) );
  XOR U16318 ( .A(n13760), .B(n13761), .Z(n13750) );
  ANDN U16319 ( .B(n13762), .A(n13763), .Z(n13760) );
  XOR U16320 ( .A(n13761), .B(n13764), .Z(n13762) );
  XOR U16321 ( .A(n13765), .B(n13766), .Z(n13749) );
  XOR U16322 ( .A(n13767), .B(n13768), .Z(n13766) );
  ANDN U16323 ( .B(n13769), .A(n13770), .Z(n13767) );
  XOR U16324 ( .A(n13771), .B(n13768), .Z(n13769) );
  IV U16325 ( .A(n13747), .Z(n13765) );
  XOR U16326 ( .A(n13772), .B(n13773), .Z(n13747) );
  ANDN U16327 ( .B(n13774), .A(n13775), .Z(n13772) );
  XOR U16328 ( .A(n13773), .B(n13776), .Z(n13774) );
  IV U16329 ( .A(n13755), .Z(n13759) );
  XOR U16330 ( .A(n13755), .B(n13737), .Z(n13757) );
  XOR U16331 ( .A(n13777), .B(n13778), .Z(n13737) );
  AND U16332 ( .A(n238), .B(n13779), .Z(n13777) );
  XOR U16333 ( .A(n13780), .B(n13778), .Z(n13779) );
  NANDN U16334 ( .A(n13739), .B(n13741), .Z(n13755) );
  XOR U16335 ( .A(n13781), .B(n13782), .Z(n13741) );
  AND U16336 ( .A(n238), .B(n13783), .Z(n13781) );
  XOR U16337 ( .A(n13782), .B(n13784), .Z(n13783) );
  XOR U16338 ( .A(n13785), .B(n13786), .Z(n238) );
  AND U16339 ( .A(n13787), .B(n13788), .Z(n13785) );
  XNOR U16340 ( .A(n13786), .B(n13752), .Z(n13788) );
  XNOR U16341 ( .A(n13789), .B(n13790), .Z(n13752) );
  ANDN U16342 ( .B(n13791), .A(n13792), .Z(n13789) );
  XOR U16343 ( .A(n13790), .B(n13793), .Z(n13791) );
  XOR U16344 ( .A(n13786), .B(n13754), .Z(n13787) );
  XOR U16345 ( .A(n13794), .B(n13795), .Z(n13754) );
  AND U16346 ( .A(n242), .B(n13796), .Z(n13794) );
  XOR U16347 ( .A(n13797), .B(n13795), .Z(n13796) );
  XNOR U16348 ( .A(n13798), .B(n13799), .Z(n13786) );
  NAND U16349 ( .A(n13800), .B(n13801), .Z(n13799) );
  XOR U16350 ( .A(n13802), .B(n13778), .Z(n13801) );
  XOR U16351 ( .A(n13792), .B(n13793), .Z(n13778) );
  XOR U16352 ( .A(n13803), .B(n13804), .Z(n13793) );
  ANDN U16353 ( .B(n13805), .A(n13806), .Z(n13803) );
  XOR U16354 ( .A(n13804), .B(n13807), .Z(n13805) );
  XOR U16355 ( .A(n13808), .B(n13809), .Z(n13792) );
  XOR U16356 ( .A(n13810), .B(n13811), .Z(n13809) );
  ANDN U16357 ( .B(n13812), .A(n13813), .Z(n13810) );
  XOR U16358 ( .A(n13814), .B(n13811), .Z(n13812) );
  IV U16359 ( .A(n13790), .Z(n13808) );
  XOR U16360 ( .A(n13815), .B(n13816), .Z(n13790) );
  ANDN U16361 ( .B(n13817), .A(n13818), .Z(n13815) );
  XOR U16362 ( .A(n13816), .B(n13819), .Z(n13817) );
  IV U16363 ( .A(n13798), .Z(n13802) );
  XOR U16364 ( .A(n13798), .B(n13780), .Z(n13800) );
  XOR U16365 ( .A(n13820), .B(n13821), .Z(n13780) );
  AND U16366 ( .A(n242), .B(n13822), .Z(n13820) );
  XOR U16367 ( .A(n13823), .B(n13821), .Z(n13822) );
  NANDN U16368 ( .A(n13782), .B(n13784), .Z(n13798) );
  XOR U16369 ( .A(n13824), .B(n13825), .Z(n13784) );
  AND U16370 ( .A(n242), .B(n13826), .Z(n13824) );
  XOR U16371 ( .A(n13825), .B(n13827), .Z(n13826) );
  XOR U16372 ( .A(n13828), .B(n13829), .Z(n242) );
  AND U16373 ( .A(n13830), .B(n13831), .Z(n13828) );
  XNOR U16374 ( .A(n13829), .B(n13795), .Z(n13831) );
  XNOR U16375 ( .A(n13832), .B(n13833), .Z(n13795) );
  ANDN U16376 ( .B(n13834), .A(n13835), .Z(n13832) );
  XOR U16377 ( .A(n13833), .B(n13836), .Z(n13834) );
  XOR U16378 ( .A(n13829), .B(n13797), .Z(n13830) );
  XOR U16379 ( .A(n13837), .B(n13838), .Z(n13797) );
  AND U16380 ( .A(n246), .B(n13839), .Z(n13837) );
  XOR U16381 ( .A(n13840), .B(n13838), .Z(n13839) );
  XNOR U16382 ( .A(n13841), .B(n13842), .Z(n13829) );
  NAND U16383 ( .A(n13843), .B(n13844), .Z(n13842) );
  XOR U16384 ( .A(n13845), .B(n13821), .Z(n13844) );
  XOR U16385 ( .A(n13835), .B(n13836), .Z(n13821) );
  XOR U16386 ( .A(n13846), .B(n13847), .Z(n13836) );
  ANDN U16387 ( .B(n13848), .A(n13849), .Z(n13846) );
  XOR U16388 ( .A(n13847), .B(n13850), .Z(n13848) );
  XOR U16389 ( .A(n13851), .B(n13852), .Z(n13835) );
  XOR U16390 ( .A(n13853), .B(n13854), .Z(n13852) );
  ANDN U16391 ( .B(n13855), .A(n13856), .Z(n13853) );
  XOR U16392 ( .A(n13857), .B(n13854), .Z(n13855) );
  IV U16393 ( .A(n13833), .Z(n13851) );
  XOR U16394 ( .A(n13858), .B(n13859), .Z(n13833) );
  ANDN U16395 ( .B(n13860), .A(n13861), .Z(n13858) );
  XOR U16396 ( .A(n13859), .B(n13862), .Z(n13860) );
  IV U16397 ( .A(n13841), .Z(n13845) );
  XOR U16398 ( .A(n13841), .B(n13823), .Z(n13843) );
  XOR U16399 ( .A(n13863), .B(n13864), .Z(n13823) );
  AND U16400 ( .A(n246), .B(n13865), .Z(n13863) );
  XOR U16401 ( .A(n13866), .B(n13864), .Z(n13865) );
  NANDN U16402 ( .A(n13825), .B(n13827), .Z(n13841) );
  XOR U16403 ( .A(n13867), .B(n13868), .Z(n13827) );
  AND U16404 ( .A(n246), .B(n13869), .Z(n13867) );
  XOR U16405 ( .A(n13868), .B(n13870), .Z(n13869) );
  XOR U16406 ( .A(n13871), .B(n13872), .Z(n246) );
  AND U16407 ( .A(n13873), .B(n13874), .Z(n13871) );
  XNOR U16408 ( .A(n13872), .B(n13838), .Z(n13874) );
  XNOR U16409 ( .A(n13875), .B(n13876), .Z(n13838) );
  ANDN U16410 ( .B(n13877), .A(n13878), .Z(n13875) );
  XOR U16411 ( .A(n13876), .B(n13879), .Z(n13877) );
  XOR U16412 ( .A(n13872), .B(n13840), .Z(n13873) );
  XOR U16413 ( .A(n13880), .B(n13881), .Z(n13840) );
  AND U16414 ( .A(n250), .B(n13882), .Z(n13880) );
  XOR U16415 ( .A(n13883), .B(n13881), .Z(n13882) );
  XNOR U16416 ( .A(n13884), .B(n13885), .Z(n13872) );
  NAND U16417 ( .A(n13886), .B(n13887), .Z(n13885) );
  XOR U16418 ( .A(n13888), .B(n13864), .Z(n13887) );
  XOR U16419 ( .A(n13878), .B(n13879), .Z(n13864) );
  XOR U16420 ( .A(n13889), .B(n13890), .Z(n13879) );
  ANDN U16421 ( .B(n13891), .A(n13892), .Z(n13889) );
  XOR U16422 ( .A(n13890), .B(n13893), .Z(n13891) );
  XOR U16423 ( .A(n13894), .B(n13895), .Z(n13878) );
  XOR U16424 ( .A(n13896), .B(n13897), .Z(n13895) );
  ANDN U16425 ( .B(n13898), .A(n13899), .Z(n13896) );
  XOR U16426 ( .A(n13900), .B(n13897), .Z(n13898) );
  IV U16427 ( .A(n13876), .Z(n13894) );
  XOR U16428 ( .A(n13901), .B(n13902), .Z(n13876) );
  ANDN U16429 ( .B(n13903), .A(n13904), .Z(n13901) );
  XOR U16430 ( .A(n13902), .B(n13905), .Z(n13903) );
  IV U16431 ( .A(n13884), .Z(n13888) );
  XOR U16432 ( .A(n13884), .B(n13866), .Z(n13886) );
  XOR U16433 ( .A(n13906), .B(n13907), .Z(n13866) );
  AND U16434 ( .A(n250), .B(n13908), .Z(n13906) );
  XOR U16435 ( .A(n13909), .B(n13907), .Z(n13908) );
  NANDN U16436 ( .A(n13868), .B(n13870), .Z(n13884) );
  XOR U16437 ( .A(n13910), .B(n13911), .Z(n13870) );
  AND U16438 ( .A(n250), .B(n13912), .Z(n13910) );
  XOR U16439 ( .A(n13911), .B(n13913), .Z(n13912) );
  XOR U16440 ( .A(n13914), .B(n13915), .Z(n250) );
  AND U16441 ( .A(n13916), .B(n13917), .Z(n13914) );
  XNOR U16442 ( .A(n13915), .B(n13881), .Z(n13917) );
  XNOR U16443 ( .A(n13918), .B(n13919), .Z(n13881) );
  ANDN U16444 ( .B(n13920), .A(n13921), .Z(n13918) );
  XOR U16445 ( .A(n13919), .B(n13922), .Z(n13920) );
  XOR U16446 ( .A(n13915), .B(n13883), .Z(n13916) );
  XOR U16447 ( .A(n13923), .B(n13924), .Z(n13883) );
  AND U16448 ( .A(n254), .B(n13925), .Z(n13923) );
  XOR U16449 ( .A(n13926), .B(n13924), .Z(n13925) );
  XNOR U16450 ( .A(n13927), .B(n13928), .Z(n13915) );
  NAND U16451 ( .A(n13929), .B(n13930), .Z(n13928) );
  XOR U16452 ( .A(n13931), .B(n13907), .Z(n13930) );
  XOR U16453 ( .A(n13921), .B(n13922), .Z(n13907) );
  XOR U16454 ( .A(n13932), .B(n13933), .Z(n13922) );
  ANDN U16455 ( .B(n13934), .A(n13935), .Z(n13932) );
  XOR U16456 ( .A(n13933), .B(n13936), .Z(n13934) );
  XOR U16457 ( .A(n13937), .B(n13938), .Z(n13921) );
  XOR U16458 ( .A(n13939), .B(n13940), .Z(n13938) );
  ANDN U16459 ( .B(n13941), .A(n13942), .Z(n13939) );
  XOR U16460 ( .A(n13943), .B(n13940), .Z(n13941) );
  IV U16461 ( .A(n13919), .Z(n13937) );
  XOR U16462 ( .A(n13944), .B(n13945), .Z(n13919) );
  ANDN U16463 ( .B(n13946), .A(n13947), .Z(n13944) );
  XOR U16464 ( .A(n13945), .B(n13948), .Z(n13946) );
  IV U16465 ( .A(n13927), .Z(n13931) );
  XOR U16466 ( .A(n13927), .B(n13909), .Z(n13929) );
  XOR U16467 ( .A(n13949), .B(n13950), .Z(n13909) );
  AND U16468 ( .A(n254), .B(n13951), .Z(n13949) );
  XOR U16469 ( .A(n13952), .B(n13950), .Z(n13951) );
  NANDN U16470 ( .A(n13911), .B(n13913), .Z(n13927) );
  XOR U16471 ( .A(n13953), .B(n13954), .Z(n13913) );
  AND U16472 ( .A(n254), .B(n13955), .Z(n13953) );
  XOR U16473 ( .A(n13954), .B(n13956), .Z(n13955) );
  XOR U16474 ( .A(n13957), .B(n13958), .Z(n254) );
  AND U16475 ( .A(n13959), .B(n13960), .Z(n13957) );
  XNOR U16476 ( .A(n13958), .B(n13924), .Z(n13960) );
  XNOR U16477 ( .A(n13961), .B(n13962), .Z(n13924) );
  ANDN U16478 ( .B(n13963), .A(n13964), .Z(n13961) );
  XOR U16479 ( .A(n13962), .B(n13965), .Z(n13963) );
  XOR U16480 ( .A(n13958), .B(n13926), .Z(n13959) );
  XOR U16481 ( .A(n13966), .B(n13967), .Z(n13926) );
  AND U16482 ( .A(n258), .B(n13968), .Z(n13966) );
  XOR U16483 ( .A(n13969), .B(n13967), .Z(n13968) );
  XNOR U16484 ( .A(n13970), .B(n13971), .Z(n13958) );
  NAND U16485 ( .A(n13972), .B(n13973), .Z(n13971) );
  XOR U16486 ( .A(n13974), .B(n13950), .Z(n13973) );
  XOR U16487 ( .A(n13964), .B(n13965), .Z(n13950) );
  XOR U16488 ( .A(n13975), .B(n13976), .Z(n13965) );
  ANDN U16489 ( .B(n13977), .A(n13978), .Z(n13975) );
  XOR U16490 ( .A(n13976), .B(n13979), .Z(n13977) );
  XOR U16491 ( .A(n13980), .B(n13981), .Z(n13964) );
  XOR U16492 ( .A(n13982), .B(n13983), .Z(n13981) );
  ANDN U16493 ( .B(n13984), .A(n13985), .Z(n13982) );
  XOR U16494 ( .A(n13986), .B(n13983), .Z(n13984) );
  IV U16495 ( .A(n13962), .Z(n13980) );
  XOR U16496 ( .A(n13987), .B(n13988), .Z(n13962) );
  ANDN U16497 ( .B(n13989), .A(n13990), .Z(n13987) );
  XOR U16498 ( .A(n13988), .B(n13991), .Z(n13989) );
  IV U16499 ( .A(n13970), .Z(n13974) );
  XOR U16500 ( .A(n13970), .B(n13952), .Z(n13972) );
  XOR U16501 ( .A(n13992), .B(n13993), .Z(n13952) );
  AND U16502 ( .A(n258), .B(n13994), .Z(n13992) );
  XOR U16503 ( .A(n13995), .B(n13993), .Z(n13994) );
  NANDN U16504 ( .A(n13954), .B(n13956), .Z(n13970) );
  XOR U16505 ( .A(n13996), .B(n13997), .Z(n13956) );
  AND U16506 ( .A(n258), .B(n13998), .Z(n13996) );
  XOR U16507 ( .A(n13997), .B(n13999), .Z(n13998) );
  XOR U16508 ( .A(n14000), .B(n14001), .Z(n258) );
  AND U16509 ( .A(n14002), .B(n14003), .Z(n14000) );
  XNOR U16510 ( .A(n14001), .B(n13967), .Z(n14003) );
  XNOR U16511 ( .A(n14004), .B(n14005), .Z(n13967) );
  ANDN U16512 ( .B(n14006), .A(n14007), .Z(n14004) );
  XOR U16513 ( .A(n14005), .B(n14008), .Z(n14006) );
  XOR U16514 ( .A(n14001), .B(n13969), .Z(n14002) );
  XOR U16515 ( .A(n14009), .B(n14010), .Z(n13969) );
  AND U16516 ( .A(n262), .B(n14011), .Z(n14009) );
  XOR U16517 ( .A(n14012), .B(n14010), .Z(n14011) );
  XNOR U16518 ( .A(n14013), .B(n14014), .Z(n14001) );
  NAND U16519 ( .A(n14015), .B(n14016), .Z(n14014) );
  XOR U16520 ( .A(n14017), .B(n13993), .Z(n14016) );
  XOR U16521 ( .A(n14007), .B(n14008), .Z(n13993) );
  XOR U16522 ( .A(n14018), .B(n14019), .Z(n14008) );
  ANDN U16523 ( .B(n14020), .A(n14021), .Z(n14018) );
  XOR U16524 ( .A(n14019), .B(n14022), .Z(n14020) );
  XOR U16525 ( .A(n14023), .B(n14024), .Z(n14007) );
  XOR U16526 ( .A(n14025), .B(n14026), .Z(n14024) );
  ANDN U16527 ( .B(n14027), .A(n14028), .Z(n14025) );
  XOR U16528 ( .A(n14029), .B(n14026), .Z(n14027) );
  IV U16529 ( .A(n14005), .Z(n14023) );
  XOR U16530 ( .A(n14030), .B(n14031), .Z(n14005) );
  ANDN U16531 ( .B(n14032), .A(n14033), .Z(n14030) );
  XOR U16532 ( .A(n14031), .B(n14034), .Z(n14032) );
  IV U16533 ( .A(n14013), .Z(n14017) );
  XOR U16534 ( .A(n14013), .B(n13995), .Z(n14015) );
  XOR U16535 ( .A(n14035), .B(n14036), .Z(n13995) );
  AND U16536 ( .A(n262), .B(n14037), .Z(n14035) );
  XOR U16537 ( .A(n14038), .B(n14036), .Z(n14037) );
  NANDN U16538 ( .A(n13997), .B(n13999), .Z(n14013) );
  XOR U16539 ( .A(n14039), .B(n14040), .Z(n13999) );
  AND U16540 ( .A(n262), .B(n14041), .Z(n14039) );
  XOR U16541 ( .A(n14040), .B(n14042), .Z(n14041) );
  XOR U16542 ( .A(n14043), .B(n14044), .Z(n262) );
  AND U16543 ( .A(n14045), .B(n14046), .Z(n14043) );
  XNOR U16544 ( .A(n14044), .B(n14010), .Z(n14046) );
  XNOR U16545 ( .A(n14047), .B(n14048), .Z(n14010) );
  ANDN U16546 ( .B(n14049), .A(n14050), .Z(n14047) );
  XOR U16547 ( .A(n14048), .B(n14051), .Z(n14049) );
  XOR U16548 ( .A(n14044), .B(n14012), .Z(n14045) );
  XOR U16549 ( .A(n14052), .B(n14053), .Z(n14012) );
  AND U16550 ( .A(n266), .B(n14054), .Z(n14052) );
  XOR U16551 ( .A(n14055), .B(n14053), .Z(n14054) );
  XNOR U16552 ( .A(n14056), .B(n14057), .Z(n14044) );
  NAND U16553 ( .A(n14058), .B(n14059), .Z(n14057) );
  XOR U16554 ( .A(n14060), .B(n14036), .Z(n14059) );
  XOR U16555 ( .A(n14050), .B(n14051), .Z(n14036) );
  XOR U16556 ( .A(n14061), .B(n14062), .Z(n14051) );
  ANDN U16557 ( .B(n14063), .A(n14064), .Z(n14061) );
  XOR U16558 ( .A(n14062), .B(n14065), .Z(n14063) );
  XOR U16559 ( .A(n14066), .B(n14067), .Z(n14050) );
  XOR U16560 ( .A(n14068), .B(n14069), .Z(n14067) );
  ANDN U16561 ( .B(n14070), .A(n14071), .Z(n14068) );
  XOR U16562 ( .A(n14072), .B(n14069), .Z(n14070) );
  IV U16563 ( .A(n14048), .Z(n14066) );
  XOR U16564 ( .A(n14073), .B(n14074), .Z(n14048) );
  ANDN U16565 ( .B(n14075), .A(n14076), .Z(n14073) );
  XOR U16566 ( .A(n14074), .B(n14077), .Z(n14075) );
  IV U16567 ( .A(n14056), .Z(n14060) );
  XOR U16568 ( .A(n14056), .B(n14038), .Z(n14058) );
  XOR U16569 ( .A(n14078), .B(n14079), .Z(n14038) );
  AND U16570 ( .A(n266), .B(n14080), .Z(n14078) );
  XOR U16571 ( .A(n14081), .B(n14079), .Z(n14080) );
  NANDN U16572 ( .A(n14040), .B(n14042), .Z(n14056) );
  XOR U16573 ( .A(n14082), .B(n14083), .Z(n14042) );
  AND U16574 ( .A(n266), .B(n14084), .Z(n14082) );
  XOR U16575 ( .A(n14083), .B(n14085), .Z(n14084) );
  XOR U16576 ( .A(n14086), .B(n14087), .Z(n266) );
  AND U16577 ( .A(n14088), .B(n14089), .Z(n14086) );
  XNOR U16578 ( .A(n14087), .B(n14053), .Z(n14089) );
  XNOR U16579 ( .A(n14090), .B(n14091), .Z(n14053) );
  ANDN U16580 ( .B(n14092), .A(n14093), .Z(n14090) );
  XOR U16581 ( .A(n14091), .B(n14094), .Z(n14092) );
  XOR U16582 ( .A(n14087), .B(n14055), .Z(n14088) );
  XOR U16583 ( .A(n14095), .B(n14096), .Z(n14055) );
  AND U16584 ( .A(n270), .B(n14097), .Z(n14095) );
  XOR U16585 ( .A(n14098), .B(n14096), .Z(n14097) );
  XNOR U16586 ( .A(n14099), .B(n14100), .Z(n14087) );
  NAND U16587 ( .A(n14101), .B(n14102), .Z(n14100) );
  XOR U16588 ( .A(n14103), .B(n14079), .Z(n14102) );
  XOR U16589 ( .A(n14093), .B(n14094), .Z(n14079) );
  XOR U16590 ( .A(n14104), .B(n14105), .Z(n14094) );
  ANDN U16591 ( .B(n14106), .A(n14107), .Z(n14104) );
  XOR U16592 ( .A(n14105), .B(n14108), .Z(n14106) );
  XOR U16593 ( .A(n14109), .B(n14110), .Z(n14093) );
  XOR U16594 ( .A(n14111), .B(n14112), .Z(n14110) );
  ANDN U16595 ( .B(n14113), .A(n14114), .Z(n14111) );
  XOR U16596 ( .A(n14115), .B(n14112), .Z(n14113) );
  IV U16597 ( .A(n14091), .Z(n14109) );
  XOR U16598 ( .A(n14116), .B(n14117), .Z(n14091) );
  ANDN U16599 ( .B(n14118), .A(n14119), .Z(n14116) );
  XOR U16600 ( .A(n14117), .B(n14120), .Z(n14118) );
  IV U16601 ( .A(n14099), .Z(n14103) );
  XOR U16602 ( .A(n14099), .B(n14081), .Z(n14101) );
  XOR U16603 ( .A(n14121), .B(n14122), .Z(n14081) );
  AND U16604 ( .A(n270), .B(n14123), .Z(n14121) );
  XOR U16605 ( .A(n14124), .B(n14122), .Z(n14123) );
  NANDN U16606 ( .A(n14083), .B(n14085), .Z(n14099) );
  XOR U16607 ( .A(n14125), .B(n14126), .Z(n14085) );
  AND U16608 ( .A(n270), .B(n14127), .Z(n14125) );
  XOR U16609 ( .A(n14126), .B(n14128), .Z(n14127) );
  XOR U16610 ( .A(n14129), .B(n14130), .Z(n270) );
  AND U16611 ( .A(n14131), .B(n14132), .Z(n14129) );
  XNOR U16612 ( .A(n14130), .B(n14096), .Z(n14132) );
  XNOR U16613 ( .A(n14133), .B(n14134), .Z(n14096) );
  ANDN U16614 ( .B(n14135), .A(n14136), .Z(n14133) );
  XOR U16615 ( .A(n14134), .B(n14137), .Z(n14135) );
  XOR U16616 ( .A(n14130), .B(n14098), .Z(n14131) );
  XOR U16617 ( .A(n14138), .B(n14139), .Z(n14098) );
  AND U16618 ( .A(n274), .B(n14140), .Z(n14138) );
  XOR U16619 ( .A(n14141), .B(n14139), .Z(n14140) );
  XNOR U16620 ( .A(n14142), .B(n14143), .Z(n14130) );
  NAND U16621 ( .A(n14144), .B(n14145), .Z(n14143) );
  XOR U16622 ( .A(n14146), .B(n14122), .Z(n14145) );
  XOR U16623 ( .A(n14136), .B(n14137), .Z(n14122) );
  XOR U16624 ( .A(n14147), .B(n14148), .Z(n14137) );
  ANDN U16625 ( .B(n14149), .A(n14150), .Z(n14147) );
  XOR U16626 ( .A(n14148), .B(n14151), .Z(n14149) );
  XOR U16627 ( .A(n14152), .B(n14153), .Z(n14136) );
  XOR U16628 ( .A(n14154), .B(n14155), .Z(n14153) );
  ANDN U16629 ( .B(n14156), .A(n14157), .Z(n14154) );
  XOR U16630 ( .A(n14158), .B(n14155), .Z(n14156) );
  IV U16631 ( .A(n14134), .Z(n14152) );
  XOR U16632 ( .A(n14159), .B(n14160), .Z(n14134) );
  ANDN U16633 ( .B(n14161), .A(n14162), .Z(n14159) );
  XOR U16634 ( .A(n14160), .B(n14163), .Z(n14161) );
  IV U16635 ( .A(n14142), .Z(n14146) );
  XOR U16636 ( .A(n14142), .B(n14124), .Z(n14144) );
  XOR U16637 ( .A(n14164), .B(n14165), .Z(n14124) );
  AND U16638 ( .A(n274), .B(n14166), .Z(n14164) );
  XOR U16639 ( .A(n14167), .B(n14165), .Z(n14166) );
  NANDN U16640 ( .A(n14126), .B(n14128), .Z(n14142) );
  XOR U16641 ( .A(n14168), .B(n14169), .Z(n14128) );
  AND U16642 ( .A(n274), .B(n14170), .Z(n14168) );
  XOR U16643 ( .A(n14169), .B(n14171), .Z(n14170) );
  XOR U16644 ( .A(n14172), .B(n14173), .Z(n274) );
  AND U16645 ( .A(n14174), .B(n14175), .Z(n14172) );
  XNOR U16646 ( .A(n14173), .B(n14139), .Z(n14175) );
  XNOR U16647 ( .A(n14176), .B(n14177), .Z(n14139) );
  ANDN U16648 ( .B(n14178), .A(n14179), .Z(n14176) );
  XOR U16649 ( .A(n14177), .B(n14180), .Z(n14178) );
  XOR U16650 ( .A(n14173), .B(n14141), .Z(n14174) );
  XOR U16651 ( .A(n14181), .B(n14182), .Z(n14141) );
  AND U16652 ( .A(n278), .B(n14183), .Z(n14181) );
  XOR U16653 ( .A(n14184), .B(n14182), .Z(n14183) );
  XNOR U16654 ( .A(n14185), .B(n14186), .Z(n14173) );
  NAND U16655 ( .A(n14187), .B(n14188), .Z(n14186) );
  XOR U16656 ( .A(n14189), .B(n14165), .Z(n14188) );
  XOR U16657 ( .A(n14179), .B(n14180), .Z(n14165) );
  XOR U16658 ( .A(n14190), .B(n14191), .Z(n14180) );
  ANDN U16659 ( .B(n14192), .A(n14193), .Z(n14190) );
  XOR U16660 ( .A(n14191), .B(n14194), .Z(n14192) );
  XOR U16661 ( .A(n14195), .B(n14196), .Z(n14179) );
  XOR U16662 ( .A(n14197), .B(n14198), .Z(n14196) );
  ANDN U16663 ( .B(n14199), .A(n14200), .Z(n14197) );
  XOR U16664 ( .A(n14201), .B(n14198), .Z(n14199) );
  IV U16665 ( .A(n14177), .Z(n14195) );
  XOR U16666 ( .A(n14202), .B(n14203), .Z(n14177) );
  ANDN U16667 ( .B(n14204), .A(n14205), .Z(n14202) );
  XOR U16668 ( .A(n14203), .B(n14206), .Z(n14204) );
  IV U16669 ( .A(n14185), .Z(n14189) );
  XOR U16670 ( .A(n14185), .B(n14167), .Z(n14187) );
  XOR U16671 ( .A(n14207), .B(n14208), .Z(n14167) );
  AND U16672 ( .A(n278), .B(n14209), .Z(n14207) );
  XOR U16673 ( .A(n14210), .B(n14208), .Z(n14209) );
  NANDN U16674 ( .A(n14169), .B(n14171), .Z(n14185) );
  XOR U16675 ( .A(n14211), .B(n14212), .Z(n14171) );
  AND U16676 ( .A(n278), .B(n14213), .Z(n14211) );
  XOR U16677 ( .A(n14212), .B(n14214), .Z(n14213) );
  XOR U16678 ( .A(n14215), .B(n14216), .Z(n278) );
  AND U16679 ( .A(n14217), .B(n14218), .Z(n14215) );
  XNOR U16680 ( .A(n14216), .B(n14182), .Z(n14218) );
  XNOR U16681 ( .A(n14219), .B(n14220), .Z(n14182) );
  ANDN U16682 ( .B(n14221), .A(n14222), .Z(n14219) );
  XOR U16683 ( .A(n14220), .B(n14223), .Z(n14221) );
  XOR U16684 ( .A(n14216), .B(n14184), .Z(n14217) );
  XOR U16685 ( .A(n14224), .B(n14225), .Z(n14184) );
  AND U16686 ( .A(n282), .B(n14226), .Z(n14224) );
  XOR U16687 ( .A(n14227), .B(n14225), .Z(n14226) );
  XNOR U16688 ( .A(n14228), .B(n14229), .Z(n14216) );
  NAND U16689 ( .A(n14230), .B(n14231), .Z(n14229) );
  XOR U16690 ( .A(n14232), .B(n14208), .Z(n14231) );
  XOR U16691 ( .A(n14222), .B(n14223), .Z(n14208) );
  XOR U16692 ( .A(n14233), .B(n14234), .Z(n14223) );
  ANDN U16693 ( .B(n14235), .A(n14236), .Z(n14233) );
  XOR U16694 ( .A(n14234), .B(n14237), .Z(n14235) );
  XOR U16695 ( .A(n14238), .B(n14239), .Z(n14222) );
  XOR U16696 ( .A(n14240), .B(n14241), .Z(n14239) );
  ANDN U16697 ( .B(n14242), .A(n14243), .Z(n14240) );
  XOR U16698 ( .A(n14244), .B(n14241), .Z(n14242) );
  IV U16699 ( .A(n14220), .Z(n14238) );
  XOR U16700 ( .A(n14245), .B(n14246), .Z(n14220) );
  ANDN U16701 ( .B(n14247), .A(n14248), .Z(n14245) );
  XOR U16702 ( .A(n14246), .B(n14249), .Z(n14247) );
  IV U16703 ( .A(n14228), .Z(n14232) );
  XOR U16704 ( .A(n14228), .B(n14210), .Z(n14230) );
  XOR U16705 ( .A(n14250), .B(n14251), .Z(n14210) );
  AND U16706 ( .A(n282), .B(n14252), .Z(n14250) );
  XOR U16707 ( .A(n14253), .B(n14251), .Z(n14252) );
  NANDN U16708 ( .A(n14212), .B(n14214), .Z(n14228) );
  XOR U16709 ( .A(n14254), .B(n14255), .Z(n14214) );
  AND U16710 ( .A(n282), .B(n14256), .Z(n14254) );
  XOR U16711 ( .A(n14255), .B(n14257), .Z(n14256) );
  XOR U16712 ( .A(n14258), .B(n14259), .Z(n282) );
  AND U16713 ( .A(n14260), .B(n14261), .Z(n14258) );
  XNOR U16714 ( .A(n14259), .B(n14225), .Z(n14261) );
  XNOR U16715 ( .A(n14262), .B(n14263), .Z(n14225) );
  ANDN U16716 ( .B(n14264), .A(n14265), .Z(n14262) );
  XOR U16717 ( .A(n14263), .B(n14266), .Z(n14264) );
  XOR U16718 ( .A(n14259), .B(n14227), .Z(n14260) );
  XOR U16719 ( .A(n14267), .B(n14268), .Z(n14227) );
  AND U16720 ( .A(n286), .B(n14269), .Z(n14267) );
  XOR U16721 ( .A(n14270), .B(n14268), .Z(n14269) );
  XNOR U16722 ( .A(n14271), .B(n14272), .Z(n14259) );
  NAND U16723 ( .A(n14273), .B(n14274), .Z(n14272) );
  XOR U16724 ( .A(n14275), .B(n14251), .Z(n14274) );
  XOR U16725 ( .A(n14265), .B(n14266), .Z(n14251) );
  XOR U16726 ( .A(n14276), .B(n14277), .Z(n14266) );
  ANDN U16727 ( .B(n14278), .A(n14279), .Z(n14276) );
  XOR U16728 ( .A(n14277), .B(n14280), .Z(n14278) );
  XOR U16729 ( .A(n14281), .B(n14282), .Z(n14265) );
  XOR U16730 ( .A(n14283), .B(n14284), .Z(n14282) );
  ANDN U16731 ( .B(n14285), .A(n14286), .Z(n14283) );
  XOR U16732 ( .A(n14287), .B(n14284), .Z(n14285) );
  IV U16733 ( .A(n14263), .Z(n14281) );
  XOR U16734 ( .A(n14288), .B(n14289), .Z(n14263) );
  ANDN U16735 ( .B(n14290), .A(n14291), .Z(n14288) );
  XOR U16736 ( .A(n14289), .B(n14292), .Z(n14290) );
  IV U16737 ( .A(n14271), .Z(n14275) );
  XOR U16738 ( .A(n14271), .B(n14253), .Z(n14273) );
  XOR U16739 ( .A(n14293), .B(n14294), .Z(n14253) );
  AND U16740 ( .A(n286), .B(n14295), .Z(n14293) );
  XOR U16741 ( .A(n14296), .B(n14294), .Z(n14295) );
  NANDN U16742 ( .A(n14255), .B(n14257), .Z(n14271) );
  XOR U16743 ( .A(n14297), .B(n14298), .Z(n14257) );
  AND U16744 ( .A(n286), .B(n14299), .Z(n14297) );
  XOR U16745 ( .A(n14298), .B(n14300), .Z(n14299) );
  XOR U16746 ( .A(n14301), .B(n14302), .Z(n286) );
  AND U16747 ( .A(n14303), .B(n14304), .Z(n14301) );
  XNOR U16748 ( .A(n14302), .B(n14268), .Z(n14304) );
  XNOR U16749 ( .A(n14305), .B(n14306), .Z(n14268) );
  ANDN U16750 ( .B(n14307), .A(n14308), .Z(n14305) );
  XOR U16751 ( .A(n14306), .B(n14309), .Z(n14307) );
  XOR U16752 ( .A(n14302), .B(n14270), .Z(n14303) );
  XOR U16753 ( .A(n14310), .B(n14311), .Z(n14270) );
  AND U16754 ( .A(n290), .B(n14312), .Z(n14310) );
  XOR U16755 ( .A(n14313), .B(n14311), .Z(n14312) );
  XNOR U16756 ( .A(n14314), .B(n14315), .Z(n14302) );
  NAND U16757 ( .A(n14316), .B(n14317), .Z(n14315) );
  XOR U16758 ( .A(n14318), .B(n14294), .Z(n14317) );
  XOR U16759 ( .A(n14308), .B(n14309), .Z(n14294) );
  XOR U16760 ( .A(n14319), .B(n14320), .Z(n14309) );
  ANDN U16761 ( .B(n14321), .A(n14322), .Z(n14319) );
  XOR U16762 ( .A(n14320), .B(n14323), .Z(n14321) );
  XOR U16763 ( .A(n14324), .B(n14325), .Z(n14308) );
  XOR U16764 ( .A(n14326), .B(n14327), .Z(n14325) );
  ANDN U16765 ( .B(n14328), .A(n14329), .Z(n14326) );
  XOR U16766 ( .A(n14330), .B(n14327), .Z(n14328) );
  IV U16767 ( .A(n14306), .Z(n14324) );
  XOR U16768 ( .A(n14331), .B(n14332), .Z(n14306) );
  ANDN U16769 ( .B(n14333), .A(n14334), .Z(n14331) );
  XOR U16770 ( .A(n14332), .B(n14335), .Z(n14333) );
  IV U16771 ( .A(n14314), .Z(n14318) );
  XOR U16772 ( .A(n14314), .B(n14296), .Z(n14316) );
  XOR U16773 ( .A(n14336), .B(n14337), .Z(n14296) );
  AND U16774 ( .A(n290), .B(n14338), .Z(n14336) );
  XOR U16775 ( .A(n14339), .B(n14337), .Z(n14338) );
  NANDN U16776 ( .A(n14298), .B(n14300), .Z(n14314) );
  XOR U16777 ( .A(n14340), .B(n14341), .Z(n14300) );
  AND U16778 ( .A(n290), .B(n14342), .Z(n14340) );
  XOR U16779 ( .A(n14341), .B(n14343), .Z(n14342) );
  XOR U16780 ( .A(n14344), .B(n14345), .Z(n290) );
  AND U16781 ( .A(n14346), .B(n14347), .Z(n14344) );
  XNOR U16782 ( .A(n14345), .B(n14311), .Z(n14347) );
  XNOR U16783 ( .A(n14348), .B(n14349), .Z(n14311) );
  ANDN U16784 ( .B(n14350), .A(n14351), .Z(n14348) );
  XOR U16785 ( .A(n14349), .B(n14352), .Z(n14350) );
  XOR U16786 ( .A(n14345), .B(n14313), .Z(n14346) );
  XOR U16787 ( .A(n14353), .B(n14354), .Z(n14313) );
  AND U16788 ( .A(n294), .B(n14355), .Z(n14353) );
  XOR U16789 ( .A(n14356), .B(n14354), .Z(n14355) );
  XNOR U16790 ( .A(n14357), .B(n14358), .Z(n14345) );
  NAND U16791 ( .A(n14359), .B(n14360), .Z(n14358) );
  XOR U16792 ( .A(n14361), .B(n14337), .Z(n14360) );
  XOR U16793 ( .A(n14351), .B(n14352), .Z(n14337) );
  XOR U16794 ( .A(n14362), .B(n14363), .Z(n14352) );
  ANDN U16795 ( .B(n14364), .A(n14365), .Z(n14362) );
  XOR U16796 ( .A(n14363), .B(n14366), .Z(n14364) );
  XOR U16797 ( .A(n14367), .B(n14368), .Z(n14351) );
  XOR U16798 ( .A(n14369), .B(n14370), .Z(n14368) );
  ANDN U16799 ( .B(n14371), .A(n14372), .Z(n14369) );
  XOR U16800 ( .A(n14373), .B(n14370), .Z(n14371) );
  IV U16801 ( .A(n14349), .Z(n14367) );
  XOR U16802 ( .A(n14374), .B(n14375), .Z(n14349) );
  ANDN U16803 ( .B(n14376), .A(n14377), .Z(n14374) );
  XOR U16804 ( .A(n14375), .B(n14378), .Z(n14376) );
  IV U16805 ( .A(n14357), .Z(n14361) );
  XOR U16806 ( .A(n14357), .B(n14339), .Z(n14359) );
  XOR U16807 ( .A(n14379), .B(n14380), .Z(n14339) );
  AND U16808 ( .A(n294), .B(n14381), .Z(n14379) );
  XOR U16809 ( .A(n14382), .B(n14380), .Z(n14381) );
  NANDN U16810 ( .A(n14341), .B(n14343), .Z(n14357) );
  XOR U16811 ( .A(n14383), .B(n14384), .Z(n14343) );
  AND U16812 ( .A(n294), .B(n14385), .Z(n14383) );
  XOR U16813 ( .A(n14384), .B(n14386), .Z(n14385) );
  XOR U16814 ( .A(n14387), .B(n14388), .Z(n294) );
  AND U16815 ( .A(n14389), .B(n14390), .Z(n14387) );
  XNOR U16816 ( .A(n14388), .B(n14354), .Z(n14390) );
  XNOR U16817 ( .A(n14391), .B(n14392), .Z(n14354) );
  ANDN U16818 ( .B(n14393), .A(n14394), .Z(n14391) );
  XOR U16819 ( .A(n14392), .B(n14395), .Z(n14393) );
  XOR U16820 ( .A(n14388), .B(n14356), .Z(n14389) );
  XOR U16821 ( .A(n14396), .B(n14397), .Z(n14356) );
  AND U16822 ( .A(n298), .B(n14398), .Z(n14396) );
  XOR U16823 ( .A(n14399), .B(n14397), .Z(n14398) );
  XNOR U16824 ( .A(n14400), .B(n14401), .Z(n14388) );
  NAND U16825 ( .A(n14402), .B(n14403), .Z(n14401) );
  XOR U16826 ( .A(n14404), .B(n14380), .Z(n14403) );
  XOR U16827 ( .A(n14394), .B(n14395), .Z(n14380) );
  XOR U16828 ( .A(n14405), .B(n14406), .Z(n14395) );
  ANDN U16829 ( .B(n14407), .A(n14408), .Z(n14405) );
  XOR U16830 ( .A(n14406), .B(n14409), .Z(n14407) );
  XOR U16831 ( .A(n14410), .B(n14411), .Z(n14394) );
  XOR U16832 ( .A(n14412), .B(n14413), .Z(n14411) );
  ANDN U16833 ( .B(n14414), .A(n14415), .Z(n14412) );
  XOR U16834 ( .A(n14416), .B(n14413), .Z(n14414) );
  IV U16835 ( .A(n14392), .Z(n14410) );
  XOR U16836 ( .A(n14417), .B(n14418), .Z(n14392) );
  ANDN U16837 ( .B(n14419), .A(n14420), .Z(n14417) );
  XOR U16838 ( .A(n14418), .B(n14421), .Z(n14419) );
  IV U16839 ( .A(n14400), .Z(n14404) );
  XOR U16840 ( .A(n14400), .B(n14382), .Z(n14402) );
  XOR U16841 ( .A(n14422), .B(n14423), .Z(n14382) );
  AND U16842 ( .A(n298), .B(n14424), .Z(n14422) );
  XOR U16843 ( .A(n14425), .B(n14423), .Z(n14424) );
  NANDN U16844 ( .A(n14384), .B(n14386), .Z(n14400) );
  XOR U16845 ( .A(n14426), .B(n14427), .Z(n14386) );
  AND U16846 ( .A(n298), .B(n14428), .Z(n14426) );
  XOR U16847 ( .A(n14427), .B(n14429), .Z(n14428) );
  XOR U16848 ( .A(n14430), .B(n14431), .Z(n298) );
  AND U16849 ( .A(n14432), .B(n14433), .Z(n14430) );
  XNOR U16850 ( .A(n14431), .B(n14397), .Z(n14433) );
  XNOR U16851 ( .A(n14434), .B(n14435), .Z(n14397) );
  ANDN U16852 ( .B(n14436), .A(n14437), .Z(n14434) );
  XOR U16853 ( .A(n14435), .B(n14438), .Z(n14436) );
  XOR U16854 ( .A(n14431), .B(n14399), .Z(n14432) );
  XOR U16855 ( .A(n14439), .B(n14440), .Z(n14399) );
  AND U16856 ( .A(n302), .B(n14441), .Z(n14439) );
  XOR U16857 ( .A(n14442), .B(n14440), .Z(n14441) );
  XNOR U16858 ( .A(n14443), .B(n14444), .Z(n14431) );
  NAND U16859 ( .A(n14445), .B(n14446), .Z(n14444) );
  XOR U16860 ( .A(n14447), .B(n14423), .Z(n14446) );
  XOR U16861 ( .A(n14437), .B(n14438), .Z(n14423) );
  XOR U16862 ( .A(n14448), .B(n14449), .Z(n14438) );
  ANDN U16863 ( .B(n14450), .A(n14451), .Z(n14448) );
  XOR U16864 ( .A(n14449), .B(n14452), .Z(n14450) );
  XOR U16865 ( .A(n14453), .B(n14454), .Z(n14437) );
  XOR U16866 ( .A(n14455), .B(n14456), .Z(n14454) );
  ANDN U16867 ( .B(n14457), .A(n14458), .Z(n14455) );
  XOR U16868 ( .A(n14459), .B(n14456), .Z(n14457) );
  IV U16869 ( .A(n14435), .Z(n14453) );
  XOR U16870 ( .A(n14460), .B(n14461), .Z(n14435) );
  ANDN U16871 ( .B(n14462), .A(n14463), .Z(n14460) );
  XOR U16872 ( .A(n14461), .B(n14464), .Z(n14462) );
  IV U16873 ( .A(n14443), .Z(n14447) );
  XOR U16874 ( .A(n14443), .B(n14425), .Z(n14445) );
  XOR U16875 ( .A(n14465), .B(n14466), .Z(n14425) );
  AND U16876 ( .A(n302), .B(n14467), .Z(n14465) );
  XOR U16877 ( .A(n14468), .B(n14466), .Z(n14467) );
  NANDN U16878 ( .A(n14427), .B(n14429), .Z(n14443) );
  XOR U16879 ( .A(n14469), .B(n14470), .Z(n14429) );
  AND U16880 ( .A(n302), .B(n14471), .Z(n14469) );
  XOR U16881 ( .A(n14470), .B(n14472), .Z(n14471) );
  XOR U16882 ( .A(n14473), .B(n14474), .Z(n302) );
  AND U16883 ( .A(n14475), .B(n14476), .Z(n14473) );
  XNOR U16884 ( .A(n14474), .B(n14440), .Z(n14476) );
  XNOR U16885 ( .A(n14477), .B(n14478), .Z(n14440) );
  ANDN U16886 ( .B(n14479), .A(n14480), .Z(n14477) );
  XOR U16887 ( .A(n14478), .B(n14481), .Z(n14479) );
  XOR U16888 ( .A(n14474), .B(n14442), .Z(n14475) );
  XOR U16889 ( .A(n14482), .B(n14483), .Z(n14442) );
  AND U16890 ( .A(n306), .B(n14484), .Z(n14482) );
  XOR U16891 ( .A(n14485), .B(n14483), .Z(n14484) );
  XNOR U16892 ( .A(n14486), .B(n14487), .Z(n14474) );
  NAND U16893 ( .A(n14488), .B(n14489), .Z(n14487) );
  XOR U16894 ( .A(n14490), .B(n14466), .Z(n14489) );
  XOR U16895 ( .A(n14480), .B(n14481), .Z(n14466) );
  XOR U16896 ( .A(n14491), .B(n14492), .Z(n14481) );
  ANDN U16897 ( .B(n14493), .A(n14494), .Z(n14491) );
  XOR U16898 ( .A(n14492), .B(n14495), .Z(n14493) );
  XOR U16899 ( .A(n14496), .B(n14497), .Z(n14480) );
  XOR U16900 ( .A(n14498), .B(n14499), .Z(n14497) );
  ANDN U16901 ( .B(n14500), .A(n14501), .Z(n14498) );
  XOR U16902 ( .A(n14502), .B(n14499), .Z(n14500) );
  IV U16903 ( .A(n14478), .Z(n14496) );
  XOR U16904 ( .A(n14503), .B(n14504), .Z(n14478) );
  ANDN U16905 ( .B(n14505), .A(n14506), .Z(n14503) );
  XOR U16906 ( .A(n14504), .B(n14507), .Z(n14505) );
  IV U16907 ( .A(n14486), .Z(n14490) );
  XOR U16908 ( .A(n14486), .B(n14468), .Z(n14488) );
  XOR U16909 ( .A(n14508), .B(n14509), .Z(n14468) );
  AND U16910 ( .A(n306), .B(n14510), .Z(n14508) );
  XOR U16911 ( .A(n14511), .B(n14509), .Z(n14510) );
  NANDN U16912 ( .A(n14470), .B(n14472), .Z(n14486) );
  XOR U16913 ( .A(n14512), .B(n14513), .Z(n14472) );
  AND U16914 ( .A(n306), .B(n14514), .Z(n14512) );
  XOR U16915 ( .A(n14513), .B(n14515), .Z(n14514) );
  XOR U16916 ( .A(n14516), .B(n14517), .Z(n306) );
  AND U16917 ( .A(n14518), .B(n14519), .Z(n14516) );
  XNOR U16918 ( .A(n14517), .B(n14483), .Z(n14519) );
  XNOR U16919 ( .A(n14520), .B(n14521), .Z(n14483) );
  ANDN U16920 ( .B(n14522), .A(n14523), .Z(n14520) );
  XOR U16921 ( .A(n14521), .B(n14524), .Z(n14522) );
  XOR U16922 ( .A(n14517), .B(n14485), .Z(n14518) );
  XOR U16923 ( .A(n14525), .B(n14526), .Z(n14485) );
  AND U16924 ( .A(n310), .B(n14527), .Z(n14525) );
  XOR U16925 ( .A(n14528), .B(n14526), .Z(n14527) );
  XNOR U16926 ( .A(n14529), .B(n14530), .Z(n14517) );
  NAND U16927 ( .A(n14531), .B(n14532), .Z(n14530) );
  XOR U16928 ( .A(n14533), .B(n14509), .Z(n14532) );
  XOR U16929 ( .A(n14523), .B(n14524), .Z(n14509) );
  XOR U16930 ( .A(n14534), .B(n14535), .Z(n14524) );
  ANDN U16931 ( .B(n14536), .A(n14537), .Z(n14534) );
  XOR U16932 ( .A(n14535), .B(n14538), .Z(n14536) );
  XOR U16933 ( .A(n14539), .B(n14540), .Z(n14523) );
  XOR U16934 ( .A(n14541), .B(n14542), .Z(n14540) );
  ANDN U16935 ( .B(n14543), .A(n14544), .Z(n14541) );
  XOR U16936 ( .A(n14545), .B(n14542), .Z(n14543) );
  IV U16937 ( .A(n14521), .Z(n14539) );
  XOR U16938 ( .A(n14546), .B(n14547), .Z(n14521) );
  ANDN U16939 ( .B(n14548), .A(n14549), .Z(n14546) );
  XOR U16940 ( .A(n14547), .B(n14550), .Z(n14548) );
  IV U16941 ( .A(n14529), .Z(n14533) );
  XOR U16942 ( .A(n14529), .B(n14511), .Z(n14531) );
  XOR U16943 ( .A(n14551), .B(n14552), .Z(n14511) );
  AND U16944 ( .A(n310), .B(n14553), .Z(n14551) );
  XOR U16945 ( .A(n14554), .B(n14552), .Z(n14553) );
  NANDN U16946 ( .A(n14513), .B(n14515), .Z(n14529) );
  XOR U16947 ( .A(n14555), .B(n14556), .Z(n14515) );
  AND U16948 ( .A(n310), .B(n14557), .Z(n14555) );
  XOR U16949 ( .A(n14556), .B(n14558), .Z(n14557) );
  XOR U16950 ( .A(n14559), .B(n14560), .Z(n310) );
  AND U16951 ( .A(n14561), .B(n14562), .Z(n14559) );
  XNOR U16952 ( .A(n14560), .B(n14526), .Z(n14562) );
  XNOR U16953 ( .A(n14563), .B(n14564), .Z(n14526) );
  ANDN U16954 ( .B(n14565), .A(n14566), .Z(n14563) );
  XOR U16955 ( .A(n14564), .B(n14567), .Z(n14565) );
  XOR U16956 ( .A(n14560), .B(n14528), .Z(n14561) );
  XOR U16957 ( .A(n14568), .B(n14569), .Z(n14528) );
  AND U16958 ( .A(n314), .B(n14570), .Z(n14568) );
  XOR U16959 ( .A(n14571), .B(n14569), .Z(n14570) );
  XNOR U16960 ( .A(n14572), .B(n14573), .Z(n14560) );
  NAND U16961 ( .A(n14574), .B(n14575), .Z(n14573) );
  XOR U16962 ( .A(n14576), .B(n14552), .Z(n14575) );
  XOR U16963 ( .A(n14566), .B(n14567), .Z(n14552) );
  XOR U16964 ( .A(n14577), .B(n14578), .Z(n14567) );
  ANDN U16965 ( .B(n14579), .A(n14580), .Z(n14577) );
  XOR U16966 ( .A(n14578), .B(n14581), .Z(n14579) );
  XOR U16967 ( .A(n14582), .B(n14583), .Z(n14566) );
  XOR U16968 ( .A(n14584), .B(n14585), .Z(n14583) );
  ANDN U16969 ( .B(n14586), .A(n14587), .Z(n14584) );
  XOR U16970 ( .A(n14588), .B(n14585), .Z(n14586) );
  IV U16971 ( .A(n14564), .Z(n14582) );
  XOR U16972 ( .A(n14589), .B(n14590), .Z(n14564) );
  ANDN U16973 ( .B(n14591), .A(n14592), .Z(n14589) );
  XOR U16974 ( .A(n14590), .B(n14593), .Z(n14591) );
  IV U16975 ( .A(n14572), .Z(n14576) );
  XOR U16976 ( .A(n14572), .B(n14554), .Z(n14574) );
  XOR U16977 ( .A(n14594), .B(n14595), .Z(n14554) );
  AND U16978 ( .A(n314), .B(n14596), .Z(n14594) );
  XOR U16979 ( .A(n14597), .B(n14595), .Z(n14596) );
  NANDN U16980 ( .A(n14556), .B(n14558), .Z(n14572) );
  XOR U16981 ( .A(n14598), .B(n14599), .Z(n14558) );
  AND U16982 ( .A(n314), .B(n14600), .Z(n14598) );
  XOR U16983 ( .A(n14599), .B(n14601), .Z(n14600) );
  XOR U16984 ( .A(n14602), .B(n14603), .Z(n314) );
  AND U16985 ( .A(n14604), .B(n14605), .Z(n14602) );
  XNOR U16986 ( .A(n14603), .B(n14569), .Z(n14605) );
  XNOR U16987 ( .A(n14606), .B(n14607), .Z(n14569) );
  ANDN U16988 ( .B(n14608), .A(n14609), .Z(n14606) );
  XOR U16989 ( .A(n14607), .B(n14610), .Z(n14608) );
  XOR U16990 ( .A(n14603), .B(n14571), .Z(n14604) );
  XOR U16991 ( .A(n14611), .B(n14612), .Z(n14571) );
  AND U16992 ( .A(n318), .B(n14613), .Z(n14611) );
  XOR U16993 ( .A(n14614), .B(n14612), .Z(n14613) );
  XNOR U16994 ( .A(n14615), .B(n14616), .Z(n14603) );
  NAND U16995 ( .A(n14617), .B(n14618), .Z(n14616) );
  XOR U16996 ( .A(n14619), .B(n14595), .Z(n14618) );
  XOR U16997 ( .A(n14609), .B(n14610), .Z(n14595) );
  XOR U16998 ( .A(n14620), .B(n14621), .Z(n14610) );
  ANDN U16999 ( .B(n14622), .A(n14623), .Z(n14620) );
  XOR U17000 ( .A(n14621), .B(n14624), .Z(n14622) );
  XOR U17001 ( .A(n14625), .B(n14626), .Z(n14609) );
  XOR U17002 ( .A(n14627), .B(n14628), .Z(n14626) );
  ANDN U17003 ( .B(n14629), .A(n14630), .Z(n14627) );
  XOR U17004 ( .A(n14631), .B(n14628), .Z(n14629) );
  IV U17005 ( .A(n14607), .Z(n14625) );
  XOR U17006 ( .A(n14632), .B(n14633), .Z(n14607) );
  ANDN U17007 ( .B(n14634), .A(n14635), .Z(n14632) );
  XOR U17008 ( .A(n14633), .B(n14636), .Z(n14634) );
  IV U17009 ( .A(n14615), .Z(n14619) );
  XOR U17010 ( .A(n14615), .B(n14597), .Z(n14617) );
  XOR U17011 ( .A(n14637), .B(n14638), .Z(n14597) );
  AND U17012 ( .A(n318), .B(n14639), .Z(n14637) );
  XOR U17013 ( .A(n14640), .B(n14638), .Z(n14639) );
  NANDN U17014 ( .A(n14599), .B(n14601), .Z(n14615) );
  XOR U17015 ( .A(n14641), .B(n14642), .Z(n14601) );
  AND U17016 ( .A(n318), .B(n14643), .Z(n14641) );
  XOR U17017 ( .A(n14642), .B(n14644), .Z(n14643) );
  XOR U17018 ( .A(n14645), .B(n14646), .Z(n318) );
  AND U17019 ( .A(n14647), .B(n14648), .Z(n14645) );
  XNOR U17020 ( .A(n14646), .B(n14612), .Z(n14648) );
  XNOR U17021 ( .A(n14649), .B(n14650), .Z(n14612) );
  ANDN U17022 ( .B(n14651), .A(n14652), .Z(n14649) );
  XOR U17023 ( .A(n14650), .B(n14653), .Z(n14651) );
  XOR U17024 ( .A(n14646), .B(n14614), .Z(n14647) );
  XOR U17025 ( .A(n14654), .B(n14655), .Z(n14614) );
  AND U17026 ( .A(n322), .B(n14656), .Z(n14654) );
  XOR U17027 ( .A(n14657), .B(n14655), .Z(n14656) );
  XNOR U17028 ( .A(n14658), .B(n14659), .Z(n14646) );
  NAND U17029 ( .A(n14660), .B(n14661), .Z(n14659) );
  XOR U17030 ( .A(n14662), .B(n14638), .Z(n14661) );
  XOR U17031 ( .A(n14652), .B(n14653), .Z(n14638) );
  XOR U17032 ( .A(n14663), .B(n14664), .Z(n14653) );
  ANDN U17033 ( .B(n14665), .A(n14666), .Z(n14663) );
  XOR U17034 ( .A(n14664), .B(n14667), .Z(n14665) );
  XOR U17035 ( .A(n14668), .B(n14669), .Z(n14652) );
  XOR U17036 ( .A(n14670), .B(n14671), .Z(n14669) );
  ANDN U17037 ( .B(n14672), .A(n14673), .Z(n14670) );
  XOR U17038 ( .A(n14674), .B(n14671), .Z(n14672) );
  IV U17039 ( .A(n14650), .Z(n14668) );
  XOR U17040 ( .A(n14675), .B(n14676), .Z(n14650) );
  ANDN U17041 ( .B(n14677), .A(n14678), .Z(n14675) );
  XOR U17042 ( .A(n14676), .B(n14679), .Z(n14677) );
  IV U17043 ( .A(n14658), .Z(n14662) );
  XOR U17044 ( .A(n14658), .B(n14640), .Z(n14660) );
  XOR U17045 ( .A(n14680), .B(n14681), .Z(n14640) );
  AND U17046 ( .A(n322), .B(n14682), .Z(n14680) );
  XOR U17047 ( .A(n14683), .B(n14681), .Z(n14682) );
  NANDN U17048 ( .A(n14642), .B(n14644), .Z(n14658) );
  XOR U17049 ( .A(n14684), .B(n14685), .Z(n14644) );
  AND U17050 ( .A(n322), .B(n14686), .Z(n14684) );
  XOR U17051 ( .A(n14685), .B(n14687), .Z(n14686) );
  XOR U17052 ( .A(n14688), .B(n14689), .Z(n322) );
  AND U17053 ( .A(n14690), .B(n14691), .Z(n14688) );
  XNOR U17054 ( .A(n14689), .B(n14655), .Z(n14691) );
  XNOR U17055 ( .A(n14692), .B(n14693), .Z(n14655) );
  ANDN U17056 ( .B(n14694), .A(n14695), .Z(n14692) );
  XOR U17057 ( .A(n14693), .B(n14696), .Z(n14694) );
  XOR U17058 ( .A(n14689), .B(n14657), .Z(n14690) );
  XOR U17059 ( .A(n14697), .B(n14698), .Z(n14657) );
  AND U17060 ( .A(n326), .B(n14699), .Z(n14697) );
  XOR U17061 ( .A(n14700), .B(n14698), .Z(n14699) );
  XNOR U17062 ( .A(n14701), .B(n14702), .Z(n14689) );
  NAND U17063 ( .A(n14703), .B(n14704), .Z(n14702) );
  XOR U17064 ( .A(n14705), .B(n14681), .Z(n14704) );
  XOR U17065 ( .A(n14695), .B(n14696), .Z(n14681) );
  XOR U17066 ( .A(n14706), .B(n14707), .Z(n14696) );
  ANDN U17067 ( .B(n14708), .A(n14709), .Z(n14706) );
  XOR U17068 ( .A(n14707), .B(n14710), .Z(n14708) );
  XOR U17069 ( .A(n14711), .B(n14712), .Z(n14695) );
  XOR U17070 ( .A(n14713), .B(n14714), .Z(n14712) );
  ANDN U17071 ( .B(n14715), .A(n14716), .Z(n14713) );
  XOR U17072 ( .A(n14717), .B(n14714), .Z(n14715) );
  IV U17073 ( .A(n14693), .Z(n14711) );
  XOR U17074 ( .A(n14718), .B(n14719), .Z(n14693) );
  ANDN U17075 ( .B(n14720), .A(n14721), .Z(n14718) );
  XOR U17076 ( .A(n14719), .B(n14722), .Z(n14720) );
  IV U17077 ( .A(n14701), .Z(n14705) );
  XOR U17078 ( .A(n14701), .B(n14683), .Z(n14703) );
  XOR U17079 ( .A(n14723), .B(n14724), .Z(n14683) );
  AND U17080 ( .A(n326), .B(n14725), .Z(n14723) );
  XOR U17081 ( .A(n14726), .B(n14724), .Z(n14725) );
  NANDN U17082 ( .A(n14685), .B(n14687), .Z(n14701) );
  XOR U17083 ( .A(n14727), .B(n14728), .Z(n14687) );
  AND U17084 ( .A(n326), .B(n14729), .Z(n14727) );
  XOR U17085 ( .A(n14728), .B(n14730), .Z(n14729) );
  XOR U17086 ( .A(n14731), .B(n14732), .Z(n326) );
  AND U17087 ( .A(n14733), .B(n14734), .Z(n14731) );
  XNOR U17088 ( .A(n14732), .B(n14698), .Z(n14734) );
  XNOR U17089 ( .A(n14735), .B(n14736), .Z(n14698) );
  ANDN U17090 ( .B(n14737), .A(n14738), .Z(n14735) );
  XOR U17091 ( .A(n14736), .B(n14739), .Z(n14737) );
  XOR U17092 ( .A(n14732), .B(n14700), .Z(n14733) );
  XOR U17093 ( .A(n14740), .B(n14741), .Z(n14700) );
  AND U17094 ( .A(n330), .B(n14742), .Z(n14740) );
  XOR U17095 ( .A(n14743), .B(n14741), .Z(n14742) );
  XNOR U17096 ( .A(n14744), .B(n14745), .Z(n14732) );
  NAND U17097 ( .A(n14746), .B(n14747), .Z(n14745) );
  XOR U17098 ( .A(n14748), .B(n14724), .Z(n14747) );
  XOR U17099 ( .A(n14738), .B(n14739), .Z(n14724) );
  XOR U17100 ( .A(n14749), .B(n14750), .Z(n14739) );
  ANDN U17101 ( .B(n14751), .A(n14752), .Z(n14749) );
  XOR U17102 ( .A(n14750), .B(n14753), .Z(n14751) );
  XOR U17103 ( .A(n14754), .B(n14755), .Z(n14738) );
  XOR U17104 ( .A(n14756), .B(n14757), .Z(n14755) );
  ANDN U17105 ( .B(n14758), .A(n14759), .Z(n14756) );
  XOR U17106 ( .A(n14760), .B(n14757), .Z(n14758) );
  IV U17107 ( .A(n14736), .Z(n14754) );
  XOR U17108 ( .A(n14761), .B(n14762), .Z(n14736) );
  ANDN U17109 ( .B(n14763), .A(n14764), .Z(n14761) );
  XOR U17110 ( .A(n14762), .B(n14765), .Z(n14763) );
  IV U17111 ( .A(n14744), .Z(n14748) );
  XOR U17112 ( .A(n14744), .B(n14726), .Z(n14746) );
  XOR U17113 ( .A(n14766), .B(n14767), .Z(n14726) );
  AND U17114 ( .A(n330), .B(n14768), .Z(n14766) );
  XOR U17115 ( .A(n14769), .B(n14767), .Z(n14768) );
  NANDN U17116 ( .A(n14728), .B(n14730), .Z(n14744) );
  XOR U17117 ( .A(n14770), .B(n14771), .Z(n14730) );
  AND U17118 ( .A(n330), .B(n14772), .Z(n14770) );
  XOR U17119 ( .A(n14771), .B(n14773), .Z(n14772) );
  XOR U17120 ( .A(n14774), .B(n14775), .Z(n330) );
  AND U17121 ( .A(n14776), .B(n14777), .Z(n14774) );
  XNOR U17122 ( .A(n14775), .B(n14741), .Z(n14777) );
  XNOR U17123 ( .A(n14778), .B(n14779), .Z(n14741) );
  ANDN U17124 ( .B(n14780), .A(n14781), .Z(n14778) );
  XOR U17125 ( .A(n14779), .B(n14782), .Z(n14780) );
  XOR U17126 ( .A(n14775), .B(n14743), .Z(n14776) );
  XOR U17127 ( .A(n14783), .B(n14784), .Z(n14743) );
  AND U17128 ( .A(n334), .B(n14785), .Z(n14783) );
  XOR U17129 ( .A(n14786), .B(n14784), .Z(n14785) );
  XNOR U17130 ( .A(n14787), .B(n14788), .Z(n14775) );
  NAND U17131 ( .A(n14789), .B(n14790), .Z(n14788) );
  XOR U17132 ( .A(n14791), .B(n14767), .Z(n14790) );
  XOR U17133 ( .A(n14781), .B(n14782), .Z(n14767) );
  XOR U17134 ( .A(n14792), .B(n14793), .Z(n14782) );
  ANDN U17135 ( .B(n14794), .A(n14795), .Z(n14792) );
  XOR U17136 ( .A(n14793), .B(n14796), .Z(n14794) );
  XOR U17137 ( .A(n14797), .B(n14798), .Z(n14781) );
  XOR U17138 ( .A(n14799), .B(n14800), .Z(n14798) );
  ANDN U17139 ( .B(n14801), .A(n14802), .Z(n14799) );
  XOR U17140 ( .A(n14803), .B(n14800), .Z(n14801) );
  IV U17141 ( .A(n14779), .Z(n14797) );
  XOR U17142 ( .A(n14804), .B(n14805), .Z(n14779) );
  ANDN U17143 ( .B(n14806), .A(n14807), .Z(n14804) );
  XOR U17144 ( .A(n14805), .B(n14808), .Z(n14806) );
  IV U17145 ( .A(n14787), .Z(n14791) );
  XOR U17146 ( .A(n14787), .B(n14769), .Z(n14789) );
  XOR U17147 ( .A(n14809), .B(n14810), .Z(n14769) );
  AND U17148 ( .A(n334), .B(n14811), .Z(n14809) );
  XOR U17149 ( .A(n14812), .B(n14810), .Z(n14811) );
  NANDN U17150 ( .A(n14771), .B(n14773), .Z(n14787) );
  XOR U17151 ( .A(n14813), .B(n14814), .Z(n14773) );
  AND U17152 ( .A(n334), .B(n14815), .Z(n14813) );
  XOR U17153 ( .A(n14814), .B(n14816), .Z(n14815) );
  XOR U17154 ( .A(n14817), .B(n14818), .Z(n334) );
  AND U17155 ( .A(n14819), .B(n14820), .Z(n14817) );
  XNOR U17156 ( .A(n14818), .B(n14784), .Z(n14820) );
  XNOR U17157 ( .A(n14821), .B(n14822), .Z(n14784) );
  ANDN U17158 ( .B(n14823), .A(n14824), .Z(n14821) );
  XOR U17159 ( .A(n14822), .B(n14825), .Z(n14823) );
  XOR U17160 ( .A(n14818), .B(n14786), .Z(n14819) );
  XOR U17161 ( .A(n14826), .B(n14827), .Z(n14786) );
  AND U17162 ( .A(n338), .B(n14828), .Z(n14826) );
  XOR U17163 ( .A(n14829), .B(n14827), .Z(n14828) );
  XNOR U17164 ( .A(n14830), .B(n14831), .Z(n14818) );
  NAND U17165 ( .A(n14832), .B(n14833), .Z(n14831) );
  XOR U17166 ( .A(n14834), .B(n14810), .Z(n14833) );
  XOR U17167 ( .A(n14824), .B(n14825), .Z(n14810) );
  XOR U17168 ( .A(n14835), .B(n14836), .Z(n14825) );
  ANDN U17169 ( .B(n14837), .A(n14838), .Z(n14835) );
  XOR U17170 ( .A(n14836), .B(n14839), .Z(n14837) );
  XOR U17171 ( .A(n14840), .B(n14841), .Z(n14824) );
  XOR U17172 ( .A(n14842), .B(n14843), .Z(n14841) );
  ANDN U17173 ( .B(n14844), .A(n14845), .Z(n14842) );
  XOR U17174 ( .A(n14846), .B(n14843), .Z(n14844) );
  IV U17175 ( .A(n14822), .Z(n14840) );
  XOR U17176 ( .A(n14847), .B(n14848), .Z(n14822) );
  ANDN U17177 ( .B(n14849), .A(n14850), .Z(n14847) );
  XOR U17178 ( .A(n14848), .B(n14851), .Z(n14849) );
  IV U17179 ( .A(n14830), .Z(n14834) );
  XOR U17180 ( .A(n14830), .B(n14812), .Z(n14832) );
  XOR U17181 ( .A(n14852), .B(n14853), .Z(n14812) );
  AND U17182 ( .A(n338), .B(n14854), .Z(n14852) );
  XOR U17183 ( .A(n14855), .B(n14853), .Z(n14854) );
  NANDN U17184 ( .A(n14814), .B(n14816), .Z(n14830) );
  XOR U17185 ( .A(n14856), .B(n14857), .Z(n14816) );
  AND U17186 ( .A(n338), .B(n14858), .Z(n14856) );
  XOR U17187 ( .A(n14857), .B(n14859), .Z(n14858) );
  XOR U17188 ( .A(n14860), .B(n14861), .Z(n338) );
  AND U17189 ( .A(n14862), .B(n14863), .Z(n14860) );
  XNOR U17190 ( .A(n14861), .B(n14827), .Z(n14863) );
  XNOR U17191 ( .A(n14864), .B(n14865), .Z(n14827) );
  ANDN U17192 ( .B(n14866), .A(n14867), .Z(n14864) );
  XOR U17193 ( .A(n14865), .B(n14868), .Z(n14866) );
  XOR U17194 ( .A(n14861), .B(n14829), .Z(n14862) );
  XOR U17195 ( .A(n14869), .B(n14870), .Z(n14829) );
  AND U17196 ( .A(n342), .B(n14871), .Z(n14869) );
  XOR U17197 ( .A(n14872), .B(n14870), .Z(n14871) );
  XNOR U17198 ( .A(n14873), .B(n14874), .Z(n14861) );
  NAND U17199 ( .A(n14875), .B(n14876), .Z(n14874) );
  XOR U17200 ( .A(n14877), .B(n14853), .Z(n14876) );
  XOR U17201 ( .A(n14867), .B(n14868), .Z(n14853) );
  XOR U17202 ( .A(n14878), .B(n14879), .Z(n14868) );
  ANDN U17203 ( .B(n14880), .A(n14881), .Z(n14878) );
  XOR U17204 ( .A(n14879), .B(n14882), .Z(n14880) );
  XOR U17205 ( .A(n14883), .B(n14884), .Z(n14867) );
  XOR U17206 ( .A(n14885), .B(n14886), .Z(n14884) );
  ANDN U17207 ( .B(n14887), .A(n14888), .Z(n14885) );
  XOR U17208 ( .A(n14889), .B(n14886), .Z(n14887) );
  IV U17209 ( .A(n14865), .Z(n14883) );
  XOR U17210 ( .A(n14890), .B(n14891), .Z(n14865) );
  ANDN U17211 ( .B(n14892), .A(n14893), .Z(n14890) );
  XOR U17212 ( .A(n14891), .B(n14894), .Z(n14892) );
  IV U17213 ( .A(n14873), .Z(n14877) );
  XOR U17214 ( .A(n14873), .B(n14855), .Z(n14875) );
  XOR U17215 ( .A(n14895), .B(n14896), .Z(n14855) );
  AND U17216 ( .A(n342), .B(n14897), .Z(n14895) );
  XOR U17217 ( .A(n14898), .B(n14896), .Z(n14897) );
  NANDN U17218 ( .A(n14857), .B(n14859), .Z(n14873) );
  XOR U17219 ( .A(n14899), .B(n14900), .Z(n14859) );
  AND U17220 ( .A(n342), .B(n14901), .Z(n14899) );
  XOR U17221 ( .A(n14900), .B(n14902), .Z(n14901) );
  XOR U17222 ( .A(n14903), .B(n14904), .Z(n342) );
  AND U17223 ( .A(n14905), .B(n14906), .Z(n14903) );
  XNOR U17224 ( .A(n14904), .B(n14870), .Z(n14906) );
  XNOR U17225 ( .A(n14907), .B(n14908), .Z(n14870) );
  ANDN U17226 ( .B(n14909), .A(n14910), .Z(n14907) );
  XOR U17227 ( .A(n14908), .B(n14911), .Z(n14909) );
  XOR U17228 ( .A(n14904), .B(n14872), .Z(n14905) );
  XOR U17229 ( .A(n14912), .B(n14913), .Z(n14872) );
  AND U17230 ( .A(n346), .B(n14914), .Z(n14912) );
  XOR U17231 ( .A(n14915), .B(n14913), .Z(n14914) );
  XNOR U17232 ( .A(n14916), .B(n14917), .Z(n14904) );
  NAND U17233 ( .A(n14918), .B(n14919), .Z(n14917) );
  XOR U17234 ( .A(n14920), .B(n14896), .Z(n14919) );
  XOR U17235 ( .A(n14910), .B(n14911), .Z(n14896) );
  XOR U17236 ( .A(n14921), .B(n14922), .Z(n14911) );
  ANDN U17237 ( .B(n14923), .A(n14924), .Z(n14921) );
  XOR U17238 ( .A(n14922), .B(n14925), .Z(n14923) );
  XOR U17239 ( .A(n14926), .B(n14927), .Z(n14910) );
  XOR U17240 ( .A(n14928), .B(n14929), .Z(n14927) );
  ANDN U17241 ( .B(n14930), .A(n14931), .Z(n14928) );
  XOR U17242 ( .A(n14932), .B(n14929), .Z(n14930) );
  IV U17243 ( .A(n14908), .Z(n14926) );
  XOR U17244 ( .A(n14933), .B(n14934), .Z(n14908) );
  ANDN U17245 ( .B(n14935), .A(n14936), .Z(n14933) );
  XOR U17246 ( .A(n14934), .B(n14937), .Z(n14935) );
  IV U17247 ( .A(n14916), .Z(n14920) );
  XOR U17248 ( .A(n14916), .B(n14898), .Z(n14918) );
  XOR U17249 ( .A(n14938), .B(n14939), .Z(n14898) );
  AND U17250 ( .A(n346), .B(n14940), .Z(n14938) );
  XOR U17251 ( .A(n14941), .B(n14939), .Z(n14940) );
  NANDN U17252 ( .A(n14900), .B(n14902), .Z(n14916) );
  XOR U17253 ( .A(n14942), .B(n14943), .Z(n14902) );
  AND U17254 ( .A(n346), .B(n14944), .Z(n14942) );
  XOR U17255 ( .A(n14943), .B(n14945), .Z(n14944) );
  XOR U17256 ( .A(n14946), .B(n14947), .Z(n346) );
  AND U17257 ( .A(n14948), .B(n14949), .Z(n14946) );
  XNOR U17258 ( .A(n14947), .B(n14913), .Z(n14949) );
  XNOR U17259 ( .A(n14950), .B(n14951), .Z(n14913) );
  ANDN U17260 ( .B(n14952), .A(n14953), .Z(n14950) );
  XOR U17261 ( .A(n14951), .B(n14954), .Z(n14952) );
  XOR U17262 ( .A(n14947), .B(n14915), .Z(n14948) );
  XOR U17263 ( .A(n14955), .B(n14956), .Z(n14915) );
  AND U17264 ( .A(n350), .B(n14957), .Z(n14955) );
  XOR U17265 ( .A(n14958), .B(n14956), .Z(n14957) );
  XNOR U17266 ( .A(n14959), .B(n14960), .Z(n14947) );
  NAND U17267 ( .A(n14961), .B(n14962), .Z(n14960) );
  XOR U17268 ( .A(n14963), .B(n14939), .Z(n14962) );
  XOR U17269 ( .A(n14953), .B(n14954), .Z(n14939) );
  XOR U17270 ( .A(n14964), .B(n14965), .Z(n14954) );
  ANDN U17271 ( .B(n14966), .A(n14967), .Z(n14964) );
  XOR U17272 ( .A(n14965), .B(n14968), .Z(n14966) );
  XOR U17273 ( .A(n14969), .B(n14970), .Z(n14953) );
  XOR U17274 ( .A(n14971), .B(n14972), .Z(n14970) );
  ANDN U17275 ( .B(n14973), .A(n14974), .Z(n14971) );
  XOR U17276 ( .A(n14975), .B(n14972), .Z(n14973) );
  IV U17277 ( .A(n14951), .Z(n14969) );
  XOR U17278 ( .A(n14976), .B(n14977), .Z(n14951) );
  ANDN U17279 ( .B(n14978), .A(n14979), .Z(n14976) );
  XOR U17280 ( .A(n14977), .B(n14980), .Z(n14978) );
  IV U17281 ( .A(n14959), .Z(n14963) );
  XOR U17282 ( .A(n14959), .B(n14941), .Z(n14961) );
  XOR U17283 ( .A(n14981), .B(n14982), .Z(n14941) );
  AND U17284 ( .A(n350), .B(n14983), .Z(n14981) );
  XOR U17285 ( .A(n14984), .B(n14982), .Z(n14983) );
  NANDN U17286 ( .A(n14943), .B(n14945), .Z(n14959) );
  XOR U17287 ( .A(n14985), .B(n14986), .Z(n14945) );
  AND U17288 ( .A(n350), .B(n14987), .Z(n14985) );
  XOR U17289 ( .A(n14986), .B(n14988), .Z(n14987) );
  XOR U17290 ( .A(n14989), .B(n14990), .Z(n350) );
  AND U17291 ( .A(n14991), .B(n14992), .Z(n14989) );
  XNOR U17292 ( .A(n14990), .B(n14956), .Z(n14992) );
  XNOR U17293 ( .A(n14993), .B(n14994), .Z(n14956) );
  ANDN U17294 ( .B(n14995), .A(n14996), .Z(n14993) );
  XOR U17295 ( .A(n14994), .B(n14997), .Z(n14995) );
  XOR U17296 ( .A(n14990), .B(n14958), .Z(n14991) );
  XOR U17297 ( .A(n14998), .B(n14999), .Z(n14958) );
  AND U17298 ( .A(n354), .B(n15000), .Z(n14998) );
  XOR U17299 ( .A(n15001), .B(n14999), .Z(n15000) );
  XNOR U17300 ( .A(n15002), .B(n15003), .Z(n14990) );
  NAND U17301 ( .A(n15004), .B(n15005), .Z(n15003) );
  XOR U17302 ( .A(n15006), .B(n14982), .Z(n15005) );
  XOR U17303 ( .A(n14996), .B(n14997), .Z(n14982) );
  XOR U17304 ( .A(n15007), .B(n15008), .Z(n14997) );
  ANDN U17305 ( .B(n15009), .A(n15010), .Z(n15007) );
  XOR U17306 ( .A(n15008), .B(n15011), .Z(n15009) );
  XOR U17307 ( .A(n15012), .B(n15013), .Z(n14996) );
  XOR U17308 ( .A(n15014), .B(n15015), .Z(n15013) );
  ANDN U17309 ( .B(n15016), .A(n15017), .Z(n15014) );
  XOR U17310 ( .A(n15018), .B(n15015), .Z(n15016) );
  IV U17311 ( .A(n14994), .Z(n15012) );
  XOR U17312 ( .A(n15019), .B(n15020), .Z(n14994) );
  ANDN U17313 ( .B(n15021), .A(n15022), .Z(n15019) );
  XOR U17314 ( .A(n15020), .B(n15023), .Z(n15021) );
  IV U17315 ( .A(n15002), .Z(n15006) );
  XOR U17316 ( .A(n15002), .B(n14984), .Z(n15004) );
  XOR U17317 ( .A(n15024), .B(n15025), .Z(n14984) );
  AND U17318 ( .A(n354), .B(n15026), .Z(n15024) );
  XOR U17319 ( .A(n15027), .B(n15025), .Z(n15026) );
  NANDN U17320 ( .A(n14986), .B(n14988), .Z(n15002) );
  XOR U17321 ( .A(n15028), .B(n15029), .Z(n14988) );
  AND U17322 ( .A(n354), .B(n15030), .Z(n15028) );
  XOR U17323 ( .A(n15029), .B(n15031), .Z(n15030) );
  XOR U17324 ( .A(n15032), .B(n15033), .Z(n354) );
  AND U17325 ( .A(n15034), .B(n15035), .Z(n15032) );
  XNOR U17326 ( .A(n15033), .B(n14999), .Z(n15035) );
  XNOR U17327 ( .A(n15036), .B(n15037), .Z(n14999) );
  ANDN U17328 ( .B(n15038), .A(n15039), .Z(n15036) );
  XOR U17329 ( .A(n15037), .B(n15040), .Z(n15038) );
  XOR U17330 ( .A(n15033), .B(n15001), .Z(n15034) );
  XOR U17331 ( .A(n15041), .B(n15042), .Z(n15001) );
  AND U17332 ( .A(n358), .B(n15043), .Z(n15041) );
  XOR U17333 ( .A(n15044), .B(n15042), .Z(n15043) );
  XNOR U17334 ( .A(n15045), .B(n15046), .Z(n15033) );
  NAND U17335 ( .A(n15047), .B(n15048), .Z(n15046) );
  XOR U17336 ( .A(n15049), .B(n15025), .Z(n15048) );
  XOR U17337 ( .A(n15039), .B(n15040), .Z(n15025) );
  XOR U17338 ( .A(n15050), .B(n15051), .Z(n15040) );
  ANDN U17339 ( .B(n15052), .A(n15053), .Z(n15050) );
  XOR U17340 ( .A(n15051), .B(n15054), .Z(n15052) );
  XOR U17341 ( .A(n15055), .B(n15056), .Z(n15039) );
  XOR U17342 ( .A(n15057), .B(n15058), .Z(n15056) );
  ANDN U17343 ( .B(n15059), .A(n15060), .Z(n15057) );
  XOR U17344 ( .A(n15061), .B(n15058), .Z(n15059) );
  IV U17345 ( .A(n15037), .Z(n15055) );
  XOR U17346 ( .A(n15062), .B(n15063), .Z(n15037) );
  ANDN U17347 ( .B(n15064), .A(n15065), .Z(n15062) );
  XOR U17348 ( .A(n15063), .B(n15066), .Z(n15064) );
  IV U17349 ( .A(n15045), .Z(n15049) );
  XOR U17350 ( .A(n15045), .B(n15027), .Z(n15047) );
  XOR U17351 ( .A(n15067), .B(n15068), .Z(n15027) );
  AND U17352 ( .A(n358), .B(n15069), .Z(n15067) );
  XOR U17353 ( .A(n15070), .B(n15068), .Z(n15069) );
  NANDN U17354 ( .A(n15029), .B(n15031), .Z(n15045) );
  XOR U17355 ( .A(n15071), .B(n15072), .Z(n15031) );
  AND U17356 ( .A(n358), .B(n15073), .Z(n15071) );
  XOR U17357 ( .A(n15072), .B(n15074), .Z(n15073) );
  XOR U17358 ( .A(n15075), .B(n15076), .Z(n358) );
  AND U17359 ( .A(n15077), .B(n15078), .Z(n15075) );
  XNOR U17360 ( .A(n15076), .B(n15042), .Z(n15078) );
  XNOR U17361 ( .A(n15079), .B(n15080), .Z(n15042) );
  ANDN U17362 ( .B(n15081), .A(n15082), .Z(n15079) );
  XOR U17363 ( .A(n15080), .B(n15083), .Z(n15081) );
  XOR U17364 ( .A(n15076), .B(n15044), .Z(n15077) );
  XOR U17365 ( .A(n15084), .B(n15085), .Z(n15044) );
  AND U17366 ( .A(n362), .B(n15086), .Z(n15084) );
  XOR U17367 ( .A(n15087), .B(n15085), .Z(n15086) );
  XNOR U17368 ( .A(n15088), .B(n15089), .Z(n15076) );
  NAND U17369 ( .A(n15090), .B(n15091), .Z(n15089) );
  XOR U17370 ( .A(n15092), .B(n15068), .Z(n15091) );
  XOR U17371 ( .A(n15082), .B(n15083), .Z(n15068) );
  XOR U17372 ( .A(n15093), .B(n15094), .Z(n15083) );
  ANDN U17373 ( .B(n15095), .A(n15096), .Z(n15093) );
  XOR U17374 ( .A(n15094), .B(n15097), .Z(n15095) );
  XOR U17375 ( .A(n15098), .B(n15099), .Z(n15082) );
  XOR U17376 ( .A(n15100), .B(n15101), .Z(n15099) );
  ANDN U17377 ( .B(n15102), .A(n15103), .Z(n15100) );
  XOR U17378 ( .A(n15104), .B(n15101), .Z(n15102) );
  IV U17379 ( .A(n15080), .Z(n15098) );
  XOR U17380 ( .A(n15105), .B(n15106), .Z(n15080) );
  ANDN U17381 ( .B(n15107), .A(n15108), .Z(n15105) );
  XOR U17382 ( .A(n15106), .B(n15109), .Z(n15107) );
  IV U17383 ( .A(n15088), .Z(n15092) );
  XOR U17384 ( .A(n15088), .B(n15070), .Z(n15090) );
  XOR U17385 ( .A(n15110), .B(n15111), .Z(n15070) );
  AND U17386 ( .A(n362), .B(n15112), .Z(n15110) );
  XOR U17387 ( .A(n15113), .B(n15111), .Z(n15112) );
  NANDN U17388 ( .A(n15072), .B(n15074), .Z(n15088) );
  XOR U17389 ( .A(n15114), .B(n15115), .Z(n15074) );
  AND U17390 ( .A(n362), .B(n15116), .Z(n15114) );
  XOR U17391 ( .A(n15115), .B(n15117), .Z(n15116) );
  XOR U17392 ( .A(n15118), .B(n15119), .Z(n362) );
  AND U17393 ( .A(n15120), .B(n15121), .Z(n15118) );
  XNOR U17394 ( .A(n15119), .B(n15085), .Z(n15121) );
  XNOR U17395 ( .A(n15122), .B(n15123), .Z(n15085) );
  ANDN U17396 ( .B(n15124), .A(n15125), .Z(n15122) );
  XOR U17397 ( .A(n15123), .B(n15126), .Z(n15124) );
  XOR U17398 ( .A(n15119), .B(n15087), .Z(n15120) );
  XOR U17399 ( .A(n15127), .B(n15128), .Z(n15087) );
  AND U17400 ( .A(n366), .B(n15129), .Z(n15127) );
  XOR U17401 ( .A(n15130), .B(n15128), .Z(n15129) );
  XNOR U17402 ( .A(n15131), .B(n15132), .Z(n15119) );
  NAND U17403 ( .A(n15133), .B(n15134), .Z(n15132) );
  XOR U17404 ( .A(n15135), .B(n15111), .Z(n15134) );
  XOR U17405 ( .A(n15125), .B(n15126), .Z(n15111) );
  XOR U17406 ( .A(n15136), .B(n15137), .Z(n15126) );
  ANDN U17407 ( .B(n15138), .A(n15139), .Z(n15136) );
  XOR U17408 ( .A(n15137), .B(n15140), .Z(n15138) );
  XOR U17409 ( .A(n15141), .B(n15142), .Z(n15125) );
  XOR U17410 ( .A(n15143), .B(n15144), .Z(n15142) );
  ANDN U17411 ( .B(n15145), .A(n15146), .Z(n15143) );
  XOR U17412 ( .A(n15147), .B(n15144), .Z(n15145) );
  IV U17413 ( .A(n15123), .Z(n15141) );
  XOR U17414 ( .A(n15148), .B(n15149), .Z(n15123) );
  ANDN U17415 ( .B(n15150), .A(n15151), .Z(n15148) );
  XOR U17416 ( .A(n15149), .B(n15152), .Z(n15150) );
  IV U17417 ( .A(n15131), .Z(n15135) );
  XOR U17418 ( .A(n15131), .B(n15113), .Z(n15133) );
  XOR U17419 ( .A(n15153), .B(n15154), .Z(n15113) );
  AND U17420 ( .A(n366), .B(n15155), .Z(n15153) );
  XOR U17421 ( .A(n15156), .B(n15154), .Z(n15155) );
  NANDN U17422 ( .A(n15115), .B(n15117), .Z(n15131) );
  XOR U17423 ( .A(n15157), .B(n15158), .Z(n15117) );
  AND U17424 ( .A(n366), .B(n15159), .Z(n15157) );
  XOR U17425 ( .A(n15158), .B(n15160), .Z(n15159) );
  XOR U17426 ( .A(n15161), .B(n15162), .Z(n366) );
  AND U17427 ( .A(n15163), .B(n15164), .Z(n15161) );
  XNOR U17428 ( .A(n15162), .B(n15128), .Z(n15164) );
  XNOR U17429 ( .A(n15165), .B(n15166), .Z(n15128) );
  ANDN U17430 ( .B(n15167), .A(n15168), .Z(n15165) );
  XOR U17431 ( .A(n15166), .B(n15169), .Z(n15167) );
  XOR U17432 ( .A(n15162), .B(n15130), .Z(n15163) );
  XOR U17433 ( .A(n15170), .B(n15171), .Z(n15130) );
  AND U17434 ( .A(n370), .B(n15172), .Z(n15170) );
  XOR U17435 ( .A(n15173), .B(n15171), .Z(n15172) );
  XNOR U17436 ( .A(n15174), .B(n15175), .Z(n15162) );
  NAND U17437 ( .A(n15176), .B(n15177), .Z(n15175) );
  XOR U17438 ( .A(n15178), .B(n15154), .Z(n15177) );
  XOR U17439 ( .A(n15168), .B(n15169), .Z(n15154) );
  XOR U17440 ( .A(n15179), .B(n15180), .Z(n15169) );
  ANDN U17441 ( .B(n15181), .A(n15182), .Z(n15179) );
  XOR U17442 ( .A(n15180), .B(n15183), .Z(n15181) );
  XOR U17443 ( .A(n15184), .B(n15185), .Z(n15168) );
  XOR U17444 ( .A(n15186), .B(n15187), .Z(n15185) );
  ANDN U17445 ( .B(n15188), .A(n15189), .Z(n15186) );
  XOR U17446 ( .A(n15190), .B(n15187), .Z(n15188) );
  IV U17447 ( .A(n15166), .Z(n15184) );
  XOR U17448 ( .A(n15191), .B(n15192), .Z(n15166) );
  ANDN U17449 ( .B(n15193), .A(n15194), .Z(n15191) );
  XOR U17450 ( .A(n15192), .B(n15195), .Z(n15193) );
  IV U17451 ( .A(n15174), .Z(n15178) );
  XOR U17452 ( .A(n15174), .B(n15156), .Z(n15176) );
  XOR U17453 ( .A(n15196), .B(n15197), .Z(n15156) );
  AND U17454 ( .A(n370), .B(n15198), .Z(n15196) );
  XOR U17455 ( .A(n15199), .B(n15197), .Z(n15198) );
  NANDN U17456 ( .A(n15158), .B(n15160), .Z(n15174) );
  XOR U17457 ( .A(n15200), .B(n15201), .Z(n15160) );
  AND U17458 ( .A(n370), .B(n15202), .Z(n15200) );
  XOR U17459 ( .A(n15201), .B(n15203), .Z(n15202) );
  XOR U17460 ( .A(n15204), .B(n15205), .Z(n370) );
  AND U17461 ( .A(n15206), .B(n15207), .Z(n15204) );
  XNOR U17462 ( .A(n15205), .B(n15171), .Z(n15207) );
  XNOR U17463 ( .A(n15208), .B(n15209), .Z(n15171) );
  ANDN U17464 ( .B(n15210), .A(n15211), .Z(n15208) );
  XOR U17465 ( .A(n15209), .B(n15212), .Z(n15210) );
  XOR U17466 ( .A(n15205), .B(n15173), .Z(n15206) );
  XOR U17467 ( .A(n15213), .B(n15214), .Z(n15173) );
  AND U17468 ( .A(n374), .B(n15215), .Z(n15213) );
  XOR U17469 ( .A(n15216), .B(n15214), .Z(n15215) );
  XNOR U17470 ( .A(n15217), .B(n15218), .Z(n15205) );
  NAND U17471 ( .A(n15219), .B(n15220), .Z(n15218) );
  XOR U17472 ( .A(n15221), .B(n15197), .Z(n15220) );
  XOR U17473 ( .A(n15211), .B(n15212), .Z(n15197) );
  XOR U17474 ( .A(n15222), .B(n15223), .Z(n15212) );
  ANDN U17475 ( .B(n15224), .A(n15225), .Z(n15222) );
  XOR U17476 ( .A(n15223), .B(n15226), .Z(n15224) );
  XOR U17477 ( .A(n15227), .B(n15228), .Z(n15211) );
  XOR U17478 ( .A(n15229), .B(n15230), .Z(n15228) );
  ANDN U17479 ( .B(n15231), .A(n15232), .Z(n15229) );
  XOR U17480 ( .A(n15233), .B(n15230), .Z(n15231) );
  IV U17481 ( .A(n15209), .Z(n15227) );
  XOR U17482 ( .A(n15234), .B(n15235), .Z(n15209) );
  ANDN U17483 ( .B(n15236), .A(n15237), .Z(n15234) );
  XOR U17484 ( .A(n15235), .B(n15238), .Z(n15236) );
  IV U17485 ( .A(n15217), .Z(n15221) );
  XOR U17486 ( .A(n15217), .B(n15199), .Z(n15219) );
  XOR U17487 ( .A(n15239), .B(n15240), .Z(n15199) );
  AND U17488 ( .A(n374), .B(n15241), .Z(n15239) );
  XOR U17489 ( .A(n15242), .B(n15240), .Z(n15241) );
  NANDN U17490 ( .A(n15201), .B(n15203), .Z(n15217) );
  XOR U17491 ( .A(n15243), .B(n15244), .Z(n15203) );
  AND U17492 ( .A(n374), .B(n15245), .Z(n15243) );
  XOR U17493 ( .A(n15244), .B(n15246), .Z(n15245) );
  XOR U17494 ( .A(n15247), .B(n15248), .Z(n374) );
  AND U17495 ( .A(n15249), .B(n15250), .Z(n15247) );
  XNOR U17496 ( .A(n15248), .B(n15214), .Z(n15250) );
  XNOR U17497 ( .A(n15251), .B(n15252), .Z(n15214) );
  ANDN U17498 ( .B(n15253), .A(n15254), .Z(n15251) );
  XOR U17499 ( .A(n15252), .B(n15255), .Z(n15253) );
  XOR U17500 ( .A(n15248), .B(n15216), .Z(n15249) );
  XOR U17501 ( .A(n15256), .B(n15257), .Z(n15216) );
  AND U17502 ( .A(n378), .B(n15258), .Z(n15256) );
  XOR U17503 ( .A(n15259), .B(n15257), .Z(n15258) );
  XNOR U17504 ( .A(n15260), .B(n15261), .Z(n15248) );
  NAND U17505 ( .A(n15262), .B(n15263), .Z(n15261) );
  XOR U17506 ( .A(n15264), .B(n15240), .Z(n15263) );
  XOR U17507 ( .A(n15254), .B(n15255), .Z(n15240) );
  XOR U17508 ( .A(n15265), .B(n15266), .Z(n15255) );
  ANDN U17509 ( .B(n15267), .A(n15268), .Z(n15265) );
  XOR U17510 ( .A(n15266), .B(n15269), .Z(n15267) );
  XOR U17511 ( .A(n15270), .B(n15271), .Z(n15254) );
  XOR U17512 ( .A(n15272), .B(n15273), .Z(n15271) );
  ANDN U17513 ( .B(n15274), .A(n15275), .Z(n15272) );
  XOR U17514 ( .A(n15276), .B(n15273), .Z(n15274) );
  IV U17515 ( .A(n15252), .Z(n15270) );
  XOR U17516 ( .A(n15277), .B(n15278), .Z(n15252) );
  ANDN U17517 ( .B(n15279), .A(n15280), .Z(n15277) );
  XOR U17518 ( .A(n15278), .B(n15281), .Z(n15279) );
  IV U17519 ( .A(n15260), .Z(n15264) );
  XOR U17520 ( .A(n15260), .B(n15242), .Z(n15262) );
  XOR U17521 ( .A(n15282), .B(n15283), .Z(n15242) );
  AND U17522 ( .A(n378), .B(n15284), .Z(n15282) );
  XOR U17523 ( .A(n15285), .B(n15283), .Z(n15284) );
  NANDN U17524 ( .A(n15244), .B(n15246), .Z(n15260) );
  XOR U17525 ( .A(n15286), .B(n15287), .Z(n15246) );
  AND U17526 ( .A(n378), .B(n15288), .Z(n15286) );
  XOR U17527 ( .A(n15287), .B(n15289), .Z(n15288) );
  XOR U17528 ( .A(n15290), .B(n15291), .Z(n378) );
  AND U17529 ( .A(n15292), .B(n15293), .Z(n15290) );
  XNOR U17530 ( .A(n15291), .B(n15257), .Z(n15293) );
  XNOR U17531 ( .A(n15294), .B(n15295), .Z(n15257) );
  ANDN U17532 ( .B(n15296), .A(n15297), .Z(n15294) );
  XOR U17533 ( .A(n15295), .B(n15298), .Z(n15296) );
  XOR U17534 ( .A(n15291), .B(n15259), .Z(n15292) );
  XOR U17535 ( .A(n15299), .B(n15300), .Z(n15259) );
  AND U17536 ( .A(n382), .B(n15301), .Z(n15299) );
  XOR U17537 ( .A(n15302), .B(n15300), .Z(n15301) );
  XNOR U17538 ( .A(n15303), .B(n15304), .Z(n15291) );
  NAND U17539 ( .A(n15305), .B(n15306), .Z(n15304) );
  XOR U17540 ( .A(n15307), .B(n15283), .Z(n15306) );
  XOR U17541 ( .A(n15297), .B(n15298), .Z(n15283) );
  XOR U17542 ( .A(n15308), .B(n15309), .Z(n15298) );
  ANDN U17543 ( .B(n15310), .A(n15311), .Z(n15308) );
  XOR U17544 ( .A(n15309), .B(n15312), .Z(n15310) );
  XOR U17545 ( .A(n15313), .B(n15314), .Z(n15297) );
  XOR U17546 ( .A(n15315), .B(n15316), .Z(n15314) );
  ANDN U17547 ( .B(n15317), .A(n15318), .Z(n15315) );
  XOR U17548 ( .A(n15319), .B(n15316), .Z(n15317) );
  IV U17549 ( .A(n15295), .Z(n15313) );
  XOR U17550 ( .A(n15320), .B(n15321), .Z(n15295) );
  ANDN U17551 ( .B(n15322), .A(n15323), .Z(n15320) );
  XOR U17552 ( .A(n15321), .B(n15324), .Z(n15322) );
  IV U17553 ( .A(n15303), .Z(n15307) );
  XOR U17554 ( .A(n15303), .B(n15285), .Z(n15305) );
  XOR U17555 ( .A(n15325), .B(n15326), .Z(n15285) );
  AND U17556 ( .A(n382), .B(n15327), .Z(n15325) );
  XOR U17557 ( .A(n15328), .B(n15326), .Z(n15327) );
  NANDN U17558 ( .A(n15287), .B(n15289), .Z(n15303) );
  XOR U17559 ( .A(n15329), .B(n15330), .Z(n15289) );
  AND U17560 ( .A(n382), .B(n15331), .Z(n15329) );
  XOR U17561 ( .A(n15330), .B(n15332), .Z(n15331) );
  XOR U17562 ( .A(n15333), .B(n15334), .Z(n382) );
  AND U17563 ( .A(n15335), .B(n15336), .Z(n15333) );
  XNOR U17564 ( .A(n15334), .B(n15300), .Z(n15336) );
  XNOR U17565 ( .A(n15337), .B(n15338), .Z(n15300) );
  ANDN U17566 ( .B(n15339), .A(n15340), .Z(n15337) );
  XOR U17567 ( .A(n15338), .B(n15341), .Z(n15339) );
  XOR U17568 ( .A(n15334), .B(n15302), .Z(n15335) );
  XOR U17569 ( .A(n15342), .B(n15343), .Z(n15302) );
  AND U17570 ( .A(n386), .B(n15344), .Z(n15342) );
  XOR U17571 ( .A(n15345), .B(n15343), .Z(n15344) );
  XNOR U17572 ( .A(n15346), .B(n15347), .Z(n15334) );
  NAND U17573 ( .A(n15348), .B(n15349), .Z(n15347) );
  XOR U17574 ( .A(n15350), .B(n15326), .Z(n15349) );
  XOR U17575 ( .A(n15340), .B(n15341), .Z(n15326) );
  XOR U17576 ( .A(n15351), .B(n15352), .Z(n15341) );
  ANDN U17577 ( .B(n15353), .A(n15354), .Z(n15351) );
  XOR U17578 ( .A(n15352), .B(n15355), .Z(n15353) );
  XOR U17579 ( .A(n15356), .B(n15357), .Z(n15340) );
  XOR U17580 ( .A(n15358), .B(n15359), .Z(n15357) );
  ANDN U17581 ( .B(n15360), .A(n15361), .Z(n15358) );
  XOR U17582 ( .A(n15362), .B(n15359), .Z(n15360) );
  IV U17583 ( .A(n15338), .Z(n15356) );
  XOR U17584 ( .A(n15363), .B(n15364), .Z(n15338) );
  ANDN U17585 ( .B(n15365), .A(n15366), .Z(n15363) );
  XOR U17586 ( .A(n15364), .B(n15367), .Z(n15365) );
  IV U17587 ( .A(n15346), .Z(n15350) );
  XOR U17588 ( .A(n15346), .B(n15328), .Z(n15348) );
  XOR U17589 ( .A(n15368), .B(n15369), .Z(n15328) );
  AND U17590 ( .A(n386), .B(n15370), .Z(n15368) );
  XOR U17591 ( .A(n15371), .B(n15369), .Z(n15370) );
  NANDN U17592 ( .A(n15330), .B(n15332), .Z(n15346) );
  XOR U17593 ( .A(n15372), .B(n15373), .Z(n15332) );
  AND U17594 ( .A(n386), .B(n15374), .Z(n15372) );
  XOR U17595 ( .A(n15373), .B(n15375), .Z(n15374) );
  XOR U17596 ( .A(n15376), .B(n15377), .Z(n386) );
  AND U17597 ( .A(n15378), .B(n15379), .Z(n15376) );
  XNOR U17598 ( .A(n15377), .B(n15343), .Z(n15379) );
  XNOR U17599 ( .A(n15380), .B(n15381), .Z(n15343) );
  ANDN U17600 ( .B(n15382), .A(n15383), .Z(n15380) );
  XOR U17601 ( .A(n15381), .B(n15384), .Z(n15382) );
  XOR U17602 ( .A(n15377), .B(n15345), .Z(n15378) );
  XOR U17603 ( .A(n15385), .B(n15386), .Z(n15345) );
  AND U17604 ( .A(n390), .B(n15387), .Z(n15385) );
  XOR U17605 ( .A(n15388), .B(n15386), .Z(n15387) );
  XNOR U17606 ( .A(n15389), .B(n15390), .Z(n15377) );
  NAND U17607 ( .A(n15391), .B(n15392), .Z(n15390) );
  XOR U17608 ( .A(n15393), .B(n15369), .Z(n15392) );
  XOR U17609 ( .A(n15383), .B(n15384), .Z(n15369) );
  XOR U17610 ( .A(n15394), .B(n15395), .Z(n15384) );
  ANDN U17611 ( .B(n15396), .A(n15397), .Z(n15394) );
  XOR U17612 ( .A(n15395), .B(n15398), .Z(n15396) );
  XOR U17613 ( .A(n15399), .B(n15400), .Z(n15383) );
  XOR U17614 ( .A(n15401), .B(n15402), .Z(n15400) );
  ANDN U17615 ( .B(n15403), .A(n15404), .Z(n15401) );
  XOR U17616 ( .A(n15405), .B(n15402), .Z(n15403) );
  IV U17617 ( .A(n15381), .Z(n15399) );
  XOR U17618 ( .A(n15406), .B(n15407), .Z(n15381) );
  ANDN U17619 ( .B(n15408), .A(n15409), .Z(n15406) );
  XOR U17620 ( .A(n15407), .B(n15410), .Z(n15408) );
  IV U17621 ( .A(n15389), .Z(n15393) );
  XOR U17622 ( .A(n15389), .B(n15371), .Z(n15391) );
  XOR U17623 ( .A(n15411), .B(n15412), .Z(n15371) );
  AND U17624 ( .A(n390), .B(n15413), .Z(n15411) );
  XOR U17625 ( .A(n15414), .B(n15412), .Z(n15413) );
  NANDN U17626 ( .A(n15373), .B(n15375), .Z(n15389) );
  XOR U17627 ( .A(n15415), .B(n15416), .Z(n15375) );
  AND U17628 ( .A(n390), .B(n15417), .Z(n15415) );
  XOR U17629 ( .A(n15416), .B(n15418), .Z(n15417) );
  XOR U17630 ( .A(n15419), .B(n15420), .Z(n390) );
  AND U17631 ( .A(n15421), .B(n15422), .Z(n15419) );
  XNOR U17632 ( .A(n15420), .B(n15386), .Z(n15422) );
  XNOR U17633 ( .A(n15423), .B(n15424), .Z(n15386) );
  ANDN U17634 ( .B(n15425), .A(n15426), .Z(n15423) );
  XOR U17635 ( .A(n15424), .B(n15427), .Z(n15425) );
  XOR U17636 ( .A(n15420), .B(n15388), .Z(n15421) );
  XOR U17637 ( .A(n15428), .B(n15429), .Z(n15388) );
  AND U17638 ( .A(n394), .B(n15430), .Z(n15428) );
  XOR U17639 ( .A(n15431), .B(n15429), .Z(n15430) );
  XNOR U17640 ( .A(n15432), .B(n15433), .Z(n15420) );
  NAND U17641 ( .A(n15434), .B(n15435), .Z(n15433) );
  XOR U17642 ( .A(n15436), .B(n15412), .Z(n15435) );
  XOR U17643 ( .A(n15426), .B(n15427), .Z(n15412) );
  XOR U17644 ( .A(n15437), .B(n15438), .Z(n15427) );
  ANDN U17645 ( .B(n15439), .A(n15440), .Z(n15437) );
  XOR U17646 ( .A(n15438), .B(n15441), .Z(n15439) );
  XOR U17647 ( .A(n15442), .B(n15443), .Z(n15426) );
  XOR U17648 ( .A(n15444), .B(n15445), .Z(n15443) );
  ANDN U17649 ( .B(n15446), .A(n15447), .Z(n15444) );
  XOR U17650 ( .A(n15448), .B(n15445), .Z(n15446) );
  IV U17651 ( .A(n15424), .Z(n15442) );
  XOR U17652 ( .A(n15449), .B(n15450), .Z(n15424) );
  ANDN U17653 ( .B(n15451), .A(n15452), .Z(n15449) );
  XOR U17654 ( .A(n15450), .B(n15453), .Z(n15451) );
  IV U17655 ( .A(n15432), .Z(n15436) );
  XOR U17656 ( .A(n15432), .B(n15414), .Z(n15434) );
  XOR U17657 ( .A(n15454), .B(n15455), .Z(n15414) );
  AND U17658 ( .A(n394), .B(n15456), .Z(n15454) );
  XOR U17659 ( .A(n15457), .B(n15455), .Z(n15456) );
  NANDN U17660 ( .A(n15416), .B(n15418), .Z(n15432) );
  XOR U17661 ( .A(n15458), .B(n15459), .Z(n15418) );
  AND U17662 ( .A(n394), .B(n15460), .Z(n15458) );
  XOR U17663 ( .A(n15459), .B(n15461), .Z(n15460) );
  XOR U17664 ( .A(n15462), .B(n15463), .Z(n394) );
  AND U17665 ( .A(n15464), .B(n15465), .Z(n15462) );
  XNOR U17666 ( .A(n15463), .B(n15429), .Z(n15465) );
  XNOR U17667 ( .A(n15466), .B(n15467), .Z(n15429) );
  ANDN U17668 ( .B(n15468), .A(n15469), .Z(n15466) );
  XOR U17669 ( .A(n15467), .B(n15470), .Z(n15468) );
  XOR U17670 ( .A(n15463), .B(n15431), .Z(n15464) );
  XOR U17671 ( .A(n15471), .B(n15472), .Z(n15431) );
  AND U17672 ( .A(n398), .B(n15473), .Z(n15471) );
  XOR U17673 ( .A(n15474), .B(n15472), .Z(n15473) );
  XNOR U17674 ( .A(n15475), .B(n15476), .Z(n15463) );
  NAND U17675 ( .A(n15477), .B(n15478), .Z(n15476) );
  XOR U17676 ( .A(n15479), .B(n15455), .Z(n15478) );
  XOR U17677 ( .A(n15469), .B(n15470), .Z(n15455) );
  XOR U17678 ( .A(n15480), .B(n15481), .Z(n15470) );
  ANDN U17679 ( .B(n15482), .A(n15483), .Z(n15480) );
  XOR U17680 ( .A(n15481), .B(n15484), .Z(n15482) );
  XOR U17681 ( .A(n15485), .B(n15486), .Z(n15469) );
  XOR U17682 ( .A(n15487), .B(n15488), .Z(n15486) );
  ANDN U17683 ( .B(n15489), .A(n15490), .Z(n15487) );
  XOR U17684 ( .A(n15491), .B(n15488), .Z(n15489) );
  IV U17685 ( .A(n15467), .Z(n15485) );
  XOR U17686 ( .A(n15492), .B(n15493), .Z(n15467) );
  ANDN U17687 ( .B(n15494), .A(n15495), .Z(n15492) );
  XOR U17688 ( .A(n15493), .B(n15496), .Z(n15494) );
  IV U17689 ( .A(n15475), .Z(n15479) );
  XOR U17690 ( .A(n15475), .B(n15457), .Z(n15477) );
  XOR U17691 ( .A(n15497), .B(n15498), .Z(n15457) );
  AND U17692 ( .A(n398), .B(n15499), .Z(n15497) );
  XOR U17693 ( .A(n15500), .B(n15498), .Z(n15499) );
  NANDN U17694 ( .A(n15459), .B(n15461), .Z(n15475) );
  XOR U17695 ( .A(n15501), .B(n15502), .Z(n15461) );
  AND U17696 ( .A(n398), .B(n15503), .Z(n15501) );
  XOR U17697 ( .A(n15502), .B(n15504), .Z(n15503) );
  XOR U17698 ( .A(n15505), .B(n15506), .Z(n398) );
  AND U17699 ( .A(n15507), .B(n15508), .Z(n15505) );
  XNOR U17700 ( .A(n15506), .B(n15472), .Z(n15508) );
  XNOR U17701 ( .A(n15509), .B(n15510), .Z(n15472) );
  ANDN U17702 ( .B(n15511), .A(n15512), .Z(n15509) );
  XOR U17703 ( .A(n15510), .B(n15513), .Z(n15511) );
  XOR U17704 ( .A(n15506), .B(n15474), .Z(n15507) );
  XOR U17705 ( .A(n15514), .B(n15515), .Z(n15474) );
  AND U17706 ( .A(n402), .B(n15516), .Z(n15514) );
  XOR U17707 ( .A(n15517), .B(n15515), .Z(n15516) );
  XNOR U17708 ( .A(n15518), .B(n15519), .Z(n15506) );
  NAND U17709 ( .A(n15520), .B(n15521), .Z(n15519) );
  XOR U17710 ( .A(n15522), .B(n15498), .Z(n15521) );
  XOR U17711 ( .A(n15512), .B(n15513), .Z(n15498) );
  XOR U17712 ( .A(n15523), .B(n15524), .Z(n15513) );
  ANDN U17713 ( .B(n15525), .A(n15526), .Z(n15523) );
  XOR U17714 ( .A(n15524), .B(n15527), .Z(n15525) );
  XOR U17715 ( .A(n15528), .B(n15529), .Z(n15512) );
  XOR U17716 ( .A(n15530), .B(n15531), .Z(n15529) );
  ANDN U17717 ( .B(n15532), .A(n15533), .Z(n15530) );
  XOR U17718 ( .A(n15534), .B(n15531), .Z(n15532) );
  IV U17719 ( .A(n15510), .Z(n15528) );
  XOR U17720 ( .A(n15535), .B(n15536), .Z(n15510) );
  ANDN U17721 ( .B(n15537), .A(n15538), .Z(n15535) );
  XOR U17722 ( .A(n15536), .B(n15539), .Z(n15537) );
  IV U17723 ( .A(n15518), .Z(n15522) );
  XOR U17724 ( .A(n15518), .B(n15500), .Z(n15520) );
  XOR U17725 ( .A(n15540), .B(n15541), .Z(n15500) );
  AND U17726 ( .A(n402), .B(n15542), .Z(n15540) );
  XOR U17727 ( .A(n15543), .B(n15541), .Z(n15542) );
  NANDN U17728 ( .A(n15502), .B(n15504), .Z(n15518) );
  XOR U17729 ( .A(n15544), .B(n15545), .Z(n15504) );
  AND U17730 ( .A(n402), .B(n15546), .Z(n15544) );
  XOR U17731 ( .A(n15545), .B(n15547), .Z(n15546) );
  XOR U17732 ( .A(n15548), .B(n15549), .Z(n402) );
  AND U17733 ( .A(n15550), .B(n15551), .Z(n15548) );
  XNOR U17734 ( .A(n15549), .B(n15515), .Z(n15551) );
  XNOR U17735 ( .A(n15552), .B(n15553), .Z(n15515) );
  ANDN U17736 ( .B(n15554), .A(n15555), .Z(n15552) );
  XOR U17737 ( .A(n15553), .B(n15556), .Z(n15554) );
  XOR U17738 ( .A(n15549), .B(n15517), .Z(n15550) );
  XOR U17739 ( .A(n15557), .B(n15558), .Z(n15517) );
  AND U17740 ( .A(n406), .B(n15559), .Z(n15557) );
  XOR U17741 ( .A(n15560), .B(n15558), .Z(n15559) );
  XNOR U17742 ( .A(n15561), .B(n15562), .Z(n15549) );
  NAND U17743 ( .A(n15563), .B(n15564), .Z(n15562) );
  XOR U17744 ( .A(n15565), .B(n15541), .Z(n15564) );
  XOR U17745 ( .A(n15555), .B(n15556), .Z(n15541) );
  XOR U17746 ( .A(n15566), .B(n15567), .Z(n15556) );
  ANDN U17747 ( .B(n15568), .A(n15569), .Z(n15566) );
  XOR U17748 ( .A(n15567), .B(n15570), .Z(n15568) );
  XOR U17749 ( .A(n15571), .B(n15572), .Z(n15555) );
  XOR U17750 ( .A(n15573), .B(n15574), .Z(n15572) );
  ANDN U17751 ( .B(n15575), .A(n15576), .Z(n15573) );
  XOR U17752 ( .A(n15577), .B(n15574), .Z(n15575) );
  IV U17753 ( .A(n15553), .Z(n15571) );
  XOR U17754 ( .A(n15578), .B(n15579), .Z(n15553) );
  ANDN U17755 ( .B(n15580), .A(n15581), .Z(n15578) );
  XOR U17756 ( .A(n15579), .B(n15582), .Z(n15580) );
  IV U17757 ( .A(n15561), .Z(n15565) );
  XOR U17758 ( .A(n15561), .B(n15543), .Z(n15563) );
  XOR U17759 ( .A(n15583), .B(n15584), .Z(n15543) );
  AND U17760 ( .A(n406), .B(n15585), .Z(n15583) );
  XOR U17761 ( .A(n15586), .B(n15584), .Z(n15585) );
  NANDN U17762 ( .A(n15545), .B(n15547), .Z(n15561) );
  XOR U17763 ( .A(n15587), .B(n15588), .Z(n15547) );
  AND U17764 ( .A(n406), .B(n15589), .Z(n15587) );
  XOR U17765 ( .A(n15588), .B(n15590), .Z(n15589) );
  XOR U17766 ( .A(n15591), .B(n15592), .Z(n406) );
  AND U17767 ( .A(n15593), .B(n15594), .Z(n15591) );
  XNOR U17768 ( .A(n15592), .B(n15558), .Z(n15594) );
  XNOR U17769 ( .A(n15595), .B(n15596), .Z(n15558) );
  ANDN U17770 ( .B(n15597), .A(n15598), .Z(n15595) );
  XOR U17771 ( .A(n15596), .B(n15599), .Z(n15597) );
  XOR U17772 ( .A(n15592), .B(n15560), .Z(n15593) );
  XOR U17773 ( .A(n15600), .B(n15601), .Z(n15560) );
  AND U17774 ( .A(n410), .B(n15602), .Z(n15600) );
  XOR U17775 ( .A(n15603), .B(n15601), .Z(n15602) );
  XNOR U17776 ( .A(n15604), .B(n15605), .Z(n15592) );
  NAND U17777 ( .A(n15606), .B(n15607), .Z(n15605) );
  XOR U17778 ( .A(n15608), .B(n15584), .Z(n15607) );
  XOR U17779 ( .A(n15598), .B(n15599), .Z(n15584) );
  XOR U17780 ( .A(n15609), .B(n15610), .Z(n15599) );
  ANDN U17781 ( .B(n15611), .A(n15612), .Z(n15609) );
  XOR U17782 ( .A(n15610), .B(n15613), .Z(n15611) );
  XOR U17783 ( .A(n15614), .B(n15615), .Z(n15598) );
  XOR U17784 ( .A(n15616), .B(n15617), .Z(n15615) );
  ANDN U17785 ( .B(n15618), .A(n15619), .Z(n15616) );
  XOR U17786 ( .A(n15620), .B(n15617), .Z(n15618) );
  IV U17787 ( .A(n15596), .Z(n15614) );
  XOR U17788 ( .A(n15621), .B(n15622), .Z(n15596) );
  ANDN U17789 ( .B(n15623), .A(n15624), .Z(n15621) );
  XOR U17790 ( .A(n15622), .B(n15625), .Z(n15623) );
  IV U17791 ( .A(n15604), .Z(n15608) );
  XOR U17792 ( .A(n15604), .B(n15586), .Z(n15606) );
  XOR U17793 ( .A(n15626), .B(n15627), .Z(n15586) );
  AND U17794 ( .A(n410), .B(n15628), .Z(n15626) );
  XOR U17795 ( .A(n15629), .B(n15627), .Z(n15628) );
  NANDN U17796 ( .A(n15588), .B(n15590), .Z(n15604) );
  XOR U17797 ( .A(n15630), .B(n15631), .Z(n15590) );
  AND U17798 ( .A(n410), .B(n15632), .Z(n15630) );
  XOR U17799 ( .A(n15631), .B(n15633), .Z(n15632) );
  XOR U17800 ( .A(n15634), .B(n15635), .Z(n410) );
  AND U17801 ( .A(n15636), .B(n15637), .Z(n15634) );
  XNOR U17802 ( .A(n15635), .B(n15601), .Z(n15637) );
  XNOR U17803 ( .A(n15638), .B(n15639), .Z(n15601) );
  ANDN U17804 ( .B(n15640), .A(n15641), .Z(n15638) );
  XOR U17805 ( .A(n15639), .B(n15642), .Z(n15640) );
  XOR U17806 ( .A(n15635), .B(n15603), .Z(n15636) );
  XOR U17807 ( .A(n15643), .B(n15644), .Z(n15603) );
  AND U17808 ( .A(n414), .B(n15645), .Z(n15643) );
  XOR U17809 ( .A(n15646), .B(n15644), .Z(n15645) );
  XNOR U17810 ( .A(n15647), .B(n15648), .Z(n15635) );
  NAND U17811 ( .A(n15649), .B(n15650), .Z(n15648) );
  XOR U17812 ( .A(n15651), .B(n15627), .Z(n15650) );
  XOR U17813 ( .A(n15641), .B(n15642), .Z(n15627) );
  XOR U17814 ( .A(n15652), .B(n15653), .Z(n15642) );
  ANDN U17815 ( .B(n15654), .A(n15655), .Z(n15652) );
  XOR U17816 ( .A(n15653), .B(n15656), .Z(n15654) );
  XOR U17817 ( .A(n15657), .B(n15658), .Z(n15641) );
  XOR U17818 ( .A(n15659), .B(n15660), .Z(n15658) );
  ANDN U17819 ( .B(n15661), .A(n15662), .Z(n15659) );
  XOR U17820 ( .A(n15663), .B(n15660), .Z(n15661) );
  IV U17821 ( .A(n15639), .Z(n15657) );
  XOR U17822 ( .A(n15664), .B(n15665), .Z(n15639) );
  ANDN U17823 ( .B(n15666), .A(n15667), .Z(n15664) );
  XOR U17824 ( .A(n15665), .B(n15668), .Z(n15666) );
  IV U17825 ( .A(n15647), .Z(n15651) );
  XOR U17826 ( .A(n15647), .B(n15629), .Z(n15649) );
  XOR U17827 ( .A(n15669), .B(n15670), .Z(n15629) );
  AND U17828 ( .A(n414), .B(n15671), .Z(n15669) );
  XOR U17829 ( .A(n15672), .B(n15670), .Z(n15671) );
  NANDN U17830 ( .A(n15631), .B(n15633), .Z(n15647) );
  XOR U17831 ( .A(n15673), .B(n15674), .Z(n15633) );
  AND U17832 ( .A(n414), .B(n15675), .Z(n15673) );
  XOR U17833 ( .A(n15674), .B(n15676), .Z(n15675) );
  XOR U17834 ( .A(n15677), .B(n15678), .Z(n414) );
  AND U17835 ( .A(n15679), .B(n15680), .Z(n15677) );
  XNOR U17836 ( .A(n15678), .B(n15644), .Z(n15680) );
  XNOR U17837 ( .A(n15681), .B(n15682), .Z(n15644) );
  ANDN U17838 ( .B(n15683), .A(n15684), .Z(n15681) );
  XOR U17839 ( .A(n15682), .B(n15685), .Z(n15683) );
  XOR U17840 ( .A(n15678), .B(n15646), .Z(n15679) );
  XOR U17841 ( .A(n15686), .B(n15687), .Z(n15646) );
  AND U17842 ( .A(n418), .B(n15688), .Z(n15686) );
  XOR U17843 ( .A(n15689), .B(n15687), .Z(n15688) );
  XNOR U17844 ( .A(n15690), .B(n15691), .Z(n15678) );
  NAND U17845 ( .A(n15692), .B(n15693), .Z(n15691) );
  XOR U17846 ( .A(n15694), .B(n15670), .Z(n15693) );
  XOR U17847 ( .A(n15684), .B(n15685), .Z(n15670) );
  XOR U17848 ( .A(n15695), .B(n15696), .Z(n15685) );
  ANDN U17849 ( .B(n15697), .A(n15698), .Z(n15695) );
  XOR U17850 ( .A(n15696), .B(n15699), .Z(n15697) );
  XOR U17851 ( .A(n15700), .B(n15701), .Z(n15684) );
  XOR U17852 ( .A(n15702), .B(n15703), .Z(n15701) );
  ANDN U17853 ( .B(n15704), .A(n15705), .Z(n15702) );
  XOR U17854 ( .A(n15706), .B(n15703), .Z(n15704) );
  IV U17855 ( .A(n15682), .Z(n15700) );
  XOR U17856 ( .A(n15707), .B(n15708), .Z(n15682) );
  ANDN U17857 ( .B(n15709), .A(n15710), .Z(n15707) );
  XOR U17858 ( .A(n15708), .B(n15711), .Z(n15709) );
  IV U17859 ( .A(n15690), .Z(n15694) );
  XOR U17860 ( .A(n15690), .B(n15672), .Z(n15692) );
  XOR U17861 ( .A(n15712), .B(n15713), .Z(n15672) );
  AND U17862 ( .A(n418), .B(n15714), .Z(n15712) );
  XOR U17863 ( .A(n15715), .B(n15713), .Z(n15714) );
  NANDN U17864 ( .A(n15674), .B(n15676), .Z(n15690) );
  XOR U17865 ( .A(n15716), .B(n15717), .Z(n15676) );
  AND U17866 ( .A(n418), .B(n15718), .Z(n15716) );
  XOR U17867 ( .A(n15717), .B(n15719), .Z(n15718) );
  XOR U17868 ( .A(n15720), .B(n15721), .Z(n418) );
  AND U17869 ( .A(n15722), .B(n15723), .Z(n15720) );
  XNOR U17870 ( .A(n15721), .B(n15687), .Z(n15723) );
  XNOR U17871 ( .A(n15724), .B(n15725), .Z(n15687) );
  ANDN U17872 ( .B(n15726), .A(n15727), .Z(n15724) );
  XOR U17873 ( .A(n15725), .B(n15728), .Z(n15726) );
  XOR U17874 ( .A(n15721), .B(n15689), .Z(n15722) );
  XOR U17875 ( .A(n15729), .B(n15730), .Z(n15689) );
  AND U17876 ( .A(n422), .B(n15731), .Z(n15729) );
  XOR U17877 ( .A(n15732), .B(n15730), .Z(n15731) );
  XNOR U17878 ( .A(n15733), .B(n15734), .Z(n15721) );
  NAND U17879 ( .A(n15735), .B(n15736), .Z(n15734) );
  XOR U17880 ( .A(n15737), .B(n15713), .Z(n15736) );
  XOR U17881 ( .A(n15727), .B(n15728), .Z(n15713) );
  XOR U17882 ( .A(n15738), .B(n15739), .Z(n15728) );
  ANDN U17883 ( .B(n15740), .A(n15741), .Z(n15738) );
  XOR U17884 ( .A(n15739), .B(n15742), .Z(n15740) );
  XOR U17885 ( .A(n15743), .B(n15744), .Z(n15727) );
  XOR U17886 ( .A(n15745), .B(n15746), .Z(n15744) );
  ANDN U17887 ( .B(n15747), .A(n15748), .Z(n15745) );
  XOR U17888 ( .A(n15749), .B(n15746), .Z(n15747) );
  IV U17889 ( .A(n15725), .Z(n15743) );
  XOR U17890 ( .A(n15750), .B(n15751), .Z(n15725) );
  ANDN U17891 ( .B(n15752), .A(n15753), .Z(n15750) );
  XOR U17892 ( .A(n15751), .B(n15754), .Z(n15752) );
  IV U17893 ( .A(n15733), .Z(n15737) );
  XOR U17894 ( .A(n15733), .B(n15715), .Z(n15735) );
  XOR U17895 ( .A(n15755), .B(n15756), .Z(n15715) );
  AND U17896 ( .A(n422), .B(n15757), .Z(n15755) );
  XOR U17897 ( .A(n15758), .B(n15756), .Z(n15757) );
  NANDN U17898 ( .A(n15717), .B(n15719), .Z(n15733) );
  XOR U17899 ( .A(n15759), .B(n15760), .Z(n15719) );
  AND U17900 ( .A(n422), .B(n15761), .Z(n15759) );
  XOR U17901 ( .A(n15760), .B(n15762), .Z(n15761) );
  XOR U17902 ( .A(n15763), .B(n15764), .Z(n422) );
  AND U17903 ( .A(n15765), .B(n15766), .Z(n15763) );
  XNOR U17904 ( .A(n15764), .B(n15730), .Z(n15766) );
  XNOR U17905 ( .A(n15767), .B(n15768), .Z(n15730) );
  ANDN U17906 ( .B(n15769), .A(n15770), .Z(n15767) );
  XOR U17907 ( .A(n15768), .B(n15771), .Z(n15769) );
  XOR U17908 ( .A(n15764), .B(n15732), .Z(n15765) );
  XOR U17909 ( .A(n15772), .B(n15773), .Z(n15732) );
  AND U17910 ( .A(n426), .B(n15774), .Z(n15772) );
  XOR U17911 ( .A(n15775), .B(n15773), .Z(n15774) );
  XNOR U17912 ( .A(n15776), .B(n15777), .Z(n15764) );
  NAND U17913 ( .A(n15778), .B(n15779), .Z(n15777) );
  XOR U17914 ( .A(n15780), .B(n15756), .Z(n15779) );
  XOR U17915 ( .A(n15770), .B(n15771), .Z(n15756) );
  XOR U17916 ( .A(n15781), .B(n15782), .Z(n15771) );
  ANDN U17917 ( .B(n15783), .A(n15784), .Z(n15781) );
  XOR U17918 ( .A(n15782), .B(n15785), .Z(n15783) );
  XOR U17919 ( .A(n15786), .B(n15787), .Z(n15770) );
  XOR U17920 ( .A(n15788), .B(n15789), .Z(n15787) );
  ANDN U17921 ( .B(n15790), .A(n15791), .Z(n15788) );
  XOR U17922 ( .A(n15792), .B(n15789), .Z(n15790) );
  IV U17923 ( .A(n15768), .Z(n15786) );
  XOR U17924 ( .A(n15793), .B(n15794), .Z(n15768) );
  ANDN U17925 ( .B(n15795), .A(n15796), .Z(n15793) );
  XOR U17926 ( .A(n15794), .B(n15797), .Z(n15795) );
  IV U17927 ( .A(n15776), .Z(n15780) );
  XOR U17928 ( .A(n15776), .B(n15758), .Z(n15778) );
  XOR U17929 ( .A(n15798), .B(n15799), .Z(n15758) );
  AND U17930 ( .A(n426), .B(n15800), .Z(n15798) );
  XOR U17931 ( .A(n15801), .B(n15799), .Z(n15800) );
  NANDN U17932 ( .A(n15760), .B(n15762), .Z(n15776) );
  XOR U17933 ( .A(n15802), .B(n15803), .Z(n15762) );
  AND U17934 ( .A(n426), .B(n15804), .Z(n15802) );
  XOR U17935 ( .A(n15803), .B(n15805), .Z(n15804) );
  XOR U17936 ( .A(n15806), .B(n15807), .Z(n426) );
  AND U17937 ( .A(n15808), .B(n15809), .Z(n15806) );
  XNOR U17938 ( .A(n15807), .B(n15773), .Z(n15809) );
  XNOR U17939 ( .A(n15810), .B(n15811), .Z(n15773) );
  ANDN U17940 ( .B(n15812), .A(n15813), .Z(n15810) );
  XOR U17941 ( .A(n15811), .B(n15814), .Z(n15812) );
  XOR U17942 ( .A(n15807), .B(n15775), .Z(n15808) );
  XOR U17943 ( .A(n15815), .B(n15816), .Z(n15775) );
  AND U17944 ( .A(n430), .B(n15817), .Z(n15815) );
  XOR U17945 ( .A(n15818), .B(n15816), .Z(n15817) );
  XNOR U17946 ( .A(n15819), .B(n15820), .Z(n15807) );
  NAND U17947 ( .A(n15821), .B(n15822), .Z(n15820) );
  XOR U17948 ( .A(n15823), .B(n15799), .Z(n15822) );
  XOR U17949 ( .A(n15813), .B(n15814), .Z(n15799) );
  XOR U17950 ( .A(n15824), .B(n15825), .Z(n15814) );
  ANDN U17951 ( .B(n15826), .A(n15827), .Z(n15824) );
  XOR U17952 ( .A(n15825), .B(n15828), .Z(n15826) );
  XOR U17953 ( .A(n15829), .B(n15830), .Z(n15813) );
  XOR U17954 ( .A(n15831), .B(n15832), .Z(n15830) );
  ANDN U17955 ( .B(n15833), .A(n15834), .Z(n15831) );
  XOR U17956 ( .A(n15835), .B(n15832), .Z(n15833) );
  IV U17957 ( .A(n15811), .Z(n15829) );
  XOR U17958 ( .A(n15836), .B(n15837), .Z(n15811) );
  ANDN U17959 ( .B(n15838), .A(n15839), .Z(n15836) );
  XOR U17960 ( .A(n15837), .B(n15840), .Z(n15838) );
  IV U17961 ( .A(n15819), .Z(n15823) );
  XOR U17962 ( .A(n15819), .B(n15801), .Z(n15821) );
  XOR U17963 ( .A(n15841), .B(n15842), .Z(n15801) );
  AND U17964 ( .A(n430), .B(n15843), .Z(n15841) );
  XOR U17965 ( .A(n15844), .B(n15842), .Z(n15843) );
  NANDN U17966 ( .A(n15803), .B(n15805), .Z(n15819) );
  XOR U17967 ( .A(n15845), .B(n15846), .Z(n15805) );
  AND U17968 ( .A(n430), .B(n15847), .Z(n15845) );
  XOR U17969 ( .A(n15846), .B(n15848), .Z(n15847) );
  XOR U17970 ( .A(n15849), .B(n15850), .Z(n430) );
  AND U17971 ( .A(n15851), .B(n15852), .Z(n15849) );
  XNOR U17972 ( .A(n15850), .B(n15816), .Z(n15852) );
  XNOR U17973 ( .A(n15853), .B(n15854), .Z(n15816) );
  ANDN U17974 ( .B(n15855), .A(n15856), .Z(n15853) );
  XOR U17975 ( .A(n15854), .B(n15857), .Z(n15855) );
  XOR U17976 ( .A(n15850), .B(n15818), .Z(n15851) );
  XOR U17977 ( .A(n15858), .B(n15859), .Z(n15818) );
  AND U17978 ( .A(n434), .B(n15860), .Z(n15858) );
  XOR U17979 ( .A(n15861), .B(n15859), .Z(n15860) );
  XNOR U17980 ( .A(n15862), .B(n15863), .Z(n15850) );
  NAND U17981 ( .A(n15864), .B(n15865), .Z(n15863) );
  XOR U17982 ( .A(n15866), .B(n15842), .Z(n15865) );
  XOR U17983 ( .A(n15856), .B(n15857), .Z(n15842) );
  XOR U17984 ( .A(n15867), .B(n15868), .Z(n15857) );
  ANDN U17985 ( .B(n15869), .A(n15870), .Z(n15867) );
  XOR U17986 ( .A(n15868), .B(n15871), .Z(n15869) );
  XOR U17987 ( .A(n15872), .B(n15873), .Z(n15856) );
  XOR U17988 ( .A(n15874), .B(n15875), .Z(n15873) );
  ANDN U17989 ( .B(n15876), .A(n15877), .Z(n15874) );
  XOR U17990 ( .A(n15878), .B(n15875), .Z(n15876) );
  IV U17991 ( .A(n15854), .Z(n15872) );
  XOR U17992 ( .A(n15879), .B(n15880), .Z(n15854) );
  ANDN U17993 ( .B(n15881), .A(n15882), .Z(n15879) );
  XOR U17994 ( .A(n15880), .B(n15883), .Z(n15881) );
  IV U17995 ( .A(n15862), .Z(n15866) );
  XOR U17996 ( .A(n15862), .B(n15844), .Z(n15864) );
  XOR U17997 ( .A(n15884), .B(n15885), .Z(n15844) );
  AND U17998 ( .A(n434), .B(n15886), .Z(n15884) );
  XOR U17999 ( .A(n15887), .B(n15885), .Z(n15886) );
  NANDN U18000 ( .A(n15846), .B(n15848), .Z(n15862) );
  XOR U18001 ( .A(n15888), .B(n15889), .Z(n15848) );
  AND U18002 ( .A(n434), .B(n15890), .Z(n15888) );
  XOR U18003 ( .A(n15889), .B(n15891), .Z(n15890) );
  XOR U18004 ( .A(n15892), .B(n15893), .Z(n434) );
  AND U18005 ( .A(n15894), .B(n15895), .Z(n15892) );
  XNOR U18006 ( .A(n15893), .B(n15859), .Z(n15895) );
  XNOR U18007 ( .A(n15896), .B(n15897), .Z(n15859) );
  ANDN U18008 ( .B(n15898), .A(n15899), .Z(n15896) );
  XOR U18009 ( .A(n15897), .B(n15900), .Z(n15898) );
  XOR U18010 ( .A(n15893), .B(n15861), .Z(n15894) );
  XOR U18011 ( .A(n15901), .B(n15902), .Z(n15861) );
  AND U18012 ( .A(n438), .B(n15903), .Z(n15901) );
  XOR U18013 ( .A(n15904), .B(n15902), .Z(n15903) );
  XNOR U18014 ( .A(n15905), .B(n15906), .Z(n15893) );
  NAND U18015 ( .A(n15907), .B(n15908), .Z(n15906) );
  XOR U18016 ( .A(n15909), .B(n15885), .Z(n15908) );
  XOR U18017 ( .A(n15899), .B(n15900), .Z(n15885) );
  XOR U18018 ( .A(n15910), .B(n15911), .Z(n15900) );
  ANDN U18019 ( .B(n15912), .A(n15913), .Z(n15910) );
  XOR U18020 ( .A(n15911), .B(n15914), .Z(n15912) );
  XOR U18021 ( .A(n15915), .B(n15916), .Z(n15899) );
  XOR U18022 ( .A(n15917), .B(n15918), .Z(n15916) );
  ANDN U18023 ( .B(n15919), .A(n15920), .Z(n15917) );
  XOR U18024 ( .A(n15921), .B(n15918), .Z(n15919) );
  IV U18025 ( .A(n15897), .Z(n15915) );
  XOR U18026 ( .A(n15922), .B(n15923), .Z(n15897) );
  ANDN U18027 ( .B(n15924), .A(n15925), .Z(n15922) );
  XOR U18028 ( .A(n15923), .B(n15926), .Z(n15924) );
  IV U18029 ( .A(n15905), .Z(n15909) );
  XOR U18030 ( .A(n15905), .B(n15887), .Z(n15907) );
  XOR U18031 ( .A(n15927), .B(n15928), .Z(n15887) );
  AND U18032 ( .A(n438), .B(n15929), .Z(n15927) );
  XOR U18033 ( .A(n15930), .B(n15928), .Z(n15929) );
  NANDN U18034 ( .A(n15889), .B(n15891), .Z(n15905) );
  XOR U18035 ( .A(n15931), .B(n15932), .Z(n15891) );
  AND U18036 ( .A(n438), .B(n15933), .Z(n15931) );
  XOR U18037 ( .A(n15932), .B(n15934), .Z(n15933) );
  XOR U18038 ( .A(n15935), .B(n15936), .Z(n438) );
  AND U18039 ( .A(n15937), .B(n15938), .Z(n15935) );
  XNOR U18040 ( .A(n15936), .B(n15902), .Z(n15938) );
  XNOR U18041 ( .A(n15939), .B(n15940), .Z(n15902) );
  ANDN U18042 ( .B(n15941), .A(n15942), .Z(n15939) );
  XOR U18043 ( .A(n15940), .B(n15943), .Z(n15941) );
  XOR U18044 ( .A(n15936), .B(n15904), .Z(n15937) );
  XOR U18045 ( .A(n15944), .B(n15945), .Z(n15904) );
  AND U18046 ( .A(n442), .B(n15946), .Z(n15944) );
  XOR U18047 ( .A(n15947), .B(n15945), .Z(n15946) );
  XNOR U18048 ( .A(n15948), .B(n15949), .Z(n15936) );
  NAND U18049 ( .A(n15950), .B(n15951), .Z(n15949) );
  XOR U18050 ( .A(n15952), .B(n15928), .Z(n15951) );
  XOR U18051 ( .A(n15942), .B(n15943), .Z(n15928) );
  XOR U18052 ( .A(n15953), .B(n15954), .Z(n15943) );
  ANDN U18053 ( .B(n15955), .A(n15956), .Z(n15953) );
  XOR U18054 ( .A(n15954), .B(n15957), .Z(n15955) );
  XOR U18055 ( .A(n15958), .B(n15959), .Z(n15942) );
  XOR U18056 ( .A(n15960), .B(n15961), .Z(n15959) );
  ANDN U18057 ( .B(n15962), .A(n15963), .Z(n15960) );
  XOR U18058 ( .A(n15964), .B(n15961), .Z(n15962) );
  IV U18059 ( .A(n15940), .Z(n15958) );
  XOR U18060 ( .A(n15965), .B(n15966), .Z(n15940) );
  ANDN U18061 ( .B(n15967), .A(n15968), .Z(n15965) );
  XOR U18062 ( .A(n15966), .B(n15969), .Z(n15967) );
  IV U18063 ( .A(n15948), .Z(n15952) );
  XOR U18064 ( .A(n15948), .B(n15930), .Z(n15950) );
  XOR U18065 ( .A(n15970), .B(n15971), .Z(n15930) );
  AND U18066 ( .A(n442), .B(n15972), .Z(n15970) );
  XOR U18067 ( .A(n15973), .B(n15971), .Z(n15972) );
  NANDN U18068 ( .A(n15932), .B(n15934), .Z(n15948) );
  XOR U18069 ( .A(n15974), .B(n15975), .Z(n15934) );
  AND U18070 ( .A(n442), .B(n15976), .Z(n15974) );
  XOR U18071 ( .A(n15975), .B(n15977), .Z(n15976) );
  XOR U18072 ( .A(n15978), .B(n15979), .Z(n442) );
  AND U18073 ( .A(n15980), .B(n15981), .Z(n15978) );
  XNOR U18074 ( .A(n15979), .B(n15945), .Z(n15981) );
  XNOR U18075 ( .A(n15982), .B(n15983), .Z(n15945) );
  ANDN U18076 ( .B(n15984), .A(n15985), .Z(n15982) );
  XOR U18077 ( .A(n15983), .B(n15986), .Z(n15984) );
  XOR U18078 ( .A(n15979), .B(n15947), .Z(n15980) );
  XOR U18079 ( .A(n15987), .B(n15988), .Z(n15947) );
  AND U18080 ( .A(n446), .B(n15989), .Z(n15987) );
  XOR U18081 ( .A(n15990), .B(n15988), .Z(n15989) );
  XNOR U18082 ( .A(n15991), .B(n15992), .Z(n15979) );
  NAND U18083 ( .A(n15993), .B(n15994), .Z(n15992) );
  XOR U18084 ( .A(n15995), .B(n15971), .Z(n15994) );
  XOR U18085 ( .A(n15985), .B(n15986), .Z(n15971) );
  XOR U18086 ( .A(n15996), .B(n15997), .Z(n15986) );
  ANDN U18087 ( .B(n15998), .A(n15999), .Z(n15996) );
  XOR U18088 ( .A(n15997), .B(n16000), .Z(n15998) );
  XOR U18089 ( .A(n16001), .B(n16002), .Z(n15985) );
  XOR U18090 ( .A(n16003), .B(n16004), .Z(n16002) );
  ANDN U18091 ( .B(n16005), .A(n16006), .Z(n16003) );
  XOR U18092 ( .A(n16007), .B(n16004), .Z(n16005) );
  IV U18093 ( .A(n15983), .Z(n16001) );
  XOR U18094 ( .A(n16008), .B(n16009), .Z(n15983) );
  ANDN U18095 ( .B(n16010), .A(n16011), .Z(n16008) );
  XOR U18096 ( .A(n16009), .B(n16012), .Z(n16010) );
  IV U18097 ( .A(n15991), .Z(n15995) );
  XOR U18098 ( .A(n15991), .B(n15973), .Z(n15993) );
  XOR U18099 ( .A(n16013), .B(n16014), .Z(n15973) );
  AND U18100 ( .A(n446), .B(n16015), .Z(n16013) );
  XOR U18101 ( .A(n16016), .B(n16014), .Z(n16015) );
  NANDN U18102 ( .A(n15975), .B(n15977), .Z(n15991) );
  XOR U18103 ( .A(n16017), .B(n16018), .Z(n15977) );
  AND U18104 ( .A(n446), .B(n16019), .Z(n16017) );
  XOR U18105 ( .A(n16018), .B(n16020), .Z(n16019) );
  XOR U18106 ( .A(n16021), .B(n16022), .Z(n446) );
  AND U18107 ( .A(n16023), .B(n16024), .Z(n16021) );
  XNOR U18108 ( .A(n16022), .B(n15988), .Z(n16024) );
  XNOR U18109 ( .A(n16025), .B(n16026), .Z(n15988) );
  ANDN U18110 ( .B(n16027), .A(n16028), .Z(n16025) );
  XOR U18111 ( .A(n16026), .B(n16029), .Z(n16027) );
  XOR U18112 ( .A(n16022), .B(n15990), .Z(n16023) );
  XOR U18113 ( .A(n16030), .B(n16031), .Z(n15990) );
  AND U18114 ( .A(n450), .B(n16032), .Z(n16030) );
  XOR U18115 ( .A(n16033), .B(n16031), .Z(n16032) );
  XNOR U18116 ( .A(n16034), .B(n16035), .Z(n16022) );
  NAND U18117 ( .A(n16036), .B(n16037), .Z(n16035) );
  XOR U18118 ( .A(n16038), .B(n16014), .Z(n16037) );
  XOR U18119 ( .A(n16028), .B(n16029), .Z(n16014) );
  XOR U18120 ( .A(n16039), .B(n16040), .Z(n16029) );
  ANDN U18121 ( .B(n16041), .A(n16042), .Z(n16039) );
  XOR U18122 ( .A(n16040), .B(n16043), .Z(n16041) );
  XOR U18123 ( .A(n16044), .B(n16045), .Z(n16028) );
  XOR U18124 ( .A(n16046), .B(n16047), .Z(n16045) );
  ANDN U18125 ( .B(n16048), .A(n16049), .Z(n16046) );
  XOR U18126 ( .A(n16050), .B(n16047), .Z(n16048) );
  IV U18127 ( .A(n16026), .Z(n16044) );
  XOR U18128 ( .A(n16051), .B(n16052), .Z(n16026) );
  ANDN U18129 ( .B(n16053), .A(n16054), .Z(n16051) );
  XOR U18130 ( .A(n16052), .B(n16055), .Z(n16053) );
  IV U18131 ( .A(n16034), .Z(n16038) );
  XOR U18132 ( .A(n16034), .B(n16016), .Z(n16036) );
  XOR U18133 ( .A(n16056), .B(n16057), .Z(n16016) );
  AND U18134 ( .A(n450), .B(n16058), .Z(n16056) );
  XOR U18135 ( .A(n16059), .B(n16057), .Z(n16058) );
  NANDN U18136 ( .A(n16018), .B(n16020), .Z(n16034) );
  XOR U18137 ( .A(n16060), .B(n16061), .Z(n16020) );
  AND U18138 ( .A(n450), .B(n16062), .Z(n16060) );
  XOR U18139 ( .A(n16061), .B(n16063), .Z(n16062) );
  XOR U18140 ( .A(n16064), .B(n16065), .Z(n450) );
  AND U18141 ( .A(n16066), .B(n16067), .Z(n16064) );
  XNOR U18142 ( .A(n16065), .B(n16031), .Z(n16067) );
  XNOR U18143 ( .A(n16068), .B(n16069), .Z(n16031) );
  ANDN U18144 ( .B(n16070), .A(n16071), .Z(n16068) );
  XOR U18145 ( .A(n16069), .B(n16072), .Z(n16070) );
  XOR U18146 ( .A(n16065), .B(n16033), .Z(n16066) );
  XOR U18147 ( .A(n16073), .B(n16074), .Z(n16033) );
  AND U18148 ( .A(n454), .B(n16075), .Z(n16073) );
  XOR U18149 ( .A(n16076), .B(n16074), .Z(n16075) );
  XNOR U18150 ( .A(n16077), .B(n16078), .Z(n16065) );
  NAND U18151 ( .A(n16079), .B(n16080), .Z(n16078) );
  XOR U18152 ( .A(n16081), .B(n16057), .Z(n16080) );
  XOR U18153 ( .A(n16071), .B(n16072), .Z(n16057) );
  XOR U18154 ( .A(n16082), .B(n16083), .Z(n16072) );
  ANDN U18155 ( .B(n16084), .A(n16085), .Z(n16082) );
  XOR U18156 ( .A(n16083), .B(n16086), .Z(n16084) );
  XOR U18157 ( .A(n16087), .B(n16088), .Z(n16071) );
  XOR U18158 ( .A(n16089), .B(n16090), .Z(n16088) );
  ANDN U18159 ( .B(n16091), .A(n16092), .Z(n16089) );
  XOR U18160 ( .A(n16093), .B(n16090), .Z(n16091) );
  IV U18161 ( .A(n16069), .Z(n16087) );
  XOR U18162 ( .A(n16094), .B(n16095), .Z(n16069) );
  ANDN U18163 ( .B(n16096), .A(n16097), .Z(n16094) );
  XOR U18164 ( .A(n16095), .B(n16098), .Z(n16096) );
  IV U18165 ( .A(n16077), .Z(n16081) );
  XOR U18166 ( .A(n16077), .B(n16059), .Z(n16079) );
  XOR U18167 ( .A(n16099), .B(n16100), .Z(n16059) );
  AND U18168 ( .A(n454), .B(n16101), .Z(n16099) );
  XOR U18169 ( .A(n16102), .B(n16100), .Z(n16101) );
  NANDN U18170 ( .A(n16061), .B(n16063), .Z(n16077) );
  XOR U18171 ( .A(n16103), .B(n16104), .Z(n16063) );
  AND U18172 ( .A(n454), .B(n16105), .Z(n16103) );
  XOR U18173 ( .A(n16104), .B(n16106), .Z(n16105) );
  XOR U18174 ( .A(n16107), .B(n16108), .Z(n454) );
  AND U18175 ( .A(n16109), .B(n16110), .Z(n16107) );
  XNOR U18176 ( .A(n16108), .B(n16074), .Z(n16110) );
  XNOR U18177 ( .A(n16111), .B(n16112), .Z(n16074) );
  ANDN U18178 ( .B(n16113), .A(n16114), .Z(n16111) );
  XOR U18179 ( .A(n16112), .B(n16115), .Z(n16113) );
  XOR U18180 ( .A(n16108), .B(n16076), .Z(n16109) );
  XOR U18181 ( .A(n16116), .B(n16117), .Z(n16076) );
  AND U18182 ( .A(n458), .B(n16118), .Z(n16116) );
  XOR U18183 ( .A(n16119), .B(n16117), .Z(n16118) );
  XNOR U18184 ( .A(n16120), .B(n16121), .Z(n16108) );
  NAND U18185 ( .A(n16122), .B(n16123), .Z(n16121) );
  XOR U18186 ( .A(n16124), .B(n16100), .Z(n16123) );
  XOR U18187 ( .A(n16114), .B(n16115), .Z(n16100) );
  XOR U18188 ( .A(n16125), .B(n16126), .Z(n16115) );
  ANDN U18189 ( .B(n16127), .A(n16128), .Z(n16125) );
  XOR U18190 ( .A(n16126), .B(n16129), .Z(n16127) );
  XOR U18191 ( .A(n16130), .B(n16131), .Z(n16114) );
  XOR U18192 ( .A(n16132), .B(n16133), .Z(n16131) );
  ANDN U18193 ( .B(n16134), .A(n16135), .Z(n16132) );
  XOR U18194 ( .A(n16136), .B(n16133), .Z(n16134) );
  IV U18195 ( .A(n16112), .Z(n16130) );
  XOR U18196 ( .A(n16137), .B(n16138), .Z(n16112) );
  ANDN U18197 ( .B(n16139), .A(n16140), .Z(n16137) );
  XOR U18198 ( .A(n16138), .B(n16141), .Z(n16139) );
  IV U18199 ( .A(n16120), .Z(n16124) );
  XOR U18200 ( .A(n16120), .B(n16102), .Z(n16122) );
  XOR U18201 ( .A(n16142), .B(n16143), .Z(n16102) );
  AND U18202 ( .A(n458), .B(n16144), .Z(n16142) );
  XOR U18203 ( .A(n16145), .B(n16143), .Z(n16144) );
  NANDN U18204 ( .A(n16104), .B(n16106), .Z(n16120) );
  XOR U18205 ( .A(n16146), .B(n16147), .Z(n16106) );
  AND U18206 ( .A(n458), .B(n16148), .Z(n16146) );
  XOR U18207 ( .A(n16147), .B(n16149), .Z(n16148) );
  XOR U18208 ( .A(n16150), .B(n16151), .Z(n458) );
  AND U18209 ( .A(n16152), .B(n16153), .Z(n16150) );
  XNOR U18210 ( .A(n16151), .B(n16117), .Z(n16153) );
  XNOR U18211 ( .A(n16154), .B(n16155), .Z(n16117) );
  ANDN U18212 ( .B(n16156), .A(n16157), .Z(n16154) );
  XOR U18213 ( .A(n16155), .B(n16158), .Z(n16156) );
  XOR U18214 ( .A(n16151), .B(n16119), .Z(n16152) );
  XOR U18215 ( .A(n16159), .B(n16160), .Z(n16119) );
  AND U18216 ( .A(n462), .B(n16161), .Z(n16159) );
  XOR U18217 ( .A(n16162), .B(n16160), .Z(n16161) );
  XNOR U18218 ( .A(n16163), .B(n16164), .Z(n16151) );
  NAND U18219 ( .A(n16165), .B(n16166), .Z(n16164) );
  XOR U18220 ( .A(n16167), .B(n16143), .Z(n16166) );
  XOR U18221 ( .A(n16157), .B(n16158), .Z(n16143) );
  XOR U18222 ( .A(n16168), .B(n16169), .Z(n16158) );
  ANDN U18223 ( .B(n16170), .A(n16171), .Z(n16168) );
  XOR U18224 ( .A(n16169), .B(n16172), .Z(n16170) );
  XOR U18225 ( .A(n16173), .B(n16174), .Z(n16157) );
  XOR U18226 ( .A(n16175), .B(n16176), .Z(n16174) );
  ANDN U18227 ( .B(n16177), .A(n16178), .Z(n16175) );
  XOR U18228 ( .A(n16179), .B(n16176), .Z(n16177) );
  IV U18229 ( .A(n16155), .Z(n16173) );
  XOR U18230 ( .A(n16180), .B(n16181), .Z(n16155) );
  ANDN U18231 ( .B(n16182), .A(n16183), .Z(n16180) );
  XOR U18232 ( .A(n16181), .B(n16184), .Z(n16182) );
  IV U18233 ( .A(n16163), .Z(n16167) );
  XOR U18234 ( .A(n16163), .B(n16145), .Z(n16165) );
  XOR U18235 ( .A(n16185), .B(n16186), .Z(n16145) );
  AND U18236 ( .A(n462), .B(n16187), .Z(n16185) );
  XOR U18237 ( .A(n16188), .B(n16186), .Z(n16187) );
  NANDN U18238 ( .A(n16147), .B(n16149), .Z(n16163) );
  XOR U18239 ( .A(n16189), .B(n16190), .Z(n16149) );
  AND U18240 ( .A(n462), .B(n16191), .Z(n16189) );
  XOR U18241 ( .A(n16190), .B(n16192), .Z(n16191) );
  XOR U18242 ( .A(n16193), .B(n16194), .Z(n462) );
  AND U18243 ( .A(n16195), .B(n16196), .Z(n16193) );
  XNOR U18244 ( .A(n16194), .B(n16160), .Z(n16196) );
  XNOR U18245 ( .A(n16197), .B(n16198), .Z(n16160) );
  ANDN U18246 ( .B(n16199), .A(n16200), .Z(n16197) );
  XOR U18247 ( .A(n16198), .B(n16201), .Z(n16199) );
  XOR U18248 ( .A(n16194), .B(n16162), .Z(n16195) );
  XOR U18249 ( .A(n16202), .B(n16203), .Z(n16162) );
  AND U18250 ( .A(n466), .B(n16204), .Z(n16202) );
  XOR U18251 ( .A(n16205), .B(n16203), .Z(n16204) );
  XNOR U18252 ( .A(n16206), .B(n16207), .Z(n16194) );
  NAND U18253 ( .A(n16208), .B(n16209), .Z(n16207) );
  XOR U18254 ( .A(n16210), .B(n16186), .Z(n16209) );
  XOR U18255 ( .A(n16200), .B(n16201), .Z(n16186) );
  XOR U18256 ( .A(n16211), .B(n16212), .Z(n16201) );
  ANDN U18257 ( .B(n16213), .A(n16214), .Z(n16211) );
  XOR U18258 ( .A(n16212), .B(n16215), .Z(n16213) );
  XOR U18259 ( .A(n16216), .B(n16217), .Z(n16200) );
  XOR U18260 ( .A(n16218), .B(n16219), .Z(n16217) );
  ANDN U18261 ( .B(n16220), .A(n16221), .Z(n16218) );
  XOR U18262 ( .A(n16222), .B(n16219), .Z(n16220) );
  IV U18263 ( .A(n16198), .Z(n16216) );
  XOR U18264 ( .A(n16223), .B(n16224), .Z(n16198) );
  ANDN U18265 ( .B(n16225), .A(n16226), .Z(n16223) );
  XOR U18266 ( .A(n16224), .B(n16227), .Z(n16225) );
  IV U18267 ( .A(n16206), .Z(n16210) );
  XOR U18268 ( .A(n16206), .B(n16188), .Z(n16208) );
  XOR U18269 ( .A(n16228), .B(n16229), .Z(n16188) );
  AND U18270 ( .A(n466), .B(n16230), .Z(n16228) );
  XOR U18271 ( .A(n16231), .B(n16229), .Z(n16230) );
  NANDN U18272 ( .A(n16190), .B(n16192), .Z(n16206) );
  XOR U18273 ( .A(n16232), .B(n16233), .Z(n16192) );
  AND U18274 ( .A(n466), .B(n16234), .Z(n16232) );
  XOR U18275 ( .A(n16233), .B(n16235), .Z(n16234) );
  XOR U18276 ( .A(n16236), .B(n16237), .Z(n466) );
  AND U18277 ( .A(n16238), .B(n16239), .Z(n16236) );
  XNOR U18278 ( .A(n16237), .B(n16203), .Z(n16239) );
  XNOR U18279 ( .A(n16240), .B(n16241), .Z(n16203) );
  ANDN U18280 ( .B(n16242), .A(n16243), .Z(n16240) );
  XOR U18281 ( .A(n16241), .B(n16244), .Z(n16242) );
  XOR U18282 ( .A(n16237), .B(n16205), .Z(n16238) );
  XOR U18283 ( .A(n16245), .B(n16246), .Z(n16205) );
  AND U18284 ( .A(n470), .B(n16247), .Z(n16245) );
  XOR U18285 ( .A(n16248), .B(n16246), .Z(n16247) );
  XNOR U18286 ( .A(n16249), .B(n16250), .Z(n16237) );
  NAND U18287 ( .A(n16251), .B(n16252), .Z(n16250) );
  XOR U18288 ( .A(n16253), .B(n16229), .Z(n16252) );
  XOR U18289 ( .A(n16243), .B(n16244), .Z(n16229) );
  XOR U18290 ( .A(n16254), .B(n16255), .Z(n16244) );
  ANDN U18291 ( .B(n16256), .A(n16257), .Z(n16254) );
  XOR U18292 ( .A(n16255), .B(n16258), .Z(n16256) );
  XOR U18293 ( .A(n16259), .B(n16260), .Z(n16243) );
  XOR U18294 ( .A(n16261), .B(n16262), .Z(n16260) );
  ANDN U18295 ( .B(n16263), .A(n16264), .Z(n16261) );
  XOR U18296 ( .A(n16265), .B(n16262), .Z(n16263) );
  IV U18297 ( .A(n16241), .Z(n16259) );
  XOR U18298 ( .A(n16266), .B(n16267), .Z(n16241) );
  ANDN U18299 ( .B(n16268), .A(n16269), .Z(n16266) );
  XOR U18300 ( .A(n16267), .B(n16270), .Z(n16268) );
  IV U18301 ( .A(n16249), .Z(n16253) );
  XOR U18302 ( .A(n16249), .B(n16231), .Z(n16251) );
  XOR U18303 ( .A(n16271), .B(n16272), .Z(n16231) );
  AND U18304 ( .A(n470), .B(n16273), .Z(n16271) );
  XOR U18305 ( .A(n16274), .B(n16272), .Z(n16273) );
  NANDN U18306 ( .A(n16233), .B(n16235), .Z(n16249) );
  XOR U18307 ( .A(n16275), .B(n16276), .Z(n16235) );
  AND U18308 ( .A(n470), .B(n16277), .Z(n16275) );
  XOR U18309 ( .A(n16276), .B(n16278), .Z(n16277) );
  XOR U18310 ( .A(n16279), .B(n16280), .Z(n470) );
  AND U18311 ( .A(n16281), .B(n16282), .Z(n16279) );
  XNOR U18312 ( .A(n16280), .B(n16246), .Z(n16282) );
  XNOR U18313 ( .A(n16283), .B(n16284), .Z(n16246) );
  ANDN U18314 ( .B(n16285), .A(n16286), .Z(n16283) );
  XOR U18315 ( .A(n16284), .B(n16287), .Z(n16285) );
  XOR U18316 ( .A(n16280), .B(n16248), .Z(n16281) );
  XOR U18317 ( .A(n16288), .B(n16289), .Z(n16248) );
  AND U18318 ( .A(n474), .B(n16290), .Z(n16288) );
  XOR U18319 ( .A(n16291), .B(n16289), .Z(n16290) );
  XNOR U18320 ( .A(n16292), .B(n16293), .Z(n16280) );
  NAND U18321 ( .A(n16294), .B(n16295), .Z(n16293) );
  XOR U18322 ( .A(n16296), .B(n16272), .Z(n16295) );
  XOR U18323 ( .A(n16286), .B(n16287), .Z(n16272) );
  XOR U18324 ( .A(n16297), .B(n16298), .Z(n16287) );
  ANDN U18325 ( .B(n16299), .A(n16300), .Z(n16297) );
  XOR U18326 ( .A(n16298), .B(n16301), .Z(n16299) );
  XOR U18327 ( .A(n16302), .B(n16303), .Z(n16286) );
  XOR U18328 ( .A(n16304), .B(n16305), .Z(n16303) );
  ANDN U18329 ( .B(n16306), .A(n16307), .Z(n16304) );
  XOR U18330 ( .A(n16308), .B(n16305), .Z(n16306) );
  IV U18331 ( .A(n16284), .Z(n16302) );
  XOR U18332 ( .A(n16309), .B(n16310), .Z(n16284) );
  ANDN U18333 ( .B(n16311), .A(n16312), .Z(n16309) );
  XOR U18334 ( .A(n16310), .B(n16313), .Z(n16311) );
  IV U18335 ( .A(n16292), .Z(n16296) );
  XOR U18336 ( .A(n16292), .B(n16274), .Z(n16294) );
  XOR U18337 ( .A(n16314), .B(n16315), .Z(n16274) );
  AND U18338 ( .A(n474), .B(n16316), .Z(n16314) );
  XOR U18339 ( .A(n16317), .B(n16315), .Z(n16316) );
  NANDN U18340 ( .A(n16276), .B(n16278), .Z(n16292) );
  XOR U18341 ( .A(n16318), .B(n16319), .Z(n16278) );
  AND U18342 ( .A(n474), .B(n16320), .Z(n16318) );
  XOR U18343 ( .A(n16319), .B(n16321), .Z(n16320) );
  XOR U18344 ( .A(n16322), .B(n16323), .Z(n474) );
  AND U18345 ( .A(n16324), .B(n16325), .Z(n16322) );
  XNOR U18346 ( .A(n16323), .B(n16289), .Z(n16325) );
  XNOR U18347 ( .A(n16326), .B(n16327), .Z(n16289) );
  ANDN U18348 ( .B(n16328), .A(n16329), .Z(n16326) );
  XOR U18349 ( .A(n16327), .B(n16330), .Z(n16328) );
  XOR U18350 ( .A(n16323), .B(n16291), .Z(n16324) );
  XOR U18351 ( .A(n16331), .B(n16332), .Z(n16291) );
  AND U18352 ( .A(n478), .B(n16333), .Z(n16331) );
  XOR U18353 ( .A(n16334), .B(n16332), .Z(n16333) );
  XNOR U18354 ( .A(n16335), .B(n16336), .Z(n16323) );
  NAND U18355 ( .A(n16337), .B(n16338), .Z(n16336) );
  XOR U18356 ( .A(n16339), .B(n16315), .Z(n16338) );
  XOR U18357 ( .A(n16329), .B(n16330), .Z(n16315) );
  XOR U18358 ( .A(n16340), .B(n16341), .Z(n16330) );
  ANDN U18359 ( .B(n16342), .A(n16343), .Z(n16340) );
  XOR U18360 ( .A(n16341), .B(n16344), .Z(n16342) );
  XOR U18361 ( .A(n16345), .B(n16346), .Z(n16329) );
  XOR U18362 ( .A(n16347), .B(n16348), .Z(n16346) );
  ANDN U18363 ( .B(n16349), .A(n16350), .Z(n16347) );
  XOR U18364 ( .A(n16351), .B(n16348), .Z(n16349) );
  IV U18365 ( .A(n16327), .Z(n16345) );
  XOR U18366 ( .A(n16352), .B(n16353), .Z(n16327) );
  ANDN U18367 ( .B(n16354), .A(n16355), .Z(n16352) );
  XOR U18368 ( .A(n16353), .B(n16356), .Z(n16354) );
  IV U18369 ( .A(n16335), .Z(n16339) );
  XOR U18370 ( .A(n16335), .B(n16317), .Z(n16337) );
  XOR U18371 ( .A(n16357), .B(n16358), .Z(n16317) );
  AND U18372 ( .A(n478), .B(n16359), .Z(n16357) );
  XOR U18373 ( .A(n16360), .B(n16358), .Z(n16359) );
  NANDN U18374 ( .A(n16319), .B(n16321), .Z(n16335) );
  XOR U18375 ( .A(n16361), .B(n16362), .Z(n16321) );
  AND U18376 ( .A(n478), .B(n16363), .Z(n16361) );
  XOR U18377 ( .A(n16362), .B(n16364), .Z(n16363) );
  XOR U18378 ( .A(n16365), .B(n16366), .Z(n478) );
  AND U18379 ( .A(n16367), .B(n16368), .Z(n16365) );
  XNOR U18380 ( .A(n16366), .B(n16332), .Z(n16368) );
  XNOR U18381 ( .A(n16369), .B(n16370), .Z(n16332) );
  ANDN U18382 ( .B(n16371), .A(n16372), .Z(n16369) );
  XOR U18383 ( .A(n16370), .B(n16373), .Z(n16371) );
  XOR U18384 ( .A(n16366), .B(n16334), .Z(n16367) );
  XOR U18385 ( .A(n16374), .B(n16375), .Z(n16334) );
  AND U18386 ( .A(n482), .B(n16376), .Z(n16374) );
  XOR U18387 ( .A(n16377), .B(n16375), .Z(n16376) );
  XNOR U18388 ( .A(n16378), .B(n16379), .Z(n16366) );
  NAND U18389 ( .A(n16380), .B(n16381), .Z(n16379) );
  XOR U18390 ( .A(n16382), .B(n16358), .Z(n16381) );
  XOR U18391 ( .A(n16372), .B(n16373), .Z(n16358) );
  XOR U18392 ( .A(n16383), .B(n16384), .Z(n16373) );
  ANDN U18393 ( .B(n16385), .A(n16386), .Z(n16383) );
  XOR U18394 ( .A(n16384), .B(n16387), .Z(n16385) );
  XOR U18395 ( .A(n16388), .B(n16389), .Z(n16372) );
  XOR U18396 ( .A(n16390), .B(n16391), .Z(n16389) );
  ANDN U18397 ( .B(n16392), .A(n16393), .Z(n16390) );
  XOR U18398 ( .A(n16394), .B(n16391), .Z(n16392) );
  IV U18399 ( .A(n16370), .Z(n16388) );
  XOR U18400 ( .A(n16395), .B(n16396), .Z(n16370) );
  ANDN U18401 ( .B(n16397), .A(n16398), .Z(n16395) );
  XOR U18402 ( .A(n16396), .B(n16399), .Z(n16397) );
  IV U18403 ( .A(n16378), .Z(n16382) );
  XOR U18404 ( .A(n16378), .B(n16360), .Z(n16380) );
  XOR U18405 ( .A(n16400), .B(n16401), .Z(n16360) );
  AND U18406 ( .A(n482), .B(n16402), .Z(n16400) );
  XOR U18407 ( .A(n16403), .B(n16401), .Z(n16402) );
  NANDN U18408 ( .A(n16362), .B(n16364), .Z(n16378) );
  XOR U18409 ( .A(n16404), .B(n16405), .Z(n16364) );
  AND U18410 ( .A(n482), .B(n16406), .Z(n16404) );
  XOR U18411 ( .A(n16405), .B(n16407), .Z(n16406) );
  XOR U18412 ( .A(n16408), .B(n16409), .Z(n482) );
  AND U18413 ( .A(n16410), .B(n16411), .Z(n16408) );
  XNOR U18414 ( .A(n16409), .B(n16375), .Z(n16411) );
  XNOR U18415 ( .A(n16412), .B(n16413), .Z(n16375) );
  ANDN U18416 ( .B(n16414), .A(n16415), .Z(n16412) );
  XOR U18417 ( .A(n16413), .B(n16416), .Z(n16414) );
  XOR U18418 ( .A(n16409), .B(n16377), .Z(n16410) );
  XOR U18419 ( .A(n16417), .B(n16418), .Z(n16377) );
  AND U18420 ( .A(n486), .B(n16419), .Z(n16417) );
  XOR U18421 ( .A(n16420), .B(n16418), .Z(n16419) );
  XNOR U18422 ( .A(n16421), .B(n16422), .Z(n16409) );
  NAND U18423 ( .A(n16423), .B(n16424), .Z(n16422) );
  XOR U18424 ( .A(n16425), .B(n16401), .Z(n16424) );
  XOR U18425 ( .A(n16415), .B(n16416), .Z(n16401) );
  XOR U18426 ( .A(n16426), .B(n16427), .Z(n16416) );
  ANDN U18427 ( .B(n16428), .A(n16429), .Z(n16426) );
  XOR U18428 ( .A(n16427), .B(n16430), .Z(n16428) );
  XOR U18429 ( .A(n16431), .B(n16432), .Z(n16415) );
  XOR U18430 ( .A(n16433), .B(n16434), .Z(n16432) );
  ANDN U18431 ( .B(n16435), .A(n16436), .Z(n16433) );
  XOR U18432 ( .A(n16437), .B(n16434), .Z(n16435) );
  IV U18433 ( .A(n16413), .Z(n16431) );
  XOR U18434 ( .A(n16438), .B(n16439), .Z(n16413) );
  ANDN U18435 ( .B(n16440), .A(n16441), .Z(n16438) );
  XOR U18436 ( .A(n16439), .B(n16442), .Z(n16440) );
  IV U18437 ( .A(n16421), .Z(n16425) );
  XOR U18438 ( .A(n16421), .B(n16403), .Z(n16423) );
  XOR U18439 ( .A(n16443), .B(n16444), .Z(n16403) );
  AND U18440 ( .A(n486), .B(n16445), .Z(n16443) );
  XOR U18441 ( .A(n16446), .B(n16444), .Z(n16445) );
  NANDN U18442 ( .A(n16405), .B(n16407), .Z(n16421) );
  XOR U18443 ( .A(n16447), .B(n16448), .Z(n16407) );
  AND U18444 ( .A(n486), .B(n16449), .Z(n16447) );
  XOR U18445 ( .A(n16448), .B(n16450), .Z(n16449) );
  XOR U18446 ( .A(n16451), .B(n16452), .Z(n486) );
  AND U18447 ( .A(n16453), .B(n16454), .Z(n16451) );
  XNOR U18448 ( .A(n16452), .B(n16418), .Z(n16454) );
  XNOR U18449 ( .A(n16455), .B(n16456), .Z(n16418) );
  ANDN U18450 ( .B(n16457), .A(n16458), .Z(n16455) );
  XOR U18451 ( .A(n16456), .B(n16459), .Z(n16457) );
  XOR U18452 ( .A(n16452), .B(n16420), .Z(n16453) );
  XOR U18453 ( .A(n16460), .B(n16461), .Z(n16420) );
  AND U18454 ( .A(n490), .B(n16462), .Z(n16460) );
  XOR U18455 ( .A(n16463), .B(n16461), .Z(n16462) );
  XNOR U18456 ( .A(n16464), .B(n16465), .Z(n16452) );
  NAND U18457 ( .A(n16466), .B(n16467), .Z(n16465) );
  XOR U18458 ( .A(n16468), .B(n16444), .Z(n16467) );
  XOR U18459 ( .A(n16458), .B(n16459), .Z(n16444) );
  XOR U18460 ( .A(n16469), .B(n16470), .Z(n16459) );
  ANDN U18461 ( .B(n16471), .A(n16472), .Z(n16469) );
  XOR U18462 ( .A(n16470), .B(n16473), .Z(n16471) );
  XOR U18463 ( .A(n16474), .B(n16475), .Z(n16458) );
  XOR U18464 ( .A(n16476), .B(n16477), .Z(n16475) );
  ANDN U18465 ( .B(n16478), .A(n16479), .Z(n16476) );
  XOR U18466 ( .A(n16480), .B(n16477), .Z(n16478) );
  IV U18467 ( .A(n16456), .Z(n16474) );
  XOR U18468 ( .A(n16481), .B(n16482), .Z(n16456) );
  ANDN U18469 ( .B(n16483), .A(n16484), .Z(n16481) );
  XOR U18470 ( .A(n16482), .B(n16485), .Z(n16483) );
  IV U18471 ( .A(n16464), .Z(n16468) );
  XOR U18472 ( .A(n16464), .B(n16446), .Z(n16466) );
  XOR U18473 ( .A(n16486), .B(n16487), .Z(n16446) );
  AND U18474 ( .A(n490), .B(n16488), .Z(n16486) );
  XOR U18475 ( .A(n16489), .B(n16487), .Z(n16488) );
  NANDN U18476 ( .A(n16448), .B(n16450), .Z(n16464) );
  XOR U18477 ( .A(n16490), .B(n16491), .Z(n16450) );
  AND U18478 ( .A(n490), .B(n16492), .Z(n16490) );
  XOR U18479 ( .A(n16491), .B(n16493), .Z(n16492) );
  XOR U18480 ( .A(n16494), .B(n16495), .Z(n490) );
  AND U18481 ( .A(n16496), .B(n16497), .Z(n16494) );
  XNOR U18482 ( .A(n16495), .B(n16461), .Z(n16497) );
  XNOR U18483 ( .A(n16498), .B(n16499), .Z(n16461) );
  ANDN U18484 ( .B(n16500), .A(n16501), .Z(n16498) );
  XOR U18485 ( .A(n16499), .B(n16502), .Z(n16500) );
  XOR U18486 ( .A(n16495), .B(n16463), .Z(n16496) );
  XOR U18487 ( .A(n16503), .B(n16504), .Z(n16463) );
  AND U18488 ( .A(n494), .B(n16505), .Z(n16503) );
  XOR U18489 ( .A(n16506), .B(n16504), .Z(n16505) );
  XNOR U18490 ( .A(n16507), .B(n16508), .Z(n16495) );
  NAND U18491 ( .A(n16509), .B(n16510), .Z(n16508) );
  XOR U18492 ( .A(n16511), .B(n16487), .Z(n16510) );
  XOR U18493 ( .A(n16501), .B(n16502), .Z(n16487) );
  XOR U18494 ( .A(n16512), .B(n16513), .Z(n16502) );
  ANDN U18495 ( .B(n16514), .A(n16515), .Z(n16512) );
  XOR U18496 ( .A(n16513), .B(n16516), .Z(n16514) );
  XOR U18497 ( .A(n16517), .B(n16518), .Z(n16501) );
  XOR U18498 ( .A(n16519), .B(n16520), .Z(n16518) );
  ANDN U18499 ( .B(n16521), .A(n16522), .Z(n16519) );
  XOR U18500 ( .A(n16523), .B(n16520), .Z(n16521) );
  IV U18501 ( .A(n16499), .Z(n16517) );
  XOR U18502 ( .A(n16524), .B(n16525), .Z(n16499) );
  ANDN U18503 ( .B(n16526), .A(n16527), .Z(n16524) );
  XOR U18504 ( .A(n16525), .B(n16528), .Z(n16526) );
  IV U18505 ( .A(n16507), .Z(n16511) );
  XOR U18506 ( .A(n16507), .B(n16489), .Z(n16509) );
  XOR U18507 ( .A(n16529), .B(n16530), .Z(n16489) );
  AND U18508 ( .A(n494), .B(n16531), .Z(n16529) );
  XOR U18509 ( .A(n16532), .B(n16530), .Z(n16531) );
  NANDN U18510 ( .A(n16491), .B(n16493), .Z(n16507) );
  XOR U18511 ( .A(n16533), .B(n16534), .Z(n16493) );
  AND U18512 ( .A(n494), .B(n16535), .Z(n16533) );
  XOR U18513 ( .A(n16534), .B(n16536), .Z(n16535) );
  XOR U18514 ( .A(n16537), .B(n16538), .Z(n494) );
  AND U18515 ( .A(n16539), .B(n16540), .Z(n16537) );
  XNOR U18516 ( .A(n16538), .B(n16504), .Z(n16540) );
  XNOR U18517 ( .A(n16541), .B(n16542), .Z(n16504) );
  ANDN U18518 ( .B(n16543), .A(n16544), .Z(n16541) );
  XOR U18519 ( .A(n16542), .B(n16545), .Z(n16543) );
  XOR U18520 ( .A(n16538), .B(n16506), .Z(n16539) );
  XOR U18521 ( .A(n16546), .B(n16547), .Z(n16506) );
  AND U18522 ( .A(n498), .B(n16548), .Z(n16546) );
  XOR U18523 ( .A(n16549), .B(n16547), .Z(n16548) );
  XNOR U18524 ( .A(n16550), .B(n16551), .Z(n16538) );
  NAND U18525 ( .A(n16552), .B(n16553), .Z(n16551) );
  XOR U18526 ( .A(n16554), .B(n16530), .Z(n16553) );
  XOR U18527 ( .A(n16544), .B(n16545), .Z(n16530) );
  XOR U18528 ( .A(n16555), .B(n16556), .Z(n16545) );
  ANDN U18529 ( .B(n16557), .A(n16558), .Z(n16555) );
  XOR U18530 ( .A(n16556), .B(n16559), .Z(n16557) );
  XOR U18531 ( .A(n16560), .B(n16561), .Z(n16544) );
  XOR U18532 ( .A(n16562), .B(n16563), .Z(n16561) );
  ANDN U18533 ( .B(n16564), .A(n16565), .Z(n16562) );
  XOR U18534 ( .A(n16566), .B(n16563), .Z(n16564) );
  IV U18535 ( .A(n16542), .Z(n16560) );
  XOR U18536 ( .A(n16567), .B(n16568), .Z(n16542) );
  ANDN U18537 ( .B(n16569), .A(n16570), .Z(n16567) );
  XOR U18538 ( .A(n16568), .B(n16571), .Z(n16569) );
  IV U18539 ( .A(n16550), .Z(n16554) );
  XOR U18540 ( .A(n16550), .B(n16532), .Z(n16552) );
  XOR U18541 ( .A(n16572), .B(n16573), .Z(n16532) );
  AND U18542 ( .A(n498), .B(n16574), .Z(n16572) );
  XOR U18543 ( .A(n16575), .B(n16573), .Z(n16574) );
  NANDN U18544 ( .A(n16534), .B(n16536), .Z(n16550) );
  XOR U18545 ( .A(n16576), .B(n16577), .Z(n16536) );
  AND U18546 ( .A(n498), .B(n16578), .Z(n16576) );
  XOR U18547 ( .A(n16577), .B(n16579), .Z(n16578) );
  XOR U18548 ( .A(n16580), .B(n16581), .Z(n498) );
  AND U18549 ( .A(n16582), .B(n16583), .Z(n16580) );
  XNOR U18550 ( .A(n16581), .B(n16547), .Z(n16583) );
  XNOR U18551 ( .A(n16584), .B(n16585), .Z(n16547) );
  ANDN U18552 ( .B(n16586), .A(n16587), .Z(n16584) );
  XOR U18553 ( .A(n16585), .B(n16588), .Z(n16586) );
  XOR U18554 ( .A(n16581), .B(n16549), .Z(n16582) );
  XOR U18555 ( .A(n16589), .B(n16590), .Z(n16549) );
  AND U18556 ( .A(n502), .B(n16591), .Z(n16589) );
  XOR U18557 ( .A(n16592), .B(n16590), .Z(n16591) );
  XNOR U18558 ( .A(n16593), .B(n16594), .Z(n16581) );
  NAND U18559 ( .A(n16595), .B(n16596), .Z(n16594) );
  XOR U18560 ( .A(n16597), .B(n16573), .Z(n16596) );
  XOR U18561 ( .A(n16587), .B(n16588), .Z(n16573) );
  XOR U18562 ( .A(n16598), .B(n16599), .Z(n16588) );
  ANDN U18563 ( .B(n16600), .A(n16601), .Z(n16598) );
  XOR U18564 ( .A(n16599), .B(n16602), .Z(n16600) );
  XOR U18565 ( .A(n16603), .B(n16604), .Z(n16587) );
  XOR U18566 ( .A(n16605), .B(n16606), .Z(n16604) );
  ANDN U18567 ( .B(n16607), .A(n16608), .Z(n16605) );
  XOR U18568 ( .A(n16609), .B(n16606), .Z(n16607) );
  IV U18569 ( .A(n16585), .Z(n16603) );
  XOR U18570 ( .A(n16610), .B(n16611), .Z(n16585) );
  ANDN U18571 ( .B(n16612), .A(n16613), .Z(n16610) );
  XOR U18572 ( .A(n16611), .B(n16614), .Z(n16612) );
  IV U18573 ( .A(n16593), .Z(n16597) );
  XOR U18574 ( .A(n16593), .B(n16575), .Z(n16595) );
  XOR U18575 ( .A(n16615), .B(n16616), .Z(n16575) );
  AND U18576 ( .A(n502), .B(n16617), .Z(n16615) );
  XOR U18577 ( .A(n16618), .B(n16616), .Z(n16617) );
  NANDN U18578 ( .A(n16577), .B(n16579), .Z(n16593) );
  XOR U18579 ( .A(n16619), .B(n16620), .Z(n16579) );
  AND U18580 ( .A(n502), .B(n16621), .Z(n16619) );
  XOR U18581 ( .A(n16620), .B(n16622), .Z(n16621) );
  XOR U18582 ( .A(n16623), .B(n16624), .Z(n502) );
  AND U18583 ( .A(n16625), .B(n16626), .Z(n16623) );
  XNOR U18584 ( .A(n16624), .B(n16590), .Z(n16626) );
  XNOR U18585 ( .A(n16627), .B(n16628), .Z(n16590) );
  ANDN U18586 ( .B(n16629), .A(n16630), .Z(n16627) );
  XOR U18587 ( .A(n16628), .B(n16631), .Z(n16629) );
  XOR U18588 ( .A(n16624), .B(n16592), .Z(n16625) );
  XOR U18589 ( .A(n16632), .B(n16633), .Z(n16592) );
  AND U18590 ( .A(n506), .B(n16634), .Z(n16632) );
  XOR U18591 ( .A(n16635), .B(n16633), .Z(n16634) );
  XNOR U18592 ( .A(n16636), .B(n16637), .Z(n16624) );
  NAND U18593 ( .A(n16638), .B(n16639), .Z(n16637) );
  XOR U18594 ( .A(n16640), .B(n16616), .Z(n16639) );
  XOR U18595 ( .A(n16630), .B(n16631), .Z(n16616) );
  XOR U18596 ( .A(n16641), .B(n16642), .Z(n16631) );
  ANDN U18597 ( .B(n16643), .A(n16644), .Z(n16641) );
  XOR U18598 ( .A(n16642), .B(n16645), .Z(n16643) );
  XOR U18599 ( .A(n16646), .B(n16647), .Z(n16630) );
  XOR U18600 ( .A(n16648), .B(n16649), .Z(n16647) );
  ANDN U18601 ( .B(n16650), .A(n16651), .Z(n16648) );
  XOR U18602 ( .A(n16652), .B(n16649), .Z(n16650) );
  IV U18603 ( .A(n16628), .Z(n16646) );
  XOR U18604 ( .A(n16653), .B(n16654), .Z(n16628) );
  ANDN U18605 ( .B(n16655), .A(n16656), .Z(n16653) );
  XOR U18606 ( .A(n16654), .B(n16657), .Z(n16655) );
  IV U18607 ( .A(n16636), .Z(n16640) );
  XOR U18608 ( .A(n16636), .B(n16618), .Z(n16638) );
  XOR U18609 ( .A(n16658), .B(n16659), .Z(n16618) );
  AND U18610 ( .A(n506), .B(n16660), .Z(n16658) );
  XOR U18611 ( .A(n16661), .B(n16659), .Z(n16660) );
  NANDN U18612 ( .A(n16620), .B(n16622), .Z(n16636) );
  XOR U18613 ( .A(n16662), .B(n16663), .Z(n16622) );
  AND U18614 ( .A(n506), .B(n16664), .Z(n16662) );
  XOR U18615 ( .A(n16663), .B(n16665), .Z(n16664) );
  XOR U18616 ( .A(n16666), .B(n16667), .Z(n506) );
  AND U18617 ( .A(n16668), .B(n16669), .Z(n16666) );
  XNOR U18618 ( .A(n16667), .B(n16633), .Z(n16669) );
  XNOR U18619 ( .A(n16670), .B(n16671), .Z(n16633) );
  ANDN U18620 ( .B(n16672), .A(n16673), .Z(n16670) );
  XOR U18621 ( .A(n16671), .B(n16674), .Z(n16672) );
  XOR U18622 ( .A(n16667), .B(n16635), .Z(n16668) );
  XOR U18623 ( .A(n16675), .B(n16676), .Z(n16635) );
  AND U18624 ( .A(n510), .B(n16677), .Z(n16675) );
  XOR U18625 ( .A(n16678), .B(n16676), .Z(n16677) );
  XNOR U18626 ( .A(n16679), .B(n16680), .Z(n16667) );
  NAND U18627 ( .A(n16681), .B(n16682), .Z(n16680) );
  XOR U18628 ( .A(n16683), .B(n16659), .Z(n16682) );
  XOR U18629 ( .A(n16673), .B(n16674), .Z(n16659) );
  XOR U18630 ( .A(n16684), .B(n16685), .Z(n16674) );
  ANDN U18631 ( .B(n16686), .A(n16687), .Z(n16684) );
  XOR U18632 ( .A(n16685), .B(n16688), .Z(n16686) );
  XOR U18633 ( .A(n16689), .B(n16690), .Z(n16673) );
  XOR U18634 ( .A(n16691), .B(n16692), .Z(n16690) );
  ANDN U18635 ( .B(n16693), .A(n16694), .Z(n16691) );
  XOR U18636 ( .A(n16695), .B(n16692), .Z(n16693) );
  IV U18637 ( .A(n16671), .Z(n16689) );
  XOR U18638 ( .A(n16696), .B(n16697), .Z(n16671) );
  ANDN U18639 ( .B(n16698), .A(n16699), .Z(n16696) );
  XOR U18640 ( .A(n16697), .B(n16700), .Z(n16698) );
  IV U18641 ( .A(n16679), .Z(n16683) );
  XOR U18642 ( .A(n16679), .B(n16661), .Z(n16681) );
  XOR U18643 ( .A(n16701), .B(n16702), .Z(n16661) );
  AND U18644 ( .A(n510), .B(n16703), .Z(n16701) );
  XOR U18645 ( .A(n16704), .B(n16702), .Z(n16703) );
  NANDN U18646 ( .A(n16663), .B(n16665), .Z(n16679) );
  XOR U18647 ( .A(n16705), .B(n16706), .Z(n16665) );
  AND U18648 ( .A(n510), .B(n16707), .Z(n16705) );
  XOR U18649 ( .A(n16706), .B(n16708), .Z(n16707) );
  XOR U18650 ( .A(n16709), .B(n16710), .Z(n510) );
  AND U18651 ( .A(n16711), .B(n16712), .Z(n16709) );
  XNOR U18652 ( .A(n16710), .B(n16676), .Z(n16712) );
  XNOR U18653 ( .A(n16713), .B(n16714), .Z(n16676) );
  ANDN U18654 ( .B(n16715), .A(n16716), .Z(n16713) );
  XOR U18655 ( .A(n16714), .B(n16717), .Z(n16715) );
  XOR U18656 ( .A(n16710), .B(n16678), .Z(n16711) );
  XOR U18657 ( .A(n16718), .B(n16719), .Z(n16678) );
  AND U18658 ( .A(n514), .B(n16720), .Z(n16718) );
  XOR U18659 ( .A(n16721), .B(n16719), .Z(n16720) );
  XNOR U18660 ( .A(n16722), .B(n16723), .Z(n16710) );
  NAND U18661 ( .A(n16724), .B(n16725), .Z(n16723) );
  XOR U18662 ( .A(n16726), .B(n16702), .Z(n16725) );
  XOR U18663 ( .A(n16716), .B(n16717), .Z(n16702) );
  XOR U18664 ( .A(n16727), .B(n16728), .Z(n16717) );
  ANDN U18665 ( .B(n16729), .A(n16730), .Z(n16727) );
  XOR U18666 ( .A(n16728), .B(n16731), .Z(n16729) );
  XOR U18667 ( .A(n16732), .B(n16733), .Z(n16716) );
  XOR U18668 ( .A(n16734), .B(n16735), .Z(n16733) );
  ANDN U18669 ( .B(n16736), .A(n16737), .Z(n16734) );
  XOR U18670 ( .A(n16738), .B(n16735), .Z(n16736) );
  IV U18671 ( .A(n16714), .Z(n16732) );
  XOR U18672 ( .A(n16739), .B(n16740), .Z(n16714) );
  ANDN U18673 ( .B(n16741), .A(n16742), .Z(n16739) );
  XOR U18674 ( .A(n16740), .B(n16743), .Z(n16741) );
  IV U18675 ( .A(n16722), .Z(n16726) );
  XOR U18676 ( .A(n16722), .B(n16704), .Z(n16724) );
  XOR U18677 ( .A(n16744), .B(n16745), .Z(n16704) );
  AND U18678 ( .A(n514), .B(n16746), .Z(n16744) );
  XOR U18679 ( .A(n16747), .B(n16745), .Z(n16746) );
  NANDN U18680 ( .A(n16706), .B(n16708), .Z(n16722) );
  XOR U18681 ( .A(n16748), .B(n16749), .Z(n16708) );
  AND U18682 ( .A(n514), .B(n16750), .Z(n16748) );
  XOR U18683 ( .A(n16749), .B(n16751), .Z(n16750) );
  XOR U18684 ( .A(n16752), .B(n16753), .Z(n514) );
  AND U18685 ( .A(n16754), .B(n16755), .Z(n16752) );
  XNOR U18686 ( .A(n16753), .B(n16719), .Z(n16755) );
  XNOR U18687 ( .A(n16756), .B(n16757), .Z(n16719) );
  ANDN U18688 ( .B(n16758), .A(n16759), .Z(n16756) );
  XOR U18689 ( .A(n16757), .B(n16760), .Z(n16758) );
  XOR U18690 ( .A(n16753), .B(n16721), .Z(n16754) );
  XOR U18691 ( .A(n16761), .B(n16762), .Z(n16721) );
  AND U18692 ( .A(n518), .B(n16763), .Z(n16761) );
  XOR U18693 ( .A(n16764), .B(n16762), .Z(n16763) );
  XNOR U18694 ( .A(n16765), .B(n16766), .Z(n16753) );
  NAND U18695 ( .A(n16767), .B(n16768), .Z(n16766) );
  XOR U18696 ( .A(n16769), .B(n16745), .Z(n16768) );
  XOR U18697 ( .A(n16759), .B(n16760), .Z(n16745) );
  XOR U18698 ( .A(n16770), .B(n16771), .Z(n16760) );
  ANDN U18699 ( .B(n16772), .A(n16773), .Z(n16770) );
  XOR U18700 ( .A(n16771), .B(n16774), .Z(n16772) );
  XOR U18701 ( .A(n16775), .B(n16776), .Z(n16759) );
  XOR U18702 ( .A(n16777), .B(n16778), .Z(n16776) );
  ANDN U18703 ( .B(n16779), .A(n16780), .Z(n16777) );
  XOR U18704 ( .A(n16781), .B(n16778), .Z(n16779) );
  IV U18705 ( .A(n16757), .Z(n16775) );
  XOR U18706 ( .A(n16782), .B(n16783), .Z(n16757) );
  ANDN U18707 ( .B(n16784), .A(n16785), .Z(n16782) );
  XOR U18708 ( .A(n16783), .B(n16786), .Z(n16784) );
  IV U18709 ( .A(n16765), .Z(n16769) );
  XOR U18710 ( .A(n16765), .B(n16747), .Z(n16767) );
  XOR U18711 ( .A(n16787), .B(n16788), .Z(n16747) );
  AND U18712 ( .A(n518), .B(n16789), .Z(n16787) );
  XOR U18713 ( .A(n16790), .B(n16788), .Z(n16789) );
  NANDN U18714 ( .A(n16749), .B(n16751), .Z(n16765) );
  XOR U18715 ( .A(n16791), .B(n16792), .Z(n16751) );
  AND U18716 ( .A(n518), .B(n16793), .Z(n16791) );
  XOR U18717 ( .A(n16792), .B(n16794), .Z(n16793) );
  XOR U18718 ( .A(n16795), .B(n16796), .Z(n518) );
  AND U18719 ( .A(n16797), .B(n16798), .Z(n16795) );
  XNOR U18720 ( .A(n16796), .B(n16762), .Z(n16798) );
  XNOR U18721 ( .A(n16799), .B(n16800), .Z(n16762) );
  ANDN U18722 ( .B(n16801), .A(n16802), .Z(n16799) );
  XOR U18723 ( .A(n16800), .B(n16803), .Z(n16801) );
  XOR U18724 ( .A(n16796), .B(n16764), .Z(n16797) );
  XOR U18725 ( .A(n16804), .B(n16805), .Z(n16764) );
  AND U18726 ( .A(n522), .B(n16806), .Z(n16804) );
  XOR U18727 ( .A(n16807), .B(n16805), .Z(n16806) );
  XNOR U18728 ( .A(n16808), .B(n16809), .Z(n16796) );
  NAND U18729 ( .A(n16810), .B(n16811), .Z(n16809) );
  XOR U18730 ( .A(n16812), .B(n16788), .Z(n16811) );
  XOR U18731 ( .A(n16802), .B(n16803), .Z(n16788) );
  XOR U18732 ( .A(n16813), .B(n16814), .Z(n16803) );
  ANDN U18733 ( .B(n16815), .A(n16816), .Z(n16813) );
  XOR U18734 ( .A(n16814), .B(n16817), .Z(n16815) );
  XOR U18735 ( .A(n16818), .B(n16819), .Z(n16802) );
  XOR U18736 ( .A(n16820), .B(n16821), .Z(n16819) );
  ANDN U18737 ( .B(n16822), .A(n16823), .Z(n16820) );
  XOR U18738 ( .A(n16824), .B(n16821), .Z(n16822) );
  IV U18739 ( .A(n16800), .Z(n16818) );
  XOR U18740 ( .A(n16825), .B(n16826), .Z(n16800) );
  ANDN U18741 ( .B(n16827), .A(n16828), .Z(n16825) );
  XOR U18742 ( .A(n16826), .B(n16829), .Z(n16827) );
  IV U18743 ( .A(n16808), .Z(n16812) );
  XOR U18744 ( .A(n16808), .B(n16790), .Z(n16810) );
  XOR U18745 ( .A(n16830), .B(n16831), .Z(n16790) );
  AND U18746 ( .A(n522), .B(n16832), .Z(n16830) );
  XOR U18747 ( .A(n16833), .B(n16831), .Z(n16832) );
  NANDN U18748 ( .A(n16792), .B(n16794), .Z(n16808) );
  XOR U18749 ( .A(n16834), .B(n16835), .Z(n16794) );
  AND U18750 ( .A(n522), .B(n16836), .Z(n16834) );
  XOR U18751 ( .A(n16835), .B(n16837), .Z(n16836) );
  XOR U18752 ( .A(n16838), .B(n16839), .Z(n522) );
  AND U18753 ( .A(n16840), .B(n16841), .Z(n16838) );
  XNOR U18754 ( .A(n16839), .B(n16805), .Z(n16841) );
  XNOR U18755 ( .A(n16842), .B(n16843), .Z(n16805) );
  ANDN U18756 ( .B(n16844), .A(n16845), .Z(n16842) );
  XOR U18757 ( .A(n16843), .B(n16846), .Z(n16844) );
  XOR U18758 ( .A(n16839), .B(n16807), .Z(n16840) );
  XOR U18759 ( .A(n16847), .B(n16848), .Z(n16807) );
  AND U18760 ( .A(n526), .B(n16849), .Z(n16847) );
  XOR U18761 ( .A(n16850), .B(n16848), .Z(n16849) );
  XNOR U18762 ( .A(n16851), .B(n16852), .Z(n16839) );
  NAND U18763 ( .A(n16853), .B(n16854), .Z(n16852) );
  XOR U18764 ( .A(n16855), .B(n16831), .Z(n16854) );
  XOR U18765 ( .A(n16845), .B(n16846), .Z(n16831) );
  XOR U18766 ( .A(n16856), .B(n16857), .Z(n16846) );
  ANDN U18767 ( .B(n16858), .A(n16859), .Z(n16856) );
  XOR U18768 ( .A(n16857), .B(n16860), .Z(n16858) );
  XOR U18769 ( .A(n16861), .B(n16862), .Z(n16845) );
  XOR U18770 ( .A(n16863), .B(n16864), .Z(n16862) );
  ANDN U18771 ( .B(n16865), .A(n16866), .Z(n16863) );
  XOR U18772 ( .A(n16867), .B(n16864), .Z(n16865) );
  IV U18773 ( .A(n16843), .Z(n16861) );
  XOR U18774 ( .A(n16868), .B(n16869), .Z(n16843) );
  ANDN U18775 ( .B(n16870), .A(n16871), .Z(n16868) );
  XOR U18776 ( .A(n16869), .B(n16872), .Z(n16870) );
  IV U18777 ( .A(n16851), .Z(n16855) );
  XOR U18778 ( .A(n16851), .B(n16833), .Z(n16853) );
  XOR U18779 ( .A(n16873), .B(n16874), .Z(n16833) );
  AND U18780 ( .A(n526), .B(n16875), .Z(n16873) );
  XOR U18781 ( .A(n16876), .B(n16874), .Z(n16875) );
  NANDN U18782 ( .A(n16835), .B(n16837), .Z(n16851) );
  XOR U18783 ( .A(n16877), .B(n16878), .Z(n16837) );
  AND U18784 ( .A(n526), .B(n16879), .Z(n16877) );
  XOR U18785 ( .A(n16878), .B(n16880), .Z(n16879) );
  XOR U18786 ( .A(n16881), .B(n16882), .Z(n526) );
  AND U18787 ( .A(n16883), .B(n16884), .Z(n16881) );
  XNOR U18788 ( .A(n16882), .B(n16848), .Z(n16884) );
  XNOR U18789 ( .A(n16885), .B(n16886), .Z(n16848) );
  ANDN U18790 ( .B(n16887), .A(n16888), .Z(n16885) );
  XOR U18791 ( .A(n16886), .B(n16889), .Z(n16887) );
  XOR U18792 ( .A(n16882), .B(n16850), .Z(n16883) );
  XOR U18793 ( .A(n16890), .B(n16891), .Z(n16850) );
  AND U18794 ( .A(n530), .B(n16892), .Z(n16890) );
  XOR U18795 ( .A(n16893), .B(n16891), .Z(n16892) );
  XNOR U18796 ( .A(n16894), .B(n16895), .Z(n16882) );
  NAND U18797 ( .A(n16896), .B(n16897), .Z(n16895) );
  XOR U18798 ( .A(n16898), .B(n16874), .Z(n16897) );
  XOR U18799 ( .A(n16888), .B(n16889), .Z(n16874) );
  XOR U18800 ( .A(n16899), .B(n16900), .Z(n16889) );
  ANDN U18801 ( .B(n16901), .A(n16902), .Z(n16899) );
  XOR U18802 ( .A(n16900), .B(n16903), .Z(n16901) );
  XOR U18803 ( .A(n16904), .B(n16905), .Z(n16888) );
  XOR U18804 ( .A(n16906), .B(n16907), .Z(n16905) );
  ANDN U18805 ( .B(n16908), .A(n16909), .Z(n16906) );
  XOR U18806 ( .A(n16910), .B(n16907), .Z(n16908) );
  IV U18807 ( .A(n16886), .Z(n16904) );
  XOR U18808 ( .A(n16911), .B(n16912), .Z(n16886) );
  ANDN U18809 ( .B(n16913), .A(n16914), .Z(n16911) );
  XOR U18810 ( .A(n16912), .B(n16915), .Z(n16913) );
  IV U18811 ( .A(n16894), .Z(n16898) );
  XOR U18812 ( .A(n16894), .B(n16876), .Z(n16896) );
  XOR U18813 ( .A(n16916), .B(n16917), .Z(n16876) );
  AND U18814 ( .A(n530), .B(n16918), .Z(n16916) );
  XOR U18815 ( .A(n16919), .B(n16917), .Z(n16918) );
  NANDN U18816 ( .A(n16878), .B(n16880), .Z(n16894) );
  XOR U18817 ( .A(n16920), .B(n16921), .Z(n16880) );
  AND U18818 ( .A(n530), .B(n16922), .Z(n16920) );
  XOR U18819 ( .A(n16921), .B(n16923), .Z(n16922) );
  XOR U18820 ( .A(n16924), .B(n16925), .Z(n530) );
  AND U18821 ( .A(n16926), .B(n16927), .Z(n16924) );
  XNOR U18822 ( .A(n16925), .B(n16891), .Z(n16927) );
  XNOR U18823 ( .A(n16928), .B(n16929), .Z(n16891) );
  ANDN U18824 ( .B(n16930), .A(n16931), .Z(n16928) );
  XOR U18825 ( .A(n16929), .B(n16932), .Z(n16930) );
  XOR U18826 ( .A(n16925), .B(n16893), .Z(n16926) );
  XOR U18827 ( .A(n16933), .B(n16934), .Z(n16893) );
  AND U18828 ( .A(n534), .B(n16935), .Z(n16933) );
  XOR U18829 ( .A(n16936), .B(n16934), .Z(n16935) );
  XNOR U18830 ( .A(n16937), .B(n16938), .Z(n16925) );
  NAND U18831 ( .A(n16939), .B(n16940), .Z(n16938) );
  XOR U18832 ( .A(n16941), .B(n16917), .Z(n16940) );
  XOR U18833 ( .A(n16931), .B(n16932), .Z(n16917) );
  XOR U18834 ( .A(n16942), .B(n16943), .Z(n16932) );
  ANDN U18835 ( .B(n16944), .A(n16945), .Z(n16942) );
  XOR U18836 ( .A(n16943), .B(n16946), .Z(n16944) );
  XOR U18837 ( .A(n16947), .B(n16948), .Z(n16931) );
  XOR U18838 ( .A(n16949), .B(n16950), .Z(n16948) );
  ANDN U18839 ( .B(n16951), .A(n16952), .Z(n16949) );
  XOR U18840 ( .A(n16953), .B(n16950), .Z(n16951) );
  IV U18841 ( .A(n16929), .Z(n16947) );
  XOR U18842 ( .A(n16954), .B(n16955), .Z(n16929) );
  ANDN U18843 ( .B(n16956), .A(n16957), .Z(n16954) );
  XOR U18844 ( .A(n16955), .B(n16958), .Z(n16956) );
  IV U18845 ( .A(n16937), .Z(n16941) );
  XOR U18846 ( .A(n16937), .B(n16919), .Z(n16939) );
  XOR U18847 ( .A(n16959), .B(n16960), .Z(n16919) );
  AND U18848 ( .A(n534), .B(n16961), .Z(n16959) );
  XOR U18849 ( .A(n16962), .B(n16960), .Z(n16961) );
  NANDN U18850 ( .A(n16921), .B(n16923), .Z(n16937) );
  XOR U18851 ( .A(n16963), .B(n16964), .Z(n16923) );
  AND U18852 ( .A(n534), .B(n16965), .Z(n16963) );
  XOR U18853 ( .A(n16964), .B(n16966), .Z(n16965) );
  XOR U18854 ( .A(n16967), .B(n16968), .Z(n534) );
  AND U18855 ( .A(n16969), .B(n16970), .Z(n16967) );
  XNOR U18856 ( .A(n16968), .B(n16934), .Z(n16970) );
  XNOR U18857 ( .A(n16971), .B(n16972), .Z(n16934) );
  ANDN U18858 ( .B(n16973), .A(n16974), .Z(n16971) );
  XOR U18859 ( .A(n16972), .B(n16975), .Z(n16973) );
  XOR U18860 ( .A(n16968), .B(n16936), .Z(n16969) );
  XOR U18861 ( .A(n16976), .B(n16977), .Z(n16936) );
  AND U18862 ( .A(n538), .B(n16978), .Z(n16976) );
  XOR U18863 ( .A(n16979), .B(n16977), .Z(n16978) );
  XNOR U18864 ( .A(n16980), .B(n16981), .Z(n16968) );
  NAND U18865 ( .A(n16982), .B(n16983), .Z(n16981) );
  XOR U18866 ( .A(n16984), .B(n16960), .Z(n16983) );
  XOR U18867 ( .A(n16974), .B(n16975), .Z(n16960) );
  XOR U18868 ( .A(n16985), .B(n16986), .Z(n16975) );
  ANDN U18869 ( .B(n16987), .A(n16988), .Z(n16985) );
  XOR U18870 ( .A(n16986), .B(n16989), .Z(n16987) );
  XOR U18871 ( .A(n16990), .B(n16991), .Z(n16974) );
  XOR U18872 ( .A(n16992), .B(n16993), .Z(n16991) );
  ANDN U18873 ( .B(n16994), .A(n16995), .Z(n16992) );
  XOR U18874 ( .A(n16996), .B(n16993), .Z(n16994) );
  IV U18875 ( .A(n16972), .Z(n16990) );
  XOR U18876 ( .A(n16997), .B(n16998), .Z(n16972) );
  ANDN U18877 ( .B(n16999), .A(n17000), .Z(n16997) );
  XOR U18878 ( .A(n16998), .B(n17001), .Z(n16999) );
  IV U18879 ( .A(n16980), .Z(n16984) );
  XOR U18880 ( .A(n16980), .B(n16962), .Z(n16982) );
  XOR U18881 ( .A(n17002), .B(n17003), .Z(n16962) );
  AND U18882 ( .A(n538), .B(n17004), .Z(n17002) );
  XOR U18883 ( .A(n17005), .B(n17003), .Z(n17004) );
  NANDN U18884 ( .A(n16964), .B(n16966), .Z(n16980) );
  XOR U18885 ( .A(n17006), .B(n17007), .Z(n16966) );
  AND U18886 ( .A(n538), .B(n17008), .Z(n17006) );
  XOR U18887 ( .A(n17007), .B(n17009), .Z(n17008) );
  XOR U18888 ( .A(n17010), .B(n17011), .Z(n538) );
  AND U18889 ( .A(n17012), .B(n17013), .Z(n17010) );
  XNOR U18890 ( .A(n17011), .B(n16977), .Z(n17013) );
  XNOR U18891 ( .A(n17014), .B(n17015), .Z(n16977) );
  ANDN U18892 ( .B(n17016), .A(n17017), .Z(n17014) );
  XOR U18893 ( .A(n17015), .B(n17018), .Z(n17016) );
  XOR U18894 ( .A(n17011), .B(n16979), .Z(n17012) );
  XOR U18895 ( .A(n17019), .B(n17020), .Z(n16979) );
  AND U18896 ( .A(n542), .B(n17021), .Z(n17019) );
  XOR U18897 ( .A(n17022), .B(n17020), .Z(n17021) );
  XNOR U18898 ( .A(n17023), .B(n17024), .Z(n17011) );
  NAND U18899 ( .A(n17025), .B(n17026), .Z(n17024) );
  XOR U18900 ( .A(n17027), .B(n17003), .Z(n17026) );
  XOR U18901 ( .A(n17017), .B(n17018), .Z(n17003) );
  XOR U18902 ( .A(n17028), .B(n17029), .Z(n17018) );
  ANDN U18903 ( .B(n17030), .A(n17031), .Z(n17028) );
  XOR U18904 ( .A(n17029), .B(n17032), .Z(n17030) );
  XOR U18905 ( .A(n17033), .B(n17034), .Z(n17017) );
  XOR U18906 ( .A(n17035), .B(n17036), .Z(n17034) );
  ANDN U18907 ( .B(n17037), .A(n17038), .Z(n17035) );
  XOR U18908 ( .A(n17039), .B(n17036), .Z(n17037) );
  IV U18909 ( .A(n17015), .Z(n17033) );
  XOR U18910 ( .A(n17040), .B(n17041), .Z(n17015) );
  ANDN U18911 ( .B(n17042), .A(n17043), .Z(n17040) );
  XOR U18912 ( .A(n17041), .B(n17044), .Z(n17042) );
  IV U18913 ( .A(n17023), .Z(n17027) );
  XOR U18914 ( .A(n17023), .B(n17005), .Z(n17025) );
  XOR U18915 ( .A(n17045), .B(n17046), .Z(n17005) );
  AND U18916 ( .A(n542), .B(n17047), .Z(n17045) );
  XOR U18917 ( .A(n17048), .B(n17046), .Z(n17047) );
  NANDN U18918 ( .A(n17007), .B(n17009), .Z(n17023) );
  XOR U18919 ( .A(n17049), .B(n17050), .Z(n17009) );
  AND U18920 ( .A(n542), .B(n17051), .Z(n17049) );
  XOR U18921 ( .A(n17050), .B(n17052), .Z(n17051) );
  XOR U18922 ( .A(n17053), .B(n17054), .Z(n542) );
  AND U18923 ( .A(n17055), .B(n17056), .Z(n17053) );
  XNOR U18924 ( .A(n17054), .B(n17020), .Z(n17056) );
  XNOR U18925 ( .A(n17057), .B(n17058), .Z(n17020) );
  ANDN U18926 ( .B(n17059), .A(n17060), .Z(n17057) );
  XOR U18927 ( .A(n17058), .B(n17061), .Z(n17059) );
  XOR U18928 ( .A(n17054), .B(n17022), .Z(n17055) );
  XOR U18929 ( .A(n17062), .B(n17063), .Z(n17022) );
  AND U18930 ( .A(n546), .B(n17064), .Z(n17062) );
  XOR U18931 ( .A(n17065), .B(n17063), .Z(n17064) );
  XNOR U18932 ( .A(n17066), .B(n17067), .Z(n17054) );
  NAND U18933 ( .A(n17068), .B(n17069), .Z(n17067) );
  XOR U18934 ( .A(n17070), .B(n17046), .Z(n17069) );
  XOR U18935 ( .A(n17060), .B(n17061), .Z(n17046) );
  XOR U18936 ( .A(n17071), .B(n17072), .Z(n17061) );
  ANDN U18937 ( .B(n17073), .A(n17074), .Z(n17071) );
  XOR U18938 ( .A(n17072), .B(n17075), .Z(n17073) );
  XOR U18939 ( .A(n17076), .B(n17077), .Z(n17060) );
  XOR U18940 ( .A(n17078), .B(n17079), .Z(n17077) );
  ANDN U18941 ( .B(n17080), .A(n17081), .Z(n17078) );
  XOR U18942 ( .A(n17082), .B(n17079), .Z(n17080) );
  IV U18943 ( .A(n17058), .Z(n17076) );
  XOR U18944 ( .A(n17083), .B(n17084), .Z(n17058) );
  ANDN U18945 ( .B(n17085), .A(n17086), .Z(n17083) );
  XOR U18946 ( .A(n17084), .B(n17087), .Z(n17085) );
  IV U18947 ( .A(n17066), .Z(n17070) );
  XOR U18948 ( .A(n17066), .B(n17048), .Z(n17068) );
  XOR U18949 ( .A(n17088), .B(n17089), .Z(n17048) );
  AND U18950 ( .A(n546), .B(n17090), .Z(n17088) );
  XOR U18951 ( .A(n17091), .B(n17089), .Z(n17090) );
  NANDN U18952 ( .A(n17050), .B(n17052), .Z(n17066) );
  XOR U18953 ( .A(n17092), .B(n17093), .Z(n17052) );
  AND U18954 ( .A(n546), .B(n17094), .Z(n17092) );
  XOR U18955 ( .A(n17093), .B(n17095), .Z(n17094) );
  XOR U18956 ( .A(n17096), .B(n17097), .Z(n546) );
  AND U18957 ( .A(n17098), .B(n17099), .Z(n17096) );
  XNOR U18958 ( .A(n17097), .B(n17063), .Z(n17099) );
  XNOR U18959 ( .A(n17100), .B(n17101), .Z(n17063) );
  ANDN U18960 ( .B(n17102), .A(n17103), .Z(n17100) );
  XOR U18961 ( .A(n17101), .B(n17104), .Z(n17102) );
  XOR U18962 ( .A(n17097), .B(n17065), .Z(n17098) );
  XOR U18963 ( .A(n17105), .B(n17106), .Z(n17065) );
  AND U18964 ( .A(n550), .B(n17107), .Z(n17105) );
  XOR U18965 ( .A(n17108), .B(n17106), .Z(n17107) );
  XNOR U18966 ( .A(n17109), .B(n17110), .Z(n17097) );
  NAND U18967 ( .A(n17111), .B(n17112), .Z(n17110) );
  XOR U18968 ( .A(n17113), .B(n17089), .Z(n17112) );
  XOR U18969 ( .A(n17103), .B(n17104), .Z(n17089) );
  XOR U18970 ( .A(n17114), .B(n17115), .Z(n17104) );
  ANDN U18971 ( .B(n17116), .A(n17117), .Z(n17114) );
  XOR U18972 ( .A(n17115), .B(n17118), .Z(n17116) );
  XOR U18973 ( .A(n17119), .B(n17120), .Z(n17103) );
  XOR U18974 ( .A(n17121), .B(n17122), .Z(n17120) );
  ANDN U18975 ( .B(n17123), .A(n17124), .Z(n17121) );
  XOR U18976 ( .A(n17125), .B(n17122), .Z(n17123) );
  IV U18977 ( .A(n17101), .Z(n17119) );
  XOR U18978 ( .A(n17126), .B(n17127), .Z(n17101) );
  ANDN U18979 ( .B(n17128), .A(n17129), .Z(n17126) );
  XOR U18980 ( .A(n17127), .B(n17130), .Z(n17128) );
  IV U18981 ( .A(n17109), .Z(n17113) );
  XOR U18982 ( .A(n17109), .B(n17091), .Z(n17111) );
  XOR U18983 ( .A(n17131), .B(n17132), .Z(n17091) );
  AND U18984 ( .A(n550), .B(n17133), .Z(n17131) );
  XOR U18985 ( .A(n17134), .B(n17132), .Z(n17133) );
  NANDN U18986 ( .A(n17093), .B(n17095), .Z(n17109) );
  XOR U18987 ( .A(n17135), .B(n17136), .Z(n17095) );
  AND U18988 ( .A(n550), .B(n17137), .Z(n17135) );
  XOR U18989 ( .A(n17136), .B(n17138), .Z(n17137) );
  XOR U18990 ( .A(n17139), .B(n17140), .Z(n550) );
  AND U18991 ( .A(n17141), .B(n17142), .Z(n17139) );
  XNOR U18992 ( .A(n17140), .B(n17106), .Z(n17142) );
  XNOR U18993 ( .A(n17143), .B(n17144), .Z(n17106) );
  ANDN U18994 ( .B(n17145), .A(n17146), .Z(n17143) );
  XOR U18995 ( .A(n17144), .B(n17147), .Z(n17145) );
  XOR U18996 ( .A(n17140), .B(n17108), .Z(n17141) );
  XOR U18997 ( .A(n17148), .B(n17149), .Z(n17108) );
  AND U18998 ( .A(n554), .B(n17150), .Z(n17148) );
  XOR U18999 ( .A(n17151), .B(n17149), .Z(n17150) );
  XNOR U19000 ( .A(n17152), .B(n17153), .Z(n17140) );
  NAND U19001 ( .A(n17154), .B(n17155), .Z(n17153) );
  XOR U19002 ( .A(n17156), .B(n17132), .Z(n17155) );
  XOR U19003 ( .A(n17146), .B(n17147), .Z(n17132) );
  XOR U19004 ( .A(n17157), .B(n17158), .Z(n17147) );
  ANDN U19005 ( .B(n17159), .A(n17160), .Z(n17157) );
  XOR U19006 ( .A(n17158), .B(n17161), .Z(n17159) );
  XOR U19007 ( .A(n17162), .B(n17163), .Z(n17146) );
  XOR U19008 ( .A(n17164), .B(n17165), .Z(n17163) );
  ANDN U19009 ( .B(n17166), .A(n17167), .Z(n17164) );
  XOR U19010 ( .A(n17168), .B(n17165), .Z(n17166) );
  IV U19011 ( .A(n17144), .Z(n17162) );
  XOR U19012 ( .A(n17169), .B(n17170), .Z(n17144) );
  ANDN U19013 ( .B(n17171), .A(n17172), .Z(n17169) );
  XOR U19014 ( .A(n17170), .B(n17173), .Z(n17171) );
  IV U19015 ( .A(n17152), .Z(n17156) );
  XOR U19016 ( .A(n17152), .B(n17134), .Z(n17154) );
  XOR U19017 ( .A(n17174), .B(n17175), .Z(n17134) );
  AND U19018 ( .A(n554), .B(n17176), .Z(n17174) );
  XOR U19019 ( .A(n17177), .B(n17175), .Z(n17176) );
  NANDN U19020 ( .A(n17136), .B(n17138), .Z(n17152) );
  XOR U19021 ( .A(n17178), .B(n17179), .Z(n17138) );
  AND U19022 ( .A(n554), .B(n17180), .Z(n17178) );
  XOR U19023 ( .A(n17179), .B(n17181), .Z(n17180) );
  XOR U19024 ( .A(n17182), .B(n17183), .Z(n554) );
  AND U19025 ( .A(n17184), .B(n17185), .Z(n17182) );
  XNOR U19026 ( .A(n17183), .B(n17149), .Z(n17185) );
  XNOR U19027 ( .A(n17186), .B(n17187), .Z(n17149) );
  ANDN U19028 ( .B(n17188), .A(n17189), .Z(n17186) );
  XOR U19029 ( .A(n17187), .B(n17190), .Z(n17188) );
  XOR U19030 ( .A(n17183), .B(n17151), .Z(n17184) );
  XOR U19031 ( .A(n17191), .B(n17192), .Z(n17151) );
  AND U19032 ( .A(n558), .B(n17193), .Z(n17191) );
  XOR U19033 ( .A(n17194), .B(n17192), .Z(n17193) );
  XNOR U19034 ( .A(n17195), .B(n17196), .Z(n17183) );
  NAND U19035 ( .A(n17197), .B(n17198), .Z(n17196) );
  XOR U19036 ( .A(n17199), .B(n17175), .Z(n17198) );
  XOR U19037 ( .A(n17189), .B(n17190), .Z(n17175) );
  XOR U19038 ( .A(n17200), .B(n17201), .Z(n17190) );
  ANDN U19039 ( .B(n17202), .A(n17203), .Z(n17200) );
  XOR U19040 ( .A(n17201), .B(n17204), .Z(n17202) );
  XOR U19041 ( .A(n17205), .B(n17206), .Z(n17189) );
  XOR U19042 ( .A(n17207), .B(n17208), .Z(n17206) );
  ANDN U19043 ( .B(n17209), .A(n17210), .Z(n17207) );
  XOR U19044 ( .A(n17211), .B(n17208), .Z(n17209) );
  IV U19045 ( .A(n17187), .Z(n17205) );
  XOR U19046 ( .A(n17212), .B(n17213), .Z(n17187) );
  ANDN U19047 ( .B(n17214), .A(n17215), .Z(n17212) );
  XOR U19048 ( .A(n17213), .B(n17216), .Z(n17214) );
  IV U19049 ( .A(n17195), .Z(n17199) );
  XOR U19050 ( .A(n17195), .B(n17177), .Z(n17197) );
  XOR U19051 ( .A(n17217), .B(n17218), .Z(n17177) );
  AND U19052 ( .A(n558), .B(n17219), .Z(n17217) );
  XOR U19053 ( .A(n17220), .B(n17218), .Z(n17219) );
  NANDN U19054 ( .A(n17179), .B(n17181), .Z(n17195) );
  XOR U19055 ( .A(n17221), .B(n17222), .Z(n17181) );
  AND U19056 ( .A(n558), .B(n17223), .Z(n17221) );
  XOR U19057 ( .A(n17222), .B(n17224), .Z(n17223) );
  XOR U19058 ( .A(n17225), .B(n17226), .Z(n558) );
  AND U19059 ( .A(n17227), .B(n17228), .Z(n17225) );
  XNOR U19060 ( .A(n17226), .B(n17192), .Z(n17228) );
  XNOR U19061 ( .A(n17229), .B(n17230), .Z(n17192) );
  ANDN U19062 ( .B(n17231), .A(n17232), .Z(n17229) );
  XOR U19063 ( .A(n17230), .B(n17233), .Z(n17231) );
  XOR U19064 ( .A(n17226), .B(n17194), .Z(n17227) );
  XOR U19065 ( .A(n17234), .B(n17235), .Z(n17194) );
  AND U19066 ( .A(n562), .B(n17236), .Z(n17234) );
  XOR U19067 ( .A(n17237), .B(n17235), .Z(n17236) );
  XNOR U19068 ( .A(n17238), .B(n17239), .Z(n17226) );
  NAND U19069 ( .A(n17240), .B(n17241), .Z(n17239) );
  XOR U19070 ( .A(n17242), .B(n17218), .Z(n17241) );
  XOR U19071 ( .A(n17232), .B(n17233), .Z(n17218) );
  XOR U19072 ( .A(n17243), .B(n17244), .Z(n17233) );
  ANDN U19073 ( .B(n17245), .A(n17246), .Z(n17243) );
  XOR U19074 ( .A(n17244), .B(n17247), .Z(n17245) );
  XOR U19075 ( .A(n17248), .B(n17249), .Z(n17232) );
  XOR U19076 ( .A(n17250), .B(n17251), .Z(n17249) );
  ANDN U19077 ( .B(n17252), .A(n17253), .Z(n17250) );
  XOR U19078 ( .A(n17254), .B(n17251), .Z(n17252) );
  IV U19079 ( .A(n17230), .Z(n17248) );
  XOR U19080 ( .A(n17255), .B(n17256), .Z(n17230) );
  ANDN U19081 ( .B(n17257), .A(n17258), .Z(n17255) );
  XOR U19082 ( .A(n17256), .B(n17259), .Z(n17257) );
  IV U19083 ( .A(n17238), .Z(n17242) );
  XOR U19084 ( .A(n17238), .B(n17220), .Z(n17240) );
  XOR U19085 ( .A(n17260), .B(n17261), .Z(n17220) );
  AND U19086 ( .A(n562), .B(n17262), .Z(n17260) );
  XOR U19087 ( .A(n17263), .B(n17261), .Z(n17262) );
  NANDN U19088 ( .A(n17222), .B(n17224), .Z(n17238) );
  XOR U19089 ( .A(n17264), .B(n17265), .Z(n17224) );
  AND U19090 ( .A(n562), .B(n17266), .Z(n17264) );
  XOR U19091 ( .A(n17265), .B(n17267), .Z(n17266) );
  XOR U19092 ( .A(n17268), .B(n17269), .Z(n562) );
  AND U19093 ( .A(n17270), .B(n17271), .Z(n17268) );
  XNOR U19094 ( .A(n17269), .B(n17235), .Z(n17271) );
  XNOR U19095 ( .A(n17272), .B(n17273), .Z(n17235) );
  ANDN U19096 ( .B(n17274), .A(n17275), .Z(n17272) );
  XOR U19097 ( .A(n17273), .B(n17276), .Z(n17274) );
  XOR U19098 ( .A(n17269), .B(n17237), .Z(n17270) );
  XOR U19099 ( .A(n17277), .B(n17278), .Z(n17237) );
  AND U19100 ( .A(n566), .B(n17279), .Z(n17277) );
  XOR U19101 ( .A(n17280), .B(n17278), .Z(n17279) );
  XNOR U19102 ( .A(n17281), .B(n17282), .Z(n17269) );
  NAND U19103 ( .A(n17283), .B(n17284), .Z(n17282) );
  XOR U19104 ( .A(n17285), .B(n17261), .Z(n17284) );
  XOR U19105 ( .A(n17275), .B(n17276), .Z(n17261) );
  XOR U19106 ( .A(n17286), .B(n17287), .Z(n17276) );
  ANDN U19107 ( .B(n17288), .A(n17289), .Z(n17286) );
  XOR U19108 ( .A(n17287), .B(n17290), .Z(n17288) );
  XOR U19109 ( .A(n17291), .B(n17292), .Z(n17275) );
  XOR U19110 ( .A(n17293), .B(n17294), .Z(n17292) );
  ANDN U19111 ( .B(n17295), .A(n17296), .Z(n17293) );
  XOR U19112 ( .A(n17297), .B(n17294), .Z(n17295) );
  IV U19113 ( .A(n17273), .Z(n17291) );
  XOR U19114 ( .A(n17298), .B(n17299), .Z(n17273) );
  ANDN U19115 ( .B(n17300), .A(n17301), .Z(n17298) );
  XOR U19116 ( .A(n17299), .B(n17302), .Z(n17300) );
  IV U19117 ( .A(n17281), .Z(n17285) );
  XOR U19118 ( .A(n17281), .B(n17263), .Z(n17283) );
  XOR U19119 ( .A(n17303), .B(n17304), .Z(n17263) );
  AND U19120 ( .A(n566), .B(n17305), .Z(n17303) );
  XOR U19121 ( .A(n17306), .B(n17304), .Z(n17305) );
  NANDN U19122 ( .A(n17265), .B(n17267), .Z(n17281) );
  XOR U19123 ( .A(n17307), .B(n17308), .Z(n17267) );
  AND U19124 ( .A(n566), .B(n17309), .Z(n17307) );
  XOR U19125 ( .A(n17308), .B(n17310), .Z(n17309) );
  XOR U19126 ( .A(n17311), .B(n17312), .Z(n566) );
  AND U19127 ( .A(n17313), .B(n17314), .Z(n17311) );
  XNOR U19128 ( .A(n17312), .B(n17278), .Z(n17314) );
  XNOR U19129 ( .A(n17315), .B(n17316), .Z(n17278) );
  ANDN U19130 ( .B(n17317), .A(n17318), .Z(n17315) );
  XOR U19131 ( .A(n17316), .B(n17319), .Z(n17317) );
  XOR U19132 ( .A(n17312), .B(n17280), .Z(n17313) );
  XOR U19133 ( .A(n17320), .B(n17321), .Z(n17280) );
  AND U19134 ( .A(n570), .B(n17322), .Z(n17320) );
  XOR U19135 ( .A(n17323), .B(n17321), .Z(n17322) );
  XNOR U19136 ( .A(n17324), .B(n17325), .Z(n17312) );
  NAND U19137 ( .A(n17326), .B(n17327), .Z(n17325) );
  XOR U19138 ( .A(n17328), .B(n17304), .Z(n17327) );
  XOR U19139 ( .A(n17318), .B(n17319), .Z(n17304) );
  XOR U19140 ( .A(n17329), .B(n17330), .Z(n17319) );
  ANDN U19141 ( .B(n17331), .A(n17332), .Z(n17329) );
  XOR U19142 ( .A(n17330), .B(n17333), .Z(n17331) );
  XOR U19143 ( .A(n17334), .B(n17335), .Z(n17318) );
  XOR U19144 ( .A(n17336), .B(n17337), .Z(n17335) );
  ANDN U19145 ( .B(n17338), .A(n17339), .Z(n17336) );
  XOR U19146 ( .A(n17340), .B(n17337), .Z(n17338) );
  IV U19147 ( .A(n17316), .Z(n17334) );
  XOR U19148 ( .A(n17341), .B(n17342), .Z(n17316) );
  ANDN U19149 ( .B(n17343), .A(n17344), .Z(n17341) );
  XOR U19150 ( .A(n17342), .B(n17345), .Z(n17343) );
  IV U19151 ( .A(n17324), .Z(n17328) );
  XOR U19152 ( .A(n17324), .B(n17306), .Z(n17326) );
  XOR U19153 ( .A(n17346), .B(n17347), .Z(n17306) );
  AND U19154 ( .A(n570), .B(n17348), .Z(n17346) );
  XOR U19155 ( .A(n17349), .B(n17347), .Z(n17348) );
  NANDN U19156 ( .A(n17308), .B(n17310), .Z(n17324) );
  XOR U19157 ( .A(n17350), .B(n17351), .Z(n17310) );
  AND U19158 ( .A(n570), .B(n17352), .Z(n17350) );
  XOR U19159 ( .A(n17351), .B(n17353), .Z(n17352) );
  XOR U19160 ( .A(n17354), .B(n17355), .Z(n570) );
  AND U19161 ( .A(n17356), .B(n17357), .Z(n17354) );
  XNOR U19162 ( .A(n17355), .B(n17321), .Z(n17357) );
  XNOR U19163 ( .A(n17358), .B(n17359), .Z(n17321) );
  ANDN U19164 ( .B(n17360), .A(n17361), .Z(n17358) );
  XOR U19165 ( .A(n17359), .B(n17362), .Z(n17360) );
  XOR U19166 ( .A(n17355), .B(n17323), .Z(n17356) );
  XOR U19167 ( .A(n17363), .B(n17364), .Z(n17323) );
  AND U19168 ( .A(n574), .B(n17365), .Z(n17363) );
  XOR U19169 ( .A(n17366), .B(n17364), .Z(n17365) );
  XNOR U19170 ( .A(n17367), .B(n17368), .Z(n17355) );
  NAND U19171 ( .A(n17369), .B(n17370), .Z(n17368) );
  XOR U19172 ( .A(n17371), .B(n17347), .Z(n17370) );
  XOR U19173 ( .A(n17361), .B(n17362), .Z(n17347) );
  XOR U19174 ( .A(n17372), .B(n17373), .Z(n17362) );
  ANDN U19175 ( .B(n17374), .A(n17375), .Z(n17372) );
  XOR U19176 ( .A(n17373), .B(n17376), .Z(n17374) );
  XOR U19177 ( .A(n17377), .B(n17378), .Z(n17361) );
  XOR U19178 ( .A(n17379), .B(n17380), .Z(n17378) );
  ANDN U19179 ( .B(n17381), .A(n17382), .Z(n17379) );
  XOR U19180 ( .A(n17383), .B(n17380), .Z(n17381) );
  IV U19181 ( .A(n17359), .Z(n17377) );
  XOR U19182 ( .A(n17384), .B(n17385), .Z(n17359) );
  ANDN U19183 ( .B(n17386), .A(n17387), .Z(n17384) );
  XOR U19184 ( .A(n17385), .B(n17388), .Z(n17386) );
  IV U19185 ( .A(n17367), .Z(n17371) );
  XOR U19186 ( .A(n17367), .B(n17349), .Z(n17369) );
  XOR U19187 ( .A(n17389), .B(n17390), .Z(n17349) );
  AND U19188 ( .A(n574), .B(n17391), .Z(n17389) );
  XOR U19189 ( .A(n17392), .B(n17390), .Z(n17391) );
  NANDN U19190 ( .A(n17351), .B(n17353), .Z(n17367) );
  XOR U19191 ( .A(n17393), .B(n17394), .Z(n17353) );
  AND U19192 ( .A(n574), .B(n17395), .Z(n17393) );
  XOR U19193 ( .A(n17394), .B(n17396), .Z(n17395) );
  XOR U19194 ( .A(n17397), .B(n17398), .Z(n574) );
  AND U19195 ( .A(n17399), .B(n17400), .Z(n17397) );
  XNOR U19196 ( .A(n17398), .B(n17364), .Z(n17400) );
  XNOR U19197 ( .A(n17401), .B(n17402), .Z(n17364) );
  ANDN U19198 ( .B(n17403), .A(n17404), .Z(n17401) );
  XOR U19199 ( .A(n17402), .B(n17405), .Z(n17403) );
  XOR U19200 ( .A(n17398), .B(n17366), .Z(n17399) );
  XOR U19201 ( .A(n17406), .B(n17407), .Z(n17366) );
  AND U19202 ( .A(n578), .B(n17408), .Z(n17406) );
  XOR U19203 ( .A(n17409), .B(n17407), .Z(n17408) );
  XNOR U19204 ( .A(n17410), .B(n17411), .Z(n17398) );
  NAND U19205 ( .A(n17412), .B(n17413), .Z(n17411) );
  XOR U19206 ( .A(n17414), .B(n17390), .Z(n17413) );
  XOR U19207 ( .A(n17404), .B(n17405), .Z(n17390) );
  XOR U19208 ( .A(n17415), .B(n17416), .Z(n17405) );
  ANDN U19209 ( .B(n17417), .A(n17418), .Z(n17415) );
  XOR U19210 ( .A(n17416), .B(n17419), .Z(n17417) );
  XOR U19211 ( .A(n17420), .B(n17421), .Z(n17404) );
  XOR U19212 ( .A(n17422), .B(n17423), .Z(n17421) );
  ANDN U19213 ( .B(n17424), .A(n17425), .Z(n17422) );
  XOR U19214 ( .A(n17426), .B(n17423), .Z(n17424) );
  IV U19215 ( .A(n17402), .Z(n17420) );
  XOR U19216 ( .A(n17427), .B(n17428), .Z(n17402) );
  ANDN U19217 ( .B(n17429), .A(n17430), .Z(n17427) );
  XOR U19218 ( .A(n17428), .B(n17431), .Z(n17429) );
  IV U19219 ( .A(n17410), .Z(n17414) );
  XOR U19220 ( .A(n17410), .B(n17392), .Z(n17412) );
  XOR U19221 ( .A(n17432), .B(n17433), .Z(n17392) );
  AND U19222 ( .A(n578), .B(n17434), .Z(n17432) );
  XOR U19223 ( .A(n17435), .B(n17433), .Z(n17434) );
  NANDN U19224 ( .A(n17394), .B(n17396), .Z(n17410) );
  XOR U19225 ( .A(n17436), .B(n17437), .Z(n17396) );
  AND U19226 ( .A(n578), .B(n17438), .Z(n17436) );
  XOR U19227 ( .A(n17437), .B(n17439), .Z(n17438) );
  XOR U19228 ( .A(n17440), .B(n17441), .Z(n578) );
  AND U19229 ( .A(n17442), .B(n17443), .Z(n17440) );
  XNOR U19230 ( .A(n17441), .B(n17407), .Z(n17443) );
  XNOR U19231 ( .A(n17444), .B(n17445), .Z(n17407) );
  ANDN U19232 ( .B(n17446), .A(n17447), .Z(n17444) );
  XOR U19233 ( .A(n17445), .B(n17448), .Z(n17446) );
  XOR U19234 ( .A(n17441), .B(n17409), .Z(n17442) );
  XOR U19235 ( .A(n17449), .B(n17450), .Z(n17409) );
  AND U19236 ( .A(n582), .B(n17451), .Z(n17449) );
  XOR U19237 ( .A(n17452), .B(n17450), .Z(n17451) );
  XNOR U19238 ( .A(n17453), .B(n17454), .Z(n17441) );
  NAND U19239 ( .A(n17455), .B(n17456), .Z(n17454) );
  XOR U19240 ( .A(n17457), .B(n17433), .Z(n17456) );
  XOR U19241 ( .A(n17447), .B(n17448), .Z(n17433) );
  XOR U19242 ( .A(n17458), .B(n17459), .Z(n17448) );
  ANDN U19243 ( .B(n17460), .A(n17461), .Z(n17458) );
  XOR U19244 ( .A(n17459), .B(n17462), .Z(n17460) );
  XOR U19245 ( .A(n17463), .B(n17464), .Z(n17447) );
  XOR U19246 ( .A(n17465), .B(n17466), .Z(n17464) );
  ANDN U19247 ( .B(n17467), .A(n17468), .Z(n17465) );
  XOR U19248 ( .A(n17469), .B(n17466), .Z(n17467) );
  IV U19249 ( .A(n17445), .Z(n17463) );
  XOR U19250 ( .A(n17470), .B(n17471), .Z(n17445) );
  ANDN U19251 ( .B(n17472), .A(n17473), .Z(n17470) );
  XOR U19252 ( .A(n17471), .B(n17474), .Z(n17472) );
  IV U19253 ( .A(n17453), .Z(n17457) );
  XOR U19254 ( .A(n17453), .B(n17435), .Z(n17455) );
  XOR U19255 ( .A(n17475), .B(n17476), .Z(n17435) );
  AND U19256 ( .A(n582), .B(n17477), .Z(n17475) );
  XOR U19257 ( .A(n17478), .B(n17476), .Z(n17477) );
  NANDN U19258 ( .A(n17437), .B(n17439), .Z(n17453) );
  XOR U19259 ( .A(n17479), .B(n17480), .Z(n17439) );
  AND U19260 ( .A(n582), .B(n17481), .Z(n17479) );
  XOR U19261 ( .A(n17480), .B(n17482), .Z(n17481) );
  XOR U19262 ( .A(n17483), .B(n17484), .Z(n582) );
  AND U19263 ( .A(n17485), .B(n17486), .Z(n17483) );
  XNOR U19264 ( .A(n17484), .B(n17450), .Z(n17486) );
  XNOR U19265 ( .A(n17487), .B(n17488), .Z(n17450) );
  ANDN U19266 ( .B(n17489), .A(n17490), .Z(n17487) );
  XOR U19267 ( .A(n17488), .B(n17491), .Z(n17489) );
  XOR U19268 ( .A(n17484), .B(n17452), .Z(n17485) );
  XOR U19269 ( .A(n17492), .B(n17493), .Z(n17452) );
  AND U19270 ( .A(n586), .B(n17494), .Z(n17492) );
  XOR U19271 ( .A(n17495), .B(n17493), .Z(n17494) );
  XNOR U19272 ( .A(n17496), .B(n17497), .Z(n17484) );
  NAND U19273 ( .A(n17498), .B(n17499), .Z(n17497) );
  XOR U19274 ( .A(n17500), .B(n17476), .Z(n17499) );
  XOR U19275 ( .A(n17490), .B(n17491), .Z(n17476) );
  XOR U19276 ( .A(n17501), .B(n17502), .Z(n17491) );
  ANDN U19277 ( .B(n17503), .A(n17504), .Z(n17501) );
  XOR U19278 ( .A(n17502), .B(n17505), .Z(n17503) );
  XOR U19279 ( .A(n17506), .B(n17507), .Z(n17490) );
  XOR U19280 ( .A(n17508), .B(n17509), .Z(n17507) );
  ANDN U19281 ( .B(n17510), .A(n17511), .Z(n17508) );
  XOR U19282 ( .A(n17512), .B(n17509), .Z(n17510) );
  IV U19283 ( .A(n17488), .Z(n17506) );
  XOR U19284 ( .A(n17513), .B(n17514), .Z(n17488) );
  ANDN U19285 ( .B(n17515), .A(n17516), .Z(n17513) );
  XOR U19286 ( .A(n17514), .B(n17517), .Z(n17515) );
  IV U19287 ( .A(n17496), .Z(n17500) );
  XOR U19288 ( .A(n17496), .B(n17478), .Z(n17498) );
  XOR U19289 ( .A(n17518), .B(n17519), .Z(n17478) );
  AND U19290 ( .A(n586), .B(n17520), .Z(n17518) );
  XOR U19291 ( .A(n17521), .B(n17519), .Z(n17520) );
  NANDN U19292 ( .A(n17480), .B(n17482), .Z(n17496) );
  XOR U19293 ( .A(n17522), .B(n17523), .Z(n17482) );
  AND U19294 ( .A(n586), .B(n17524), .Z(n17522) );
  XOR U19295 ( .A(n17523), .B(n17525), .Z(n17524) );
  XOR U19296 ( .A(n17526), .B(n17527), .Z(n586) );
  AND U19297 ( .A(n17528), .B(n17529), .Z(n17526) );
  XNOR U19298 ( .A(n17527), .B(n17493), .Z(n17529) );
  XNOR U19299 ( .A(n17530), .B(n17531), .Z(n17493) );
  ANDN U19300 ( .B(n17532), .A(n17533), .Z(n17530) );
  XOR U19301 ( .A(n17531), .B(n17534), .Z(n17532) );
  XOR U19302 ( .A(n17527), .B(n17495), .Z(n17528) );
  XOR U19303 ( .A(n17535), .B(n17536), .Z(n17495) );
  AND U19304 ( .A(n590), .B(n17537), .Z(n17535) );
  XOR U19305 ( .A(n17538), .B(n17536), .Z(n17537) );
  XNOR U19306 ( .A(n17539), .B(n17540), .Z(n17527) );
  NAND U19307 ( .A(n17541), .B(n17542), .Z(n17540) );
  XOR U19308 ( .A(n17543), .B(n17519), .Z(n17542) );
  XOR U19309 ( .A(n17533), .B(n17534), .Z(n17519) );
  XOR U19310 ( .A(n17544), .B(n17545), .Z(n17534) );
  ANDN U19311 ( .B(n17546), .A(n17547), .Z(n17544) );
  XOR U19312 ( .A(n17545), .B(n17548), .Z(n17546) );
  XOR U19313 ( .A(n17549), .B(n17550), .Z(n17533) );
  XOR U19314 ( .A(n17551), .B(n17552), .Z(n17550) );
  ANDN U19315 ( .B(n17553), .A(n17554), .Z(n17551) );
  XOR U19316 ( .A(n17555), .B(n17552), .Z(n17553) );
  IV U19317 ( .A(n17531), .Z(n17549) );
  XOR U19318 ( .A(n17556), .B(n17557), .Z(n17531) );
  ANDN U19319 ( .B(n17558), .A(n17559), .Z(n17556) );
  XOR U19320 ( .A(n17557), .B(n17560), .Z(n17558) );
  IV U19321 ( .A(n17539), .Z(n17543) );
  XOR U19322 ( .A(n17539), .B(n17521), .Z(n17541) );
  XOR U19323 ( .A(n17561), .B(n17562), .Z(n17521) );
  AND U19324 ( .A(n590), .B(n17563), .Z(n17561) );
  XOR U19325 ( .A(n17564), .B(n17562), .Z(n17563) );
  NANDN U19326 ( .A(n17523), .B(n17525), .Z(n17539) );
  XOR U19327 ( .A(n17565), .B(n17566), .Z(n17525) );
  AND U19328 ( .A(n590), .B(n17567), .Z(n17565) );
  XOR U19329 ( .A(n17566), .B(n17568), .Z(n17567) );
  XOR U19330 ( .A(n17569), .B(n17570), .Z(n590) );
  AND U19331 ( .A(n17571), .B(n17572), .Z(n17569) );
  XNOR U19332 ( .A(n17570), .B(n17536), .Z(n17572) );
  XNOR U19333 ( .A(n17573), .B(n17574), .Z(n17536) );
  ANDN U19334 ( .B(n17575), .A(n17576), .Z(n17573) );
  XOR U19335 ( .A(n17574), .B(n17577), .Z(n17575) );
  XOR U19336 ( .A(n17570), .B(n17538), .Z(n17571) );
  XOR U19337 ( .A(n17578), .B(n17579), .Z(n17538) );
  AND U19338 ( .A(n594), .B(n17580), .Z(n17578) );
  XOR U19339 ( .A(n17581), .B(n17579), .Z(n17580) );
  XNOR U19340 ( .A(n17582), .B(n17583), .Z(n17570) );
  NAND U19341 ( .A(n17584), .B(n17585), .Z(n17583) );
  XOR U19342 ( .A(n17586), .B(n17562), .Z(n17585) );
  XOR U19343 ( .A(n17576), .B(n17577), .Z(n17562) );
  XOR U19344 ( .A(n17587), .B(n17588), .Z(n17577) );
  ANDN U19345 ( .B(n17589), .A(n17590), .Z(n17587) );
  XOR U19346 ( .A(n17588), .B(n17591), .Z(n17589) );
  XOR U19347 ( .A(n17592), .B(n17593), .Z(n17576) );
  XOR U19348 ( .A(n17594), .B(n17595), .Z(n17593) );
  ANDN U19349 ( .B(n17596), .A(n17597), .Z(n17594) );
  XOR U19350 ( .A(n17598), .B(n17595), .Z(n17596) );
  IV U19351 ( .A(n17574), .Z(n17592) );
  XOR U19352 ( .A(n17599), .B(n17600), .Z(n17574) );
  ANDN U19353 ( .B(n17601), .A(n17602), .Z(n17599) );
  XOR U19354 ( .A(n17600), .B(n17603), .Z(n17601) );
  IV U19355 ( .A(n17582), .Z(n17586) );
  XOR U19356 ( .A(n17582), .B(n17564), .Z(n17584) );
  XOR U19357 ( .A(n17604), .B(n17605), .Z(n17564) );
  AND U19358 ( .A(n594), .B(n17606), .Z(n17604) );
  XOR U19359 ( .A(n17607), .B(n17605), .Z(n17606) );
  NANDN U19360 ( .A(n17566), .B(n17568), .Z(n17582) );
  XOR U19361 ( .A(n17608), .B(n17609), .Z(n17568) );
  AND U19362 ( .A(n594), .B(n17610), .Z(n17608) );
  XOR U19363 ( .A(n17609), .B(n17611), .Z(n17610) );
  XOR U19364 ( .A(n17612), .B(n17613), .Z(n594) );
  AND U19365 ( .A(n17614), .B(n17615), .Z(n17612) );
  XNOR U19366 ( .A(n17613), .B(n17579), .Z(n17615) );
  XNOR U19367 ( .A(n17616), .B(n17617), .Z(n17579) );
  ANDN U19368 ( .B(n17618), .A(n17619), .Z(n17616) );
  XOR U19369 ( .A(n17617), .B(n17620), .Z(n17618) );
  XOR U19370 ( .A(n17613), .B(n17581), .Z(n17614) );
  XOR U19371 ( .A(n17621), .B(n17622), .Z(n17581) );
  AND U19372 ( .A(n598), .B(n17623), .Z(n17621) );
  XOR U19373 ( .A(n17624), .B(n17622), .Z(n17623) );
  XNOR U19374 ( .A(n17625), .B(n17626), .Z(n17613) );
  NAND U19375 ( .A(n17627), .B(n17628), .Z(n17626) );
  XOR U19376 ( .A(n17629), .B(n17605), .Z(n17628) );
  XOR U19377 ( .A(n17619), .B(n17620), .Z(n17605) );
  XOR U19378 ( .A(n17630), .B(n17631), .Z(n17620) );
  ANDN U19379 ( .B(n17632), .A(n17633), .Z(n17630) );
  XOR U19380 ( .A(n17631), .B(n17634), .Z(n17632) );
  XOR U19381 ( .A(n17635), .B(n17636), .Z(n17619) );
  XOR U19382 ( .A(n17637), .B(n17638), .Z(n17636) );
  ANDN U19383 ( .B(n17639), .A(n17640), .Z(n17637) );
  XOR U19384 ( .A(n17641), .B(n17638), .Z(n17639) );
  IV U19385 ( .A(n17617), .Z(n17635) );
  XOR U19386 ( .A(n17642), .B(n17643), .Z(n17617) );
  ANDN U19387 ( .B(n17644), .A(n17645), .Z(n17642) );
  XOR U19388 ( .A(n17643), .B(n17646), .Z(n17644) );
  IV U19389 ( .A(n17625), .Z(n17629) );
  XOR U19390 ( .A(n17625), .B(n17607), .Z(n17627) );
  XOR U19391 ( .A(n17647), .B(n17648), .Z(n17607) );
  AND U19392 ( .A(n598), .B(n17649), .Z(n17647) );
  XOR U19393 ( .A(n17650), .B(n17648), .Z(n17649) );
  NANDN U19394 ( .A(n17609), .B(n17611), .Z(n17625) );
  XOR U19395 ( .A(n17651), .B(n17652), .Z(n17611) );
  AND U19396 ( .A(n598), .B(n17653), .Z(n17651) );
  XOR U19397 ( .A(n17652), .B(n17654), .Z(n17653) );
  XOR U19398 ( .A(n17655), .B(n17656), .Z(n598) );
  AND U19399 ( .A(n17657), .B(n17658), .Z(n17655) );
  XNOR U19400 ( .A(n17656), .B(n17622), .Z(n17658) );
  XNOR U19401 ( .A(n17659), .B(n17660), .Z(n17622) );
  ANDN U19402 ( .B(n17661), .A(n17662), .Z(n17659) );
  XOR U19403 ( .A(n17660), .B(n17663), .Z(n17661) );
  XOR U19404 ( .A(n17656), .B(n17624), .Z(n17657) );
  XOR U19405 ( .A(n17664), .B(n17665), .Z(n17624) );
  AND U19406 ( .A(n602), .B(n17666), .Z(n17664) );
  XOR U19407 ( .A(n17667), .B(n17665), .Z(n17666) );
  XNOR U19408 ( .A(n17668), .B(n17669), .Z(n17656) );
  NAND U19409 ( .A(n17670), .B(n17671), .Z(n17669) );
  XOR U19410 ( .A(n17672), .B(n17648), .Z(n17671) );
  XOR U19411 ( .A(n17662), .B(n17663), .Z(n17648) );
  XOR U19412 ( .A(n17673), .B(n17674), .Z(n17663) );
  ANDN U19413 ( .B(n17675), .A(n17676), .Z(n17673) );
  XOR U19414 ( .A(n17674), .B(n17677), .Z(n17675) );
  XOR U19415 ( .A(n17678), .B(n17679), .Z(n17662) );
  XOR U19416 ( .A(n17680), .B(n17681), .Z(n17679) );
  ANDN U19417 ( .B(n17682), .A(n17683), .Z(n17680) );
  XOR U19418 ( .A(n17684), .B(n17681), .Z(n17682) );
  IV U19419 ( .A(n17660), .Z(n17678) );
  XOR U19420 ( .A(n17685), .B(n17686), .Z(n17660) );
  ANDN U19421 ( .B(n17687), .A(n17688), .Z(n17685) );
  XOR U19422 ( .A(n17686), .B(n17689), .Z(n17687) );
  IV U19423 ( .A(n17668), .Z(n17672) );
  XOR U19424 ( .A(n17668), .B(n17650), .Z(n17670) );
  XOR U19425 ( .A(n17690), .B(n17691), .Z(n17650) );
  AND U19426 ( .A(n602), .B(n17692), .Z(n17690) );
  XOR U19427 ( .A(n17693), .B(n17691), .Z(n17692) );
  NANDN U19428 ( .A(n17652), .B(n17654), .Z(n17668) );
  XOR U19429 ( .A(n17694), .B(n17695), .Z(n17654) );
  AND U19430 ( .A(n602), .B(n17696), .Z(n17694) );
  XOR U19431 ( .A(n17695), .B(n17697), .Z(n17696) );
  XOR U19432 ( .A(n17698), .B(n17699), .Z(n602) );
  AND U19433 ( .A(n17700), .B(n17701), .Z(n17698) );
  XNOR U19434 ( .A(n17699), .B(n17665), .Z(n17701) );
  XNOR U19435 ( .A(n17702), .B(n17703), .Z(n17665) );
  ANDN U19436 ( .B(n17704), .A(n17705), .Z(n17702) );
  XOR U19437 ( .A(n17703), .B(n17706), .Z(n17704) );
  XOR U19438 ( .A(n17699), .B(n17667), .Z(n17700) );
  XOR U19439 ( .A(n17707), .B(n17708), .Z(n17667) );
  AND U19440 ( .A(n606), .B(n17709), .Z(n17707) );
  XOR U19441 ( .A(n17710), .B(n17708), .Z(n17709) );
  XNOR U19442 ( .A(n17711), .B(n17712), .Z(n17699) );
  NAND U19443 ( .A(n17713), .B(n17714), .Z(n17712) );
  XOR U19444 ( .A(n17715), .B(n17691), .Z(n17714) );
  XOR U19445 ( .A(n17705), .B(n17706), .Z(n17691) );
  XOR U19446 ( .A(n17716), .B(n17717), .Z(n17706) );
  ANDN U19447 ( .B(n17718), .A(n17719), .Z(n17716) );
  XOR U19448 ( .A(n17717), .B(n17720), .Z(n17718) );
  XOR U19449 ( .A(n17721), .B(n17722), .Z(n17705) );
  XOR U19450 ( .A(n17723), .B(n17724), .Z(n17722) );
  ANDN U19451 ( .B(n17725), .A(n17726), .Z(n17723) );
  XOR U19452 ( .A(n17727), .B(n17724), .Z(n17725) );
  IV U19453 ( .A(n17703), .Z(n17721) );
  XOR U19454 ( .A(n17728), .B(n17729), .Z(n17703) );
  ANDN U19455 ( .B(n17730), .A(n17731), .Z(n17728) );
  XOR U19456 ( .A(n17729), .B(n17732), .Z(n17730) );
  IV U19457 ( .A(n17711), .Z(n17715) );
  XOR U19458 ( .A(n17711), .B(n17693), .Z(n17713) );
  XOR U19459 ( .A(n17733), .B(n17734), .Z(n17693) );
  AND U19460 ( .A(n606), .B(n17735), .Z(n17733) );
  XOR U19461 ( .A(n17736), .B(n17734), .Z(n17735) );
  NANDN U19462 ( .A(n17695), .B(n17697), .Z(n17711) );
  XOR U19463 ( .A(n17737), .B(n17738), .Z(n17697) );
  AND U19464 ( .A(n606), .B(n17739), .Z(n17737) );
  XOR U19465 ( .A(n17738), .B(n17740), .Z(n17739) );
  XOR U19466 ( .A(n17741), .B(n17742), .Z(n606) );
  AND U19467 ( .A(n17743), .B(n17744), .Z(n17741) );
  XNOR U19468 ( .A(n17742), .B(n17708), .Z(n17744) );
  XNOR U19469 ( .A(n17745), .B(n17746), .Z(n17708) );
  ANDN U19470 ( .B(n17747), .A(n17748), .Z(n17745) );
  XOR U19471 ( .A(n17746), .B(n17749), .Z(n17747) );
  XOR U19472 ( .A(n17742), .B(n17710), .Z(n17743) );
  XOR U19473 ( .A(n17750), .B(n17751), .Z(n17710) );
  AND U19474 ( .A(n610), .B(n17752), .Z(n17750) );
  XOR U19475 ( .A(n17753), .B(n17751), .Z(n17752) );
  XNOR U19476 ( .A(n17754), .B(n17755), .Z(n17742) );
  NAND U19477 ( .A(n17756), .B(n17757), .Z(n17755) );
  XOR U19478 ( .A(n17758), .B(n17734), .Z(n17757) );
  XOR U19479 ( .A(n17748), .B(n17749), .Z(n17734) );
  XOR U19480 ( .A(n17759), .B(n17760), .Z(n17749) );
  ANDN U19481 ( .B(n17761), .A(n17762), .Z(n17759) );
  XOR U19482 ( .A(n17760), .B(n17763), .Z(n17761) );
  XOR U19483 ( .A(n17764), .B(n17765), .Z(n17748) );
  XOR U19484 ( .A(n17766), .B(n17767), .Z(n17765) );
  ANDN U19485 ( .B(n17768), .A(n17769), .Z(n17766) );
  XOR U19486 ( .A(n17770), .B(n17767), .Z(n17768) );
  IV U19487 ( .A(n17746), .Z(n17764) );
  XOR U19488 ( .A(n17771), .B(n17772), .Z(n17746) );
  ANDN U19489 ( .B(n17773), .A(n17774), .Z(n17771) );
  XOR U19490 ( .A(n17772), .B(n17775), .Z(n17773) );
  IV U19491 ( .A(n17754), .Z(n17758) );
  XOR U19492 ( .A(n17754), .B(n17736), .Z(n17756) );
  XOR U19493 ( .A(n17776), .B(n17777), .Z(n17736) );
  AND U19494 ( .A(n610), .B(n17778), .Z(n17776) );
  XOR U19495 ( .A(n17779), .B(n17777), .Z(n17778) );
  NANDN U19496 ( .A(n17738), .B(n17740), .Z(n17754) );
  XOR U19497 ( .A(n17780), .B(n17781), .Z(n17740) );
  AND U19498 ( .A(n610), .B(n17782), .Z(n17780) );
  XOR U19499 ( .A(n17781), .B(n17783), .Z(n17782) );
  XOR U19500 ( .A(n17784), .B(n17785), .Z(n610) );
  AND U19501 ( .A(n17786), .B(n17787), .Z(n17784) );
  XNOR U19502 ( .A(n17785), .B(n17751), .Z(n17787) );
  XNOR U19503 ( .A(n17788), .B(n17789), .Z(n17751) );
  ANDN U19504 ( .B(n17790), .A(n17791), .Z(n17788) );
  XOR U19505 ( .A(n17789), .B(n17792), .Z(n17790) );
  XOR U19506 ( .A(n17785), .B(n17753), .Z(n17786) );
  XOR U19507 ( .A(n17793), .B(n17794), .Z(n17753) );
  AND U19508 ( .A(n614), .B(n17795), .Z(n17793) );
  XOR U19509 ( .A(n17796), .B(n17794), .Z(n17795) );
  XNOR U19510 ( .A(n17797), .B(n17798), .Z(n17785) );
  NAND U19511 ( .A(n17799), .B(n17800), .Z(n17798) );
  XOR U19512 ( .A(n17801), .B(n17777), .Z(n17800) );
  XOR U19513 ( .A(n17791), .B(n17792), .Z(n17777) );
  XOR U19514 ( .A(n17802), .B(n17803), .Z(n17792) );
  ANDN U19515 ( .B(n17804), .A(n17805), .Z(n17802) );
  XOR U19516 ( .A(n17803), .B(n17806), .Z(n17804) );
  XOR U19517 ( .A(n17807), .B(n17808), .Z(n17791) );
  XOR U19518 ( .A(n17809), .B(n17810), .Z(n17808) );
  ANDN U19519 ( .B(n17811), .A(n17812), .Z(n17809) );
  XOR U19520 ( .A(n17813), .B(n17810), .Z(n17811) );
  IV U19521 ( .A(n17789), .Z(n17807) );
  XOR U19522 ( .A(n17814), .B(n17815), .Z(n17789) );
  ANDN U19523 ( .B(n17816), .A(n17817), .Z(n17814) );
  XOR U19524 ( .A(n17815), .B(n17818), .Z(n17816) );
  IV U19525 ( .A(n17797), .Z(n17801) );
  XOR U19526 ( .A(n17797), .B(n17779), .Z(n17799) );
  XOR U19527 ( .A(n17819), .B(n17820), .Z(n17779) );
  AND U19528 ( .A(n614), .B(n17821), .Z(n17819) );
  XOR U19529 ( .A(n17822), .B(n17820), .Z(n17821) );
  NANDN U19530 ( .A(n17781), .B(n17783), .Z(n17797) );
  XOR U19531 ( .A(n17823), .B(n17824), .Z(n17783) );
  AND U19532 ( .A(n614), .B(n17825), .Z(n17823) );
  XOR U19533 ( .A(n17824), .B(n17826), .Z(n17825) );
  XOR U19534 ( .A(n17827), .B(n17828), .Z(n614) );
  AND U19535 ( .A(n17829), .B(n17830), .Z(n17827) );
  XNOR U19536 ( .A(n17828), .B(n17794), .Z(n17830) );
  XNOR U19537 ( .A(n17831), .B(n17832), .Z(n17794) );
  ANDN U19538 ( .B(n17833), .A(n17834), .Z(n17831) );
  XOR U19539 ( .A(n17832), .B(n17835), .Z(n17833) );
  XOR U19540 ( .A(n17828), .B(n17796), .Z(n17829) );
  XOR U19541 ( .A(n17836), .B(n17837), .Z(n17796) );
  AND U19542 ( .A(n618), .B(n17838), .Z(n17836) );
  XOR U19543 ( .A(n17839), .B(n17837), .Z(n17838) );
  XNOR U19544 ( .A(n17840), .B(n17841), .Z(n17828) );
  NAND U19545 ( .A(n17842), .B(n17843), .Z(n17841) );
  XOR U19546 ( .A(n17844), .B(n17820), .Z(n17843) );
  XOR U19547 ( .A(n17834), .B(n17835), .Z(n17820) );
  XOR U19548 ( .A(n17845), .B(n17846), .Z(n17835) );
  ANDN U19549 ( .B(n17847), .A(n17848), .Z(n17845) );
  XOR U19550 ( .A(n17846), .B(n17849), .Z(n17847) );
  XOR U19551 ( .A(n17850), .B(n17851), .Z(n17834) );
  XOR U19552 ( .A(n17852), .B(n17853), .Z(n17851) );
  ANDN U19553 ( .B(n17854), .A(n17855), .Z(n17852) );
  XOR U19554 ( .A(n17856), .B(n17853), .Z(n17854) );
  IV U19555 ( .A(n17832), .Z(n17850) );
  XOR U19556 ( .A(n17857), .B(n17858), .Z(n17832) );
  ANDN U19557 ( .B(n17859), .A(n17860), .Z(n17857) );
  XOR U19558 ( .A(n17858), .B(n17861), .Z(n17859) );
  IV U19559 ( .A(n17840), .Z(n17844) );
  XOR U19560 ( .A(n17840), .B(n17822), .Z(n17842) );
  XOR U19561 ( .A(n17862), .B(n17863), .Z(n17822) );
  AND U19562 ( .A(n618), .B(n17864), .Z(n17862) );
  XOR U19563 ( .A(n17865), .B(n17863), .Z(n17864) );
  NANDN U19564 ( .A(n17824), .B(n17826), .Z(n17840) );
  XOR U19565 ( .A(n17866), .B(n17867), .Z(n17826) );
  AND U19566 ( .A(n618), .B(n17868), .Z(n17866) );
  XOR U19567 ( .A(n17867), .B(n17869), .Z(n17868) );
  XOR U19568 ( .A(n17870), .B(n17871), .Z(n618) );
  AND U19569 ( .A(n17872), .B(n17873), .Z(n17870) );
  XNOR U19570 ( .A(n17871), .B(n17837), .Z(n17873) );
  XNOR U19571 ( .A(n17874), .B(n17875), .Z(n17837) );
  ANDN U19572 ( .B(n17876), .A(n17877), .Z(n17874) );
  XOR U19573 ( .A(n17875), .B(n17878), .Z(n17876) );
  XOR U19574 ( .A(n17871), .B(n17839), .Z(n17872) );
  XOR U19575 ( .A(n17879), .B(n17880), .Z(n17839) );
  AND U19576 ( .A(n622), .B(n17881), .Z(n17879) );
  XOR U19577 ( .A(n17882), .B(n17880), .Z(n17881) );
  XNOR U19578 ( .A(n17883), .B(n17884), .Z(n17871) );
  NAND U19579 ( .A(n17885), .B(n17886), .Z(n17884) );
  XOR U19580 ( .A(n17887), .B(n17863), .Z(n17886) );
  XOR U19581 ( .A(n17877), .B(n17878), .Z(n17863) );
  XOR U19582 ( .A(n17888), .B(n17889), .Z(n17878) );
  ANDN U19583 ( .B(n17890), .A(n17891), .Z(n17888) );
  XOR U19584 ( .A(n17889), .B(n17892), .Z(n17890) );
  XOR U19585 ( .A(n17893), .B(n17894), .Z(n17877) );
  XOR U19586 ( .A(n17895), .B(n17896), .Z(n17894) );
  ANDN U19587 ( .B(n17897), .A(n17898), .Z(n17895) );
  XOR U19588 ( .A(n17899), .B(n17896), .Z(n17897) );
  IV U19589 ( .A(n17875), .Z(n17893) );
  XOR U19590 ( .A(n17900), .B(n17901), .Z(n17875) );
  ANDN U19591 ( .B(n17902), .A(n17903), .Z(n17900) );
  XOR U19592 ( .A(n17901), .B(n17904), .Z(n17902) );
  IV U19593 ( .A(n17883), .Z(n17887) );
  XOR U19594 ( .A(n17883), .B(n17865), .Z(n17885) );
  XOR U19595 ( .A(n17905), .B(n17906), .Z(n17865) );
  AND U19596 ( .A(n622), .B(n17907), .Z(n17905) );
  XOR U19597 ( .A(n17908), .B(n17906), .Z(n17907) );
  NANDN U19598 ( .A(n17867), .B(n17869), .Z(n17883) );
  XOR U19599 ( .A(n17909), .B(n17910), .Z(n17869) );
  AND U19600 ( .A(n622), .B(n17911), .Z(n17909) );
  XOR U19601 ( .A(n17910), .B(n17912), .Z(n17911) );
  XOR U19602 ( .A(n17913), .B(n17914), .Z(n622) );
  AND U19603 ( .A(n17915), .B(n17916), .Z(n17913) );
  XNOR U19604 ( .A(n17914), .B(n17880), .Z(n17916) );
  XNOR U19605 ( .A(n17917), .B(n17918), .Z(n17880) );
  ANDN U19606 ( .B(n17919), .A(n17920), .Z(n17917) );
  XOR U19607 ( .A(n17918), .B(n17921), .Z(n17919) );
  XOR U19608 ( .A(n17914), .B(n17882), .Z(n17915) );
  XOR U19609 ( .A(n17922), .B(n17923), .Z(n17882) );
  AND U19610 ( .A(n626), .B(n17924), .Z(n17922) );
  XOR U19611 ( .A(n17925), .B(n17923), .Z(n17924) );
  XNOR U19612 ( .A(n17926), .B(n17927), .Z(n17914) );
  NAND U19613 ( .A(n17928), .B(n17929), .Z(n17927) );
  XOR U19614 ( .A(n17930), .B(n17906), .Z(n17929) );
  XOR U19615 ( .A(n17920), .B(n17921), .Z(n17906) );
  XOR U19616 ( .A(n17931), .B(n17932), .Z(n17921) );
  ANDN U19617 ( .B(n17933), .A(n17934), .Z(n17931) );
  XOR U19618 ( .A(n17932), .B(n17935), .Z(n17933) );
  XOR U19619 ( .A(n17936), .B(n17937), .Z(n17920) );
  XOR U19620 ( .A(n17938), .B(n17939), .Z(n17937) );
  ANDN U19621 ( .B(n17940), .A(n17941), .Z(n17938) );
  XOR U19622 ( .A(n17942), .B(n17939), .Z(n17940) );
  IV U19623 ( .A(n17918), .Z(n17936) );
  XOR U19624 ( .A(n17943), .B(n17944), .Z(n17918) );
  ANDN U19625 ( .B(n17945), .A(n17946), .Z(n17943) );
  XOR U19626 ( .A(n17944), .B(n17947), .Z(n17945) );
  IV U19627 ( .A(n17926), .Z(n17930) );
  XOR U19628 ( .A(n17926), .B(n17908), .Z(n17928) );
  XOR U19629 ( .A(n17948), .B(n17949), .Z(n17908) );
  AND U19630 ( .A(n626), .B(n17950), .Z(n17948) );
  XOR U19631 ( .A(n17951), .B(n17949), .Z(n17950) );
  NANDN U19632 ( .A(n17910), .B(n17912), .Z(n17926) );
  XOR U19633 ( .A(n17952), .B(n17953), .Z(n17912) );
  AND U19634 ( .A(n626), .B(n17954), .Z(n17952) );
  XOR U19635 ( .A(n17953), .B(n17955), .Z(n17954) );
  XOR U19636 ( .A(n17956), .B(n17957), .Z(n626) );
  AND U19637 ( .A(n17958), .B(n17959), .Z(n17956) );
  XNOR U19638 ( .A(n17957), .B(n17923), .Z(n17959) );
  XNOR U19639 ( .A(n17960), .B(n17961), .Z(n17923) );
  ANDN U19640 ( .B(n17962), .A(n17963), .Z(n17960) );
  XOR U19641 ( .A(n17961), .B(n17964), .Z(n17962) );
  XOR U19642 ( .A(n17957), .B(n17925), .Z(n17958) );
  XOR U19643 ( .A(n17965), .B(n17966), .Z(n17925) );
  AND U19644 ( .A(n630), .B(n17967), .Z(n17965) );
  XOR U19645 ( .A(n17968), .B(n17966), .Z(n17967) );
  XNOR U19646 ( .A(n17969), .B(n17970), .Z(n17957) );
  NAND U19647 ( .A(n17971), .B(n17972), .Z(n17970) );
  XOR U19648 ( .A(n17973), .B(n17949), .Z(n17972) );
  XOR U19649 ( .A(n17963), .B(n17964), .Z(n17949) );
  XOR U19650 ( .A(n17974), .B(n17975), .Z(n17964) );
  ANDN U19651 ( .B(n17976), .A(n17977), .Z(n17974) );
  XOR U19652 ( .A(n17975), .B(n17978), .Z(n17976) );
  XOR U19653 ( .A(n17979), .B(n17980), .Z(n17963) );
  XOR U19654 ( .A(n17981), .B(n17982), .Z(n17980) );
  ANDN U19655 ( .B(n17983), .A(n17984), .Z(n17981) );
  XOR U19656 ( .A(n17985), .B(n17982), .Z(n17983) );
  IV U19657 ( .A(n17961), .Z(n17979) );
  XOR U19658 ( .A(n17986), .B(n17987), .Z(n17961) );
  ANDN U19659 ( .B(n17988), .A(n17989), .Z(n17986) );
  XOR U19660 ( .A(n17987), .B(n17990), .Z(n17988) );
  IV U19661 ( .A(n17969), .Z(n17973) );
  XOR U19662 ( .A(n17969), .B(n17951), .Z(n17971) );
  XOR U19663 ( .A(n17991), .B(n17992), .Z(n17951) );
  AND U19664 ( .A(n630), .B(n17993), .Z(n17991) );
  XOR U19665 ( .A(n17994), .B(n17992), .Z(n17993) );
  NANDN U19666 ( .A(n17953), .B(n17955), .Z(n17969) );
  XOR U19667 ( .A(n17995), .B(n17996), .Z(n17955) );
  AND U19668 ( .A(n630), .B(n17997), .Z(n17995) );
  XOR U19669 ( .A(n17996), .B(n17998), .Z(n17997) );
  XOR U19670 ( .A(n17999), .B(n18000), .Z(n630) );
  AND U19671 ( .A(n18001), .B(n18002), .Z(n17999) );
  XNOR U19672 ( .A(n18000), .B(n17966), .Z(n18002) );
  XNOR U19673 ( .A(n18003), .B(n18004), .Z(n17966) );
  ANDN U19674 ( .B(n18005), .A(n18006), .Z(n18003) );
  XOR U19675 ( .A(n18004), .B(n18007), .Z(n18005) );
  XOR U19676 ( .A(n18000), .B(n17968), .Z(n18001) );
  XOR U19677 ( .A(n18008), .B(n18009), .Z(n17968) );
  AND U19678 ( .A(n634), .B(n18010), .Z(n18008) );
  XOR U19679 ( .A(n18011), .B(n18009), .Z(n18010) );
  XNOR U19680 ( .A(n18012), .B(n18013), .Z(n18000) );
  NAND U19681 ( .A(n18014), .B(n18015), .Z(n18013) );
  XOR U19682 ( .A(n18016), .B(n17992), .Z(n18015) );
  XOR U19683 ( .A(n18006), .B(n18007), .Z(n17992) );
  XOR U19684 ( .A(n18017), .B(n18018), .Z(n18007) );
  ANDN U19685 ( .B(n18019), .A(n18020), .Z(n18017) );
  XOR U19686 ( .A(n18018), .B(n18021), .Z(n18019) );
  XOR U19687 ( .A(n18022), .B(n18023), .Z(n18006) );
  XOR U19688 ( .A(n18024), .B(n18025), .Z(n18023) );
  ANDN U19689 ( .B(n18026), .A(n18027), .Z(n18024) );
  XOR U19690 ( .A(n18028), .B(n18025), .Z(n18026) );
  IV U19691 ( .A(n18004), .Z(n18022) );
  XOR U19692 ( .A(n18029), .B(n18030), .Z(n18004) );
  ANDN U19693 ( .B(n18031), .A(n18032), .Z(n18029) );
  XOR U19694 ( .A(n18030), .B(n18033), .Z(n18031) );
  IV U19695 ( .A(n18012), .Z(n18016) );
  XOR U19696 ( .A(n18012), .B(n17994), .Z(n18014) );
  XOR U19697 ( .A(n18034), .B(n18035), .Z(n17994) );
  AND U19698 ( .A(n634), .B(n18036), .Z(n18034) );
  XOR U19699 ( .A(n18037), .B(n18035), .Z(n18036) );
  NANDN U19700 ( .A(n17996), .B(n17998), .Z(n18012) );
  XOR U19701 ( .A(n18038), .B(n18039), .Z(n17998) );
  AND U19702 ( .A(n634), .B(n18040), .Z(n18038) );
  XOR U19703 ( .A(n18039), .B(n18041), .Z(n18040) );
  XOR U19704 ( .A(n18042), .B(n18043), .Z(n634) );
  AND U19705 ( .A(n18044), .B(n18045), .Z(n18042) );
  XNOR U19706 ( .A(n18043), .B(n18009), .Z(n18045) );
  XNOR U19707 ( .A(n18046), .B(n18047), .Z(n18009) );
  ANDN U19708 ( .B(n18048), .A(n18049), .Z(n18046) );
  XOR U19709 ( .A(n18047), .B(n18050), .Z(n18048) );
  XOR U19710 ( .A(n18043), .B(n18011), .Z(n18044) );
  XOR U19711 ( .A(n18051), .B(n18052), .Z(n18011) );
  AND U19712 ( .A(n638), .B(n18053), .Z(n18051) );
  XOR U19713 ( .A(n18054), .B(n18052), .Z(n18053) );
  XNOR U19714 ( .A(n18055), .B(n18056), .Z(n18043) );
  NAND U19715 ( .A(n18057), .B(n18058), .Z(n18056) );
  XOR U19716 ( .A(n18059), .B(n18035), .Z(n18058) );
  XOR U19717 ( .A(n18049), .B(n18050), .Z(n18035) );
  XOR U19718 ( .A(n18060), .B(n18061), .Z(n18050) );
  ANDN U19719 ( .B(n18062), .A(n18063), .Z(n18060) );
  XOR U19720 ( .A(n18061), .B(n18064), .Z(n18062) );
  XOR U19721 ( .A(n18065), .B(n18066), .Z(n18049) );
  XOR U19722 ( .A(n18067), .B(n18068), .Z(n18066) );
  ANDN U19723 ( .B(n18069), .A(n18070), .Z(n18067) );
  XOR U19724 ( .A(n18071), .B(n18068), .Z(n18069) );
  IV U19725 ( .A(n18047), .Z(n18065) );
  XOR U19726 ( .A(n18072), .B(n18073), .Z(n18047) );
  ANDN U19727 ( .B(n18074), .A(n18075), .Z(n18072) );
  XOR U19728 ( .A(n18073), .B(n18076), .Z(n18074) );
  IV U19729 ( .A(n18055), .Z(n18059) );
  XOR U19730 ( .A(n18055), .B(n18037), .Z(n18057) );
  XOR U19731 ( .A(n18077), .B(n18078), .Z(n18037) );
  AND U19732 ( .A(n638), .B(n18079), .Z(n18077) );
  XOR U19733 ( .A(n18080), .B(n18078), .Z(n18079) );
  NANDN U19734 ( .A(n18039), .B(n18041), .Z(n18055) );
  XOR U19735 ( .A(n18081), .B(n18082), .Z(n18041) );
  AND U19736 ( .A(n638), .B(n18083), .Z(n18081) );
  XOR U19737 ( .A(n18082), .B(n18084), .Z(n18083) );
  XOR U19738 ( .A(n18085), .B(n18086), .Z(n638) );
  AND U19739 ( .A(n18087), .B(n18088), .Z(n18085) );
  XNOR U19740 ( .A(n18086), .B(n18052), .Z(n18088) );
  XNOR U19741 ( .A(n18089), .B(n18090), .Z(n18052) );
  ANDN U19742 ( .B(n18091), .A(n18092), .Z(n18089) );
  XOR U19743 ( .A(n18090), .B(n18093), .Z(n18091) );
  XOR U19744 ( .A(n18086), .B(n18054), .Z(n18087) );
  XOR U19745 ( .A(n18094), .B(n18095), .Z(n18054) );
  AND U19746 ( .A(n642), .B(n18096), .Z(n18094) );
  XOR U19747 ( .A(n18097), .B(n18095), .Z(n18096) );
  XNOR U19748 ( .A(n18098), .B(n18099), .Z(n18086) );
  NAND U19749 ( .A(n18100), .B(n18101), .Z(n18099) );
  XOR U19750 ( .A(n18102), .B(n18078), .Z(n18101) );
  XOR U19751 ( .A(n18092), .B(n18093), .Z(n18078) );
  XOR U19752 ( .A(n18103), .B(n18104), .Z(n18093) );
  ANDN U19753 ( .B(n18105), .A(n18106), .Z(n18103) );
  XOR U19754 ( .A(n18104), .B(n18107), .Z(n18105) );
  XOR U19755 ( .A(n18108), .B(n18109), .Z(n18092) );
  XOR U19756 ( .A(n18110), .B(n18111), .Z(n18109) );
  ANDN U19757 ( .B(n18112), .A(n18113), .Z(n18110) );
  XOR U19758 ( .A(n18114), .B(n18111), .Z(n18112) );
  IV U19759 ( .A(n18090), .Z(n18108) );
  XOR U19760 ( .A(n18115), .B(n18116), .Z(n18090) );
  ANDN U19761 ( .B(n18117), .A(n18118), .Z(n18115) );
  XOR U19762 ( .A(n18116), .B(n18119), .Z(n18117) );
  IV U19763 ( .A(n18098), .Z(n18102) );
  XOR U19764 ( .A(n18098), .B(n18080), .Z(n18100) );
  XOR U19765 ( .A(n18120), .B(n18121), .Z(n18080) );
  AND U19766 ( .A(n642), .B(n18122), .Z(n18120) );
  XOR U19767 ( .A(n18123), .B(n18121), .Z(n18122) );
  NANDN U19768 ( .A(n18082), .B(n18084), .Z(n18098) );
  XOR U19769 ( .A(n18124), .B(n18125), .Z(n18084) );
  AND U19770 ( .A(n642), .B(n18126), .Z(n18124) );
  XOR U19771 ( .A(n18125), .B(n18127), .Z(n18126) );
  XOR U19772 ( .A(n18128), .B(n18129), .Z(n642) );
  AND U19773 ( .A(n18130), .B(n18131), .Z(n18128) );
  XNOR U19774 ( .A(n18129), .B(n18095), .Z(n18131) );
  XNOR U19775 ( .A(n18132), .B(n18133), .Z(n18095) );
  ANDN U19776 ( .B(n18134), .A(n18135), .Z(n18132) );
  XOR U19777 ( .A(n18133), .B(n18136), .Z(n18134) );
  XOR U19778 ( .A(n18129), .B(n18097), .Z(n18130) );
  XOR U19779 ( .A(n18137), .B(n18138), .Z(n18097) );
  AND U19780 ( .A(n646), .B(n18139), .Z(n18137) );
  XOR U19781 ( .A(n18140), .B(n18138), .Z(n18139) );
  XNOR U19782 ( .A(n18141), .B(n18142), .Z(n18129) );
  NAND U19783 ( .A(n18143), .B(n18144), .Z(n18142) );
  XOR U19784 ( .A(n18145), .B(n18121), .Z(n18144) );
  XOR U19785 ( .A(n18135), .B(n18136), .Z(n18121) );
  XOR U19786 ( .A(n18146), .B(n18147), .Z(n18136) );
  ANDN U19787 ( .B(n18148), .A(n18149), .Z(n18146) );
  XOR U19788 ( .A(n18147), .B(n18150), .Z(n18148) );
  XOR U19789 ( .A(n18151), .B(n18152), .Z(n18135) );
  XOR U19790 ( .A(n18153), .B(n18154), .Z(n18152) );
  ANDN U19791 ( .B(n18155), .A(n18156), .Z(n18153) );
  XOR U19792 ( .A(n18157), .B(n18154), .Z(n18155) );
  IV U19793 ( .A(n18133), .Z(n18151) );
  XOR U19794 ( .A(n18158), .B(n18159), .Z(n18133) );
  ANDN U19795 ( .B(n18160), .A(n18161), .Z(n18158) );
  XOR U19796 ( .A(n18159), .B(n18162), .Z(n18160) );
  IV U19797 ( .A(n18141), .Z(n18145) );
  XOR U19798 ( .A(n18141), .B(n18123), .Z(n18143) );
  XOR U19799 ( .A(n18163), .B(n18164), .Z(n18123) );
  AND U19800 ( .A(n646), .B(n18165), .Z(n18163) );
  XOR U19801 ( .A(n18166), .B(n18164), .Z(n18165) );
  NANDN U19802 ( .A(n18125), .B(n18127), .Z(n18141) );
  XOR U19803 ( .A(n18167), .B(n18168), .Z(n18127) );
  AND U19804 ( .A(n646), .B(n18169), .Z(n18167) );
  XOR U19805 ( .A(n18168), .B(n18170), .Z(n18169) );
  XOR U19806 ( .A(n18171), .B(n18172), .Z(n646) );
  AND U19807 ( .A(n18173), .B(n18174), .Z(n18171) );
  XNOR U19808 ( .A(n18172), .B(n18138), .Z(n18174) );
  XNOR U19809 ( .A(n18175), .B(n18176), .Z(n18138) );
  ANDN U19810 ( .B(n18177), .A(n18178), .Z(n18175) );
  XOR U19811 ( .A(n18176), .B(n18179), .Z(n18177) );
  XOR U19812 ( .A(n18172), .B(n18140), .Z(n18173) );
  XOR U19813 ( .A(n18180), .B(n18181), .Z(n18140) );
  AND U19814 ( .A(n650), .B(n18182), .Z(n18180) );
  XOR U19815 ( .A(n18183), .B(n18181), .Z(n18182) );
  XNOR U19816 ( .A(n18184), .B(n18185), .Z(n18172) );
  NAND U19817 ( .A(n18186), .B(n18187), .Z(n18185) );
  XOR U19818 ( .A(n18188), .B(n18164), .Z(n18187) );
  XOR U19819 ( .A(n18178), .B(n18179), .Z(n18164) );
  XOR U19820 ( .A(n18189), .B(n18190), .Z(n18179) );
  ANDN U19821 ( .B(n18191), .A(n18192), .Z(n18189) );
  XOR U19822 ( .A(n18190), .B(n18193), .Z(n18191) );
  XOR U19823 ( .A(n18194), .B(n18195), .Z(n18178) );
  XOR U19824 ( .A(n18196), .B(n18197), .Z(n18195) );
  ANDN U19825 ( .B(n18198), .A(n18199), .Z(n18196) );
  XOR U19826 ( .A(n18200), .B(n18197), .Z(n18198) );
  IV U19827 ( .A(n18176), .Z(n18194) );
  XOR U19828 ( .A(n18201), .B(n18202), .Z(n18176) );
  ANDN U19829 ( .B(n18203), .A(n18204), .Z(n18201) );
  XOR U19830 ( .A(n18202), .B(n18205), .Z(n18203) );
  IV U19831 ( .A(n18184), .Z(n18188) );
  XOR U19832 ( .A(n18184), .B(n18166), .Z(n18186) );
  XOR U19833 ( .A(n18206), .B(n18207), .Z(n18166) );
  AND U19834 ( .A(n650), .B(n18208), .Z(n18206) );
  XOR U19835 ( .A(n18209), .B(n18207), .Z(n18208) );
  NANDN U19836 ( .A(n18168), .B(n18170), .Z(n18184) );
  XOR U19837 ( .A(n18210), .B(n18211), .Z(n18170) );
  AND U19838 ( .A(n650), .B(n18212), .Z(n18210) );
  XOR U19839 ( .A(n18211), .B(n18213), .Z(n18212) );
  XOR U19840 ( .A(n18214), .B(n18215), .Z(n650) );
  AND U19841 ( .A(n18216), .B(n18217), .Z(n18214) );
  XNOR U19842 ( .A(n18215), .B(n18181), .Z(n18217) );
  XNOR U19843 ( .A(n18218), .B(n18219), .Z(n18181) );
  ANDN U19844 ( .B(n18220), .A(n18221), .Z(n18218) );
  XOR U19845 ( .A(n18219), .B(n18222), .Z(n18220) );
  XOR U19846 ( .A(n18215), .B(n18183), .Z(n18216) );
  XOR U19847 ( .A(n18223), .B(n18224), .Z(n18183) );
  AND U19848 ( .A(n654), .B(n18225), .Z(n18223) );
  XOR U19849 ( .A(n18226), .B(n18224), .Z(n18225) );
  XNOR U19850 ( .A(n18227), .B(n18228), .Z(n18215) );
  NAND U19851 ( .A(n18229), .B(n18230), .Z(n18228) );
  XOR U19852 ( .A(n18231), .B(n18207), .Z(n18230) );
  XOR U19853 ( .A(n18221), .B(n18222), .Z(n18207) );
  XOR U19854 ( .A(n18232), .B(n18233), .Z(n18222) );
  ANDN U19855 ( .B(n18234), .A(n18235), .Z(n18232) );
  XOR U19856 ( .A(n18233), .B(n18236), .Z(n18234) );
  XOR U19857 ( .A(n18237), .B(n18238), .Z(n18221) );
  XOR U19858 ( .A(n18239), .B(n18240), .Z(n18238) );
  ANDN U19859 ( .B(n18241), .A(n18242), .Z(n18239) );
  XOR U19860 ( .A(n18243), .B(n18240), .Z(n18241) );
  IV U19861 ( .A(n18219), .Z(n18237) );
  XOR U19862 ( .A(n18244), .B(n18245), .Z(n18219) );
  ANDN U19863 ( .B(n18246), .A(n18247), .Z(n18244) );
  XOR U19864 ( .A(n18245), .B(n18248), .Z(n18246) );
  IV U19865 ( .A(n18227), .Z(n18231) );
  XOR U19866 ( .A(n18227), .B(n18209), .Z(n18229) );
  XOR U19867 ( .A(n18249), .B(n18250), .Z(n18209) );
  AND U19868 ( .A(n654), .B(n18251), .Z(n18249) );
  XOR U19869 ( .A(n18252), .B(n18250), .Z(n18251) );
  NANDN U19870 ( .A(n18211), .B(n18213), .Z(n18227) );
  XOR U19871 ( .A(n18253), .B(n18254), .Z(n18213) );
  AND U19872 ( .A(n654), .B(n18255), .Z(n18253) );
  XOR U19873 ( .A(n18254), .B(n18256), .Z(n18255) );
  XOR U19874 ( .A(n18257), .B(n18258), .Z(n654) );
  AND U19875 ( .A(n18259), .B(n18260), .Z(n18257) );
  XNOR U19876 ( .A(n18258), .B(n18224), .Z(n18260) );
  XNOR U19877 ( .A(n18261), .B(n18262), .Z(n18224) );
  ANDN U19878 ( .B(n18263), .A(n18264), .Z(n18261) );
  XOR U19879 ( .A(n18262), .B(n18265), .Z(n18263) );
  XOR U19880 ( .A(n18258), .B(n18226), .Z(n18259) );
  XOR U19881 ( .A(n18266), .B(n18267), .Z(n18226) );
  AND U19882 ( .A(n658), .B(n18268), .Z(n18266) );
  XOR U19883 ( .A(n18269), .B(n18267), .Z(n18268) );
  XNOR U19884 ( .A(n18270), .B(n18271), .Z(n18258) );
  NAND U19885 ( .A(n18272), .B(n18273), .Z(n18271) );
  XOR U19886 ( .A(n18274), .B(n18250), .Z(n18273) );
  XOR U19887 ( .A(n18264), .B(n18265), .Z(n18250) );
  XOR U19888 ( .A(n18275), .B(n18276), .Z(n18265) );
  ANDN U19889 ( .B(n18277), .A(n18278), .Z(n18275) );
  XOR U19890 ( .A(n18276), .B(n18279), .Z(n18277) );
  XOR U19891 ( .A(n18280), .B(n18281), .Z(n18264) );
  XOR U19892 ( .A(n18282), .B(n18283), .Z(n18281) );
  ANDN U19893 ( .B(n18284), .A(n18285), .Z(n18282) );
  XOR U19894 ( .A(n18286), .B(n18283), .Z(n18284) );
  IV U19895 ( .A(n18262), .Z(n18280) );
  XOR U19896 ( .A(n18287), .B(n18288), .Z(n18262) );
  ANDN U19897 ( .B(n18289), .A(n18290), .Z(n18287) );
  XOR U19898 ( .A(n18288), .B(n18291), .Z(n18289) );
  IV U19899 ( .A(n18270), .Z(n18274) );
  XOR U19900 ( .A(n18270), .B(n18252), .Z(n18272) );
  XOR U19901 ( .A(n18292), .B(n18293), .Z(n18252) );
  AND U19902 ( .A(n658), .B(n18294), .Z(n18292) );
  XOR U19903 ( .A(n18295), .B(n18293), .Z(n18294) );
  NANDN U19904 ( .A(n18254), .B(n18256), .Z(n18270) );
  XOR U19905 ( .A(n18296), .B(n18297), .Z(n18256) );
  AND U19906 ( .A(n658), .B(n18298), .Z(n18296) );
  XOR U19907 ( .A(n18297), .B(n18299), .Z(n18298) );
  XOR U19908 ( .A(n18300), .B(n18301), .Z(n658) );
  AND U19909 ( .A(n18302), .B(n18303), .Z(n18300) );
  XNOR U19910 ( .A(n18301), .B(n18267), .Z(n18303) );
  XNOR U19911 ( .A(n18304), .B(n18305), .Z(n18267) );
  ANDN U19912 ( .B(n18306), .A(n18307), .Z(n18304) );
  XOR U19913 ( .A(n18305), .B(n18308), .Z(n18306) );
  XOR U19914 ( .A(n18301), .B(n18269), .Z(n18302) );
  XOR U19915 ( .A(n18309), .B(n18310), .Z(n18269) );
  AND U19916 ( .A(n662), .B(n18311), .Z(n18309) );
  XOR U19917 ( .A(n18312), .B(n18310), .Z(n18311) );
  XNOR U19918 ( .A(n18313), .B(n18314), .Z(n18301) );
  NAND U19919 ( .A(n18315), .B(n18316), .Z(n18314) );
  XOR U19920 ( .A(n18317), .B(n18293), .Z(n18316) );
  XOR U19921 ( .A(n18307), .B(n18308), .Z(n18293) );
  XOR U19922 ( .A(n18318), .B(n18319), .Z(n18308) );
  ANDN U19923 ( .B(n18320), .A(n18321), .Z(n18318) );
  XOR U19924 ( .A(n18319), .B(n18322), .Z(n18320) );
  XOR U19925 ( .A(n18323), .B(n18324), .Z(n18307) );
  XOR U19926 ( .A(n18325), .B(n18326), .Z(n18324) );
  ANDN U19927 ( .B(n18327), .A(n18328), .Z(n18325) );
  XOR U19928 ( .A(n18329), .B(n18326), .Z(n18327) );
  IV U19929 ( .A(n18305), .Z(n18323) );
  XOR U19930 ( .A(n18330), .B(n18331), .Z(n18305) );
  ANDN U19931 ( .B(n18332), .A(n18333), .Z(n18330) );
  XOR U19932 ( .A(n18331), .B(n18334), .Z(n18332) );
  IV U19933 ( .A(n18313), .Z(n18317) );
  XOR U19934 ( .A(n18313), .B(n18295), .Z(n18315) );
  XOR U19935 ( .A(n18335), .B(n18336), .Z(n18295) );
  AND U19936 ( .A(n662), .B(n18337), .Z(n18335) );
  XOR U19937 ( .A(n18338), .B(n18336), .Z(n18337) );
  NANDN U19938 ( .A(n18297), .B(n18299), .Z(n18313) );
  XOR U19939 ( .A(n18339), .B(n18340), .Z(n18299) );
  AND U19940 ( .A(n662), .B(n18341), .Z(n18339) );
  XOR U19941 ( .A(n18340), .B(n18342), .Z(n18341) );
  XOR U19942 ( .A(n18343), .B(n18344), .Z(n662) );
  AND U19943 ( .A(n18345), .B(n18346), .Z(n18343) );
  XNOR U19944 ( .A(n18344), .B(n18310), .Z(n18346) );
  XNOR U19945 ( .A(n18347), .B(n18348), .Z(n18310) );
  ANDN U19946 ( .B(n18349), .A(n18350), .Z(n18347) );
  XOR U19947 ( .A(n18348), .B(n18351), .Z(n18349) );
  XOR U19948 ( .A(n18344), .B(n18312), .Z(n18345) );
  XOR U19949 ( .A(n18352), .B(n18353), .Z(n18312) );
  AND U19950 ( .A(n666), .B(n18354), .Z(n18352) );
  XOR U19951 ( .A(n18355), .B(n18353), .Z(n18354) );
  XNOR U19952 ( .A(n18356), .B(n18357), .Z(n18344) );
  NAND U19953 ( .A(n18358), .B(n18359), .Z(n18357) );
  XOR U19954 ( .A(n18360), .B(n18336), .Z(n18359) );
  XOR U19955 ( .A(n18350), .B(n18351), .Z(n18336) );
  XOR U19956 ( .A(n18361), .B(n18362), .Z(n18351) );
  ANDN U19957 ( .B(n18363), .A(n18364), .Z(n18361) );
  XOR U19958 ( .A(n18362), .B(n18365), .Z(n18363) );
  XOR U19959 ( .A(n18366), .B(n18367), .Z(n18350) );
  XOR U19960 ( .A(n18368), .B(n18369), .Z(n18367) );
  ANDN U19961 ( .B(n18370), .A(n18371), .Z(n18368) );
  XOR U19962 ( .A(n18372), .B(n18369), .Z(n18370) );
  IV U19963 ( .A(n18348), .Z(n18366) );
  XOR U19964 ( .A(n18373), .B(n18374), .Z(n18348) );
  ANDN U19965 ( .B(n18375), .A(n18376), .Z(n18373) );
  XOR U19966 ( .A(n18374), .B(n18377), .Z(n18375) );
  IV U19967 ( .A(n18356), .Z(n18360) );
  XOR U19968 ( .A(n18356), .B(n18338), .Z(n18358) );
  XOR U19969 ( .A(n18378), .B(n18379), .Z(n18338) );
  AND U19970 ( .A(n666), .B(n18380), .Z(n18378) );
  XOR U19971 ( .A(n18381), .B(n18379), .Z(n18380) );
  NANDN U19972 ( .A(n18340), .B(n18342), .Z(n18356) );
  XOR U19973 ( .A(n18382), .B(n18383), .Z(n18342) );
  AND U19974 ( .A(n666), .B(n18384), .Z(n18382) );
  XOR U19975 ( .A(n18383), .B(n18385), .Z(n18384) );
  XOR U19976 ( .A(n18386), .B(n18387), .Z(n666) );
  AND U19977 ( .A(n18388), .B(n18389), .Z(n18386) );
  XNOR U19978 ( .A(n18387), .B(n18353), .Z(n18389) );
  XNOR U19979 ( .A(n18390), .B(n18391), .Z(n18353) );
  ANDN U19980 ( .B(n18392), .A(n18393), .Z(n18390) );
  XOR U19981 ( .A(n18391), .B(n18394), .Z(n18392) );
  XOR U19982 ( .A(n18387), .B(n18355), .Z(n18388) );
  XOR U19983 ( .A(n18395), .B(n18396), .Z(n18355) );
  AND U19984 ( .A(n670), .B(n18397), .Z(n18395) );
  XOR U19985 ( .A(n18398), .B(n18396), .Z(n18397) );
  XNOR U19986 ( .A(n18399), .B(n18400), .Z(n18387) );
  NAND U19987 ( .A(n18401), .B(n18402), .Z(n18400) );
  XOR U19988 ( .A(n18403), .B(n18379), .Z(n18402) );
  XOR U19989 ( .A(n18393), .B(n18394), .Z(n18379) );
  XOR U19990 ( .A(n18404), .B(n18405), .Z(n18394) );
  ANDN U19991 ( .B(n18406), .A(n18407), .Z(n18404) );
  XOR U19992 ( .A(n18405), .B(n18408), .Z(n18406) );
  XOR U19993 ( .A(n18409), .B(n18410), .Z(n18393) );
  XOR U19994 ( .A(n18411), .B(n18412), .Z(n18410) );
  ANDN U19995 ( .B(n18413), .A(n18414), .Z(n18411) );
  XOR U19996 ( .A(n18415), .B(n18412), .Z(n18413) );
  IV U19997 ( .A(n18391), .Z(n18409) );
  XOR U19998 ( .A(n18416), .B(n18417), .Z(n18391) );
  ANDN U19999 ( .B(n18418), .A(n18419), .Z(n18416) );
  XOR U20000 ( .A(n18417), .B(n18420), .Z(n18418) );
  IV U20001 ( .A(n18399), .Z(n18403) );
  XOR U20002 ( .A(n18399), .B(n18381), .Z(n18401) );
  XOR U20003 ( .A(n18421), .B(n18422), .Z(n18381) );
  AND U20004 ( .A(n670), .B(n18423), .Z(n18421) );
  XOR U20005 ( .A(n18424), .B(n18422), .Z(n18423) );
  NANDN U20006 ( .A(n18383), .B(n18385), .Z(n18399) );
  XOR U20007 ( .A(n18425), .B(n18426), .Z(n18385) );
  AND U20008 ( .A(n670), .B(n18427), .Z(n18425) );
  XOR U20009 ( .A(n18426), .B(n18428), .Z(n18427) );
  XOR U20010 ( .A(n18429), .B(n18430), .Z(n670) );
  AND U20011 ( .A(n18431), .B(n18432), .Z(n18429) );
  XNOR U20012 ( .A(n18430), .B(n18396), .Z(n18432) );
  XNOR U20013 ( .A(n18433), .B(n18434), .Z(n18396) );
  ANDN U20014 ( .B(n18435), .A(n18436), .Z(n18433) );
  XOR U20015 ( .A(n18434), .B(n18437), .Z(n18435) );
  XOR U20016 ( .A(n18430), .B(n18398), .Z(n18431) );
  XOR U20017 ( .A(n18438), .B(n18439), .Z(n18398) );
  AND U20018 ( .A(n674), .B(n18440), .Z(n18438) );
  XOR U20019 ( .A(n18441), .B(n18439), .Z(n18440) );
  XNOR U20020 ( .A(n18442), .B(n18443), .Z(n18430) );
  NAND U20021 ( .A(n18444), .B(n18445), .Z(n18443) );
  XOR U20022 ( .A(n18446), .B(n18422), .Z(n18445) );
  XOR U20023 ( .A(n18436), .B(n18437), .Z(n18422) );
  XOR U20024 ( .A(n18447), .B(n18448), .Z(n18437) );
  ANDN U20025 ( .B(n18449), .A(n18450), .Z(n18447) );
  XOR U20026 ( .A(n18448), .B(n18451), .Z(n18449) );
  XOR U20027 ( .A(n18452), .B(n18453), .Z(n18436) );
  XOR U20028 ( .A(n18454), .B(n18455), .Z(n18453) );
  ANDN U20029 ( .B(n18456), .A(n18457), .Z(n18454) );
  XOR U20030 ( .A(n18458), .B(n18455), .Z(n18456) );
  IV U20031 ( .A(n18434), .Z(n18452) );
  XOR U20032 ( .A(n18459), .B(n18460), .Z(n18434) );
  ANDN U20033 ( .B(n18461), .A(n18462), .Z(n18459) );
  XOR U20034 ( .A(n18460), .B(n18463), .Z(n18461) );
  IV U20035 ( .A(n18442), .Z(n18446) );
  XOR U20036 ( .A(n18442), .B(n18424), .Z(n18444) );
  XOR U20037 ( .A(n18464), .B(n18465), .Z(n18424) );
  AND U20038 ( .A(n674), .B(n18466), .Z(n18464) );
  XOR U20039 ( .A(n18467), .B(n18465), .Z(n18466) );
  NANDN U20040 ( .A(n18426), .B(n18428), .Z(n18442) );
  XOR U20041 ( .A(n18468), .B(n18469), .Z(n18428) );
  AND U20042 ( .A(n674), .B(n18470), .Z(n18468) );
  XOR U20043 ( .A(n18469), .B(n18471), .Z(n18470) );
  XOR U20044 ( .A(n18472), .B(n18473), .Z(n674) );
  AND U20045 ( .A(n18474), .B(n18475), .Z(n18472) );
  XNOR U20046 ( .A(n18473), .B(n18439), .Z(n18475) );
  XNOR U20047 ( .A(n18476), .B(n18477), .Z(n18439) );
  ANDN U20048 ( .B(n18478), .A(n18479), .Z(n18476) );
  XOR U20049 ( .A(n18477), .B(n18480), .Z(n18478) );
  XOR U20050 ( .A(n18473), .B(n18441), .Z(n18474) );
  XOR U20051 ( .A(n18481), .B(n18482), .Z(n18441) );
  AND U20052 ( .A(n678), .B(n18483), .Z(n18481) );
  XOR U20053 ( .A(n18484), .B(n18482), .Z(n18483) );
  XNOR U20054 ( .A(n18485), .B(n18486), .Z(n18473) );
  NAND U20055 ( .A(n18487), .B(n18488), .Z(n18486) );
  XOR U20056 ( .A(n18489), .B(n18465), .Z(n18488) );
  XOR U20057 ( .A(n18479), .B(n18480), .Z(n18465) );
  XOR U20058 ( .A(n18490), .B(n18491), .Z(n18480) );
  ANDN U20059 ( .B(n18492), .A(n18493), .Z(n18490) );
  XOR U20060 ( .A(n18491), .B(n18494), .Z(n18492) );
  XOR U20061 ( .A(n18495), .B(n18496), .Z(n18479) );
  XOR U20062 ( .A(n18497), .B(n18498), .Z(n18496) );
  ANDN U20063 ( .B(n18499), .A(n18500), .Z(n18497) );
  XOR U20064 ( .A(n18501), .B(n18498), .Z(n18499) );
  IV U20065 ( .A(n18477), .Z(n18495) );
  XOR U20066 ( .A(n18502), .B(n18503), .Z(n18477) );
  ANDN U20067 ( .B(n18504), .A(n18505), .Z(n18502) );
  XOR U20068 ( .A(n18503), .B(n18506), .Z(n18504) );
  IV U20069 ( .A(n18485), .Z(n18489) );
  XOR U20070 ( .A(n18485), .B(n18467), .Z(n18487) );
  XOR U20071 ( .A(n18507), .B(n18508), .Z(n18467) );
  AND U20072 ( .A(n678), .B(n18509), .Z(n18507) );
  XOR U20073 ( .A(n18510), .B(n18508), .Z(n18509) );
  NANDN U20074 ( .A(n18469), .B(n18471), .Z(n18485) );
  XOR U20075 ( .A(n18511), .B(n18512), .Z(n18471) );
  AND U20076 ( .A(n678), .B(n18513), .Z(n18511) );
  XOR U20077 ( .A(n18512), .B(n18514), .Z(n18513) );
  XOR U20078 ( .A(n18515), .B(n18516), .Z(n678) );
  AND U20079 ( .A(n18517), .B(n18518), .Z(n18515) );
  XNOR U20080 ( .A(n18516), .B(n18482), .Z(n18518) );
  XNOR U20081 ( .A(n18519), .B(n18520), .Z(n18482) );
  ANDN U20082 ( .B(n18521), .A(n18522), .Z(n18519) );
  XOR U20083 ( .A(n18520), .B(n18523), .Z(n18521) );
  XOR U20084 ( .A(n18516), .B(n18484), .Z(n18517) );
  XOR U20085 ( .A(n18524), .B(n18525), .Z(n18484) );
  AND U20086 ( .A(n682), .B(n18526), .Z(n18524) );
  XOR U20087 ( .A(n18527), .B(n18525), .Z(n18526) );
  XNOR U20088 ( .A(n18528), .B(n18529), .Z(n18516) );
  NAND U20089 ( .A(n18530), .B(n18531), .Z(n18529) );
  XOR U20090 ( .A(n18532), .B(n18508), .Z(n18531) );
  XOR U20091 ( .A(n18522), .B(n18523), .Z(n18508) );
  XOR U20092 ( .A(n18533), .B(n18534), .Z(n18523) );
  ANDN U20093 ( .B(n18535), .A(n18536), .Z(n18533) );
  XOR U20094 ( .A(n18534), .B(n18537), .Z(n18535) );
  XOR U20095 ( .A(n18538), .B(n18539), .Z(n18522) );
  XOR U20096 ( .A(n18540), .B(n18541), .Z(n18539) );
  ANDN U20097 ( .B(n18542), .A(n18543), .Z(n18540) );
  XOR U20098 ( .A(n18544), .B(n18541), .Z(n18542) );
  IV U20099 ( .A(n18520), .Z(n18538) );
  XOR U20100 ( .A(n18545), .B(n18546), .Z(n18520) );
  ANDN U20101 ( .B(n18547), .A(n18548), .Z(n18545) );
  XOR U20102 ( .A(n18546), .B(n18549), .Z(n18547) );
  IV U20103 ( .A(n18528), .Z(n18532) );
  XOR U20104 ( .A(n18528), .B(n18510), .Z(n18530) );
  XOR U20105 ( .A(n18550), .B(n18551), .Z(n18510) );
  AND U20106 ( .A(n682), .B(n18552), .Z(n18550) );
  XOR U20107 ( .A(n18553), .B(n18551), .Z(n18552) );
  NANDN U20108 ( .A(n18512), .B(n18514), .Z(n18528) );
  XOR U20109 ( .A(n18554), .B(n18555), .Z(n18514) );
  AND U20110 ( .A(n682), .B(n18556), .Z(n18554) );
  XOR U20111 ( .A(n18555), .B(n18557), .Z(n18556) );
  XOR U20112 ( .A(n18558), .B(n18559), .Z(n682) );
  AND U20113 ( .A(n18560), .B(n18561), .Z(n18558) );
  XNOR U20114 ( .A(n18559), .B(n18525), .Z(n18561) );
  XNOR U20115 ( .A(n18562), .B(n18563), .Z(n18525) );
  ANDN U20116 ( .B(n18564), .A(n18565), .Z(n18562) );
  XOR U20117 ( .A(n18563), .B(n18566), .Z(n18564) );
  XOR U20118 ( .A(n18559), .B(n18527), .Z(n18560) );
  XOR U20119 ( .A(n18567), .B(n18568), .Z(n18527) );
  AND U20120 ( .A(n686), .B(n18569), .Z(n18567) );
  XOR U20121 ( .A(n18570), .B(n18568), .Z(n18569) );
  XNOR U20122 ( .A(n18571), .B(n18572), .Z(n18559) );
  NAND U20123 ( .A(n18573), .B(n18574), .Z(n18572) );
  XOR U20124 ( .A(n18575), .B(n18551), .Z(n18574) );
  XOR U20125 ( .A(n18565), .B(n18566), .Z(n18551) );
  XOR U20126 ( .A(n18576), .B(n18577), .Z(n18566) );
  ANDN U20127 ( .B(n18578), .A(n18579), .Z(n18576) );
  XOR U20128 ( .A(n18577), .B(n18580), .Z(n18578) );
  XOR U20129 ( .A(n18581), .B(n18582), .Z(n18565) );
  XOR U20130 ( .A(n18583), .B(n18584), .Z(n18582) );
  ANDN U20131 ( .B(n18585), .A(n18586), .Z(n18583) );
  XOR U20132 ( .A(n18587), .B(n18584), .Z(n18585) );
  IV U20133 ( .A(n18563), .Z(n18581) );
  XOR U20134 ( .A(n18588), .B(n18589), .Z(n18563) );
  ANDN U20135 ( .B(n18590), .A(n18591), .Z(n18588) );
  XOR U20136 ( .A(n18589), .B(n18592), .Z(n18590) );
  IV U20137 ( .A(n18571), .Z(n18575) );
  XOR U20138 ( .A(n18571), .B(n18553), .Z(n18573) );
  XOR U20139 ( .A(n18593), .B(n18594), .Z(n18553) );
  AND U20140 ( .A(n686), .B(n18595), .Z(n18593) );
  XOR U20141 ( .A(n18596), .B(n18594), .Z(n18595) );
  NANDN U20142 ( .A(n18555), .B(n18557), .Z(n18571) );
  XOR U20143 ( .A(n18597), .B(n18598), .Z(n18557) );
  AND U20144 ( .A(n686), .B(n18599), .Z(n18597) );
  XOR U20145 ( .A(n18598), .B(n18600), .Z(n18599) );
  XOR U20146 ( .A(n18601), .B(n18602), .Z(n686) );
  AND U20147 ( .A(n18603), .B(n18604), .Z(n18601) );
  XNOR U20148 ( .A(n18602), .B(n18568), .Z(n18604) );
  XNOR U20149 ( .A(n18605), .B(n18606), .Z(n18568) );
  ANDN U20150 ( .B(n18607), .A(n18608), .Z(n18605) );
  XOR U20151 ( .A(n18606), .B(n18609), .Z(n18607) );
  XOR U20152 ( .A(n18602), .B(n18570), .Z(n18603) );
  XOR U20153 ( .A(n18610), .B(n18611), .Z(n18570) );
  AND U20154 ( .A(n690), .B(n18612), .Z(n18610) );
  XOR U20155 ( .A(n18613), .B(n18611), .Z(n18612) );
  XNOR U20156 ( .A(n18614), .B(n18615), .Z(n18602) );
  NAND U20157 ( .A(n18616), .B(n18617), .Z(n18615) );
  XOR U20158 ( .A(n18618), .B(n18594), .Z(n18617) );
  XOR U20159 ( .A(n18608), .B(n18609), .Z(n18594) );
  XOR U20160 ( .A(n18619), .B(n18620), .Z(n18609) );
  ANDN U20161 ( .B(n18621), .A(n18622), .Z(n18619) );
  XOR U20162 ( .A(n18620), .B(n18623), .Z(n18621) );
  XOR U20163 ( .A(n18624), .B(n18625), .Z(n18608) );
  XOR U20164 ( .A(n18626), .B(n18627), .Z(n18625) );
  ANDN U20165 ( .B(n18628), .A(n18629), .Z(n18626) );
  XOR U20166 ( .A(n18630), .B(n18627), .Z(n18628) );
  IV U20167 ( .A(n18606), .Z(n18624) );
  XOR U20168 ( .A(n18631), .B(n18632), .Z(n18606) );
  ANDN U20169 ( .B(n18633), .A(n18634), .Z(n18631) );
  XOR U20170 ( .A(n18632), .B(n18635), .Z(n18633) );
  IV U20171 ( .A(n18614), .Z(n18618) );
  XOR U20172 ( .A(n18614), .B(n18596), .Z(n18616) );
  XOR U20173 ( .A(n18636), .B(n18637), .Z(n18596) );
  AND U20174 ( .A(n690), .B(n18638), .Z(n18636) );
  XOR U20175 ( .A(n18639), .B(n18637), .Z(n18638) );
  NANDN U20176 ( .A(n18598), .B(n18600), .Z(n18614) );
  XOR U20177 ( .A(n18640), .B(n18641), .Z(n18600) );
  AND U20178 ( .A(n690), .B(n18642), .Z(n18640) );
  XOR U20179 ( .A(n18641), .B(n18643), .Z(n18642) );
  XOR U20180 ( .A(n18644), .B(n18645), .Z(n690) );
  AND U20181 ( .A(n18646), .B(n18647), .Z(n18644) );
  XNOR U20182 ( .A(n18645), .B(n18611), .Z(n18647) );
  XNOR U20183 ( .A(n18648), .B(n18649), .Z(n18611) );
  ANDN U20184 ( .B(n18650), .A(n18651), .Z(n18648) );
  XOR U20185 ( .A(n18649), .B(n18652), .Z(n18650) );
  XOR U20186 ( .A(n18645), .B(n18613), .Z(n18646) );
  XOR U20187 ( .A(n18653), .B(n18654), .Z(n18613) );
  AND U20188 ( .A(n694), .B(n18655), .Z(n18653) );
  XOR U20189 ( .A(n18656), .B(n18654), .Z(n18655) );
  XNOR U20190 ( .A(n18657), .B(n18658), .Z(n18645) );
  NAND U20191 ( .A(n18659), .B(n18660), .Z(n18658) );
  XOR U20192 ( .A(n18661), .B(n18637), .Z(n18660) );
  XOR U20193 ( .A(n18651), .B(n18652), .Z(n18637) );
  XOR U20194 ( .A(n18662), .B(n18663), .Z(n18652) );
  ANDN U20195 ( .B(n18664), .A(n18665), .Z(n18662) );
  XOR U20196 ( .A(n18663), .B(n18666), .Z(n18664) );
  XOR U20197 ( .A(n18667), .B(n18668), .Z(n18651) );
  XOR U20198 ( .A(n18669), .B(n18670), .Z(n18668) );
  ANDN U20199 ( .B(n18671), .A(n18672), .Z(n18669) );
  XOR U20200 ( .A(n18673), .B(n18670), .Z(n18671) );
  IV U20201 ( .A(n18649), .Z(n18667) );
  XOR U20202 ( .A(n18674), .B(n18675), .Z(n18649) );
  ANDN U20203 ( .B(n18676), .A(n18677), .Z(n18674) );
  XOR U20204 ( .A(n18675), .B(n18678), .Z(n18676) );
  IV U20205 ( .A(n18657), .Z(n18661) );
  XOR U20206 ( .A(n18657), .B(n18639), .Z(n18659) );
  XOR U20207 ( .A(n18679), .B(n18680), .Z(n18639) );
  AND U20208 ( .A(n694), .B(n18681), .Z(n18679) );
  XOR U20209 ( .A(n18682), .B(n18680), .Z(n18681) );
  NANDN U20210 ( .A(n18641), .B(n18643), .Z(n18657) );
  XOR U20211 ( .A(n18683), .B(n18684), .Z(n18643) );
  AND U20212 ( .A(n694), .B(n18685), .Z(n18683) );
  XOR U20213 ( .A(n18684), .B(n18686), .Z(n18685) );
  XOR U20214 ( .A(n18687), .B(n18688), .Z(n694) );
  AND U20215 ( .A(n18689), .B(n18690), .Z(n18687) );
  XNOR U20216 ( .A(n18688), .B(n18654), .Z(n18690) );
  XNOR U20217 ( .A(n18691), .B(n18692), .Z(n18654) );
  ANDN U20218 ( .B(n18693), .A(n18694), .Z(n18691) );
  XOR U20219 ( .A(n18692), .B(n18695), .Z(n18693) );
  XOR U20220 ( .A(n18688), .B(n18656), .Z(n18689) );
  XOR U20221 ( .A(n18696), .B(n18697), .Z(n18656) );
  AND U20222 ( .A(n698), .B(n18698), .Z(n18696) );
  XOR U20223 ( .A(n18699), .B(n18697), .Z(n18698) );
  XNOR U20224 ( .A(n18700), .B(n18701), .Z(n18688) );
  NAND U20225 ( .A(n18702), .B(n18703), .Z(n18701) );
  XOR U20226 ( .A(n18704), .B(n18680), .Z(n18703) );
  XOR U20227 ( .A(n18694), .B(n18695), .Z(n18680) );
  XOR U20228 ( .A(n18705), .B(n18706), .Z(n18695) );
  ANDN U20229 ( .B(n18707), .A(n18708), .Z(n18705) );
  XOR U20230 ( .A(n18706), .B(n18709), .Z(n18707) );
  XOR U20231 ( .A(n18710), .B(n18711), .Z(n18694) );
  XOR U20232 ( .A(n18712), .B(n18713), .Z(n18711) );
  ANDN U20233 ( .B(n18714), .A(n18715), .Z(n18712) );
  XOR U20234 ( .A(n18716), .B(n18713), .Z(n18714) );
  IV U20235 ( .A(n18692), .Z(n18710) );
  XOR U20236 ( .A(n18717), .B(n18718), .Z(n18692) );
  ANDN U20237 ( .B(n18719), .A(n18720), .Z(n18717) );
  XOR U20238 ( .A(n18718), .B(n18721), .Z(n18719) );
  IV U20239 ( .A(n18700), .Z(n18704) );
  XOR U20240 ( .A(n18700), .B(n18682), .Z(n18702) );
  XOR U20241 ( .A(n18722), .B(n18723), .Z(n18682) );
  AND U20242 ( .A(n698), .B(n18724), .Z(n18722) );
  XOR U20243 ( .A(n18725), .B(n18723), .Z(n18724) );
  NANDN U20244 ( .A(n18684), .B(n18686), .Z(n18700) );
  XOR U20245 ( .A(n18726), .B(n18727), .Z(n18686) );
  AND U20246 ( .A(n698), .B(n18728), .Z(n18726) );
  XOR U20247 ( .A(n18727), .B(n18729), .Z(n18728) );
  XOR U20248 ( .A(n18730), .B(n18731), .Z(n698) );
  AND U20249 ( .A(n18732), .B(n18733), .Z(n18730) );
  XNOR U20250 ( .A(n18731), .B(n18697), .Z(n18733) );
  XNOR U20251 ( .A(n18734), .B(n18735), .Z(n18697) );
  ANDN U20252 ( .B(n18736), .A(n18737), .Z(n18734) );
  XOR U20253 ( .A(n18735), .B(n18738), .Z(n18736) );
  XOR U20254 ( .A(n18731), .B(n18699), .Z(n18732) );
  XOR U20255 ( .A(n18739), .B(n18740), .Z(n18699) );
  AND U20256 ( .A(n702), .B(n18741), .Z(n18739) );
  XOR U20257 ( .A(n18742), .B(n18740), .Z(n18741) );
  XNOR U20258 ( .A(n18743), .B(n18744), .Z(n18731) );
  NAND U20259 ( .A(n18745), .B(n18746), .Z(n18744) );
  XOR U20260 ( .A(n18747), .B(n18723), .Z(n18746) );
  XOR U20261 ( .A(n18737), .B(n18738), .Z(n18723) );
  XOR U20262 ( .A(n18748), .B(n18749), .Z(n18738) );
  ANDN U20263 ( .B(n18750), .A(n18751), .Z(n18748) );
  XOR U20264 ( .A(n18749), .B(n18752), .Z(n18750) );
  XOR U20265 ( .A(n18753), .B(n18754), .Z(n18737) );
  XOR U20266 ( .A(n18755), .B(n18756), .Z(n18754) );
  ANDN U20267 ( .B(n18757), .A(n18758), .Z(n18755) );
  XOR U20268 ( .A(n18759), .B(n18756), .Z(n18757) );
  IV U20269 ( .A(n18735), .Z(n18753) );
  XOR U20270 ( .A(n18760), .B(n18761), .Z(n18735) );
  ANDN U20271 ( .B(n18762), .A(n18763), .Z(n18760) );
  XOR U20272 ( .A(n18761), .B(n18764), .Z(n18762) );
  IV U20273 ( .A(n18743), .Z(n18747) );
  XOR U20274 ( .A(n18743), .B(n18725), .Z(n18745) );
  XOR U20275 ( .A(n18765), .B(n18766), .Z(n18725) );
  AND U20276 ( .A(n702), .B(n18767), .Z(n18765) );
  XOR U20277 ( .A(n18768), .B(n18766), .Z(n18767) );
  NANDN U20278 ( .A(n18727), .B(n18729), .Z(n18743) );
  XOR U20279 ( .A(n18769), .B(n18770), .Z(n18729) );
  AND U20280 ( .A(n702), .B(n18771), .Z(n18769) );
  XOR U20281 ( .A(n18770), .B(n18772), .Z(n18771) );
  XOR U20282 ( .A(n18773), .B(n18774), .Z(n702) );
  AND U20283 ( .A(n18775), .B(n18776), .Z(n18773) );
  XNOR U20284 ( .A(n18774), .B(n18740), .Z(n18776) );
  XNOR U20285 ( .A(n18777), .B(n18778), .Z(n18740) );
  ANDN U20286 ( .B(n18779), .A(n18780), .Z(n18777) );
  XOR U20287 ( .A(n18778), .B(n18781), .Z(n18779) );
  XOR U20288 ( .A(n18774), .B(n18742), .Z(n18775) );
  XOR U20289 ( .A(n18782), .B(n18783), .Z(n18742) );
  AND U20290 ( .A(n706), .B(n18784), .Z(n18782) );
  XOR U20291 ( .A(n18785), .B(n18783), .Z(n18784) );
  XNOR U20292 ( .A(n18786), .B(n18787), .Z(n18774) );
  NAND U20293 ( .A(n18788), .B(n18789), .Z(n18787) );
  XOR U20294 ( .A(n18790), .B(n18766), .Z(n18789) );
  XOR U20295 ( .A(n18780), .B(n18781), .Z(n18766) );
  XOR U20296 ( .A(n18791), .B(n18792), .Z(n18781) );
  ANDN U20297 ( .B(n18793), .A(n18794), .Z(n18791) );
  XOR U20298 ( .A(n18792), .B(n18795), .Z(n18793) );
  XOR U20299 ( .A(n18796), .B(n18797), .Z(n18780) );
  XOR U20300 ( .A(n18798), .B(n18799), .Z(n18797) );
  ANDN U20301 ( .B(n18800), .A(n18801), .Z(n18798) );
  XOR U20302 ( .A(n18802), .B(n18799), .Z(n18800) );
  IV U20303 ( .A(n18778), .Z(n18796) );
  XOR U20304 ( .A(n18803), .B(n18804), .Z(n18778) );
  ANDN U20305 ( .B(n18805), .A(n18806), .Z(n18803) );
  XOR U20306 ( .A(n18804), .B(n18807), .Z(n18805) );
  IV U20307 ( .A(n18786), .Z(n18790) );
  XOR U20308 ( .A(n18786), .B(n18768), .Z(n18788) );
  XOR U20309 ( .A(n18808), .B(n18809), .Z(n18768) );
  AND U20310 ( .A(n706), .B(n18810), .Z(n18808) );
  XOR U20311 ( .A(n18811), .B(n18809), .Z(n18810) );
  NANDN U20312 ( .A(n18770), .B(n18772), .Z(n18786) );
  XOR U20313 ( .A(n18812), .B(n18813), .Z(n18772) );
  AND U20314 ( .A(n706), .B(n18814), .Z(n18812) );
  XOR U20315 ( .A(n18813), .B(n18815), .Z(n18814) );
  XOR U20316 ( .A(n18816), .B(n18817), .Z(n706) );
  AND U20317 ( .A(n18818), .B(n18819), .Z(n18816) );
  XNOR U20318 ( .A(n18817), .B(n18783), .Z(n18819) );
  XNOR U20319 ( .A(n18820), .B(n18821), .Z(n18783) );
  ANDN U20320 ( .B(n18822), .A(n18823), .Z(n18820) );
  XOR U20321 ( .A(n18821), .B(n18824), .Z(n18822) );
  XOR U20322 ( .A(n18817), .B(n18785), .Z(n18818) );
  XOR U20323 ( .A(n18825), .B(n18826), .Z(n18785) );
  AND U20324 ( .A(n710), .B(n18827), .Z(n18825) );
  XOR U20325 ( .A(n18828), .B(n18826), .Z(n18827) );
  XNOR U20326 ( .A(n18829), .B(n18830), .Z(n18817) );
  NAND U20327 ( .A(n18831), .B(n18832), .Z(n18830) );
  XOR U20328 ( .A(n18833), .B(n18809), .Z(n18832) );
  XOR U20329 ( .A(n18823), .B(n18824), .Z(n18809) );
  XOR U20330 ( .A(n18834), .B(n18835), .Z(n18824) );
  ANDN U20331 ( .B(n18836), .A(n18837), .Z(n18834) );
  XOR U20332 ( .A(n18835), .B(n18838), .Z(n18836) );
  XOR U20333 ( .A(n18839), .B(n18840), .Z(n18823) );
  XOR U20334 ( .A(n18841), .B(n18842), .Z(n18840) );
  ANDN U20335 ( .B(n18843), .A(n18844), .Z(n18841) );
  XOR U20336 ( .A(n18845), .B(n18842), .Z(n18843) );
  IV U20337 ( .A(n18821), .Z(n18839) );
  XOR U20338 ( .A(n18846), .B(n18847), .Z(n18821) );
  ANDN U20339 ( .B(n18848), .A(n18849), .Z(n18846) );
  XOR U20340 ( .A(n18847), .B(n18850), .Z(n18848) );
  IV U20341 ( .A(n18829), .Z(n18833) );
  XOR U20342 ( .A(n18829), .B(n18811), .Z(n18831) );
  XOR U20343 ( .A(n18851), .B(n18852), .Z(n18811) );
  AND U20344 ( .A(n710), .B(n18853), .Z(n18851) );
  XOR U20345 ( .A(n18854), .B(n18852), .Z(n18853) );
  NANDN U20346 ( .A(n18813), .B(n18815), .Z(n18829) );
  XOR U20347 ( .A(n18855), .B(n18856), .Z(n18815) );
  AND U20348 ( .A(n710), .B(n18857), .Z(n18855) );
  XOR U20349 ( .A(n18856), .B(n18858), .Z(n18857) );
  XOR U20350 ( .A(n18859), .B(n18860), .Z(n710) );
  AND U20351 ( .A(n18861), .B(n18862), .Z(n18859) );
  XNOR U20352 ( .A(n18860), .B(n18826), .Z(n18862) );
  XNOR U20353 ( .A(n18863), .B(n18864), .Z(n18826) );
  ANDN U20354 ( .B(n18865), .A(n18866), .Z(n18863) );
  XOR U20355 ( .A(n18864), .B(n18867), .Z(n18865) );
  XOR U20356 ( .A(n18860), .B(n18828), .Z(n18861) );
  XOR U20357 ( .A(n18868), .B(n18869), .Z(n18828) );
  AND U20358 ( .A(n714), .B(n18870), .Z(n18868) );
  XOR U20359 ( .A(n18871), .B(n18869), .Z(n18870) );
  XNOR U20360 ( .A(n18872), .B(n18873), .Z(n18860) );
  NAND U20361 ( .A(n18874), .B(n18875), .Z(n18873) );
  XOR U20362 ( .A(n18876), .B(n18852), .Z(n18875) );
  XOR U20363 ( .A(n18866), .B(n18867), .Z(n18852) );
  XOR U20364 ( .A(n18877), .B(n18878), .Z(n18867) );
  ANDN U20365 ( .B(n18879), .A(n18880), .Z(n18877) );
  XOR U20366 ( .A(n18878), .B(n18881), .Z(n18879) );
  XOR U20367 ( .A(n18882), .B(n18883), .Z(n18866) );
  XOR U20368 ( .A(n18884), .B(n18885), .Z(n18883) );
  ANDN U20369 ( .B(n18886), .A(n18887), .Z(n18884) );
  XOR U20370 ( .A(n18888), .B(n18885), .Z(n18886) );
  IV U20371 ( .A(n18864), .Z(n18882) );
  XOR U20372 ( .A(n18889), .B(n18890), .Z(n18864) );
  ANDN U20373 ( .B(n18891), .A(n18892), .Z(n18889) );
  XOR U20374 ( .A(n18890), .B(n18893), .Z(n18891) );
  IV U20375 ( .A(n18872), .Z(n18876) );
  XOR U20376 ( .A(n18872), .B(n18854), .Z(n18874) );
  XOR U20377 ( .A(n18894), .B(n18895), .Z(n18854) );
  AND U20378 ( .A(n714), .B(n18896), .Z(n18894) );
  XOR U20379 ( .A(n18897), .B(n18895), .Z(n18896) );
  NANDN U20380 ( .A(n18856), .B(n18858), .Z(n18872) );
  XOR U20381 ( .A(n18898), .B(n18899), .Z(n18858) );
  AND U20382 ( .A(n714), .B(n18900), .Z(n18898) );
  XOR U20383 ( .A(n18899), .B(n18901), .Z(n18900) );
  XOR U20384 ( .A(n18902), .B(n18903), .Z(n714) );
  AND U20385 ( .A(n18904), .B(n18905), .Z(n18902) );
  XNOR U20386 ( .A(n18903), .B(n18869), .Z(n18905) );
  XNOR U20387 ( .A(n18906), .B(n18907), .Z(n18869) );
  ANDN U20388 ( .B(n18908), .A(n18909), .Z(n18906) );
  XOR U20389 ( .A(n18907), .B(n18910), .Z(n18908) );
  XOR U20390 ( .A(n18903), .B(n18871), .Z(n18904) );
  XOR U20391 ( .A(n18911), .B(n18912), .Z(n18871) );
  AND U20392 ( .A(n718), .B(n18913), .Z(n18911) );
  XOR U20393 ( .A(n18914), .B(n18912), .Z(n18913) );
  XNOR U20394 ( .A(n18915), .B(n18916), .Z(n18903) );
  NAND U20395 ( .A(n18917), .B(n18918), .Z(n18916) );
  XOR U20396 ( .A(n18919), .B(n18895), .Z(n18918) );
  XOR U20397 ( .A(n18909), .B(n18910), .Z(n18895) );
  XOR U20398 ( .A(n18920), .B(n18921), .Z(n18910) );
  ANDN U20399 ( .B(n18922), .A(n18923), .Z(n18920) );
  XOR U20400 ( .A(n18921), .B(n18924), .Z(n18922) );
  XOR U20401 ( .A(n18925), .B(n18926), .Z(n18909) );
  XOR U20402 ( .A(n18927), .B(n18928), .Z(n18926) );
  ANDN U20403 ( .B(n18929), .A(n18930), .Z(n18927) );
  XOR U20404 ( .A(n18931), .B(n18928), .Z(n18929) );
  IV U20405 ( .A(n18907), .Z(n18925) );
  XOR U20406 ( .A(n18932), .B(n18933), .Z(n18907) );
  ANDN U20407 ( .B(n18934), .A(n18935), .Z(n18932) );
  XOR U20408 ( .A(n18933), .B(n18936), .Z(n18934) );
  IV U20409 ( .A(n18915), .Z(n18919) );
  XOR U20410 ( .A(n18915), .B(n18897), .Z(n18917) );
  XOR U20411 ( .A(n18937), .B(n18938), .Z(n18897) );
  AND U20412 ( .A(n718), .B(n18939), .Z(n18937) );
  XOR U20413 ( .A(n18940), .B(n18938), .Z(n18939) );
  NANDN U20414 ( .A(n18899), .B(n18901), .Z(n18915) );
  XOR U20415 ( .A(n18941), .B(n18942), .Z(n18901) );
  AND U20416 ( .A(n718), .B(n18943), .Z(n18941) );
  XOR U20417 ( .A(n18942), .B(n18944), .Z(n18943) );
  XOR U20418 ( .A(n18945), .B(n18946), .Z(n718) );
  AND U20419 ( .A(n18947), .B(n18948), .Z(n18945) );
  XNOR U20420 ( .A(n18946), .B(n18912), .Z(n18948) );
  XNOR U20421 ( .A(n18949), .B(n18950), .Z(n18912) );
  ANDN U20422 ( .B(n18951), .A(n18952), .Z(n18949) );
  XOR U20423 ( .A(n18950), .B(n18953), .Z(n18951) );
  XOR U20424 ( .A(n18946), .B(n18914), .Z(n18947) );
  XOR U20425 ( .A(n18954), .B(n18955), .Z(n18914) );
  AND U20426 ( .A(n722), .B(n18956), .Z(n18954) );
  XOR U20427 ( .A(n18957), .B(n18955), .Z(n18956) );
  XNOR U20428 ( .A(n18958), .B(n18959), .Z(n18946) );
  NAND U20429 ( .A(n18960), .B(n18961), .Z(n18959) );
  XOR U20430 ( .A(n18962), .B(n18938), .Z(n18961) );
  XOR U20431 ( .A(n18952), .B(n18953), .Z(n18938) );
  XOR U20432 ( .A(n18963), .B(n18964), .Z(n18953) );
  ANDN U20433 ( .B(n18965), .A(n18966), .Z(n18963) );
  XOR U20434 ( .A(n18964), .B(n18967), .Z(n18965) );
  XOR U20435 ( .A(n18968), .B(n18969), .Z(n18952) );
  XOR U20436 ( .A(n18970), .B(n18971), .Z(n18969) );
  ANDN U20437 ( .B(n18972), .A(n18973), .Z(n18970) );
  XOR U20438 ( .A(n18974), .B(n18971), .Z(n18972) );
  IV U20439 ( .A(n18950), .Z(n18968) );
  XOR U20440 ( .A(n18975), .B(n18976), .Z(n18950) );
  ANDN U20441 ( .B(n18977), .A(n18978), .Z(n18975) );
  XOR U20442 ( .A(n18976), .B(n18979), .Z(n18977) );
  IV U20443 ( .A(n18958), .Z(n18962) );
  XOR U20444 ( .A(n18958), .B(n18940), .Z(n18960) );
  XOR U20445 ( .A(n18980), .B(n18981), .Z(n18940) );
  AND U20446 ( .A(n722), .B(n18982), .Z(n18980) );
  XOR U20447 ( .A(n18983), .B(n18981), .Z(n18982) );
  NANDN U20448 ( .A(n18942), .B(n18944), .Z(n18958) );
  XOR U20449 ( .A(n18984), .B(n18985), .Z(n18944) );
  AND U20450 ( .A(n722), .B(n18986), .Z(n18984) );
  XOR U20451 ( .A(n18985), .B(n18987), .Z(n18986) );
  XOR U20452 ( .A(n18988), .B(n18989), .Z(n722) );
  AND U20453 ( .A(n18990), .B(n18991), .Z(n18988) );
  XNOR U20454 ( .A(n18989), .B(n18955), .Z(n18991) );
  XNOR U20455 ( .A(n18992), .B(n18993), .Z(n18955) );
  ANDN U20456 ( .B(n18994), .A(n18995), .Z(n18992) );
  XOR U20457 ( .A(n18993), .B(n18996), .Z(n18994) );
  XOR U20458 ( .A(n18989), .B(n18957), .Z(n18990) );
  XOR U20459 ( .A(n18997), .B(n18998), .Z(n18957) );
  AND U20460 ( .A(n726), .B(n18999), .Z(n18997) );
  XOR U20461 ( .A(n19000), .B(n18998), .Z(n18999) );
  XNOR U20462 ( .A(n19001), .B(n19002), .Z(n18989) );
  NAND U20463 ( .A(n19003), .B(n19004), .Z(n19002) );
  XOR U20464 ( .A(n19005), .B(n18981), .Z(n19004) );
  XOR U20465 ( .A(n18995), .B(n18996), .Z(n18981) );
  XOR U20466 ( .A(n19006), .B(n19007), .Z(n18996) );
  ANDN U20467 ( .B(n19008), .A(n19009), .Z(n19006) );
  XOR U20468 ( .A(n19007), .B(n19010), .Z(n19008) );
  XOR U20469 ( .A(n19011), .B(n19012), .Z(n18995) );
  XOR U20470 ( .A(n19013), .B(n19014), .Z(n19012) );
  ANDN U20471 ( .B(n19015), .A(n19016), .Z(n19013) );
  XOR U20472 ( .A(n19017), .B(n19014), .Z(n19015) );
  IV U20473 ( .A(n18993), .Z(n19011) );
  XOR U20474 ( .A(n19018), .B(n19019), .Z(n18993) );
  ANDN U20475 ( .B(n19020), .A(n19021), .Z(n19018) );
  XOR U20476 ( .A(n19019), .B(n19022), .Z(n19020) );
  IV U20477 ( .A(n19001), .Z(n19005) );
  XOR U20478 ( .A(n19001), .B(n18983), .Z(n19003) );
  XOR U20479 ( .A(n19023), .B(n19024), .Z(n18983) );
  AND U20480 ( .A(n726), .B(n19025), .Z(n19023) );
  XOR U20481 ( .A(n19026), .B(n19024), .Z(n19025) );
  NANDN U20482 ( .A(n18985), .B(n18987), .Z(n19001) );
  XOR U20483 ( .A(n19027), .B(n19028), .Z(n18987) );
  AND U20484 ( .A(n726), .B(n19029), .Z(n19027) );
  XOR U20485 ( .A(n19028), .B(n19030), .Z(n19029) );
  XOR U20486 ( .A(n19031), .B(n19032), .Z(n726) );
  AND U20487 ( .A(n19033), .B(n19034), .Z(n19031) );
  XNOR U20488 ( .A(n19032), .B(n18998), .Z(n19034) );
  XNOR U20489 ( .A(n19035), .B(n19036), .Z(n18998) );
  ANDN U20490 ( .B(n19037), .A(n19038), .Z(n19035) );
  XOR U20491 ( .A(n19036), .B(n19039), .Z(n19037) );
  XOR U20492 ( .A(n19032), .B(n19000), .Z(n19033) );
  XOR U20493 ( .A(n19040), .B(n19041), .Z(n19000) );
  AND U20494 ( .A(n730), .B(n19042), .Z(n19040) );
  XOR U20495 ( .A(n19043), .B(n19041), .Z(n19042) );
  XNOR U20496 ( .A(n19044), .B(n19045), .Z(n19032) );
  NAND U20497 ( .A(n19046), .B(n19047), .Z(n19045) );
  XOR U20498 ( .A(n19048), .B(n19024), .Z(n19047) );
  XOR U20499 ( .A(n19038), .B(n19039), .Z(n19024) );
  XOR U20500 ( .A(n19049), .B(n19050), .Z(n19039) );
  ANDN U20501 ( .B(n19051), .A(n19052), .Z(n19049) );
  XOR U20502 ( .A(n19050), .B(n19053), .Z(n19051) );
  XOR U20503 ( .A(n19054), .B(n19055), .Z(n19038) );
  XOR U20504 ( .A(n19056), .B(n19057), .Z(n19055) );
  ANDN U20505 ( .B(n19058), .A(n19059), .Z(n19056) );
  XOR U20506 ( .A(n19060), .B(n19057), .Z(n19058) );
  IV U20507 ( .A(n19036), .Z(n19054) );
  XOR U20508 ( .A(n19061), .B(n19062), .Z(n19036) );
  ANDN U20509 ( .B(n19063), .A(n19064), .Z(n19061) );
  XOR U20510 ( .A(n19062), .B(n19065), .Z(n19063) );
  IV U20511 ( .A(n19044), .Z(n19048) );
  XOR U20512 ( .A(n19044), .B(n19026), .Z(n19046) );
  XOR U20513 ( .A(n19066), .B(n19067), .Z(n19026) );
  AND U20514 ( .A(n730), .B(n19068), .Z(n19066) );
  XOR U20515 ( .A(n19069), .B(n19067), .Z(n19068) );
  NANDN U20516 ( .A(n19028), .B(n19030), .Z(n19044) );
  XOR U20517 ( .A(n19070), .B(n19071), .Z(n19030) );
  AND U20518 ( .A(n730), .B(n19072), .Z(n19070) );
  XOR U20519 ( .A(n19071), .B(n19073), .Z(n19072) );
  XOR U20520 ( .A(n19074), .B(n19075), .Z(n730) );
  AND U20521 ( .A(n19076), .B(n19077), .Z(n19074) );
  XNOR U20522 ( .A(n19075), .B(n19041), .Z(n19077) );
  XNOR U20523 ( .A(n19078), .B(n19079), .Z(n19041) );
  ANDN U20524 ( .B(n19080), .A(n19081), .Z(n19078) );
  XOR U20525 ( .A(n19079), .B(n19082), .Z(n19080) );
  XOR U20526 ( .A(n19075), .B(n19043), .Z(n19076) );
  XOR U20527 ( .A(n19083), .B(n19084), .Z(n19043) );
  AND U20528 ( .A(n734), .B(n19085), .Z(n19083) );
  XOR U20529 ( .A(n19086), .B(n19084), .Z(n19085) );
  XNOR U20530 ( .A(n19087), .B(n19088), .Z(n19075) );
  NAND U20531 ( .A(n19089), .B(n19090), .Z(n19088) );
  XOR U20532 ( .A(n19091), .B(n19067), .Z(n19090) );
  XOR U20533 ( .A(n19081), .B(n19082), .Z(n19067) );
  XOR U20534 ( .A(n19092), .B(n19093), .Z(n19082) );
  ANDN U20535 ( .B(n19094), .A(n19095), .Z(n19092) );
  XOR U20536 ( .A(n19093), .B(n19096), .Z(n19094) );
  XOR U20537 ( .A(n19097), .B(n19098), .Z(n19081) );
  XOR U20538 ( .A(n19099), .B(n19100), .Z(n19098) );
  ANDN U20539 ( .B(n19101), .A(n19102), .Z(n19099) );
  XOR U20540 ( .A(n19103), .B(n19100), .Z(n19101) );
  IV U20541 ( .A(n19079), .Z(n19097) );
  XOR U20542 ( .A(n19104), .B(n19105), .Z(n19079) );
  ANDN U20543 ( .B(n19106), .A(n19107), .Z(n19104) );
  XOR U20544 ( .A(n19105), .B(n19108), .Z(n19106) );
  IV U20545 ( .A(n19087), .Z(n19091) );
  XOR U20546 ( .A(n19087), .B(n19069), .Z(n19089) );
  XOR U20547 ( .A(n19109), .B(n19110), .Z(n19069) );
  AND U20548 ( .A(n734), .B(n19111), .Z(n19109) );
  XOR U20549 ( .A(n19112), .B(n19110), .Z(n19111) );
  NANDN U20550 ( .A(n19071), .B(n19073), .Z(n19087) );
  XOR U20551 ( .A(n19113), .B(n19114), .Z(n19073) );
  AND U20552 ( .A(n734), .B(n19115), .Z(n19113) );
  XOR U20553 ( .A(n19114), .B(n19116), .Z(n19115) );
  XOR U20554 ( .A(n19117), .B(n19118), .Z(n734) );
  AND U20555 ( .A(n19119), .B(n19120), .Z(n19117) );
  XNOR U20556 ( .A(n19118), .B(n19084), .Z(n19120) );
  XNOR U20557 ( .A(n19121), .B(n19122), .Z(n19084) );
  ANDN U20558 ( .B(n19123), .A(n19124), .Z(n19121) );
  XOR U20559 ( .A(n19122), .B(n19125), .Z(n19123) );
  XOR U20560 ( .A(n19118), .B(n19086), .Z(n19119) );
  XOR U20561 ( .A(n19126), .B(n19127), .Z(n19086) );
  AND U20562 ( .A(n738), .B(n19128), .Z(n19126) );
  XOR U20563 ( .A(n19129), .B(n19127), .Z(n19128) );
  XNOR U20564 ( .A(n19130), .B(n19131), .Z(n19118) );
  NAND U20565 ( .A(n19132), .B(n19133), .Z(n19131) );
  XOR U20566 ( .A(n19134), .B(n19110), .Z(n19133) );
  XOR U20567 ( .A(n19124), .B(n19125), .Z(n19110) );
  XOR U20568 ( .A(n19135), .B(n19136), .Z(n19125) );
  ANDN U20569 ( .B(n19137), .A(n19138), .Z(n19135) );
  XOR U20570 ( .A(n19136), .B(n19139), .Z(n19137) );
  XOR U20571 ( .A(n19140), .B(n19141), .Z(n19124) );
  XOR U20572 ( .A(n19142), .B(n19143), .Z(n19141) );
  ANDN U20573 ( .B(n19144), .A(n19145), .Z(n19142) );
  XOR U20574 ( .A(n19146), .B(n19143), .Z(n19144) );
  IV U20575 ( .A(n19122), .Z(n19140) );
  XOR U20576 ( .A(n19147), .B(n19148), .Z(n19122) );
  ANDN U20577 ( .B(n19149), .A(n19150), .Z(n19147) );
  XOR U20578 ( .A(n19148), .B(n19151), .Z(n19149) );
  IV U20579 ( .A(n19130), .Z(n19134) );
  XOR U20580 ( .A(n19130), .B(n19112), .Z(n19132) );
  XOR U20581 ( .A(n19152), .B(n19153), .Z(n19112) );
  AND U20582 ( .A(n738), .B(n19154), .Z(n19152) );
  XOR U20583 ( .A(n19155), .B(n19153), .Z(n19154) );
  NANDN U20584 ( .A(n19114), .B(n19116), .Z(n19130) );
  XOR U20585 ( .A(n19156), .B(n19157), .Z(n19116) );
  AND U20586 ( .A(n738), .B(n19158), .Z(n19156) );
  XOR U20587 ( .A(n19157), .B(n19159), .Z(n19158) );
  XOR U20588 ( .A(n19160), .B(n19161), .Z(n738) );
  AND U20589 ( .A(n19162), .B(n19163), .Z(n19160) );
  XNOR U20590 ( .A(n19161), .B(n19127), .Z(n19163) );
  XNOR U20591 ( .A(n19164), .B(n19165), .Z(n19127) );
  ANDN U20592 ( .B(n19166), .A(n19167), .Z(n19164) );
  XOR U20593 ( .A(n19165), .B(n19168), .Z(n19166) );
  XOR U20594 ( .A(n19161), .B(n19129), .Z(n19162) );
  XOR U20595 ( .A(n19169), .B(n19170), .Z(n19129) );
  AND U20596 ( .A(n742), .B(n19171), .Z(n19169) );
  XOR U20597 ( .A(n19172), .B(n19170), .Z(n19171) );
  XNOR U20598 ( .A(n19173), .B(n19174), .Z(n19161) );
  NAND U20599 ( .A(n19175), .B(n19176), .Z(n19174) );
  XOR U20600 ( .A(n19177), .B(n19153), .Z(n19176) );
  XOR U20601 ( .A(n19167), .B(n19168), .Z(n19153) );
  XOR U20602 ( .A(n19178), .B(n19179), .Z(n19168) );
  ANDN U20603 ( .B(n19180), .A(n19181), .Z(n19178) );
  XOR U20604 ( .A(n19179), .B(n19182), .Z(n19180) );
  XOR U20605 ( .A(n19183), .B(n19184), .Z(n19167) );
  XOR U20606 ( .A(n19185), .B(n19186), .Z(n19184) );
  ANDN U20607 ( .B(n19187), .A(n19188), .Z(n19185) );
  XOR U20608 ( .A(n19189), .B(n19186), .Z(n19187) );
  IV U20609 ( .A(n19165), .Z(n19183) );
  XOR U20610 ( .A(n19190), .B(n19191), .Z(n19165) );
  ANDN U20611 ( .B(n19192), .A(n19193), .Z(n19190) );
  XOR U20612 ( .A(n19191), .B(n19194), .Z(n19192) );
  IV U20613 ( .A(n19173), .Z(n19177) );
  XOR U20614 ( .A(n19173), .B(n19155), .Z(n19175) );
  XOR U20615 ( .A(n19195), .B(n19196), .Z(n19155) );
  AND U20616 ( .A(n742), .B(n19197), .Z(n19195) );
  XOR U20617 ( .A(n19198), .B(n19196), .Z(n19197) );
  NANDN U20618 ( .A(n19157), .B(n19159), .Z(n19173) );
  XOR U20619 ( .A(n19199), .B(n19200), .Z(n19159) );
  AND U20620 ( .A(n742), .B(n19201), .Z(n19199) );
  XOR U20621 ( .A(n19200), .B(n19202), .Z(n19201) );
  XOR U20622 ( .A(n19203), .B(n19204), .Z(n742) );
  AND U20623 ( .A(n19205), .B(n19206), .Z(n19203) );
  XNOR U20624 ( .A(n19204), .B(n19170), .Z(n19206) );
  XNOR U20625 ( .A(n19207), .B(n19208), .Z(n19170) );
  ANDN U20626 ( .B(n19209), .A(n19210), .Z(n19207) );
  XOR U20627 ( .A(n19208), .B(n19211), .Z(n19209) );
  XOR U20628 ( .A(n19204), .B(n19172), .Z(n19205) );
  XOR U20629 ( .A(n19212), .B(n19213), .Z(n19172) );
  AND U20630 ( .A(n746), .B(n19214), .Z(n19212) );
  XOR U20631 ( .A(n19215), .B(n19213), .Z(n19214) );
  XNOR U20632 ( .A(n19216), .B(n19217), .Z(n19204) );
  NAND U20633 ( .A(n19218), .B(n19219), .Z(n19217) );
  XOR U20634 ( .A(n19220), .B(n19196), .Z(n19219) );
  XOR U20635 ( .A(n19210), .B(n19211), .Z(n19196) );
  XOR U20636 ( .A(n19221), .B(n19222), .Z(n19211) );
  ANDN U20637 ( .B(n19223), .A(n19224), .Z(n19221) );
  XOR U20638 ( .A(n19222), .B(n19225), .Z(n19223) );
  XOR U20639 ( .A(n19226), .B(n19227), .Z(n19210) );
  XOR U20640 ( .A(n19228), .B(n19229), .Z(n19227) );
  ANDN U20641 ( .B(n19230), .A(n19231), .Z(n19228) );
  XOR U20642 ( .A(n19232), .B(n19229), .Z(n19230) );
  IV U20643 ( .A(n19208), .Z(n19226) );
  XOR U20644 ( .A(n19233), .B(n19234), .Z(n19208) );
  ANDN U20645 ( .B(n19235), .A(n19236), .Z(n19233) );
  XOR U20646 ( .A(n19234), .B(n19237), .Z(n19235) );
  IV U20647 ( .A(n19216), .Z(n19220) );
  XOR U20648 ( .A(n19216), .B(n19198), .Z(n19218) );
  XOR U20649 ( .A(n19238), .B(n19239), .Z(n19198) );
  AND U20650 ( .A(n746), .B(n19240), .Z(n19238) );
  XOR U20651 ( .A(n19241), .B(n19239), .Z(n19240) );
  NANDN U20652 ( .A(n19200), .B(n19202), .Z(n19216) );
  XOR U20653 ( .A(n19242), .B(n19243), .Z(n19202) );
  AND U20654 ( .A(n746), .B(n19244), .Z(n19242) );
  XOR U20655 ( .A(n19243), .B(n19245), .Z(n19244) );
  XOR U20656 ( .A(n19246), .B(n19247), .Z(n746) );
  AND U20657 ( .A(n19248), .B(n19249), .Z(n19246) );
  XNOR U20658 ( .A(n19247), .B(n19213), .Z(n19249) );
  XNOR U20659 ( .A(n19250), .B(n19251), .Z(n19213) );
  ANDN U20660 ( .B(n19252), .A(n19253), .Z(n19250) );
  XOR U20661 ( .A(n19251), .B(n19254), .Z(n19252) );
  XOR U20662 ( .A(n19247), .B(n19215), .Z(n19248) );
  XOR U20663 ( .A(n19255), .B(n19256), .Z(n19215) );
  AND U20664 ( .A(n750), .B(n19257), .Z(n19255) );
  XOR U20665 ( .A(n19258), .B(n19256), .Z(n19257) );
  XNOR U20666 ( .A(n19259), .B(n19260), .Z(n19247) );
  NAND U20667 ( .A(n19261), .B(n19262), .Z(n19260) );
  XOR U20668 ( .A(n19263), .B(n19239), .Z(n19262) );
  XOR U20669 ( .A(n19253), .B(n19254), .Z(n19239) );
  XOR U20670 ( .A(n19264), .B(n19265), .Z(n19254) );
  ANDN U20671 ( .B(n19266), .A(n19267), .Z(n19264) );
  XOR U20672 ( .A(n19265), .B(n19268), .Z(n19266) );
  XOR U20673 ( .A(n19269), .B(n19270), .Z(n19253) );
  XOR U20674 ( .A(n19271), .B(n19272), .Z(n19270) );
  ANDN U20675 ( .B(n19273), .A(n19274), .Z(n19271) );
  XOR U20676 ( .A(n19275), .B(n19272), .Z(n19273) );
  IV U20677 ( .A(n19251), .Z(n19269) );
  XOR U20678 ( .A(n19276), .B(n19277), .Z(n19251) );
  ANDN U20679 ( .B(n19278), .A(n19279), .Z(n19276) );
  XOR U20680 ( .A(n19277), .B(n19280), .Z(n19278) );
  IV U20681 ( .A(n19259), .Z(n19263) );
  XOR U20682 ( .A(n19259), .B(n19241), .Z(n19261) );
  XOR U20683 ( .A(n19281), .B(n19282), .Z(n19241) );
  AND U20684 ( .A(n750), .B(n19283), .Z(n19281) );
  XOR U20685 ( .A(n19284), .B(n19282), .Z(n19283) );
  NANDN U20686 ( .A(n19243), .B(n19245), .Z(n19259) );
  XOR U20687 ( .A(n19285), .B(n19286), .Z(n19245) );
  AND U20688 ( .A(n750), .B(n19287), .Z(n19285) );
  XOR U20689 ( .A(n19286), .B(n19288), .Z(n19287) );
  XOR U20690 ( .A(n19289), .B(n19290), .Z(n750) );
  AND U20691 ( .A(n19291), .B(n19292), .Z(n19289) );
  XNOR U20692 ( .A(n19290), .B(n19256), .Z(n19292) );
  XNOR U20693 ( .A(n19293), .B(n19294), .Z(n19256) );
  ANDN U20694 ( .B(n19295), .A(n19296), .Z(n19293) );
  XOR U20695 ( .A(n19294), .B(n19297), .Z(n19295) );
  XOR U20696 ( .A(n19290), .B(n19258), .Z(n19291) );
  XOR U20697 ( .A(n19298), .B(n19299), .Z(n19258) );
  AND U20698 ( .A(n754), .B(n19300), .Z(n19298) );
  XOR U20699 ( .A(n19301), .B(n19299), .Z(n19300) );
  XNOR U20700 ( .A(n19302), .B(n19303), .Z(n19290) );
  NAND U20701 ( .A(n19304), .B(n19305), .Z(n19303) );
  XOR U20702 ( .A(n19306), .B(n19282), .Z(n19305) );
  XOR U20703 ( .A(n19296), .B(n19297), .Z(n19282) );
  XOR U20704 ( .A(n19307), .B(n19308), .Z(n19297) );
  ANDN U20705 ( .B(n19309), .A(n19310), .Z(n19307) );
  XOR U20706 ( .A(n19308), .B(n19311), .Z(n19309) );
  XOR U20707 ( .A(n19312), .B(n19313), .Z(n19296) );
  XOR U20708 ( .A(n19314), .B(n19315), .Z(n19313) );
  ANDN U20709 ( .B(n19316), .A(n19317), .Z(n19314) );
  XOR U20710 ( .A(n19318), .B(n19315), .Z(n19316) );
  IV U20711 ( .A(n19294), .Z(n19312) );
  XOR U20712 ( .A(n19319), .B(n19320), .Z(n19294) );
  ANDN U20713 ( .B(n19321), .A(n19322), .Z(n19319) );
  XOR U20714 ( .A(n19320), .B(n19323), .Z(n19321) );
  IV U20715 ( .A(n19302), .Z(n19306) );
  XOR U20716 ( .A(n19302), .B(n19284), .Z(n19304) );
  XOR U20717 ( .A(n19324), .B(n19325), .Z(n19284) );
  AND U20718 ( .A(n754), .B(n19326), .Z(n19324) );
  XOR U20719 ( .A(n19327), .B(n19325), .Z(n19326) );
  NANDN U20720 ( .A(n19286), .B(n19288), .Z(n19302) );
  XOR U20721 ( .A(n19328), .B(n19329), .Z(n19288) );
  AND U20722 ( .A(n754), .B(n19330), .Z(n19328) );
  XOR U20723 ( .A(n19329), .B(n19331), .Z(n19330) );
  XOR U20724 ( .A(n19332), .B(n19333), .Z(n754) );
  AND U20725 ( .A(n19334), .B(n19335), .Z(n19332) );
  XNOR U20726 ( .A(n19333), .B(n19299), .Z(n19335) );
  XNOR U20727 ( .A(n19336), .B(n19337), .Z(n19299) );
  ANDN U20728 ( .B(n19338), .A(n19339), .Z(n19336) );
  XOR U20729 ( .A(n19337), .B(n19340), .Z(n19338) );
  XOR U20730 ( .A(n19333), .B(n19301), .Z(n19334) );
  XOR U20731 ( .A(n19341), .B(n19342), .Z(n19301) );
  AND U20732 ( .A(n758), .B(n19343), .Z(n19341) );
  XOR U20733 ( .A(n19344), .B(n19342), .Z(n19343) );
  XNOR U20734 ( .A(n19345), .B(n19346), .Z(n19333) );
  NAND U20735 ( .A(n19347), .B(n19348), .Z(n19346) );
  XOR U20736 ( .A(n19349), .B(n19325), .Z(n19348) );
  XOR U20737 ( .A(n19339), .B(n19340), .Z(n19325) );
  XOR U20738 ( .A(n19350), .B(n19351), .Z(n19340) );
  ANDN U20739 ( .B(n19352), .A(n19353), .Z(n19350) );
  XOR U20740 ( .A(n19351), .B(n19354), .Z(n19352) );
  XOR U20741 ( .A(n19355), .B(n19356), .Z(n19339) );
  XOR U20742 ( .A(n19357), .B(n19358), .Z(n19356) );
  ANDN U20743 ( .B(n19359), .A(n19360), .Z(n19357) );
  XOR U20744 ( .A(n19361), .B(n19358), .Z(n19359) );
  IV U20745 ( .A(n19337), .Z(n19355) );
  XOR U20746 ( .A(n19362), .B(n19363), .Z(n19337) );
  ANDN U20747 ( .B(n19364), .A(n19365), .Z(n19362) );
  XOR U20748 ( .A(n19363), .B(n19366), .Z(n19364) );
  IV U20749 ( .A(n19345), .Z(n19349) );
  XOR U20750 ( .A(n19345), .B(n19327), .Z(n19347) );
  XOR U20751 ( .A(n19367), .B(n19368), .Z(n19327) );
  AND U20752 ( .A(n758), .B(n19369), .Z(n19367) );
  XOR U20753 ( .A(n19370), .B(n19368), .Z(n19369) );
  NANDN U20754 ( .A(n19329), .B(n19331), .Z(n19345) );
  XOR U20755 ( .A(n19371), .B(n19372), .Z(n19331) );
  AND U20756 ( .A(n758), .B(n19373), .Z(n19371) );
  XOR U20757 ( .A(n19372), .B(n19374), .Z(n19373) );
  XOR U20758 ( .A(n19375), .B(n19376), .Z(n758) );
  AND U20759 ( .A(n19377), .B(n19378), .Z(n19375) );
  XNOR U20760 ( .A(n19376), .B(n19342), .Z(n19378) );
  XNOR U20761 ( .A(n19379), .B(n19380), .Z(n19342) );
  ANDN U20762 ( .B(n19381), .A(n19382), .Z(n19379) );
  XOR U20763 ( .A(n19380), .B(n19383), .Z(n19381) );
  XOR U20764 ( .A(n19376), .B(n19344), .Z(n19377) );
  XOR U20765 ( .A(n19384), .B(n19385), .Z(n19344) );
  AND U20766 ( .A(n762), .B(n19386), .Z(n19384) );
  XOR U20767 ( .A(n19387), .B(n19385), .Z(n19386) );
  XNOR U20768 ( .A(n19388), .B(n19389), .Z(n19376) );
  NAND U20769 ( .A(n19390), .B(n19391), .Z(n19389) );
  XOR U20770 ( .A(n19392), .B(n19368), .Z(n19391) );
  XOR U20771 ( .A(n19382), .B(n19383), .Z(n19368) );
  XOR U20772 ( .A(n19393), .B(n19394), .Z(n19383) );
  ANDN U20773 ( .B(n19395), .A(n19396), .Z(n19393) );
  XOR U20774 ( .A(n19394), .B(n19397), .Z(n19395) );
  XOR U20775 ( .A(n19398), .B(n19399), .Z(n19382) );
  XOR U20776 ( .A(n19400), .B(n19401), .Z(n19399) );
  ANDN U20777 ( .B(n19402), .A(n19403), .Z(n19400) );
  XOR U20778 ( .A(n19404), .B(n19401), .Z(n19402) );
  IV U20779 ( .A(n19380), .Z(n19398) );
  XOR U20780 ( .A(n19405), .B(n19406), .Z(n19380) );
  ANDN U20781 ( .B(n19407), .A(n19408), .Z(n19405) );
  XOR U20782 ( .A(n19406), .B(n19409), .Z(n19407) );
  IV U20783 ( .A(n19388), .Z(n19392) );
  XOR U20784 ( .A(n19388), .B(n19370), .Z(n19390) );
  XOR U20785 ( .A(n19410), .B(n19411), .Z(n19370) );
  AND U20786 ( .A(n762), .B(n19412), .Z(n19410) );
  XOR U20787 ( .A(n19413), .B(n19411), .Z(n19412) );
  NANDN U20788 ( .A(n19372), .B(n19374), .Z(n19388) );
  XOR U20789 ( .A(n19414), .B(n19415), .Z(n19374) );
  AND U20790 ( .A(n762), .B(n19416), .Z(n19414) );
  XOR U20791 ( .A(n19415), .B(n19417), .Z(n19416) );
  XOR U20792 ( .A(n19418), .B(n19419), .Z(n762) );
  AND U20793 ( .A(n19420), .B(n19421), .Z(n19418) );
  XNOR U20794 ( .A(n19419), .B(n19385), .Z(n19421) );
  XNOR U20795 ( .A(n19422), .B(n19423), .Z(n19385) );
  ANDN U20796 ( .B(n19424), .A(n19425), .Z(n19422) );
  XOR U20797 ( .A(n19423), .B(n19426), .Z(n19424) );
  XOR U20798 ( .A(n19419), .B(n19387), .Z(n19420) );
  XOR U20799 ( .A(n19427), .B(n19428), .Z(n19387) );
  AND U20800 ( .A(n766), .B(n19429), .Z(n19427) );
  XOR U20801 ( .A(n19430), .B(n19428), .Z(n19429) );
  XNOR U20802 ( .A(n19431), .B(n19432), .Z(n19419) );
  NAND U20803 ( .A(n19433), .B(n19434), .Z(n19432) );
  XOR U20804 ( .A(n19435), .B(n19411), .Z(n19434) );
  XOR U20805 ( .A(n19425), .B(n19426), .Z(n19411) );
  XOR U20806 ( .A(n19436), .B(n19437), .Z(n19426) );
  ANDN U20807 ( .B(n19438), .A(n19439), .Z(n19436) );
  XOR U20808 ( .A(n19437), .B(n19440), .Z(n19438) );
  XOR U20809 ( .A(n19441), .B(n19442), .Z(n19425) );
  XOR U20810 ( .A(n19443), .B(n19444), .Z(n19442) );
  ANDN U20811 ( .B(n19445), .A(n19446), .Z(n19443) );
  XOR U20812 ( .A(n19447), .B(n19444), .Z(n19445) );
  IV U20813 ( .A(n19423), .Z(n19441) );
  XOR U20814 ( .A(n19448), .B(n19449), .Z(n19423) );
  ANDN U20815 ( .B(n19450), .A(n19451), .Z(n19448) );
  XOR U20816 ( .A(n19449), .B(n19452), .Z(n19450) );
  IV U20817 ( .A(n19431), .Z(n19435) );
  XOR U20818 ( .A(n19431), .B(n19413), .Z(n19433) );
  XOR U20819 ( .A(n19453), .B(n19454), .Z(n19413) );
  AND U20820 ( .A(n766), .B(n19455), .Z(n19453) );
  XOR U20821 ( .A(n19456), .B(n19454), .Z(n19455) );
  NANDN U20822 ( .A(n19415), .B(n19417), .Z(n19431) );
  XOR U20823 ( .A(n19457), .B(n19458), .Z(n19417) );
  AND U20824 ( .A(n766), .B(n19459), .Z(n19457) );
  XOR U20825 ( .A(n19458), .B(n19460), .Z(n19459) );
  XOR U20826 ( .A(n19461), .B(n19462), .Z(n766) );
  AND U20827 ( .A(n19463), .B(n19464), .Z(n19461) );
  XNOR U20828 ( .A(n19462), .B(n19428), .Z(n19464) );
  XNOR U20829 ( .A(n19465), .B(n19466), .Z(n19428) );
  ANDN U20830 ( .B(n19467), .A(n19468), .Z(n19465) );
  XOR U20831 ( .A(n19466), .B(n19469), .Z(n19467) );
  XOR U20832 ( .A(n19462), .B(n19430), .Z(n19463) );
  XOR U20833 ( .A(n19470), .B(n19471), .Z(n19430) );
  AND U20834 ( .A(n770), .B(n19472), .Z(n19470) );
  XOR U20835 ( .A(n19473), .B(n19471), .Z(n19472) );
  XNOR U20836 ( .A(n19474), .B(n19475), .Z(n19462) );
  NAND U20837 ( .A(n19476), .B(n19477), .Z(n19475) );
  XOR U20838 ( .A(n19478), .B(n19454), .Z(n19477) );
  XOR U20839 ( .A(n19468), .B(n19469), .Z(n19454) );
  XOR U20840 ( .A(n19479), .B(n19480), .Z(n19469) );
  ANDN U20841 ( .B(n19481), .A(n19482), .Z(n19479) );
  XOR U20842 ( .A(n19480), .B(n19483), .Z(n19481) );
  XOR U20843 ( .A(n19484), .B(n19485), .Z(n19468) );
  XOR U20844 ( .A(n19486), .B(n19487), .Z(n19485) );
  ANDN U20845 ( .B(n19488), .A(n19489), .Z(n19486) );
  XOR U20846 ( .A(n19490), .B(n19487), .Z(n19488) );
  IV U20847 ( .A(n19466), .Z(n19484) );
  XOR U20848 ( .A(n19491), .B(n19492), .Z(n19466) );
  ANDN U20849 ( .B(n19493), .A(n19494), .Z(n19491) );
  XOR U20850 ( .A(n19492), .B(n19495), .Z(n19493) );
  IV U20851 ( .A(n19474), .Z(n19478) );
  XOR U20852 ( .A(n19474), .B(n19456), .Z(n19476) );
  XOR U20853 ( .A(n19496), .B(n19497), .Z(n19456) );
  AND U20854 ( .A(n770), .B(n19498), .Z(n19496) );
  XOR U20855 ( .A(n19499), .B(n19497), .Z(n19498) );
  NANDN U20856 ( .A(n19458), .B(n19460), .Z(n19474) );
  XOR U20857 ( .A(n19500), .B(n19501), .Z(n19460) );
  AND U20858 ( .A(n770), .B(n19502), .Z(n19500) );
  XOR U20859 ( .A(n19501), .B(n19503), .Z(n19502) );
  XOR U20860 ( .A(n19504), .B(n19505), .Z(n770) );
  AND U20861 ( .A(n19506), .B(n19507), .Z(n19504) );
  XNOR U20862 ( .A(n19505), .B(n19471), .Z(n19507) );
  XNOR U20863 ( .A(n19508), .B(n19509), .Z(n19471) );
  ANDN U20864 ( .B(n19510), .A(n19511), .Z(n19508) );
  XOR U20865 ( .A(n19509), .B(n19512), .Z(n19510) );
  XOR U20866 ( .A(n19505), .B(n19473), .Z(n19506) );
  XOR U20867 ( .A(n19513), .B(n19514), .Z(n19473) );
  AND U20868 ( .A(n774), .B(n19515), .Z(n19513) );
  XOR U20869 ( .A(n19516), .B(n19514), .Z(n19515) );
  XNOR U20870 ( .A(n19517), .B(n19518), .Z(n19505) );
  NAND U20871 ( .A(n19519), .B(n19520), .Z(n19518) );
  XOR U20872 ( .A(n19521), .B(n19497), .Z(n19520) );
  XOR U20873 ( .A(n19511), .B(n19512), .Z(n19497) );
  XOR U20874 ( .A(n19522), .B(n19523), .Z(n19512) );
  ANDN U20875 ( .B(n19524), .A(n19525), .Z(n19522) );
  XOR U20876 ( .A(n19523), .B(n19526), .Z(n19524) );
  XOR U20877 ( .A(n19527), .B(n19528), .Z(n19511) );
  XOR U20878 ( .A(n19529), .B(n19530), .Z(n19528) );
  ANDN U20879 ( .B(n19531), .A(n19532), .Z(n19529) );
  XOR U20880 ( .A(n19533), .B(n19530), .Z(n19531) );
  IV U20881 ( .A(n19509), .Z(n19527) );
  XOR U20882 ( .A(n19534), .B(n19535), .Z(n19509) );
  ANDN U20883 ( .B(n19536), .A(n19537), .Z(n19534) );
  XOR U20884 ( .A(n19535), .B(n19538), .Z(n19536) );
  IV U20885 ( .A(n19517), .Z(n19521) );
  XOR U20886 ( .A(n19517), .B(n19499), .Z(n19519) );
  XOR U20887 ( .A(n19539), .B(n19540), .Z(n19499) );
  AND U20888 ( .A(n774), .B(n19541), .Z(n19539) );
  XOR U20889 ( .A(n19542), .B(n19540), .Z(n19541) );
  NANDN U20890 ( .A(n19501), .B(n19503), .Z(n19517) );
  XOR U20891 ( .A(n19543), .B(n19544), .Z(n19503) );
  AND U20892 ( .A(n774), .B(n19545), .Z(n19543) );
  XOR U20893 ( .A(n19544), .B(n19546), .Z(n19545) );
  XOR U20894 ( .A(n19547), .B(n19548), .Z(n774) );
  AND U20895 ( .A(n19549), .B(n19550), .Z(n19547) );
  XNOR U20896 ( .A(n19548), .B(n19514), .Z(n19550) );
  XNOR U20897 ( .A(n19551), .B(n19552), .Z(n19514) );
  ANDN U20898 ( .B(n19553), .A(n19554), .Z(n19551) );
  XOR U20899 ( .A(n19552), .B(n19555), .Z(n19553) );
  XOR U20900 ( .A(n19548), .B(n19516), .Z(n19549) );
  XOR U20901 ( .A(n19556), .B(n19557), .Z(n19516) );
  AND U20902 ( .A(n778), .B(n19558), .Z(n19556) );
  XOR U20903 ( .A(n19559), .B(n19557), .Z(n19558) );
  XNOR U20904 ( .A(n19560), .B(n19561), .Z(n19548) );
  NAND U20905 ( .A(n19562), .B(n19563), .Z(n19561) );
  XOR U20906 ( .A(n19564), .B(n19540), .Z(n19563) );
  XOR U20907 ( .A(n19554), .B(n19555), .Z(n19540) );
  XOR U20908 ( .A(n19565), .B(n19566), .Z(n19555) );
  ANDN U20909 ( .B(n19567), .A(n19568), .Z(n19565) );
  XOR U20910 ( .A(n19566), .B(n19569), .Z(n19567) );
  XOR U20911 ( .A(n19570), .B(n19571), .Z(n19554) );
  XOR U20912 ( .A(n19572), .B(n19573), .Z(n19571) );
  ANDN U20913 ( .B(n19574), .A(n19575), .Z(n19572) );
  XOR U20914 ( .A(n19576), .B(n19573), .Z(n19574) );
  IV U20915 ( .A(n19552), .Z(n19570) );
  XOR U20916 ( .A(n19577), .B(n19578), .Z(n19552) );
  ANDN U20917 ( .B(n19579), .A(n19580), .Z(n19577) );
  XOR U20918 ( .A(n19578), .B(n19581), .Z(n19579) );
  IV U20919 ( .A(n19560), .Z(n19564) );
  XOR U20920 ( .A(n19560), .B(n19542), .Z(n19562) );
  XOR U20921 ( .A(n19582), .B(n19583), .Z(n19542) );
  AND U20922 ( .A(n778), .B(n19584), .Z(n19582) );
  XOR U20923 ( .A(n19585), .B(n19583), .Z(n19584) );
  NANDN U20924 ( .A(n19544), .B(n19546), .Z(n19560) );
  XOR U20925 ( .A(n19586), .B(n19587), .Z(n19546) );
  AND U20926 ( .A(n778), .B(n19588), .Z(n19586) );
  XOR U20927 ( .A(n19587), .B(n19589), .Z(n19588) );
  XOR U20928 ( .A(n19590), .B(n19591), .Z(n778) );
  AND U20929 ( .A(n19592), .B(n19593), .Z(n19590) );
  XNOR U20930 ( .A(n19591), .B(n19557), .Z(n19593) );
  XNOR U20931 ( .A(n19594), .B(n19595), .Z(n19557) );
  ANDN U20932 ( .B(n19596), .A(n19597), .Z(n19594) );
  XOR U20933 ( .A(n19595), .B(n19598), .Z(n19596) );
  XOR U20934 ( .A(n19591), .B(n19559), .Z(n19592) );
  XOR U20935 ( .A(n19599), .B(n19600), .Z(n19559) );
  AND U20936 ( .A(n782), .B(n19601), .Z(n19599) );
  XOR U20937 ( .A(n19602), .B(n19600), .Z(n19601) );
  XNOR U20938 ( .A(n19603), .B(n19604), .Z(n19591) );
  NAND U20939 ( .A(n19605), .B(n19606), .Z(n19604) );
  XOR U20940 ( .A(n19607), .B(n19583), .Z(n19606) );
  XOR U20941 ( .A(n19597), .B(n19598), .Z(n19583) );
  XOR U20942 ( .A(n19608), .B(n19609), .Z(n19598) );
  ANDN U20943 ( .B(n19610), .A(n19611), .Z(n19608) );
  XOR U20944 ( .A(n19609), .B(n19612), .Z(n19610) );
  XOR U20945 ( .A(n19613), .B(n19614), .Z(n19597) );
  XOR U20946 ( .A(n19615), .B(n19616), .Z(n19614) );
  ANDN U20947 ( .B(n19617), .A(n19618), .Z(n19615) );
  XOR U20948 ( .A(n19619), .B(n19616), .Z(n19617) );
  IV U20949 ( .A(n19595), .Z(n19613) );
  XOR U20950 ( .A(n19620), .B(n19621), .Z(n19595) );
  ANDN U20951 ( .B(n19622), .A(n19623), .Z(n19620) );
  XOR U20952 ( .A(n19621), .B(n19624), .Z(n19622) );
  IV U20953 ( .A(n19603), .Z(n19607) );
  XOR U20954 ( .A(n19603), .B(n19585), .Z(n19605) );
  XOR U20955 ( .A(n19625), .B(n19626), .Z(n19585) );
  AND U20956 ( .A(n782), .B(n19627), .Z(n19625) );
  XOR U20957 ( .A(n19628), .B(n19626), .Z(n19627) );
  NANDN U20958 ( .A(n19587), .B(n19589), .Z(n19603) );
  XOR U20959 ( .A(n19629), .B(n19630), .Z(n19589) );
  AND U20960 ( .A(n782), .B(n19631), .Z(n19629) );
  XOR U20961 ( .A(n19630), .B(n19632), .Z(n19631) );
  XOR U20962 ( .A(n19633), .B(n19634), .Z(n782) );
  AND U20963 ( .A(n19635), .B(n19636), .Z(n19633) );
  XNOR U20964 ( .A(n19634), .B(n19600), .Z(n19636) );
  XNOR U20965 ( .A(n19637), .B(n19638), .Z(n19600) );
  ANDN U20966 ( .B(n19639), .A(n19640), .Z(n19637) );
  XOR U20967 ( .A(n19638), .B(n19641), .Z(n19639) );
  XOR U20968 ( .A(n19634), .B(n19602), .Z(n19635) );
  XOR U20969 ( .A(n19642), .B(n19643), .Z(n19602) );
  AND U20970 ( .A(n786), .B(n19644), .Z(n19642) );
  XOR U20971 ( .A(n19645), .B(n19643), .Z(n19644) );
  XNOR U20972 ( .A(n19646), .B(n19647), .Z(n19634) );
  NAND U20973 ( .A(n19648), .B(n19649), .Z(n19647) );
  XOR U20974 ( .A(n19650), .B(n19626), .Z(n19649) );
  XOR U20975 ( .A(n19640), .B(n19641), .Z(n19626) );
  XOR U20976 ( .A(n19651), .B(n19652), .Z(n19641) );
  ANDN U20977 ( .B(n19653), .A(n19654), .Z(n19651) );
  XOR U20978 ( .A(n19652), .B(n19655), .Z(n19653) );
  XOR U20979 ( .A(n19656), .B(n19657), .Z(n19640) );
  XOR U20980 ( .A(n19658), .B(n19659), .Z(n19657) );
  ANDN U20981 ( .B(n19660), .A(n19661), .Z(n19658) );
  XOR U20982 ( .A(n19662), .B(n19659), .Z(n19660) );
  IV U20983 ( .A(n19638), .Z(n19656) );
  XOR U20984 ( .A(n19663), .B(n19664), .Z(n19638) );
  ANDN U20985 ( .B(n19665), .A(n19666), .Z(n19663) );
  XOR U20986 ( .A(n19664), .B(n19667), .Z(n19665) );
  IV U20987 ( .A(n19646), .Z(n19650) );
  XOR U20988 ( .A(n19646), .B(n19628), .Z(n19648) );
  XOR U20989 ( .A(n19668), .B(n19669), .Z(n19628) );
  AND U20990 ( .A(n786), .B(n19670), .Z(n19668) );
  XOR U20991 ( .A(n19671), .B(n19669), .Z(n19670) );
  NANDN U20992 ( .A(n19630), .B(n19632), .Z(n19646) );
  XOR U20993 ( .A(n19672), .B(n19673), .Z(n19632) );
  AND U20994 ( .A(n786), .B(n19674), .Z(n19672) );
  XOR U20995 ( .A(n19673), .B(n19675), .Z(n19674) );
  XOR U20996 ( .A(n19676), .B(n19677), .Z(n786) );
  AND U20997 ( .A(n19678), .B(n19679), .Z(n19676) );
  XNOR U20998 ( .A(n19677), .B(n19643), .Z(n19679) );
  XNOR U20999 ( .A(n19680), .B(n19681), .Z(n19643) );
  ANDN U21000 ( .B(n19682), .A(n19683), .Z(n19680) );
  XOR U21001 ( .A(n19681), .B(n19684), .Z(n19682) );
  XOR U21002 ( .A(n19677), .B(n19645), .Z(n19678) );
  XOR U21003 ( .A(n19685), .B(n19686), .Z(n19645) );
  AND U21004 ( .A(n790), .B(n19687), .Z(n19685) );
  XOR U21005 ( .A(n19688), .B(n19686), .Z(n19687) );
  XNOR U21006 ( .A(n19689), .B(n19690), .Z(n19677) );
  NAND U21007 ( .A(n19691), .B(n19692), .Z(n19690) );
  XOR U21008 ( .A(n19693), .B(n19669), .Z(n19692) );
  XOR U21009 ( .A(n19683), .B(n19684), .Z(n19669) );
  XOR U21010 ( .A(n19694), .B(n19695), .Z(n19684) );
  ANDN U21011 ( .B(n19696), .A(n19697), .Z(n19694) );
  XOR U21012 ( .A(n19695), .B(n19698), .Z(n19696) );
  XOR U21013 ( .A(n19699), .B(n19700), .Z(n19683) );
  XOR U21014 ( .A(n19701), .B(n19702), .Z(n19700) );
  ANDN U21015 ( .B(n19703), .A(n19704), .Z(n19701) );
  XOR U21016 ( .A(n19705), .B(n19702), .Z(n19703) );
  IV U21017 ( .A(n19681), .Z(n19699) );
  XOR U21018 ( .A(n19706), .B(n19707), .Z(n19681) );
  ANDN U21019 ( .B(n19708), .A(n19709), .Z(n19706) );
  XOR U21020 ( .A(n19707), .B(n19710), .Z(n19708) );
  IV U21021 ( .A(n19689), .Z(n19693) );
  XOR U21022 ( .A(n19689), .B(n19671), .Z(n19691) );
  XOR U21023 ( .A(n19711), .B(n19712), .Z(n19671) );
  AND U21024 ( .A(n790), .B(n19713), .Z(n19711) );
  XOR U21025 ( .A(n19714), .B(n19712), .Z(n19713) );
  NANDN U21026 ( .A(n19673), .B(n19675), .Z(n19689) );
  XOR U21027 ( .A(n19715), .B(n19716), .Z(n19675) );
  AND U21028 ( .A(n790), .B(n19717), .Z(n19715) );
  XOR U21029 ( .A(n19716), .B(n19718), .Z(n19717) );
  XOR U21030 ( .A(n19719), .B(n19720), .Z(n790) );
  AND U21031 ( .A(n19721), .B(n19722), .Z(n19719) );
  XNOR U21032 ( .A(n19720), .B(n19686), .Z(n19722) );
  XNOR U21033 ( .A(n19723), .B(n19724), .Z(n19686) );
  ANDN U21034 ( .B(n19725), .A(n19726), .Z(n19723) );
  XOR U21035 ( .A(n19724), .B(n19727), .Z(n19725) );
  XOR U21036 ( .A(n19720), .B(n19688), .Z(n19721) );
  XOR U21037 ( .A(n19728), .B(n19729), .Z(n19688) );
  AND U21038 ( .A(n794), .B(n19730), .Z(n19728) );
  XOR U21039 ( .A(n19731), .B(n19729), .Z(n19730) );
  XNOR U21040 ( .A(n19732), .B(n19733), .Z(n19720) );
  NAND U21041 ( .A(n19734), .B(n19735), .Z(n19733) );
  XOR U21042 ( .A(n19736), .B(n19712), .Z(n19735) );
  XOR U21043 ( .A(n19726), .B(n19727), .Z(n19712) );
  XOR U21044 ( .A(n19737), .B(n19738), .Z(n19727) );
  ANDN U21045 ( .B(n19739), .A(n19740), .Z(n19737) );
  XOR U21046 ( .A(n19738), .B(n19741), .Z(n19739) );
  XOR U21047 ( .A(n19742), .B(n19743), .Z(n19726) );
  XOR U21048 ( .A(n19744), .B(n19745), .Z(n19743) );
  ANDN U21049 ( .B(n19746), .A(n19747), .Z(n19744) );
  XOR U21050 ( .A(n19748), .B(n19745), .Z(n19746) );
  IV U21051 ( .A(n19724), .Z(n19742) );
  XOR U21052 ( .A(n19749), .B(n19750), .Z(n19724) );
  ANDN U21053 ( .B(n19751), .A(n19752), .Z(n19749) );
  XOR U21054 ( .A(n19750), .B(n19753), .Z(n19751) );
  IV U21055 ( .A(n19732), .Z(n19736) );
  XOR U21056 ( .A(n19732), .B(n19714), .Z(n19734) );
  XOR U21057 ( .A(n19754), .B(n19755), .Z(n19714) );
  AND U21058 ( .A(n794), .B(n19756), .Z(n19754) );
  XOR U21059 ( .A(n19757), .B(n19755), .Z(n19756) );
  NANDN U21060 ( .A(n19716), .B(n19718), .Z(n19732) );
  XOR U21061 ( .A(n19758), .B(n19759), .Z(n19718) );
  AND U21062 ( .A(n794), .B(n19760), .Z(n19758) );
  XOR U21063 ( .A(n19759), .B(n19761), .Z(n19760) );
  XOR U21064 ( .A(n19762), .B(n19763), .Z(n794) );
  AND U21065 ( .A(n19764), .B(n19765), .Z(n19762) );
  XNOR U21066 ( .A(n19763), .B(n19729), .Z(n19765) );
  XNOR U21067 ( .A(n19766), .B(n19767), .Z(n19729) );
  ANDN U21068 ( .B(n19768), .A(n19769), .Z(n19766) );
  XOR U21069 ( .A(n19767), .B(n19770), .Z(n19768) );
  XOR U21070 ( .A(n19763), .B(n19731), .Z(n19764) );
  XOR U21071 ( .A(n19771), .B(n19772), .Z(n19731) );
  AND U21072 ( .A(n798), .B(n19773), .Z(n19771) );
  XOR U21073 ( .A(n19774), .B(n19772), .Z(n19773) );
  XNOR U21074 ( .A(n19775), .B(n19776), .Z(n19763) );
  NAND U21075 ( .A(n19777), .B(n19778), .Z(n19776) );
  XOR U21076 ( .A(n19779), .B(n19755), .Z(n19778) );
  XOR U21077 ( .A(n19769), .B(n19770), .Z(n19755) );
  XOR U21078 ( .A(n19780), .B(n19781), .Z(n19770) );
  ANDN U21079 ( .B(n19782), .A(n19783), .Z(n19780) );
  XOR U21080 ( .A(n19781), .B(n19784), .Z(n19782) );
  XOR U21081 ( .A(n19785), .B(n19786), .Z(n19769) );
  XOR U21082 ( .A(n19787), .B(n19788), .Z(n19786) );
  ANDN U21083 ( .B(n19789), .A(n19790), .Z(n19787) );
  XOR U21084 ( .A(n19791), .B(n19788), .Z(n19789) );
  IV U21085 ( .A(n19767), .Z(n19785) );
  XOR U21086 ( .A(n19792), .B(n19793), .Z(n19767) );
  ANDN U21087 ( .B(n19794), .A(n19795), .Z(n19792) );
  XOR U21088 ( .A(n19793), .B(n19796), .Z(n19794) );
  IV U21089 ( .A(n19775), .Z(n19779) );
  XOR U21090 ( .A(n19775), .B(n19757), .Z(n19777) );
  XOR U21091 ( .A(n19797), .B(n19798), .Z(n19757) );
  AND U21092 ( .A(n798), .B(n19799), .Z(n19797) );
  XOR U21093 ( .A(n19800), .B(n19798), .Z(n19799) );
  NANDN U21094 ( .A(n19759), .B(n19761), .Z(n19775) );
  XOR U21095 ( .A(n19801), .B(n19802), .Z(n19761) );
  AND U21096 ( .A(n798), .B(n19803), .Z(n19801) );
  XOR U21097 ( .A(n19802), .B(n19804), .Z(n19803) );
  XOR U21098 ( .A(n19805), .B(n19806), .Z(n798) );
  AND U21099 ( .A(n19807), .B(n19808), .Z(n19805) );
  XNOR U21100 ( .A(n19806), .B(n19772), .Z(n19808) );
  XNOR U21101 ( .A(n19809), .B(n19810), .Z(n19772) );
  ANDN U21102 ( .B(n19811), .A(n19812), .Z(n19809) );
  XOR U21103 ( .A(n19810), .B(n19813), .Z(n19811) );
  XOR U21104 ( .A(n19806), .B(n19774), .Z(n19807) );
  XOR U21105 ( .A(n19814), .B(n19815), .Z(n19774) );
  AND U21106 ( .A(n802), .B(n19816), .Z(n19814) );
  XOR U21107 ( .A(n19817), .B(n19815), .Z(n19816) );
  XNOR U21108 ( .A(n19818), .B(n19819), .Z(n19806) );
  NAND U21109 ( .A(n19820), .B(n19821), .Z(n19819) );
  XOR U21110 ( .A(n19822), .B(n19798), .Z(n19821) );
  XOR U21111 ( .A(n19812), .B(n19813), .Z(n19798) );
  XOR U21112 ( .A(n19823), .B(n19824), .Z(n19813) );
  ANDN U21113 ( .B(n19825), .A(n19826), .Z(n19823) );
  XOR U21114 ( .A(n19824), .B(n19827), .Z(n19825) );
  XOR U21115 ( .A(n19828), .B(n19829), .Z(n19812) );
  XOR U21116 ( .A(n19830), .B(n19831), .Z(n19829) );
  ANDN U21117 ( .B(n19832), .A(n19833), .Z(n19830) );
  XOR U21118 ( .A(n19834), .B(n19831), .Z(n19832) );
  IV U21119 ( .A(n19810), .Z(n19828) );
  XOR U21120 ( .A(n19835), .B(n19836), .Z(n19810) );
  ANDN U21121 ( .B(n19837), .A(n19838), .Z(n19835) );
  XOR U21122 ( .A(n19836), .B(n19839), .Z(n19837) );
  IV U21123 ( .A(n19818), .Z(n19822) );
  XOR U21124 ( .A(n19818), .B(n19800), .Z(n19820) );
  XOR U21125 ( .A(n19840), .B(n19841), .Z(n19800) );
  AND U21126 ( .A(n802), .B(n19842), .Z(n19840) );
  XOR U21127 ( .A(n19843), .B(n19841), .Z(n19842) );
  NANDN U21128 ( .A(n19802), .B(n19804), .Z(n19818) );
  XOR U21129 ( .A(n19844), .B(n19845), .Z(n19804) );
  AND U21130 ( .A(n802), .B(n19846), .Z(n19844) );
  XOR U21131 ( .A(n19845), .B(n19847), .Z(n19846) );
  XOR U21132 ( .A(n19848), .B(n19849), .Z(n802) );
  AND U21133 ( .A(n19850), .B(n19851), .Z(n19848) );
  XNOR U21134 ( .A(n19849), .B(n19815), .Z(n19851) );
  XNOR U21135 ( .A(n19852), .B(n19853), .Z(n19815) );
  ANDN U21136 ( .B(n19854), .A(n19855), .Z(n19852) );
  XOR U21137 ( .A(n19853), .B(n19856), .Z(n19854) );
  XOR U21138 ( .A(n19849), .B(n19817), .Z(n19850) );
  XOR U21139 ( .A(n19857), .B(n19858), .Z(n19817) );
  AND U21140 ( .A(n806), .B(n19859), .Z(n19857) );
  XOR U21141 ( .A(n19860), .B(n19858), .Z(n19859) );
  XNOR U21142 ( .A(n19861), .B(n19862), .Z(n19849) );
  NAND U21143 ( .A(n19863), .B(n19864), .Z(n19862) );
  XOR U21144 ( .A(n19865), .B(n19841), .Z(n19864) );
  XOR U21145 ( .A(n19855), .B(n19856), .Z(n19841) );
  XOR U21146 ( .A(n19866), .B(n19867), .Z(n19856) );
  ANDN U21147 ( .B(n19868), .A(n19869), .Z(n19866) );
  XOR U21148 ( .A(n19867), .B(n19870), .Z(n19868) );
  XOR U21149 ( .A(n19871), .B(n19872), .Z(n19855) );
  XOR U21150 ( .A(n19873), .B(n19874), .Z(n19872) );
  ANDN U21151 ( .B(n19875), .A(n19876), .Z(n19873) );
  XOR U21152 ( .A(n19877), .B(n19874), .Z(n19875) );
  IV U21153 ( .A(n19853), .Z(n19871) );
  XOR U21154 ( .A(n19878), .B(n19879), .Z(n19853) );
  ANDN U21155 ( .B(n19880), .A(n19881), .Z(n19878) );
  XOR U21156 ( .A(n19879), .B(n19882), .Z(n19880) );
  IV U21157 ( .A(n19861), .Z(n19865) );
  XOR U21158 ( .A(n19861), .B(n19843), .Z(n19863) );
  XOR U21159 ( .A(n19883), .B(n19884), .Z(n19843) );
  AND U21160 ( .A(n806), .B(n19885), .Z(n19883) );
  XOR U21161 ( .A(n19886), .B(n19884), .Z(n19885) );
  NANDN U21162 ( .A(n19845), .B(n19847), .Z(n19861) );
  XOR U21163 ( .A(n19887), .B(n19888), .Z(n19847) );
  AND U21164 ( .A(n806), .B(n19889), .Z(n19887) );
  XOR U21165 ( .A(n19888), .B(n19890), .Z(n19889) );
  XOR U21166 ( .A(n19891), .B(n19892), .Z(n806) );
  AND U21167 ( .A(n19893), .B(n19894), .Z(n19891) );
  XNOR U21168 ( .A(n19892), .B(n19858), .Z(n19894) );
  XNOR U21169 ( .A(n19895), .B(n19896), .Z(n19858) );
  ANDN U21170 ( .B(n19897), .A(n19898), .Z(n19895) );
  XOR U21171 ( .A(n19896), .B(n19899), .Z(n19897) );
  XOR U21172 ( .A(n19892), .B(n19860), .Z(n19893) );
  XOR U21173 ( .A(n19900), .B(n19901), .Z(n19860) );
  AND U21174 ( .A(n810), .B(n19902), .Z(n19900) );
  XOR U21175 ( .A(n19903), .B(n19901), .Z(n19902) );
  XNOR U21176 ( .A(n19904), .B(n19905), .Z(n19892) );
  NAND U21177 ( .A(n19906), .B(n19907), .Z(n19905) );
  XOR U21178 ( .A(n19908), .B(n19884), .Z(n19907) );
  XOR U21179 ( .A(n19898), .B(n19899), .Z(n19884) );
  XOR U21180 ( .A(n19909), .B(n19910), .Z(n19899) );
  ANDN U21181 ( .B(n19911), .A(n19912), .Z(n19909) );
  XOR U21182 ( .A(n19910), .B(n19913), .Z(n19911) );
  XOR U21183 ( .A(n19914), .B(n19915), .Z(n19898) );
  XOR U21184 ( .A(n19916), .B(n19917), .Z(n19915) );
  ANDN U21185 ( .B(n19918), .A(n19919), .Z(n19916) );
  XOR U21186 ( .A(n19920), .B(n19917), .Z(n19918) );
  IV U21187 ( .A(n19896), .Z(n19914) );
  XOR U21188 ( .A(n19921), .B(n19922), .Z(n19896) );
  ANDN U21189 ( .B(n19923), .A(n19924), .Z(n19921) );
  XOR U21190 ( .A(n19922), .B(n19925), .Z(n19923) );
  IV U21191 ( .A(n19904), .Z(n19908) );
  XOR U21192 ( .A(n19904), .B(n19886), .Z(n19906) );
  XOR U21193 ( .A(n19926), .B(n19927), .Z(n19886) );
  AND U21194 ( .A(n810), .B(n19928), .Z(n19926) );
  XOR U21195 ( .A(n19929), .B(n19927), .Z(n19928) );
  NANDN U21196 ( .A(n19888), .B(n19890), .Z(n19904) );
  XOR U21197 ( .A(n19930), .B(n19931), .Z(n19890) );
  AND U21198 ( .A(n810), .B(n19932), .Z(n19930) );
  XOR U21199 ( .A(n19931), .B(n19933), .Z(n19932) );
  XOR U21200 ( .A(n19934), .B(n19935), .Z(n810) );
  AND U21201 ( .A(n19936), .B(n19937), .Z(n19934) );
  XNOR U21202 ( .A(n19935), .B(n19901), .Z(n19937) );
  XNOR U21203 ( .A(n19938), .B(n19939), .Z(n19901) );
  ANDN U21204 ( .B(n19940), .A(n19941), .Z(n19938) );
  XOR U21205 ( .A(n19939), .B(n19942), .Z(n19940) );
  XOR U21206 ( .A(n19935), .B(n19903), .Z(n19936) );
  XOR U21207 ( .A(n19943), .B(n19944), .Z(n19903) );
  AND U21208 ( .A(n814), .B(n19945), .Z(n19943) );
  XOR U21209 ( .A(n19946), .B(n19944), .Z(n19945) );
  XNOR U21210 ( .A(n19947), .B(n19948), .Z(n19935) );
  NAND U21211 ( .A(n19949), .B(n19950), .Z(n19948) );
  XOR U21212 ( .A(n19951), .B(n19927), .Z(n19950) );
  XOR U21213 ( .A(n19941), .B(n19942), .Z(n19927) );
  XOR U21214 ( .A(n19952), .B(n19953), .Z(n19942) );
  ANDN U21215 ( .B(n19954), .A(n19955), .Z(n19952) );
  XOR U21216 ( .A(n19953), .B(n19956), .Z(n19954) );
  XOR U21217 ( .A(n19957), .B(n19958), .Z(n19941) );
  XOR U21218 ( .A(n19959), .B(n19960), .Z(n19958) );
  ANDN U21219 ( .B(n19961), .A(n19962), .Z(n19959) );
  XOR U21220 ( .A(n19963), .B(n19960), .Z(n19961) );
  IV U21221 ( .A(n19939), .Z(n19957) );
  XOR U21222 ( .A(n19964), .B(n19965), .Z(n19939) );
  ANDN U21223 ( .B(n19966), .A(n19967), .Z(n19964) );
  XOR U21224 ( .A(n19965), .B(n19968), .Z(n19966) );
  IV U21225 ( .A(n19947), .Z(n19951) );
  XOR U21226 ( .A(n19947), .B(n19929), .Z(n19949) );
  XOR U21227 ( .A(n19969), .B(n19970), .Z(n19929) );
  AND U21228 ( .A(n814), .B(n19971), .Z(n19969) );
  XOR U21229 ( .A(n19972), .B(n19970), .Z(n19971) );
  NANDN U21230 ( .A(n19931), .B(n19933), .Z(n19947) );
  XOR U21231 ( .A(n19973), .B(n19974), .Z(n19933) );
  AND U21232 ( .A(n814), .B(n19975), .Z(n19973) );
  XOR U21233 ( .A(n19974), .B(n19976), .Z(n19975) );
  XOR U21234 ( .A(n19977), .B(n19978), .Z(n814) );
  AND U21235 ( .A(n19979), .B(n19980), .Z(n19977) );
  XNOR U21236 ( .A(n19978), .B(n19944), .Z(n19980) );
  XNOR U21237 ( .A(n19981), .B(n19982), .Z(n19944) );
  ANDN U21238 ( .B(n19983), .A(n19984), .Z(n19981) );
  XOR U21239 ( .A(n19982), .B(n19985), .Z(n19983) );
  XOR U21240 ( .A(n19978), .B(n19946), .Z(n19979) );
  XOR U21241 ( .A(n19986), .B(n19987), .Z(n19946) );
  AND U21242 ( .A(n818), .B(n19988), .Z(n19986) );
  XOR U21243 ( .A(n19989), .B(n19987), .Z(n19988) );
  XNOR U21244 ( .A(n19990), .B(n19991), .Z(n19978) );
  NAND U21245 ( .A(n19992), .B(n19993), .Z(n19991) );
  XOR U21246 ( .A(n19994), .B(n19970), .Z(n19993) );
  XOR U21247 ( .A(n19984), .B(n19985), .Z(n19970) );
  XOR U21248 ( .A(n19995), .B(n19996), .Z(n19985) );
  ANDN U21249 ( .B(n19997), .A(n19998), .Z(n19995) );
  XOR U21250 ( .A(n19996), .B(n19999), .Z(n19997) );
  XOR U21251 ( .A(n20000), .B(n20001), .Z(n19984) );
  XOR U21252 ( .A(n20002), .B(n20003), .Z(n20001) );
  ANDN U21253 ( .B(n20004), .A(n20005), .Z(n20002) );
  XOR U21254 ( .A(n20006), .B(n20003), .Z(n20004) );
  IV U21255 ( .A(n19982), .Z(n20000) );
  XOR U21256 ( .A(n20007), .B(n20008), .Z(n19982) );
  ANDN U21257 ( .B(n20009), .A(n20010), .Z(n20007) );
  XOR U21258 ( .A(n20008), .B(n20011), .Z(n20009) );
  IV U21259 ( .A(n19990), .Z(n19994) );
  XOR U21260 ( .A(n19990), .B(n19972), .Z(n19992) );
  XOR U21261 ( .A(n20012), .B(n20013), .Z(n19972) );
  AND U21262 ( .A(n818), .B(n20014), .Z(n20012) );
  XOR U21263 ( .A(n20015), .B(n20013), .Z(n20014) );
  NANDN U21264 ( .A(n19974), .B(n19976), .Z(n19990) );
  XOR U21265 ( .A(n20016), .B(n20017), .Z(n19976) );
  AND U21266 ( .A(n818), .B(n20018), .Z(n20016) );
  XOR U21267 ( .A(n20017), .B(n20019), .Z(n20018) );
  XOR U21268 ( .A(n20020), .B(n20021), .Z(n818) );
  AND U21269 ( .A(n20022), .B(n20023), .Z(n20020) );
  XNOR U21270 ( .A(n20021), .B(n19987), .Z(n20023) );
  XNOR U21271 ( .A(n20024), .B(n20025), .Z(n19987) );
  ANDN U21272 ( .B(n20026), .A(n20027), .Z(n20024) );
  XOR U21273 ( .A(n20025), .B(n20028), .Z(n20026) );
  XOR U21274 ( .A(n20021), .B(n19989), .Z(n20022) );
  XOR U21275 ( .A(n20029), .B(n20030), .Z(n19989) );
  AND U21276 ( .A(n822), .B(n20031), .Z(n20029) );
  XOR U21277 ( .A(n20032), .B(n20030), .Z(n20031) );
  XNOR U21278 ( .A(n20033), .B(n20034), .Z(n20021) );
  NAND U21279 ( .A(n20035), .B(n20036), .Z(n20034) );
  XOR U21280 ( .A(n20037), .B(n20013), .Z(n20036) );
  XOR U21281 ( .A(n20027), .B(n20028), .Z(n20013) );
  XOR U21282 ( .A(n20038), .B(n20039), .Z(n20028) );
  ANDN U21283 ( .B(n20040), .A(n20041), .Z(n20038) );
  XOR U21284 ( .A(n20039), .B(n20042), .Z(n20040) );
  XOR U21285 ( .A(n20043), .B(n20044), .Z(n20027) );
  XOR U21286 ( .A(n20045), .B(n20046), .Z(n20044) );
  ANDN U21287 ( .B(n20047), .A(n20048), .Z(n20045) );
  XOR U21288 ( .A(n20049), .B(n20046), .Z(n20047) );
  IV U21289 ( .A(n20025), .Z(n20043) );
  XOR U21290 ( .A(n20050), .B(n20051), .Z(n20025) );
  ANDN U21291 ( .B(n20052), .A(n20053), .Z(n20050) );
  XOR U21292 ( .A(n20051), .B(n20054), .Z(n20052) );
  IV U21293 ( .A(n20033), .Z(n20037) );
  XOR U21294 ( .A(n20033), .B(n20015), .Z(n20035) );
  XOR U21295 ( .A(n20055), .B(n20056), .Z(n20015) );
  AND U21296 ( .A(n822), .B(n20057), .Z(n20055) );
  XOR U21297 ( .A(n20058), .B(n20056), .Z(n20057) );
  NANDN U21298 ( .A(n20017), .B(n20019), .Z(n20033) );
  XOR U21299 ( .A(n20059), .B(n20060), .Z(n20019) );
  AND U21300 ( .A(n822), .B(n20061), .Z(n20059) );
  XOR U21301 ( .A(n20060), .B(n20062), .Z(n20061) );
  XOR U21302 ( .A(n20063), .B(n20064), .Z(n822) );
  AND U21303 ( .A(n20065), .B(n20066), .Z(n20063) );
  XNOR U21304 ( .A(n20064), .B(n20030), .Z(n20066) );
  XNOR U21305 ( .A(n20067), .B(n20068), .Z(n20030) );
  ANDN U21306 ( .B(n20069), .A(n20070), .Z(n20067) );
  XOR U21307 ( .A(n20068), .B(n20071), .Z(n20069) );
  XOR U21308 ( .A(n20064), .B(n20032), .Z(n20065) );
  XOR U21309 ( .A(n20072), .B(n20073), .Z(n20032) );
  AND U21310 ( .A(n826), .B(n20074), .Z(n20072) );
  XOR U21311 ( .A(n20075), .B(n20073), .Z(n20074) );
  XNOR U21312 ( .A(n20076), .B(n20077), .Z(n20064) );
  NAND U21313 ( .A(n20078), .B(n20079), .Z(n20077) );
  XOR U21314 ( .A(n20080), .B(n20056), .Z(n20079) );
  XOR U21315 ( .A(n20070), .B(n20071), .Z(n20056) );
  XOR U21316 ( .A(n20081), .B(n20082), .Z(n20071) );
  ANDN U21317 ( .B(n20083), .A(n20084), .Z(n20081) );
  XOR U21318 ( .A(n20082), .B(n20085), .Z(n20083) );
  XOR U21319 ( .A(n20086), .B(n20087), .Z(n20070) );
  XOR U21320 ( .A(n20088), .B(n20089), .Z(n20087) );
  ANDN U21321 ( .B(n20090), .A(n20091), .Z(n20088) );
  XOR U21322 ( .A(n20092), .B(n20089), .Z(n20090) );
  IV U21323 ( .A(n20068), .Z(n20086) );
  XOR U21324 ( .A(n20093), .B(n20094), .Z(n20068) );
  ANDN U21325 ( .B(n20095), .A(n20096), .Z(n20093) );
  XOR U21326 ( .A(n20094), .B(n20097), .Z(n20095) );
  IV U21327 ( .A(n20076), .Z(n20080) );
  XOR U21328 ( .A(n20076), .B(n20058), .Z(n20078) );
  XOR U21329 ( .A(n20098), .B(n20099), .Z(n20058) );
  AND U21330 ( .A(n826), .B(n20100), .Z(n20098) );
  XOR U21331 ( .A(n20101), .B(n20099), .Z(n20100) );
  NANDN U21332 ( .A(n20060), .B(n20062), .Z(n20076) );
  XOR U21333 ( .A(n20102), .B(n20103), .Z(n20062) );
  AND U21334 ( .A(n826), .B(n20104), .Z(n20102) );
  XOR U21335 ( .A(n20103), .B(n20105), .Z(n20104) );
  XOR U21336 ( .A(n20106), .B(n20107), .Z(n826) );
  AND U21337 ( .A(n20108), .B(n20109), .Z(n20106) );
  XNOR U21338 ( .A(n20107), .B(n20073), .Z(n20109) );
  XNOR U21339 ( .A(n20110), .B(n20111), .Z(n20073) );
  ANDN U21340 ( .B(n20112), .A(n20113), .Z(n20110) );
  XOR U21341 ( .A(n20111), .B(n20114), .Z(n20112) );
  XOR U21342 ( .A(n20107), .B(n20075), .Z(n20108) );
  XOR U21343 ( .A(n20115), .B(n20116), .Z(n20075) );
  AND U21344 ( .A(n830), .B(n20117), .Z(n20115) );
  XOR U21345 ( .A(n20118), .B(n20116), .Z(n20117) );
  XNOR U21346 ( .A(n20119), .B(n20120), .Z(n20107) );
  NAND U21347 ( .A(n20121), .B(n20122), .Z(n20120) );
  XOR U21348 ( .A(n20123), .B(n20099), .Z(n20122) );
  XOR U21349 ( .A(n20113), .B(n20114), .Z(n20099) );
  XOR U21350 ( .A(n20124), .B(n20125), .Z(n20114) );
  ANDN U21351 ( .B(n20126), .A(n20127), .Z(n20124) );
  XOR U21352 ( .A(n20125), .B(n20128), .Z(n20126) );
  XOR U21353 ( .A(n20129), .B(n20130), .Z(n20113) );
  XOR U21354 ( .A(n20131), .B(n20132), .Z(n20130) );
  ANDN U21355 ( .B(n20133), .A(n20134), .Z(n20131) );
  XOR U21356 ( .A(n20135), .B(n20132), .Z(n20133) );
  IV U21357 ( .A(n20111), .Z(n20129) );
  XOR U21358 ( .A(n20136), .B(n20137), .Z(n20111) );
  ANDN U21359 ( .B(n20138), .A(n20139), .Z(n20136) );
  XOR U21360 ( .A(n20137), .B(n20140), .Z(n20138) );
  IV U21361 ( .A(n20119), .Z(n20123) );
  XOR U21362 ( .A(n20119), .B(n20101), .Z(n20121) );
  XOR U21363 ( .A(n20141), .B(n20142), .Z(n20101) );
  AND U21364 ( .A(n830), .B(n20143), .Z(n20141) );
  XOR U21365 ( .A(n20144), .B(n20142), .Z(n20143) );
  NANDN U21366 ( .A(n20103), .B(n20105), .Z(n20119) );
  XOR U21367 ( .A(n20145), .B(n20146), .Z(n20105) );
  AND U21368 ( .A(n830), .B(n20147), .Z(n20145) );
  XOR U21369 ( .A(n20146), .B(n20148), .Z(n20147) );
  XOR U21370 ( .A(n20149), .B(n20150), .Z(n830) );
  AND U21371 ( .A(n20151), .B(n20152), .Z(n20149) );
  XNOR U21372 ( .A(n20150), .B(n20116), .Z(n20152) );
  XNOR U21373 ( .A(n20153), .B(n20154), .Z(n20116) );
  ANDN U21374 ( .B(n20155), .A(n20156), .Z(n20153) );
  XOR U21375 ( .A(n20154), .B(n20157), .Z(n20155) );
  XOR U21376 ( .A(n20150), .B(n20118), .Z(n20151) );
  XOR U21377 ( .A(n20158), .B(n20159), .Z(n20118) );
  AND U21378 ( .A(n834), .B(n20160), .Z(n20158) );
  XOR U21379 ( .A(n20161), .B(n20159), .Z(n20160) );
  XNOR U21380 ( .A(n20162), .B(n20163), .Z(n20150) );
  NAND U21381 ( .A(n20164), .B(n20165), .Z(n20163) );
  XOR U21382 ( .A(n20166), .B(n20142), .Z(n20165) );
  XOR U21383 ( .A(n20156), .B(n20157), .Z(n20142) );
  XOR U21384 ( .A(n20167), .B(n20168), .Z(n20157) );
  ANDN U21385 ( .B(n20169), .A(n20170), .Z(n20167) );
  XOR U21386 ( .A(n20168), .B(n20171), .Z(n20169) );
  XOR U21387 ( .A(n20172), .B(n20173), .Z(n20156) );
  XOR U21388 ( .A(n20174), .B(n20175), .Z(n20173) );
  ANDN U21389 ( .B(n20176), .A(n20177), .Z(n20174) );
  XOR U21390 ( .A(n20178), .B(n20175), .Z(n20176) );
  IV U21391 ( .A(n20154), .Z(n20172) );
  XOR U21392 ( .A(n20179), .B(n20180), .Z(n20154) );
  ANDN U21393 ( .B(n20181), .A(n20182), .Z(n20179) );
  XOR U21394 ( .A(n20180), .B(n20183), .Z(n20181) );
  IV U21395 ( .A(n20162), .Z(n20166) );
  XOR U21396 ( .A(n20162), .B(n20144), .Z(n20164) );
  XOR U21397 ( .A(n20184), .B(n20185), .Z(n20144) );
  AND U21398 ( .A(n834), .B(n20186), .Z(n20184) );
  XOR U21399 ( .A(n20187), .B(n20185), .Z(n20186) );
  NANDN U21400 ( .A(n20146), .B(n20148), .Z(n20162) );
  XOR U21401 ( .A(n20188), .B(n20189), .Z(n20148) );
  AND U21402 ( .A(n834), .B(n20190), .Z(n20188) );
  XOR U21403 ( .A(n20189), .B(n20191), .Z(n20190) );
  XOR U21404 ( .A(n20192), .B(n20193), .Z(n834) );
  AND U21405 ( .A(n20194), .B(n20195), .Z(n20192) );
  XNOR U21406 ( .A(n20193), .B(n20159), .Z(n20195) );
  XNOR U21407 ( .A(n20196), .B(n20197), .Z(n20159) );
  ANDN U21408 ( .B(n20198), .A(n20199), .Z(n20196) );
  XOR U21409 ( .A(n20197), .B(n20200), .Z(n20198) );
  XOR U21410 ( .A(n20193), .B(n20161), .Z(n20194) );
  XOR U21411 ( .A(n20201), .B(n20202), .Z(n20161) );
  AND U21412 ( .A(n838), .B(n20203), .Z(n20201) );
  XOR U21413 ( .A(n20204), .B(n20202), .Z(n20203) );
  XNOR U21414 ( .A(n20205), .B(n20206), .Z(n20193) );
  NAND U21415 ( .A(n20207), .B(n20208), .Z(n20206) );
  XOR U21416 ( .A(n20209), .B(n20185), .Z(n20208) );
  XOR U21417 ( .A(n20199), .B(n20200), .Z(n20185) );
  XOR U21418 ( .A(n20210), .B(n20211), .Z(n20200) );
  ANDN U21419 ( .B(n20212), .A(n20213), .Z(n20210) );
  XOR U21420 ( .A(n20211), .B(n20214), .Z(n20212) );
  XOR U21421 ( .A(n20215), .B(n20216), .Z(n20199) );
  XOR U21422 ( .A(n20217), .B(n20218), .Z(n20216) );
  ANDN U21423 ( .B(n20219), .A(n20220), .Z(n20217) );
  XOR U21424 ( .A(n20221), .B(n20218), .Z(n20219) );
  IV U21425 ( .A(n20197), .Z(n20215) );
  XOR U21426 ( .A(n20222), .B(n20223), .Z(n20197) );
  ANDN U21427 ( .B(n20224), .A(n20225), .Z(n20222) );
  XOR U21428 ( .A(n20223), .B(n20226), .Z(n20224) );
  IV U21429 ( .A(n20205), .Z(n20209) );
  XOR U21430 ( .A(n20205), .B(n20187), .Z(n20207) );
  XOR U21431 ( .A(n20227), .B(n20228), .Z(n20187) );
  AND U21432 ( .A(n838), .B(n20229), .Z(n20227) );
  XOR U21433 ( .A(n20230), .B(n20228), .Z(n20229) );
  NANDN U21434 ( .A(n20189), .B(n20191), .Z(n20205) );
  XOR U21435 ( .A(n20231), .B(n20232), .Z(n20191) );
  AND U21436 ( .A(n838), .B(n20233), .Z(n20231) );
  XOR U21437 ( .A(n20232), .B(n20234), .Z(n20233) );
  XOR U21438 ( .A(n20235), .B(n20236), .Z(n838) );
  AND U21439 ( .A(n20237), .B(n20238), .Z(n20235) );
  XNOR U21440 ( .A(n20236), .B(n20202), .Z(n20238) );
  XNOR U21441 ( .A(n20239), .B(n20240), .Z(n20202) );
  ANDN U21442 ( .B(n20241), .A(n20242), .Z(n20239) );
  XOR U21443 ( .A(n20240), .B(n20243), .Z(n20241) );
  XOR U21444 ( .A(n20236), .B(n20204), .Z(n20237) );
  XOR U21445 ( .A(n20244), .B(n20245), .Z(n20204) );
  AND U21446 ( .A(n842), .B(n20246), .Z(n20244) );
  XOR U21447 ( .A(n20247), .B(n20245), .Z(n20246) );
  XNOR U21448 ( .A(n20248), .B(n20249), .Z(n20236) );
  NAND U21449 ( .A(n20250), .B(n20251), .Z(n20249) );
  XOR U21450 ( .A(n20252), .B(n20228), .Z(n20251) );
  XOR U21451 ( .A(n20242), .B(n20243), .Z(n20228) );
  XOR U21452 ( .A(n20253), .B(n20254), .Z(n20243) );
  ANDN U21453 ( .B(n20255), .A(n20256), .Z(n20253) );
  XOR U21454 ( .A(n20254), .B(n20257), .Z(n20255) );
  XOR U21455 ( .A(n20258), .B(n20259), .Z(n20242) );
  XOR U21456 ( .A(n20260), .B(n20261), .Z(n20259) );
  ANDN U21457 ( .B(n20262), .A(n20263), .Z(n20260) );
  XOR U21458 ( .A(n20264), .B(n20261), .Z(n20262) );
  IV U21459 ( .A(n20240), .Z(n20258) );
  XOR U21460 ( .A(n20265), .B(n20266), .Z(n20240) );
  ANDN U21461 ( .B(n20267), .A(n20268), .Z(n20265) );
  XOR U21462 ( .A(n20266), .B(n20269), .Z(n20267) );
  IV U21463 ( .A(n20248), .Z(n20252) );
  XOR U21464 ( .A(n20248), .B(n20230), .Z(n20250) );
  XOR U21465 ( .A(n20270), .B(n20271), .Z(n20230) );
  AND U21466 ( .A(n842), .B(n20272), .Z(n20270) );
  XOR U21467 ( .A(n20273), .B(n20271), .Z(n20272) );
  NANDN U21468 ( .A(n20232), .B(n20234), .Z(n20248) );
  XOR U21469 ( .A(n20274), .B(n20275), .Z(n20234) );
  AND U21470 ( .A(n842), .B(n20276), .Z(n20274) );
  XOR U21471 ( .A(n20275), .B(n20277), .Z(n20276) );
  XOR U21472 ( .A(n20278), .B(n20279), .Z(n842) );
  AND U21473 ( .A(n20280), .B(n20281), .Z(n20278) );
  XNOR U21474 ( .A(n20279), .B(n20245), .Z(n20281) );
  XNOR U21475 ( .A(n20282), .B(n20283), .Z(n20245) );
  ANDN U21476 ( .B(n20284), .A(n20285), .Z(n20282) );
  XOR U21477 ( .A(n20283), .B(n20286), .Z(n20284) );
  XOR U21478 ( .A(n20279), .B(n20247), .Z(n20280) );
  XOR U21479 ( .A(n20287), .B(n20288), .Z(n20247) );
  AND U21480 ( .A(n846), .B(n20289), .Z(n20287) );
  XOR U21481 ( .A(n20290), .B(n20288), .Z(n20289) );
  XNOR U21482 ( .A(n20291), .B(n20292), .Z(n20279) );
  NAND U21483 ( .A(n20293), .B(n20294), .Z(n20292) );
  XOR U21484 ( .A(n20295), .B(n20271), .Z(n20294) );
  XOR U21485 ( .A(n20285), .B(n20286), .Z(n20271) );
  XOR U21486 ( .A(n20296), .B(n20297), .Z(n20286) );
  ANDN U21487 ( .B(n20298), .A(n20299), .Z(n20296) );
  XOR U21488 ( .A(n20297), .B(n20300), .Z(n20298) );
  XOR U21489 ( .A(n20301), .B(n20302), .Z(n20285) );
  XOR U21490 ( .A(n20303), .B(n20304), .Z(n20302) );
  ANDN U21491 ( .B(n20305), .A(n20306), .Z(n20303) );
  XOR U21492 ( .A(n20307), .B(n20304), .Z(n20305) );
  IV U21493 ( .A(n20283), .Z(n20301) );
  XOR U21494 ( .A(n20308), .B(n20309), .Z(n20283) );
  ANDN U21495 ( .B(n20310), .A(n20311), .Z(n20308) );
  XOR U21496 ( .A(n20309), .B(n20312), .Z(n20310) );
  IV U21497 ( .A(n20291), .Z(n20295) );
  XOR U21498 ( .A(n20291), .B(n20273), .Z(n20293) );
  XOR U21499 ( .A(n20313), .B(n20314), .Z(n20273) );
  AND U21500 ( .A(n846), .B(n20315), .Z(n20313) );
  XOR U21501 ( .A(n20316), .B(n20314), .Z(n20315) );
  NANDN U21502 ( .A(n20275), .B(n20277), .Z(n20291) );
  XOR U21503 ( .A(n20317), .B(n20318), .Z(n20277) );
  AND U21504 ( .A(n846), .B(n20319), .Z(n20317) );
  XOR U21505 ( .A(n20318), .B(n20320), .Z(n20319) );
  XOR U21506 ( .A(n20321), .B(n20322), .Z(n846) );
  AND U21507 ( .A(n20323), .B(n20324), .Z(n20321) );
  XNOR U21508 ( .A(n20322), .B(n20288), .Z(n20324) );
  XNOR U21509 ( .A(n20325), .B(n20326), .Z(n20288) );
  ANDN U21510 ( .B(n20327), .A(n20328), .Z(n20325) );
  XOR U21511 ( .A(n20326), .B(n20329), .Z(n20327) );
  XOR U21512 ( .A(n20322), .B(n20290), .Z(n20323) );
  XOR U21513 ( .A(n20330), .B(n20331), .Z(n20290) );
  AND U21514 ( .A(n850), .B(n20332), .Z(n20330) );
  XOR U21515 ( .A(n20333), .B(n20331), .Z(n20332) );
  XNOR U21516 ( .A(n20334), .B(n20335), .Z(n20322) );
  NAND U21517 ( .A(n20336), .B(n20337), .Z(n20335) );
  XOR U21518 ( .A(n20338), .B(n20314), .Z(n20337) );
  XOR U21519 ( .A(n20328), .B(n20329), .Z(n20314) );
  XOR U21520 ( .A(n20339), .B(n20340), .Z(n20329) );
  ANDN U21521 ( .B(n20341), .A(n20342), .Z(n20339) );
  XOR U21522 ( .A(n20340), .B(n20343), .Z(n20341) );
  XOR U21523 ( .A(n20344), .B(n20345), .Z(n20328) );
  XOR U21524 ( .A(n20346), .B(n20347), .Z(n20345) );
  ANDN U21525 ( .B(n20348), .A(n20349), .Z(n20346) );
  XOR U21526 ( .A(n20350), .B(n20347), .Z(n20348) );
  IV U21527 ( .A(n20326), .Z(n20344) );
  XOR U21528 ( .A(n20351), .B(n20352), .Z(n20326) );
  ANDN U21529 ( .B(n20353), .A(n20354), .Z(n20351) );
  XOR U21530 ( .A(n20352), .B(n20355), .Z(n20353) );
  IV U21531 ( .A(n20334), .Z(n20338) );
  XOR U21532 ( .A(n20334), .B(n20316), .Z(n20336) );
  XOR U21533 ( .A(n20356), .B(n20357), .Z(n20316) );
  AND U21534 ( .A(n850), .B(n20358), .Z(n20356) );
  XOR U21535 ( .A(n20359), .B(n20357), .Z(n20358) );
  NANDN U21536 ( .A(n20318), .B(n20320), .Z(n20334) );
  XOR U21537 ( .A(n20360), .B(n20361), .Z(n20320) );
  AND U21538 ( .A(n850), .B(n20362), .Z(n20360) );
  XOR U21539 ( .A(n20361), .B(n20363), .Z(n20362) );
  XOR U21540 ( .A(n20364), .B(n20365), .Z(n850) );
  AND U21541 ( .A(n20366), .B(n20367), .Z(n20364) );
  XNOR U21542 ( .A(n20365), .B(n20331), .Z(n20367) );
  XNOR U21543 ( .A(n20368), .B(n20369), .Z(n20331) );
  ANDN U21544 ( .B(n20370), .A(n20371), .Z(n20368) );
  XOR U21545 ( .A(n20369), .B(n20372), .Z(n20370) );
  XOR U21546 ( .A(n20365), .B(n20333), .Z(n20366) );
  XOR U21547 ( .A(n20373), .B(n20374), .Z(n20333) );
  AND U21548 ( .A(n854), .B(n20375), .Z(n20373) );
  XOR U21549 ( .A(n20376), .B(n20374), .Z(n20375) );
  XNOR U21550 ( .A(n20377), .B(n20378), .Z(n20365) );
  NAND U21551 ( .A(n20379), .B(n20380), .Z(n20378) );
  XOR U21552 ( .A(n20381), .B(n20357), .Z(n20380) );
  XOR U21553 ( .A(n20371), .B(n20372), .Z(n20357) );
  XOR U21554 ( .A(n20382), .B(n20383), .Z(n20372) );
  ANDN U21555 ( .B(n20384), .A(n20385), .Z(n20382) );
  XOR U21556 ( .A(n20383), .B(n20386), .Z(n20384) );
  XOR U21557 ( .A(n20387), .B(n20388), .Z(n20371) );
  XOR U21558 ( .A(n20389), .B(n20390), .Z(n20388) );
  ANDN U21559 ( .B(n20391), .A(n20392), .Z(n20389) );
  XOR U21560 ( .A(n20393), .B(n20390), .Z(n20391) );
  IV U21561 ( .A(n20369), .Z(n20387) );
  XOR U21562 ( .A(n20394), .B(n20395), .Z(n20369) );
  ANDN U21563 ( .B(n20396), .A(n20397), .Z(n20394) );
  XOR U21564 ( .A(n20395), .B(n20398), .Z(n20396) );
  IV U21565 ( .A(n20377), .Z(n20381) );
  XOR U21566 ( .A(n20377), .B(n20359), .Z(n20379) );
  XOR U21567 ( .A(n20399), .B(n20400), .Z(n20359) );
  AND U21568 ( .A(n854), .B(n20401), .Z(n20399) );
  XOR U21569 ( .A(n20402), .B(n20400), .Z(n20401) );
  NANDN U21570 ( .A(n20361), .B(n20363), .Z(n20377) );
  XOR U21571 ( .A(n20403), .B(n20404), .Z(n20363) );
  AND U21572 ( .A(n854), .B(n20405), .Z(n20403) );
  XOR U21573 ( .A(n20404), .B(n20406), .Z(n20405) );
  XOR U21574 ( .A(n20407), .B(n20408), .Z(n854) );
  AND U21575 ( .A(n20409), .B(n20410), .Z(n20407) );
  XNOR U21576 ( .A(n20408), .B(n20374), .Z(n20410) );
  XNOR U21577 ( .A(n20411), .B(n20412), .Z(n20374) );
  ANDN U21578 ( .B(n20413), .A(n20414), .Z(n20411) );
  XOR U21579 ( .A(n20412), .B(n20415), .Z(n20413) );
  XOR U21580 ( .A(n20408), .B(n20376), .Z(n20409) );
  XOR U21581 ( .A(n20416), .B(n20417), .Z(n20376) );
  AND U21582 ( .A(n858), .B(n20418), .Z(n20416) );
  XOR U21583 ( .A(n20419), .B(n20417), .Z(n20418) );
  XNOR U21584 ( .A(n20420), .B(n20421), .Z(n20408) );
  NAND U21585 ( .A(n20422), .B(n20423), .Z(n20421) );
  XOR U21586 ( .A(n20424), .B(n20400), .Z(n20423) );
  XOR U21587 ( .A(n20414), .B(n20415), .Z(n20400) );
  XOR U21588 ( .A(n20425), .B(n20426), .Z(n20415) );
  ANDN U21589 ( .B(n20427), .A(n20428), .Z(n20425) );
  XOR U21590 ( .A(n20426), .B(n20429), .Z(n20427) );
  XOR U21591 ( .A(n20430), .B(n20431), .Z(n20414) );
  XOR U21592 ( .A(n20432), .B(n20433), .Z(n20431) );
  ANDN U21593 ( .B(n20434), .A(n20435), .Z(n20432) );
  XOR U21594 ( .A(n20436), .B(n20433), .Z(n20434) );
  IV U21595 ( .A(n20412), .Z(n20430) );
  XOR U21596 ( .A(n20437), .B(n20438), .Z(n20412) );
  ANDN U21597 ( .B(n20439), .A(n20440), .Z(n20437) );
  XOR U21598 ( .A(n20438), .B(n20441), .Z(n20439) );
  IV U21599 ( .A(n20420), .Z(n20424) );
  XOR U21600 ( .A(n20420), .B(n20402), .Z(n20422) );
  XOR U21601 ( .A(n20442), .B(n20443), .Z(n20402) );
  AND U21602 ( .A(n858), .B(n20444), .Z(n20442) );
  XOR U21603 ( .A(n20445), .B(n20443), .Z(n20444) );
  NANDN U21604 ( .A(n20404), .B(n20406), .Z(n20420) );
  XOR U21605 ( .A(n20446), .B(n20447), .Z(n20406) );
  AND U21606 ( .A(n858), .B(n20448), .Z(n20446) );
  XOR U21607 ( .A(n20447), .B(n20449), .Z(n20448) );
  XOR U21608 ( .A(n20450), .B(n20451), .Z(n858) );
  AND U21609 ( .A(n20452), .B(n20453), .Z(n20450) );
  XNOR U21610 ( .A(n20451), .B(n20417), .Z(n20453) );
  XNOR U21611 ( .A(n20454), .B(n20455), .Z(n20417) );
  ANDN U21612 ( .B(n20456), .A(n20457), .Z(n20454) );
  XOR U21613 ( .A(n20455), .B(n20458), .Z(n20456) );
  XOR U21614 ( .A(n20451), .B(n20419), .Z(n20452) );
  XOR U21615 ( .A(n20459), .B(n20460), .Z(n20419) );
  AND U21616 ( .A(n862), .B(n20461), .Z(n20459) );
  XOR U21617 ( .A(n20462), .B(n20460), .Z(n20461) );
  XNOR U21618 ( .A(n20463), .B(n20464), .Z(n20451) );
  NAND U21619 ( .A(n20465), .B(n20466), .Z(n20464) );
  XOR U21620 ( .A(n20467), .B(n20443), .Z(n20466) );
  XOR U21621 ( .A(n20457), .B(n20458), .Z(n20443) );
  XOR U21622 ( .A(n20468), .B(n20469), .Z(n20458) );
  ANDN U21623 ( .B(n20470), .A(n20471), .Z(n20468) );
  XOR U21624 ( .A(n20469), .B(n20472), .Z(n20470) );
  XOR U21625 ( .A(n20473), .B(n20474), .Z(n20457) );
  XOR U21626 ( .A(n20475), .B(n20476), .Z(n20474) );
  ANDN U21627 ( .B(n20477), .A(n20478), .Z(n20475) );
  XOR U21628 ( .A(n20479), .B(n20476), .Z(n20477) );
  IV U21629 ( .A(n20455), .Z(n20473) );
  XOR U21630 ( .A(n20480), .B(n20481), .Z(n20455) );
  ANDN U21631 ( .B(n20482), .A(n20483), .Z(n20480) );
  XOR U21632 ( .A(n20481), .B(n20484), .Z(n20482) );
  IV U21633 ( .A(n20463), .Z(n20467) );
  XOR U21634 ( .A(n20463), .B(n20445), .Z(n20465) );
  XOR U21635 ( .A(n20485), .B(n20486), .Z(n20445) );
  AND U21636 ( .A(n862), .B(n20487), .Z(n20485) );
  XOR U21637 ( .A(n20488), .B(n20486), .Z(n20487) );
  NANDN U21638 ( .A(n20447), .B(n20449), .Z(n20463) );
  XOR U21639 ( .A(n20489), .B(n20490), .Z(n20449) );
  AND U21640 ( .A(n862), .B(n20491), .Z(n20489) );
  XOR U21641 ( .A(n20490), .B(n20492), .Z(n20491) );
  XOR U21642 ( .A(n20493), .B(n20494), .Z(n862) );
  AND U21643 ( .A(n20495), .B(n20496), .Z(n20493) );
  XNOR U21644 ( .A(n20494), .B(n20460), .Z(n20496) );
  XNOR U21645 ( .A(n20497), .B(n20498), .Z(n20460) );
  ANDN U21646 ( .B(n20499), .A(n20500), .Z(n20497) );
  XOR U21647 ( .A(n20498), .B(n20501), .Z(n20499) );
  XOR U21648 ( .A(n20494), .B(n20462), .Z(n20495) );
  XOR U21649 ( .A(n20502), .B(n20503), .Z(n20462) );
  AND U21650 ( .A(n866), .B(n20504), .Z(n20502) );
  XOR U21651 ( .A(n20505), .B(n20503), .Z(n20504) );
  XNOR U21652 ( .A(n20506), .B(n20507), .Z(n20494) );
  NAND U21653 ( .A(n20508), .B(n20509), .Z(n20507) );
  XOR U21654 ( .A(n20510), .B(n20486), .Z(n20509) );
  XOR U21655 ( .A(n20500), .B(n20501), .Z(n20486) );
  XOR U21656 ( .A(n20511), .B(n20512), .Z(n20501) );
  ANDN U21657 ( .B(n20513), .A(n20514), .Z(n20511) );
  XOR U21658 ( .A(n20512), .B(n20515), .Z(n20513) );
  XOR U21659 ( .A(n20516), .B(n20517), .Z(n20500) );
  XOR U21660 ( .A(n20518), .B(n20519), .Z(n20517) );
  ANDN U21661 ( .B(n20520), .A(n20521), .Z(n20518) );
  XOR U21662 ( .A(n20522), .B(n20519), .Z(n20520) );
  IV U21663 ( .A(n20498), .Z(n20516) );
  XOR U21664 ( .A(n20523), .B(n20524), .Z(n20498) );
  ANDN U21665 ( .B(n20525), .A(n20526), .Z(n20523) );
  XOR U21666 ( .A(n20524), .B(n20527), .Z(n20525) );
  IV U21667 ( .A(n20506), .Z(n20510) );
  XOR U21668 ( .A(n20506), .B(n20488), .Z(n20508) );
  XOR U21669 ( .A(n20528), .B(n20529), .Z(n20488) );
  AND U21670 ( .A(n866), .B(n20530), .Z(n20528) );
  XOR U21671 ( .A(n20531), .B(n20529), .Z(n20530) );
  NANDN U21672 ( .A(n20490), .B(n20492), .Z(n20506) );
  XOR U21673 ( .A(n20532), .B(n20533), .Z(n20492) );
  AND U21674 ( .A(n866), .B(n20534), .Z(n20532) );
  XOR U21675 ( .A(n20533), .B(n20535), .Z(n20534) );
  XOR U21676 ( .A(n20536), .B(n20537), .Z(n866) );
  AND U21677 ( .A(n20538), .B(n20539), .Z(n20536) );
  XNOR U21678 ( .A(n20537), .B(n20503), .Z(n20539) );
  XNOR U21679 ( .A(n20540), .B(n20541), .Z(n20503) );
  ANDN U21680 ( .B(n20542), .A(n20543), .Z(n20540) );
  XOR U21681 ( .A(n20541), .B(n20544), .Z(n20542) );
  XOR U21682 ( .A(n20537), .B(n20505), .Z(n20538) );
  XOR U21683 ( .A(n20545), .B(n20546), .Z(n20505) );
  AND U21684 ( .A(n870), .B(n20547), .Z(n20545) );
  XOR U21685 ( .A(n20548), .B(n20546), .Z(n20547) );
  XNOR U21686 ( .A(n20549), .B(n20550), .Z(n20537) );
  NAND U21687 ( .A(n20551), .B(n20552), .Z(n20550) );
  XOR U21688 ( .A(n20553), .B(n20529), .Z(n20552) );
  XOR U21689 ( .A(n20543), .B(n20544), .Z(n20529) );
  XOR U21690 ( .A(n20554), .B(n20555), .Z(n20544) );
  ANDN U21691 ( .B(n20556), .A(n20557), .Z(n20554) );
  XOR U21692 ( .A(n20555), .B(n20558), .Z(n20556) );
  XOR U21693 ( .A(n20559), .B(n20560), .Z(n20543) );
  XOR U21694 ( .A(n20561), .B(n20562), .Z(n20560) );
  ANDN U21695 ( .B(n20563), .A(n20564), .Z(n20561) );
  XOR U21696 ( .A(n20565), .B(n20562), .Z(n20563) );
  IV U21697 ( .A(n20541), .Z(n20559) );
  XOR U21698 ( .A(n20566), .B(n20567), .Z(n20541) );
  ANDN U21699 ( .B(n20568), .A(n20569), .Z(n20566) );
  XOR U21700 ( .A(n20567), .B(n20570), .Z(n20568) );
  IV U21701 ( .A(n20549), .Z(n20553) );
  XOR U21702 ( .A(n20549), .B(n20531), .Z(n20551) );
  XOR U21703 ( .A(n20571), .B(n20572), .Z(n20531) );
  AND U21704 ( .A(n870), .B(n20573), .Z(n20571) );
  XOR U21705 ( .A(n20574), .B(n20572), .Z(n20573) );
  NANDN U21706 ( .A(n20533), .B(n20535), .Z(n20549) );
  XOR U21707 ( .A(n20575), .B(n20576), .Z(n20535) );
  AND U21708 ( .A(n870), .B(n20577), .Z(n20575) );
  XOR U21709 ( .A(n20576), .B(n20578), .Z(n20577) );
  XOR U21710 ( .A(n20579), .B(n20580), .Z(n870) );
  AND U21711 ( .A(n20581), .B(n20582), .Z(n20579) );
  XNOR U21712 ( .A(n20580), .B(n20546), .Z(n20582) );
  XNOR U21713 ( .A(n20583), .B(n20584), .Z(n20546) );
  ANDN U21714 ( .B(n20585), .A(n20586), .Z(n20583) );
  XOR U21715 ( .A(n20584), .B(n20587), .Z(n20585) );
  XOR U21716 ( .A(n20580), .B(n20548), .Z(n20581) );
  XOR U21717 ( .A(n20588), .B(n20589), .Z(n20548) );
  AND U21718 ( .A(n874), .B(n20590), .Z(n20588) );
  XOR U21719 ( .A(n20591), .B(n20589), .Z(n20590) );
  XNOR U21720 ( .A(n20592), .B(n20593), .Z(n20580) );
  NAND U21721 ( .A(n20594), .B(n20595), .Z(n20593) );
  XOR U21722 ( .A(n20596), .B(n20572), .Z(n20595) );
  XOR U21723 ( .A(n20586), .B(n20587), .Z(n20572) );
  XOR U21724 ( .A(n20597), .B(n20598), .Z(n20587) );
  ANDN U21725 ( .B(n20599), .A(n20600), .Z(n20597) );
  XOR U21726 ( .A(n20598), .B(n20601), .Z(n20599) );
  XOR U21727 ( .A(n20602), .B(n20603), .Z(n20586) );
  XOR U21728 ( .A(n20604), .B(n20605), .Z(n20603) );
  ANDN U21729 ( .B(n20606), .A(n20607), .Z(n20604) );
  XOR U21730 ( .A(n20608), .B(n20605), .Z(n20606) );
  IV U21731 ( .A(n20584), .Z(n20602) );
  XOR U21732 ( .A(n20609), .B(n20610), .Z(n20584) );
  ANDN U21733 ( .B(n20611), .A(n20612), .Z(n20609) );
  XOR U21734 ( .A(n20610), .B(n20613), .Z(n20611) );
  IV U21735 ( .A(n20592), .Z(n20596) );
  XOR U21736 ( .A(n20592), .B(n20574), .Z(n20594) );
  XOR U21737 ( .A(n20614), .B(n20615), .Z(n20574) );
  AND U21738 ( .A(n874), .B(n20616), .Z(n20614) );
  XOR U21739 ( .A(n20617), .B(n20615), .Z(n20616) );
  NANDN U21740 ( .A(n20576), .B(n20578), .Z(n20592) );
  XOR U21741 ( .A(n20618), .B(n20619), .Z(n20578) );
  AND U21742 ( .A(n874), .B(n20620), .Z(n20618) );
  XOR U21743 ( .A(n20619), .B(n20621), .Z(n20620) );
  XOR U21744 ( .A(n20622), .B(n20623), .Z(n874) );
  AND U21745 ( .A(n20624), .B(n20625), .Z(n20622) );
  XNOR U21746 ( .A(n20623), .B(n20589), .Z(n20625) );
  XNOR U21747 ( .A(n20626), .B(n20627), .Z(n20589) );
  ANDN U21748 ( .B(n20628), .A(n20629), .Z(n20626) );
  XOR U21749 ( .A(n20627), .B(n20630), .Z(n20628) );
  XOR U21750 ( .A(n20623), .B(n20591), .Z(n20624) );
  XOR U21751 ( .A(n20631), .B(n20632), .Z(n20591) );
  AND U21752 ( .A(n878), .B(n20633), .Z(n20631) );
  XOR U21753 ( .A(n20634), .B(n20632), .Z(n20633) );
  XNOR U21754 ( .A(n20635), .B(n20636), .Z(n20623) );
  NAND U21755 ( .A(n20637), .B(n20638), .Z(n20636) );
  XOR U21756 ( .A(n20639), .B(n20615), .Z(n20638) );
  XOR U21757 ( .A(n20629), .B(n20630), .Z(n20615) );
  XOR U21758 ( .A(n20640), .B(n20641), .Z(n20630) );
  ANDN U21759 ( .B(n20642), .A(n20643), .Z(n20640) );
  XOR U21760 ( .A(n20641), .B(n20644), .Z(n20642) );
  XOR U21761 ( .A(n20645), .B(n20646), .Z(n20629) );
  XOR U21762 ( .A(n20647), .B(n20648), .Z(n20646) );
  ANDN U21763 ( .B(n20649), .A(n20650), .Z(n20647) );
  XOR U21764 ( .A(n20651), .B(n20648), .Z(n20649) );
  IV U21765 ( .A(n20627), .Z(n20645) );
  XOR U21766 ( .A(n20652), .B(n20653), .Z(n20627) );
  ANDN U21767 ( .B(n20654), .A(n20655), .Z(n20652) );
  XOR U21768 ( .A(n20653), .B(n20656), .Z(n20654) );
  IV U21769 ( .A(n20635), .Z(n20639) );
  XOR U21770 ( .A(n20635), .B(n20617), .Z(n20637) );
  XOR U21771 ( .A(n20657), .B(n20658), .Z(n20617) );
  AND U21772 ( .A(n878), .B(n20659), .Z(n20657) );
  XOR U21773 ( .A(n20660), .B(n20658), .Z(n20659) );
  NANDN U21774 ( .A(n20619), .B(n20621), .Z(n20635) );
  XOR U21775 ( .A(n20661), .B(n20662), .Z(n20621) );
  AND U21776 ( .A(n878), .B(n20663), .Z(n20661) );
  XOR U21777 ( .A(n20662), .B(n20664), .Z(n20663) );
  XOR U21778 ( .A(n20665), .B(n20666), .Z(n878) );
  AND U21779 ( .A(n20667), .B(n20668), .Z(n20665) );
  XNOR U21780 ( .A(n20666), .B(n20632), .Z(n20668) );
  XNOR U21781 ( .A(n20669), .B(n20670), .Z(n20632) );
  ANDN U21782 ( .B(n20671), .A(n20672), .Z(n20669) );
  XOR U21783 ( .A(n20670), .B(n20673), .Z(n20671) );
  XOR U21784 ( .A(n20666), .B(n20634), .Z(n20667) );
  XOR U21785 ( .A(n20674), .B(n20675), .Z(n20634) );
  AND U21786 ( .A(n882), .B(n20676), .Z(n20674) );
  XOR U21787 ( .A(n20677), .B(n20675), .Z(n20676) );
  XNOR U21788 ( .A(n20678), .B(n20679), .Z(n20666) );
  NAND U21789 ( .A(n20680), .B(n20681), .Z(n20679) );
  XOR U21790 ( .A(n20682), .B(n20658), .Z(n20681) );
  XOR U21791 ( .A(n20672), .B(n20673), .Z(n20658) );
  XOR U21792 ( .A(n20683), .B(n20684), .Z(n20673) );
  ANDN U21793 ( .B(n20685), .A(n20686), .Z(n20683) );
  XOR U21794 ( .A(n20684), .B(n20687), .Z(n20685) );
  XOR U21795 ( .A(n20688), .B(n20689), .Z(n20672) );
  XOR U21796 ( .A(n20690), .B(n20691), .Z(n20689) );
  ANDN U21797 ( .B(n20692), .A(n20693), .Z(n20690) );
  XOR U21798 ( .A(n20694), .B(n20691), .Z(n20692) );
  IV U21799 ( .A(n20670), .Z(n20688) );
  XOR U21800 ( .A(n20695), .B(n20696), .Z(n20670) );
  ANDN U21801 ( .B(n20697), .A(n20698), .Z(n20695) );
  XOR U21802 ( .A(n20696), .B(n20699), .Z(n20697) );
  IV U21803 ( .A(n20678), .Z(n20682) );
  XOR U21804 ( .A(n20678), .B(n20660), .Z(n20680) );
  XOR U21805 ( .A(n20700), .B(n20701), .Z(n20660) );
  AND U21806 ( .A(n882), .B(n20702), .Z(n20700) );
  XOR U21807 ( .A(n20703), .B(n20701), .Z(n20702) );
  NANDN U21808 ( .A(n20662), .B(n20664), .Z(n20678) );
  XOR U21809 ( .A(n20704), .B(n20705), .Z(n20664) );
  AND U21810 ( .A(n882), .B(n20706), .Z(n20704) );
  XOR U21811 ( .A(n20705), .B(n20707), .Z(n20706) );
  XOR U21812 ( .A(n20708), .B(n20709), .Z(n882) );
  AND U21813 ( .A(n20710), .B(n20711), .Z(n20708) );
  XNOR U21814 ( .A(n20709), .B(n20675), .Z(n20711) );
  XNOR U21815 ( .A(n20712), .B(n20713), .Z(n20675) );
  ANDN U21816 ( .B(n20714), .A(n20715), .Z(n20712) );
  XOR U21817 ( .A(n20713), .B(n20716), .Z(n20714) );
  XOR U21818 ( .A(n20709), .B(n20677), .Z(n20710) );
  XOR U21819 ( .A(n20717), .B(n20718), .Z(n20677) );
  AND U21820 ( .A(n886), .B(n20719), .Z(n20717) );
  XOR U21821 ( .A(n20720), .B(n20718), .Z(n20719) );
  XNOR U21822 ( .A(n20721), .B(n20722), .Z(n20709) );
  NAND U21823 ( .A(n20723), .B(n20724), .Z(n20722) );
  XOR U21824 ( .A(n20725), .B(n20701), .Z(n20724) );
  XOR U21825 ( .A(n20715), .B(n20716), .Z(n20701) );
  XOR U21826 ( .A(n20726), .B(n20727), .Z(n20716) );
  ANDN U21827 ( .B(n20728), .A(n20729), .Z(n20726) );
  XOR U21828 ( .A(n20727), .B(n20730), .Z(n20728) );
  XOR U21829 ( .A(n20731), .B(n20732), .Z(n20715) );
  XOR U21830 ( .A(n20733), .B(n20734), .Z(n20732) );
  ANDN U21831 ( .B(n20735), .A(n20736), .Z(n20733) );
  XOR U21832 ( .A(n20737), .B(n20734), .Z(n20735) );
  IV U21833 ( .A(n20713), .Z(n20731) );
  XOR U21834 ( .A(n20738), .B(n20739), .Z(n20713) );
  ANDN U21835 ( .B(n20740), .A(n20741), .Z(n20738) );
  XOR U21836 ( .A(n20739), .B(n20742), .Z(n20740) );
  IV U21837 ( .A(n20721), .Z(n20725) );
  XOR U21838 ( .A(n20721), .B(n20703), .Z(n20723) );
  XOR U21839 ( .A(n20743), .B(n20744), .Z(n20703) );
  AND U21840 ( .A(n886), .B(n20745), .Z(n20743) );
  XOR U21841 ( .A(n20746), .B(n20744), .Z(n20745) );
  NANDN U21842 ( .A(n20705), .B(n20707), .Z(n20721) );
  XOR U21843 ( .A(n20747), .B(n20748), .Z(n20707) );
  AND U21844 ( .A(n886), .B(n20749), .Z(n20747) );
  XOR U21845 ( .A(n20748), .B(n20750), .Z(n20749) );
  XOR U21846 ( .A(n20751), .B(n20752), .Z(n886) );
  AND U21847 ( .A(n20753), .B(n20754), .Z(n20751) );
  XNOR U21848 ( .A(n20752), .B(n20718), .Z(n20754) );
  XNOR U21849 ( .A(n20755), .B(n20756), .Z(n20718) );
  ANDN U21850 ( .B(n20757), .A(n20758), .Z(n20755) );
  XOR U21851 ( .A(n20756), .B(n20759), .Z(n20757) );
  XOR U21852 ( .A(n20752), .B(n20720), .Z(n20753) );
  XOR U21853 ( .A(n20760), .B(n20761), .Z(n20720) );
  AND U21854 ( .A(n890), .B(n20762), .Z(n20760) );
  XOR U21855 ( .A(n20763), .B(n20761), .Z(n20762) );
  XNOR U21856 ( .A(n20764), .B(n20765), .Z(n20752) );
  NAND U21857 ( .A(n20766), .B(n20767), .Z(n20765) );
  XOR U21858 ( .A(n20768), .B(n20744), .Z(n20767) );
  XOR U21859 ( .A(n20758), .B(n20759), .Z(n20744) );
  XOR U21860 ( .A(n20769), .B(n20770), .Z(n20759) );
  ANDN U21861 ( .B(n20771), .A(n20772), .Z(n20769) );
  XOR U21862 ( .A(n20770), .B(n20773), .Z(n20771) );
  XOR U21863 ( .A(n20774), .B(n20775), .Z(n20758) );
  XOR U21864 ( .A(n20776), .B(n20777), .Z(n20775) );
  ANDN U21865 ( .B(n20778), .A(n20779), .Z(n20776) );
  XOR U21866 ( .A(n20780), .B(n20777), .Z(n20778) );
  IV U21867 ( .A(n20756), .Z(n20774) );
  XOR U21868 ( .A(n20781), .B(n20782), .Z(n20756) );
  ANDN U21869 ( .B(n20783), .A(n20784), .Z(n20781) );
  XOR U21870 ( .A(n20782), .B(n20785), .Z(n20783) );
  IV U21871 ( .A(n20764), .Z(n20768) );
  XOR U21872 ( .A(n20764), .B(n20746), .Z(n20766) );
  XOR U21873 ( .A(n20786), .B(n20787), .Z(n20746) );
  AND U21874 ( .A(n890), .B(n20788), .Z(n20786) );
  XOR U21875 ( .A(n20789), .B(n20787), .Z(n20788) );
  NANDN U21876 ( .A(n20748), .B(n20750), .Z(n20764) );
  XOR U21877 ( .A(n20790), .B(n20791), .Z(n20750) );
  AND U21878 ( .A(n890), .B(n20792), .Z(n20790) );
  XOR U21879 ( .A(n20791), .B(n20793), .Z(n20792) );
  XOR U21880 ( .A(n20794), .B(n20795), .Z(n890) );
  AND U21881 ( .A(n20796), .B(n20797), .Z(n20794) );
  XNOR U21882 ( .A(n20795), .B(n20761), .Z(n20797) );
  XNOR U21883 ( .A(n20798), .B(n20799), .Z(n20761) );
  ANDN U21884 ( .B(n20800), .A(n20801), .Z(n20798) );
  XOR U21885 ( .A(n20799), .B(n20802), .Z(n20800) );
  XOR U21886 ( .A(n20795), .B(n20763), .Z(n20796) );
  XOR U21887 ( .A(n20803), .B(n20804), .Z(n20763) );
  AND U21888 ( .A(n894), .B(n20805), .Z(n20803) );
  XOR U21889 ( .A(n20806), .B(n20804), .Z(n20805) );
  XNOR U21890 ( .A(n20807), .B(n20808), .Z(n20795) );
  NAND U21891 ( .A(n20809), .B(n20810), .Z(n20808) );
  XOR U21892 ( .A(n20811), .B(n20787), .Z(n20810) );
  XOR U21893 ( .A(n20801), .B(n20802), .Z(n20787) );
  XOR U21894 ( .A(n20812), .B(n20813), .Z(n20802) );
  ANDN U21895 ( .B(n20814), .A(n20815), .Z(n20812) );
  XOR U21896 ( .A(n20813), .B(n20816), .Z(n20814) );
  XOR U21897 ( .A(n20817), .B(n20818), .Z(n20801) );
  XOR U21898 ( .A(n20819), .B(n20820), .Z(n20818) );
  ANDN U21899 ( .B(n20821), .A(n20822), .Z(n20819) );
  XOR U21900 ( .A(n20823), .B(n20820), .Z(n20821) );
  IV U21901 ( .A(n20799), .Z(n20817) );
  XOR U21902 ( .A(n20824), .B(n20825), .Z(n20799) );
  ANDN U21903 ( .B(n20826), .A(n20827), .Z(n20824) );
  XOR U21904 ( .A(n20825), .B(n20828), .Z(n20826) );
  IV U21905 ( .A(n20807), .Z(n20811) );
  XOR U21906 ( .A(n20807), .B(n20789), .Z(n20809) );
  XOR U21907 ( .A(n20829), .B(n20830), .Z(n20789) );
  AND U21908 ( .A(n894), .B(n20831), .Z(n20829) );
  XOR U21909 ( .A(n20832), .B(n20830), .Z(n20831) );
  NANDN U21910 ( .A(n20791), .B(n20793), .Z(n20807) );
  XOR U21911 ( .A(n20833), .B(n20834), .Z(n20793) );
  AND U21912 ( .A(n894), .B(n20835), .Z(n20833) );
  XOR U21913 ( .A(n20834), .B(n20836), .Z(n20835) );
  XOR U21914 ( .A(n20837), .B(n20838), .Z(n894) );
  AND U21915 ( .A(n20839), .B(n20840), .Z(n20837) );
  XNOR U21916 ( .A(n20838), .B(n20804), .Z(n20840) );
  XNOR U21917 ( .A(n20841), .B(n20842), .Z(n20804) );
  ANDN U21918 ( .B(n20843), .A(n20844), .Z(n20841) );
  XOR U21919 ( .A(n20842), .B(n20845), .Z(n20843) );
  XOR U21920 ( .A(n20838), .B(n20806), .Z(n20839) );
  XOR U21921 ( .A(n20846), .B(n20847), .Z(n20806) );
  AND U21922 ( .A(n898), .B(n20848), .Z(n20846) );
  XOR U21923 ( .A(n20849), .B(n20847), .Z(n20848) );
  XNOR U21924 ( .A(n20850), .B(n20851), .Z(n20838) );
  NAND U21925 ( .A(n20852), .B(n20853), .Z(n20851) );
  XOR U21926 ( .A(n20854), .B(n20830), .Z(n20853) );
  XOR U21927 ( .A(n20844), .B(n20845), .Z(n20830) );
  XOR U21928 ( .A(n20855), .B(n20856), .Z(n20845) );
  ANDN U21929 ( .B(n20857), .A(n20858), .Z(n20855) );
  XOR U21930 ( .A(n20856), .B(n20859), .Z(n20857) );
  XOR U21931 ( .A(n20860), .B(n20861), .Z(n20844) );
  XOR U21932 ( .A(n20862), .B(n20863), .Z(n20861) );
  ANDN U21933 ( .B(n20864), .A(n20865), .Z(n20862) );
  XOR U21934 ( .A(n20866), .B(n20863), .Z(n20864) );
  IV U21935 ( .A(n20842), .Z(n20860) );
  XOR U21936 ( .A(n20867), .B(n20868), .Z(n20842) );
  ANDN U21937 ( .B(n20869), .A(n20870), .Z(n20867) );
  XOR U21938 ( .A(n20868), .B(n20871), .Z(n20869) );
  IV U21939 ( .A(n20850), .Z(n20854) );
  XOR U21940 ( .A(n20850), .B(n20832), .Z(n20852) );
  XOR U21941 ( .A(n20872), .B(n20873), .Z(n20832) );
  AND U21942 ( .A(n898), .B(n20874), .Z(n20872) );
  XOR U21943 ( .A(n20875), .B(n20873), .Z(n20874) );
  NANDN U21944 ( .A(n20834), .B(n20836), .Z(n20850) );
  XOR U21945 ( .A(n20876), .B(n20877), .Z(n20836) );
  AND U21946 ( .A(n898), .B(n20878), .Z(n20876) );
  XOR U21947 ( .A(n20877), .B(n20879), .Z(n20878) );
  XOR U21948 ( .A(n20880), .B(n20881), .Z(n898) );
  AND U21949 ( .A(n20882), .B(n20883), .Z(n20880) );
  XNOR U21950 ( .A(n20881), .B(n20847), .Z(n20883) );
  XNOR U21951 ( .A(n20884), .B(n20885), .Z(n20847) );
  ANDN U21952 ( .B(n20886), .A(n20887), .Z(n20884) );
  XOR U21953 ( .A(n20885), .B(n20888), .Z(n20886) );
  XOR U21954 ( .A(n20881), .B(n20849), .Z(n20882) );
  XOR U21955 ( .A(n20889), .B(n20890), .Z(n20849) );
  AND U21956 ( .A(n902), .B(n20891), .Z(n20889) );
  XOR U21957 ( .A(n20892), .B(n20890), .Z(n20891) );
  XNOR U21958 ( .A(n20893), .B(n20894), .Z(n20881) );
  NAND U21959 ( .A(n20895), .B(n20896), .Z(n20894) );
  XOR U21960 ( .A(n20897), .B(n20873), .Z(n20896) );
  XOR U21961 ( .A(n20887), .B(n20888), .Z(n20873) );
  XOR U21962 ( .A(n20898), .B(n20899), .Z(n20888) );
  ANDN U21963 ( .B(n20900), .A(n20901), .Z(n20898) );
  XOR U21964 ( .A(n20899), .B(n20902), .Z(n20900) );
  XOR U21965 ( .A(n20903), .B(n20904), .Z(n20887) );
  XOR U21966 ( .A(n20905), .B(n20906), .Z(n20904) );
  ANDN U21967 ( .B(n20907), .A(n20908), .Z(n20905) );
  XOR U21968 ( .A(n20909), .B(n20906), .Z(n20907) );
  IV U21969 ( .A(n20885), .Z(n20903) );
  XOR U21970 ( .A(n20910), .B(n20911), .Z(n20885) );
  ANDN U21971 ( .B(n20912), .A(n20913), .Z(n20910) );
  XOR U21972 ( .A(n20911), .B(n20914), .Z(n20912) );
  IV U21973 ( .A(n20893), .Z(n20897) );
  XOR U21974 ( .A(n20893), .B(n20875), .Z(n20895) );
  XOR U21975 ( .A(n20915), .B(n20916), .Z(n20875) );
  AND U21976 ( .A(n902), .B(n20917), .Z(n20915) );
  XOR U21977 ( .A(n20918), .B(n20916), .Z(n20917) );
  NANDN U21978 ( .A(n20877), .B(n20879), .Z(n20893) );
  XOR U21979 ( .A(n20919), .B(n20920), .Z(n20879) );
  AND U21980 ( .A(n902), .B(n20921), .Z(n20919) );
  XOR U21981 ( .A(n20920), .B(n20922), .Z(n20921) );
  XOR U21982 ( .A(n20923), .B(n20924), .Z(n902) );
  AND U21983 ( .A(n20925), .B(n20926), .Z(n20923) );
  XNOR U21984 ( .A(n20924), .B(n20890), .Z(n20926) );
  XNOR U21985 ( .A(n20927), .B(n20928), .Z(n20890) );
  ANDN U21986 ( .B(n20929), .A(n20930), .Z(n20927) );
  XOR U21987 ( .A(n20928), .B(n20931), .Z(n20929) );
  XOR U21988 ( .A(n20924), .B(n20892), .Z(n20925) );
  XOR U21989 ( .A(n20932), .B(n20933), .Z(n20892) );
  AND U21990 ( .A(n906), .B(n20934), .Z(n20932) );
  XOR U21991 ( .A(n20935), .B(n20933), .Z(n20934) );
  XNOR U21992 ( .A(n20936), .B(n20937), .Z(n20924) );
  NAND U21993 ( .A(n20938), .B(n20939), .Z(n20937) );
  XOR U21994 ( .A(n20940), .B(n20916), .Z(n20939) );
  XOR U21995 ( .A(n20930), .B(n20931), .Z(n20916) );
  XOR U21996 ( .A(n20941), .B(n20942), .Z(n20931) );
  ANDN U21997 ( .B(n20943), .A(n20944), .Z(n20941) );
  XOR U21998 ( .A(n20942), .B(n20945), .Z(n20943) );
  XOR U21999 ( .A(n20946), .B(n20947), .Z(n20930) );
  XOR U22000 ( .A(n20948), .B(n20949), .Z(n20947) );
  ANDN U22001 ( .B(n20950), .A(n20951), .Z(n20948) );
  XOR U22002 ( .A(n20952), .B(n20949), .Z(n20950) );
  IV U22003 ( .A(n20928), .Z(n20946) );
  XOR U22004 ( .A(n20953), .B(n20954), .Z(n20928) );
  ANDN U22005 ( .B(n20955), .A(n20956), .Z(n20953) );
  XOR U22006 ( .A(n20954), .B(n20957), .Z(n20955) );
  IV U22007 ( .A(n20936), .Z(n20940) );
  XOR U22008 ( .A(n20936), .B(n20918), .Z(n20938) );
  XOR U22009 ( .A(n20958), .B(n20959), .Z(n20918) );
  AND U22010 ( .A(n906), .B(n20960), .Z(n20958) );
  XOR U22011 ( .A(n20961), .B(n20959), .Z(n20960) );
  NANDN U22012 ( .A(n20920), .B(n20922), .Z(n20936) );
  XOR U22013 ( .A(n20962), .B(n20963), .Z(n20922) );
  AND U22014 ( .A(n906), .B(n20964), .Z(n20962) );
  XOR U22015 ( .A(n20963), .B(n20965), .Z(n20964) );
  XOR U22016 ( .A(n20966), .B(n20967), .Z(n906) );
  AND U22017 ( .A(n20968), .B(n20969), .Z(n20966) );
  XNOR U22018 ( .A(n20967), .B(n20933), .Z(n20969) );
  XNOR U22019 ( .A(n20970), .B(n20971), .Z(n20933) );
  ANDN U22020 ( .B(n20972), .A(n20973), .Z(n20970) );
  XOR U22021 ( .A(n20971), .B(n20974), .Z(n20972) );
  XOR U22022 ( .A(n20967), .B(n20935), .Z(n20968) );
  XOR U22023 ( .A(n20975), .B(n20976), .Z(n20935) );
  AND U22024 ( .A(n910), .B(n20977), .Z(n20975) );
  XOR U22025 ( .A(n20978), .B(n20976), .Z(n20977) );
  XNOR U22026 ( .A(n20979), .B(n20980), .Z(n20967) );
  NAND U22027 ( .A(n20981), .B(n20982), .Z(n20980) );
  XOR U22028 ( .A(n20983), .B(n20959), .Z(n20982) );
  XOR U22029 ( .A(n20973), .B(n20974), .Z(n20959) );
  XOR U22030 ( .A(n20984), .B(n20985), .Z(n20974) );
  ANDN U22031 ( .B(n20986), .A(n20987), .Z(n20984) );
  XOR U22032 ( .A(n20985), .B(n20988), .Z(n20986) );
  XOR U22033 ( .A(n20989), .B(n20990), .Z(n20973) );
  XOR U22034 ( .A(n20991), .B(n20992), .Z(n20990) );
  ANDN U22035 ( .B(n20993), .A(n20994), .Z(n20991) );
  XOR U22036 ( .A(n20995), .B(n20992), .Z(n20993) );
  IV U22037 ( .A(n20971), .Z(n20989) );
  XOR U22038 ( .A(n20996), .B(n20997), .Z(n20971) );
  ANDN U22039 ( .B(n20998), .A(n20999), .Z(n20996) );
  XOR U22040 ( .A(n20997), .B(n21000), .Z(n20998) );
  IV U22041 ( .A(n20979), .Z(n20983) );
  XOR U22042 ( .A(n20979), .B(n20961), .Z(n20981) );
  XOR U22043 ( .A(n21001), .B(n21002), .Z(n20961) );
  AND U22044 ( .A(n910), .B(n21003), .Z(n21001) );
  XOR U22045 ( .A(n21004), .B(n21002), .Z(n21003) );
  NANDN U22046 ( .A(n20963), .B(n20965), .Z(n20979) );
  XOR U22047 ( .A(n21005), .B(n21006), .Z(n20965) );
  AND U22048 ( .A(n910), .B(n21007), .Z(n21005) );
  XOR U22049 ( .A(n21006), .B(n21008), .Z(n21007) );
  XOR U22050 ( .A(n21009), .B(n21010), .Z(n910) );
  AND U22051 ( .A(n21011), .B(n21012), .Z(n21009) );
  XNOR U22052 ( .A(n21010), .B(n20976), .Z(n21012) );
  XNOR U22053 ( .A(n21013), .B(n21014), .Z(n20976) );
  ANDN U22054 ( .B(n21015), .A(n21016), .Z(n21013) );
  XOR U22055 ( .A(n21014), .B(n21017), .Z(n21015) );
  XOR U22056 ( .A(n21010), .B(n20978), .Z(n21011) );
  XOR U22057 ( .A(n21018), .B(n21019), .Z(n20978) );
  AND U22058 ( .A(n914), .B(n21020), .Z(n21018) );
  XOR U22059 ( .A(n21021), .B(n21019), .Z(n21020) );
  XNOR U22060 ( .A(n21022), .B(n21023), .Z(n21010) );
  NAND U22061 ( .A(n21024), .B(n21025), .Z(n21023) );
  XOR U22062 ( .A(n21026), .B(n21002), .Z(n21025) );
  XOR U22063 ( .A(n21016), .B(n21017), .Z(n21002) );
  XOR U22064 ( .A(n21027), .B(n21028), .Z(n21017) );
  ANDN U22065 ( .B(n21029), .A(n21030), .Z(n21027) );
  XOR U22066 ( .A(n21028), .B(n21031), .Z(n21029) );
  XOR U22067 ( .A(n21032), .B(n21033), .Z(n21016) );
  XOR U22068 ( .A(n21034), .B(n21035), .Z(n21033) );
  ANDN U22069 ( .B(n21036), .A(n21037), .Z(n21034) );
  XOR U22070 ( .A(n21038), .B(n21035), .Z(n21036) );
  IV U22071 ( .A(n21014), .Z(n21032) );
  XOR U22072 ( .A(n21039), .B(n21040), .Z(n21014) );
  ANDN U22073 ( .B(n21041), .A(n21042), .Z(n21039) );
  XOR U22074 ( .A(n21040), .B(n21043), .Z(n21041) );
  IV U22075 ( .A(n21022), .Z(n21026) );
  XOR U22076 ( .A(n21022), .B(n21004), .Z(n21024) );
  XOR U22077 ( .A(n21044), .B(n21045), .Z(n21004) );
  AND U22078 ( .A(n914), .B(n21046), .Z(n21044) );
  XOR U22079 ( .A(n21047), .B(n21045), .Z(n21046) );
  NANDN U22080 ( .A(n21006), .B(n21008), .Z(n21022) );
  XOR U22081 ( .A(n21048), .B(n21049), .Z(n21008) );
  AND U22082 ( .A(n914), .B(n21050), .Z(n21048) );
  XOR U22083 ( .A(n21049), .B(n21051), .Z(n21050) );
  XOR U22084 ( .A(n21052), .B(n21053), .Z(n914) );
  AND U22085 ( .A(n21054), .B(n21055), .Z(n21052) );
  XNOR U22086 ( .A(n21053), .B(n21019), .Z(n21055) );
  XNOR U22087 ( .A(n21056), .B(n21057), .Z(n21019) );
  ANDN U22088 ( .B(n21058), .A(n21059), .Z(n21056) );
  XOR U22089 ( .A(n21057), .B(n21060), .Z(n21058) );
  XOR U22090 ( .A(n21053), .B(n21021), .Z(n21054) );
  XOR U22091 ( .A(n21061), .B(n21062), .Z(n21021) );
  AND U22092 ( .A(n918), .B(n21063), .Z(n21061) );
  XOR U22093 ( .A(n21064), .B(n21062), .Z(n21063) );
  XNOR U22094 ( .A(n21065), .B(n21066), .Z(n21053) );
  NAND U22095 ( .A(n21067), .B(n21068), .Z(n21066) );
  XOR U22096 ( .A(n21069), .B(n21045), .Z(n21068) );
  XOR U22097 ( .A(n21059), .B(n21060), .Z(n21045) );
  XOR U22098 ( .A(n21070), .B(n21071), .Z(n21060) );
  ANDN U22099 ( .B(n21072), .A(n21073), .Z(n21070) );
  XOR U22100 ( .A(n21071), .B(n21074), .Z(n21072) );
  XOR U22101 ( .A(n21075), .B(n21076), .Z(n21059) );
  XOR U22102 ( .A(n21077), .B(n21078), .Z(n21076) );
  ANDN U22103 ( .B(n21079), .A(n21080), .Z(n21077) );
  XOR U22104 ( .A(n21081), .B(n21078), .Z(n21079) );
  IV U22105 ( .A(n21057), .Z(n21075) );
  XOR U22106 ( .A(n21082), .B(n21083), .Z(n21057) );
  ANDN U22107 ( .B(n21084), .A(n21085), .Z(n21082) );
  XOR U22108 ( .A(n21083), .B(n21086), .Z(n21084) );
  IV U22109 ( .A(n21065), .Z(n21069) );
  XOR U22110 ( .A(n21065), .B(n21047), .Z(n21067) );
  XOR U22111 ( .A(n21087), .B(n21088), .Z(n21047) );
  AND U22112 ( .A(n918), .B(n21089), .Z(n21087) );
  XOR U22113 ( .A(n21090), .B(n21088), .Z(n21089) );
  NANDN U22114 ( .A(n21049), .B(n21051), .Z(n21065) );
  XOR U22115 ( .A(n21091), .B(n21092), .Z(n21051) );
  AND U22116 ( .A(n918), .B(n21093), .Z(n21091) );
  XOR U22117 ( .A(n21092), .B(n21094), .Z(n21093) );
  XOR U22118 ( .A(n21095), .B(n21096), .Z(n918) );
  AND U22119 ( .A(n21097), .B(n21098), .Z(n21095) );
  XNOR U22120 ( .A(n21096), .B(n21062), .Z(n21098) );
  XNOR U22121 ( .A(n21099), .B(n21100), .Z(n21062) );
  ANDN U22122 ( .B(n21101), .A(n21102), .Z(n21099) );
  XOR U22123 ( .A(n21100), .B(n21103), .Z(n21101) );
  XOR U22124 ( .A(n21096), .B(n21064), .Z(n21097) );
  XOR U22125 ( .A(n21104), .B(n21105), .Z(n21064) );
  AND U22126 ( .A(n922), .B(n21106), .Z(n21104) );
  XOR U22127 ( .A(n21107), .B(n21105), .Z(n21106) );
  XNOR U22128 ( .A(n21108), .B(n21109), .Z(n21096) );
  NAND U22129 ( .A(n21110), .B(n21111), .Z(n21109) );
  XOR U22130 ( .A(n21112), .B(n21088), .Z(n21111) );
  XOR U22131 ( .A(n21102), .B(n21103), .Z(n21088) );
  XOR U22132 ( .A(n21113), .B(n21114), .Z(n21103) );
  ANDN U22133 ( .B(n21115), .A(n21116), .Z(n21113) );
  XOR U22134 ( .A(n21114), .B(n21117), .Z(n21115) );
  XOR U22135 ( .A(n21118), .B(n21119), .Z(n21102) );
  XOR U22136 ( .A(n21120), .B(n21121), .Z(n21119) );
  ANDN U22137 ( .B(n21122), .A(n21123), .Z(n21120) );
  XOR U22138 ( .A(n21124), .B(n21121), .Z(n21122) );
  IV U22139 ( .A(n21100), .Z(n21118) );
  XOR U22140 ( .A(n21125), .B(n21126), .Z(n21100) );
  ANDN U22141 ( .B(n21127), .A(n21128), .Z(n21125) );
  XOR U22142 ( .A(n21126), .B(n21129), .Z(n21127) );
  IV U22143 ( .A(n21108), .Z(n21112) );
  XOR U22144 ( .A(n21108), .B(n21090), .Z(n21110) );
  XOR U22145 ( .A(n21130), .B(n21131), .Z(n21090) );
  AND U22146 ( .A(n922), .B(n21132), .Z(n21130) );
  XOR U22147 ( .A(n21133), .B(n21131), .Z(n21132) );
  NANDN U22148 ( .A(n21092), .B(n21094), .Z(n21108) );
  XOR U22149 ( .A(n21134), .B(n21135), .Z(n21094) );
  AND U22150 ( .A(n922), .B(n21136), .Z(n21134) );
  XOR U22151 ( .A(n21135), .B(n21137), .Z(n21136) );
  XOR U22152 ( .A(n21138), .B(n21139), .Z(n922) );
  AND U22153 ( .A(n21140), .B(n21141), .Z(n21138) );
  XNOR U22154 ( .A(n21139), .B(n21105), .Z(n21141) );
  XNOR U22155 ( .A(n21142), .B(n21143), .Z(n21105) );
  ANDN U22156 ( .B(n21144), .A(n21145), .Z(n21142) );
  XOR U22157 ( .A(n21143), .B(n21146), .Z(n21144) );
  XOR U22158 ( .A(n21139), .B(n21107), .Z(n21140) );
  XOR U22159 ( .A(n21147), .B(n21148), .Z(n21107) );
  AND U22160 ( .A(n926), .B(n21149), .Z(n21147) );
  XOR U22161 ( .A(n21150), .B(n21148), .Z(n21149) );
  XNOR U22162 ( .A(n21151), .B(n21152), .Z(n21139) );
  NAND U22163 ( .A(n21153), .B(n21154), .Z(n21152) );
  XOR U22164 ( .A(n21155), .B(n21131), .Z(n21154) );
  XOR U22165 ( .A(n21145), .B(n21146), .Z(n21131) );
  XOR U22166 ( .A(n21156), .B(n21157), .Z(n21146) );
  ANDN U22167 ( .B(n21158), .A(n21159), .Z(n21156) );
  XOR U22168 ( .A(n21157), .B(n21160), .Z(n21158) );
  XOR U22169 ( .A(n21161), .B(n21162), .Z(n21145) );
  XOR U22170 ( .A(n21163), .B(n21164), .Z(n21162) );
  ANDN U22171 ( .B(n21165), .A(n21166), .Z(n21163) );
  XOR U22172 ( .A(n21167), .B(n21164), .Z(n21165) );
  IV U22173 ( .A(n21143), .Z(n21161) );
  XOR U22174 ( .A(n21168), .B(n21169), .Z(n21143) );
  ANDN U22175 ( .B(n21170), .A(n21171), .Z(n21168) );
  XOR U22176 ( .A(n21169), .B(n21172), .Z(n21170) );
  IV U22177 ( .A(n21151), .Z(n21155) );
  XOR U22178 ( .A(n21151), .B(n21133), .Z(n21153) );
  XOR U22179 ( .A(n21173), .B(n21174), .Z(n21133) );
  AND U22180 ( .A(n926), .B(n21175), .Z(n21173) );
  XOR U22181 ( .A(n21176), .B(n21174), .Z(n21175) );
  NANDN U22182 ( .A(n21135), .B(n21137), .Z(n21151) );
  XOR U22183 ( .A(n21177), .B(n21178), .Z(n21137) );
  AND U22184 ( .A(n926), .B(n21179), .Z(n21177) );
  XOR U22185 ( .A(n21178), .B(n21180), .Z(n21179) );
  XOR U22186 ( .A(n21181), .B(n21182), .Z(n926) );
  AND U22187 ( .A(n21183), .B(n21184), .Z(n21181) );
  XNOR U22188 ( .A(n21182), .B(n21148), .Z(n21184) );
  XNOR U22189 ( .A(n21185), .B(n21186), .Z(n21148) );
  ANDN U22190 ( .B(n21187), .A(n21188), .Z(n21185) );
  XOR U22191 ( .A(n21186), .B(n21189), .Z(n21187) );
  XOR U22192 ( .A(n21182), .B(n21150), .Z(n21183) );
  XOR U22193 ( .A(n21190), .B(n21191), .Z(n21150) );
  AND U22194 ( .A(n930), .B(n21192), .Z(n21190) );
  XOR U22195 ( .A(n21193), .B(n21191), .Z(n21192) );
  XNOR U22196 ( .A(n21194), .B(n21195), .Z(n21182) );
  NAND U22197 ( .A(n21196), .B(n21197), .Z(n21195) );
  XOR U22198 ( .A(n21198), .B(n21174), .Z(n21197) );
  XOR U22199 ( .A(n21188), .B(n21189), .Z(n21174) );
  XOR U22200 ( .A(n21199), .B(n21200), .Z(n21189) );
  ANDN U22201 ( .B(n21201), .A(n21202), .Z(n21199) );
  XOR U22202 ( .A(n21200), .B(n21203), .Z(n21201) );
  XOR U22203 ( .A(n21204), .B(n21205), .Z(n21188) );
  XOR U22204 ( .A(n21206), .B(n21207), .Z(n21205) );
  ANDN U22205 ( .B(n21208), .A(n21209), .Z(n21206) );
  XOR U22206 ( .A(n21210), .B(n21207), .Z(n21208) );
  IV U22207 ( .A(n21186), .Z(n21204) );
  XOR U22208 ( .A(n21211), .B(n21212), .Z(n21186) );
  ANDN U22209 ( .B(n21213), .A(n21214), .Z(n21211) );
  XOR U22210 ( .A(n21212), .B(n21215), .Z(n21213) );
  IV U22211 ( .A(n21194), .Z(n21198) );
  XOR U22212 ( .A(n21194), .B(n21176), .Z(n21196) );
  XOR U22213 ( .A(n21216), .B(n21217), .Z(n21176) );
  AND U22214 ( .A(n930), .B(n21218), .Z(n21216) );
  XOR U22215 ( .A(n21219), .B(n21217), .Z(n21218) );
  NANDN U22216 ( .A(n21178), .B(n21180), .Z(n21194) );
  XOR U22217 ( .A(n21220), .B(n21221), .Z(n21180) );
  AND U22218 ( .A(n930), .B(n21222), .Z(n21220) );
  XOR U22219 ( .A(n21221), .B(n21223), .Z(n21222) );
  XOR U22220 ( .A(n21224), .B(n21225), .Z(n930) );
  AND U22221 ( .A(n21226), .B(n21227), .Z(n21224) );
  XNOR U22222 ( .A(n21225), .B(n21191), .Z(n21227) );
  XNOR U22223 ( .A(n21228), .B(n21229), .Z(n21191) );
  ANDN U22224 ( .B(n21230), .A(n21231), .Z(n21228) );
  XOR U22225 ( .A(n21229), .B(n21232), .Z(n21230) );
  XOR U22226 ( .A(n21225), .B(n21193), .Z(n21226) );
  XOR U22227 ( .A(n21233), .B(n21234), .Z(n21193) );
  AND U22228 ( .A(n934), .B(n21235), .Z(n21233) );
  XOR U22229 ( .A(n21236), .B(n21234), .Z(n21235) );
  XNOR U22230 ( .A(n21237), .B(n21238), .Z(n21225) );
  NAND U22231 ( .A(n21239), .B(n21240), .Z(n21238) );
  XOR U22232 ( .A(n21241), .B(n21217), .Z(n21240) );
  XOR U22233 ( .A(n21231), .B(n21232), .Z(n21217) );
  XOR U22234 ( .A(n21242), .B(n21243), .Z(n21232) );
  ANDN U22235 ( .B(n21244), .A(n21245), .Z(n21242) );
  XOR U22236 ( .A(n21243), .B(n21246), .Z(n21244) );
  XOR U22237 ( .A(n21247), .B(n21248), .Z(n21231) );
  XOR U22238 ( .A(n21249), .B(n21250), .Z(n21248) );
  ANDN U22239 ( .B(n21251), .A(n21252), .Z(n21249) );
  XOR U22240 ( .A(n21253), .B(n21250), .Z(n21251) );
  IV U22241 ( .A(n21229), .Z(n21247) );
  XOR U22242 ( .A(n21254), .B(n21255), .Z(n21229) );
  ANDN U22243 ( .B(n21256), .A(n21257), .Z(n21254) );
  XOR U22244 ( .A(n21255), .B(n21258), .Z(n21256) );
  IV U22245 ( .A(n21237), .Z(n21241) );
  XOR U22246 ( .A(n21237), .B(n21219), .Z(n21239) );
  XOR U22247 ( .A(n21259), .B(n21260), .Z(n21219) );
  AND U22248 ( .A(n934), .B(n21261), .Z(n21259) );
  XOR U22249 ( .A(n21262), .B(n21260), .Z(n21261) );
  NANDN U22250 ( .A(n21221), .B(n21223), .Z(n21237) );
  XOR U22251 ( .A(n21263), .B(n21264), .Z(n21223) );
  AND U22252 ( .A(n934), .B(n21265), .Z(n21263) );
  XOR U22253 ( .A(n21264), .B(n21266), .Z(n21265) );
  XOR U22254 ( .A(n21267), .B(n21268), .Z(n934) );
  AND U22255 ( .A(n21269), .B(n21270), .Z(n21267) );
  XNOR U22256 ( .A(n21268), .B(n21234), .Z(n21270) );
  XNOR U22257 ( .A(n21271), .B(n21272), .Z(n21234) );
  ANDN U22258 ( .B(n21273), .A(n21274), .Z(n21271) );
  XOR U22259 ( .A(n21272), .B(n21275), .Z(n21273) );
  XOR U22260 ( .A(n21268), .B(n21236), .Z(n21269) );
  XOR U22261 ( .A(n21276), .B(n21277), .Z(n21236) );
  AND U22262 ( .A(n938), .B(n21278), .Z(n21276) );
  XOR U22263 ( .A(n21279), .B(n21277), .Z(n21278) );
  XNOR U22264 ( .A(n21280), .B(n21281), .Z(n21268) );
  NAND U22265 ( .A(n21282), .B(n21283), .Z(n21281) );
  XOR U22266 ( .A(n21284), .B(n21260), .Z(n21283) );
  XOR U22267 ( .A(n21274), .B(n21275), .Z(n21260) );
  XOR U22268 ( .A(n21285), .B(n21286), .Z(n21275) );
  ANDN U22269 ( .B(n21287), .A(n21288), .Z(n21285) );
  XOR U22270 ( .A(n21286), .B(n21289), .Z(n21287) );
  XOR U22271 ( .A(n21290), .B(n21291), .Z(n21274) );
  XOR U22272 ( .A(n21292), .B(n21293), .Z(n21291) );
  ANDN U22273 ( .B(n21294), .A(n21295), .Z(n21292) );
  XOR U22274 ( .A(n21296), .B(n21293), .Z(n21294) );
  IV U22275 ( .A(n21272), .Z(n21290) );
  XOR U22276 ( .A(n21297), .B(n21298), .Z(n21272) );
  ANDN U22277 ( .B(n21299), .A(n21300), .Z(n21297) );
  XOR U22278 ( .A(n21298), .B(n21301), .Z(n21299) );
  IV U22279 ( .A(n21280), .Z(n21284) );
  XOR U22280 ( .A(n21280), .B(n21262), .Z(n21282) );
  XOR U22281 ( .A(n21302), .B(n21303), .Z(n21262) );
  AND U22282 ( .A(n938), .B(n21304), .Z(n21302) );
  XOR U22283 ( .A(n21305), .B(n21303), .Z(n21304) );
  NANDN U22284 ( .A(n21264), .B(n21266), .Z(n21280) );
  XOR U22285 ( .A(n21306), .B(n21307), .Z(n21266) );
  AND U22286 ( .A(n938), .B(n21308), .Z(n21306) );
  XOR U22287 ( .A(n21307), .B(n21309), .Z(n21308) );
  XOR U22288 ( .A(n21310), .B(n21311), .Z(n938) );
  AND U22289 ( .A(n21312), .B(n21313), .Z(n21310) );
  XNOR U22290 ( .A(n21311), .B(n21277), .Z(n21313) );
  XNOR U22291 ( .A(n21314), .B(n21315), .Z(n21277) );
  ANDN U22292 ( .B(n21316), .A(n21317), .Z(n21314) );
  XOR U22293 ( .A(n21315), .B(n21318), .Z(n21316) );
  XOR U22294 ( .A(n21311), .B(n21279), .Z(n21312) );
  XOR U22295 ( .A(n21319), .B(n21320), .Z(n21279) );
  AND U22296 ( .A(n942), .B(n21321), .Z(n21319) );
  XOR U22297 ( .A(n21322), .B(n21320), .Z(n21321) );
  XNOR U22298 ( .A(n21323), .B(n21324), .Z(n21311) );
  NAND U22299 ( .A(n21325), .B(n21326), .Z(n21324) );
  XOR U22300 ( .A(n21327), .B(n21303), .Z(n21326) );
  XOR U22301 ( .A(n21317), .B(n21318), .Z(n21303) );
  XOR U22302 ( .A(n21328), .B(n21329), .Z(n21318) );
  ANDN U22303 ( .B(n21330), .A(n21331), .Z(n21328) );
  XOR U22304 ( .A(n21329), .B(n21332), .Z(n21330) );
  XOR U22305 ( .A(n21333), .B(n21334), .Z(n21317) );
  XOR U22306 ( .A(n21335), .B(n21336), .Z(n21334) );
  ANDN U22307 ( .B(n21337), .A(n21338), .Z(n21335) );
  XOR U22308 ( .A(n21339), .B(n21336), .Z(n21337) );
  IV U22309 ( .A(n21315), .Z(n21333) );
  XOR U22310 ( .A(n21340), .B(n21341), .Z(n21315) );
  ANDN U22311 ( .B(n21342), .A(n21343), .Z(n21340) );
  XOR U22312 ( .A(n21341), .B(n21344), .Z(n21342) );
  IV U22313 ( .A(n21323), .Z(n21327) );
  XOR U22314 ( .A(n21323), .B(n21305), .Z(n21325) );
  XOR U22315 ( .A(n21345), .B(n21346), .Z(n21305) );
  AND U22316 ( .A(n942), .B(n21347), .Z(n21345) );
  XOR U22317 ( .A(n21348), .B(n21346), .Z(n21347) );
  NANDN U22318 ( .A(n21307), .B(n21309), .Z(n21323) );
  XOR U22319 ( .A(n21349), .B(n21350), .Z(n21309) );
  AND U22320 ( .A(n942), .B(n21351), .Z(n21349) );
  XOR U22321 ( .A(n21350), .B(n21352), .Z(n21351) );
  XOR U22322 ( .A(n21353), .B(n21354), .Z(n942) );
  AND U22323 ( .A(n21355), .B(n21356), .Z(n21353) );
  XNOR U22324 ( .A(n21354), .B(n21320), .Z(n21356) );
  XNOR U22325 ( .A(n21357), .B(n21358), .Z(n21320) );
  ANDN U22326 ( .B(n21359), .A(n21360), .Z(n21357) );
  XOR U22327 ( .A(n21358), .B(n21361), .Z(n21359) );
  XOR U22328 ( .A(n21354), .B(n21322), .Z(n21355) );
  XOR U22329 ( .A(n21362), .B(n21363), .Z(n21322) );
  AND U22330 ( .A(n946), .B(n21364), .Z(n21362) );
  XOR U22331 ( .A(n21365), .B(n21363), .Z(n21364) );
  XNOR U22332 ( .A(n21366), .B(n21367), .Z(n21354) );
  NAND U22333 ( .A(n21368), .B(n21369), .Z(n21367) );
  XOR U22334 ( .A(n21370), .B(n21346), .Z(n21369) );
  XOR U22335 ( .A(n21360), .B(n21361), .Z(n21346) );
  XOR U22336 ( .A(n21371), .B(n21372), .Z(n21361) );
  ANDN U22337 ( .B(n21373), .A(n21374), .Z(n21371) );
  XOR U22338 ( .A(n21372), .B(n21375), .Z(n21373) );
  XOR U22339 ( .A(n21376), .B(n21377), .Z(n21360) );
  XOR U22340 ( .A(n21378), .B(n21379), .Z(n21377) );
  ANDN U22341 ( .B(n21380), .A(n21381), .Z(n21378) );
  XOR U22342 ( .A(n21382), .B(n21379), .Z(n21380) );
  IV U22343 ( .A(n21358), .Z(n21376) );
  XOR U22344 ( .A(n21383), .B(n21384), .Z(n21358) );
  ANDN U22345 ( .B(n21385), .A(n21386), .Z(n21383) );
  XOR U22346 ( .A(n21384), .B(n21387), .Z(n21385) );
  IV U22347 ( .A(n21366), .Z(n21370) );
  XOR U22348 ( .A(n21366), .B(n21348), .Z(n21368) );
  XOR U22349 ( .A(n21388), .B(n21389), .Z(n21348) );
  AND U22350 ( .A(n946), .B(n21390), .Z(n21388) );
  XOR U22351 ( .A(n21391), .B(n21389), .Z(n21390) );
  NANDN U22352 ( .A(n21350), .B(n21352), .Z(n21366) );
  XOR U22353 ( .A(n21392), .B(n21393), .Z(n21352) );
  AND U22354 ( .A(n946), .B(n21394), .Z(n21392) );
  XOR U22355 ( .A(n21393), .B(n21395), .Z(n21394) );
  XOR U22356 ( .A(n21396), .B(n21397), .Z(n946) );
  AND U22357 ( .A(n21398), .B(n21399), .Z(n21396) );
  XNOR U22358 ( .A(n21397), .B(n21363), .Z(n21399) );
  XNOR U22359 ( .A(n21400), .B(n21401), .Z(n21363) );
  ANDN U22360 ( .B(n21402), .A(n21403), .Z(n21400) );
  XOR U22361 ( .A(n21401), .B(n21404), .Z(n21402) );
  XOR U22362 ( .A(n21397), .B(n21365), .Z(n21398) );
  XOR U22363 ( .A(n21405), .B(n21406), .Z(n21365) );
  AND U22364 ( .A(n950), .B(n21407), .Z(n21405) );
  XOR U22365 ( .A(n21408), .B(n21406), .Z(n21407) );
  XNOR U22366 ( .A(n21409), .B(n21410), .Z(n21397) );
  NAND U22367 ( .A(n21411), .B(n21412), .Z(n21410) );
  XOR U22368 ( .A(n21413), .B(n21389), .Z(n21412) );
  XOR U22369 ( .A(n21403), .B(n21404), .Z(n21389) );
  XOR U22370 ( .A(n21414), .B(n21415), .Z(n21404) );
  ANDN U22371 ( .B(n21416), .A(n21417), .Z(n21414) );
  XOR U22372 ( .A(n21415), .B(n21418), .Z(n21416) );
  XOR U22373 ( .A(n21419), .B(n21420), .Z(n21403) );
  XOR U22374 ( .A(n21421), .B(n21422), .Z(n21420) );
  ANDN U22375 ( .B(n21423), .A(n21424), .Z(n21421) );
  XOR U22376 ( .A(n21425), .B(n21422), .Z(n21423) );
  IV U22377 ( .A(n21401), .Z(n21419) );
  XOR U22378 ( .A(n21426), .B(n21427), .Z(n21401) );
  ANDN U22379 ( .B(n21428), .A(n21429), .Z(n21426) );
  XOR U22380 ( .A(n21427), .B(n21430), .Z(n21428) );
  IV U22381 ( .A(n21409), .Z(n21413) );
  XOR U22382 ( .A(n21409), .B(n21391), .Z(n21411) );
  XOR U22383 ( .A(n21431), .B(n21432), .Z(n21391) );
  AND U22384 ( .A(n950), .B(n21433), .Z(n21431) );
  XOR U22385 ( .A(n21434), .B(n21432), .Z(n21433) );
  NANDN U22386 ( .A(n21393), .B(n21395), .Z(n21409) );
  XOR U22387 ( .A(n21435), .B(n21436), .Z(n21395) );
  AND U22388 ( .A(n950), .B(n21437), .Z(n21435) );
  XOR U22389 ( .A(n21436), .B(n21438), .Z(n21437) );
  XOR U22390 ( .A(n21439), .B(n21440), .Z(n950) );
  AND U22391 ( .A(n21441), .B(n21442), .Z(n21439) );
  XNOR U22392 ( .A(n21440), .B(n21406), .Z(n21442) );
  XNOR U22393 ( .A(n21443), .B(n21444), .Z(n21406) );
  ANDN U22394 ( .B(n21445), .A(n21446), .Z(n21443) );
  XOR U22395 ( .A(n21444), .B(n21447), .Z(n21445) );
  XOR U22396 ( .A(n21440), .B(n21408), .Z(n21441) );
  XOR U22397 ( .A(n21448), .B(n21449), .Z(n21408) );
  AND U22398 ( .A(n954), .B(n21450), .Z(n21448) );
  XOR U22399 ( .A(n21451), .B(n21449), .Z(n21450) );
  XNOR U22400 ( .A(n21452), .B(n21453), .Z(n21440) );
  NAND U22401 ( .A(n21454), .B(n21455), .Z(n21453) );
  XOR U22402 ( .A(n21456), .B(n21432), .Z(n21455) );
  XOR U22403 ( .A(n21446), .B(n21447), .Z(n21432) );
  XOR U22404 ( .A(n21457), .B(n21458), .Z(n21447) );
  ANDN U22405 ( .B(n21459), .A(n21460), .Z(n21457) );
  XOR U22406 ( .A(n21458), .B(n21461), .Z(n21459) );
  XOR U22407 ( .A(n21462), .B(n21463), .Z(n21446) );
  XOR U22408 ( .A(n21464), .B(n21465), .Z(n21463) );
  ANDN U22409 ( .B(n21466), .A(n21467), .Z(n21464) );
  XOR U22410 ( .A(n21468), .B(n21465), .Z(n21466) );
  IV U22411 ( .A(n21444), .Z(n21462) );
  XOR U22412 ( .A(n21469), .B(n21470), .Z(n21444) );
  ANDN U22413 ( .B(n21471), .A(n21472), .Z(n21469) );
  XOR U22414 ( .A(n21470), .B(n21473), .Z(n21471) );
  IV U22415 ( .A(n21452), .Z(n21456) );
  XOR U22416 ( .A(n21452), .B(n21434), .Z(n21454) );
  XOR U22417 ( .A(n21474), .B(n21475), .Z(n21434) );
  AND U22418 ( .A(n954), .B(n21476), .Z(n21474) );
  XOR U22419 ( .A(n21477), .B(n21475), .Z(n21476) );
  NANDN U22420 ( .A(n21436), .B(n21438), .Z(n21452) );
  XOR U22421 ( .A(n21478), .B(n21479), .Z(n21438) );
  AND U22422 ( .A(n954), .B(n21480), .Z(n21478) );
  XOR U22423 ( .A(n21479), .B(n21481), .Z(n21480) );
  XOR U22424 ( .A(n21482), .B(n21483), .Z(n954) );
  AND U22425 ( .A(n21484), .B(n21485), .Z(n21482) );
  XNOR U22426 ( .A(n21483), .B(n21449), .Z(n21485) );
  XNOR U22427 ( .A(n21486), .B(n21487), .Z(n21449) );
  ANDN U22428 ( .B(n21488), .A(n21489), .Z(n21486) );
  XOR U22429 ( .A(n21487), .B(n21490), .Z(n21488) );
  XOR U22430 ( .A(n21483), .B(n21451), .Z(n21484) );
  XOR U22431 ( .A(n21491), .B(n21492), .Z(n21451) );
  AND U22432 ( .A(n958), .B(n21493), .Z(n21491) );
  XOR U22433 ( .A(n21494), .B(n21492), .Z(n21493) );
  XNOR U22434 ( .A(n21495), .B(n21496), .Z(n21483) );
  NAND U22435 ( .A(n21497), .B(n21498), .Z(n21496) );
  XOR U22436 ( .A(n21499), .B(n21475), .Z(n21498) );
  XOR U22437 ( .A(n21489), .B(n21490), .Z(n21475) );
  XOR U22438 ( .A(n21500), .B(n21501), .Z(n21490) );
  ANDN U22439 ( .B(n21502), .A(n21503), .Z(n21500) );
  XOR U22440 ( .A(n21501), .B(n21504), .Z(n21502) );
  XOR U22441 ( .A(n21505), .B(n21506), .Z(n21489) );
  XOR U22442 ( .A(n21507), .B(n21508), .Z(n21506) );
  ANDN U22443 ( .B(n21509), .A(n21510), .Z(n21507) );
  XOR U22444 ( .A(n21511), .B(n21508), .Z(n21509) );
  IV U22445 ( .A(n21487), .Z(n21505) );
  XOR U22446 ( .A(n21512), .B(n21513), .Z(n21487) );
  ANDN U22447 ( .B(n21514), .A(n21515), .Z(n21512) );
  XOR U22448 ( .A(n21513), .B(n21516), .Z(n21514) );
  IV U22449 ( .A(n21495), .Z(n21499) );
  XOR U22450 ( .A(n21495), .B(n21477), .Z(n21497) );
  XOR U22451 ( .A(n21517), .B(n21518), .Z(n21477) );
  AND U22452 ( .A(n958), .B(n21519), .Z(n21517) );
  XOR U22453 ( .A(n21520), .B(n21518), .Z(n21519) );
  NANDN U22454 ( .A(n21479), .B(n21481), .Z(n21495) );
  XOR U22455 ( .A(n21521), .B(n21522), .Z(n21481) );
  AND U22456 ( .A(n958), .B(n21523), .Z(n21521) );
  XOR U22457 ( .A(n21522), .B(n21524), .Z(n21523) );
  XOR U22458 ( .A(n21525), .B(n21526), .Z(n958) );
  AND U22459 ( .A(n21527), .B(n21528), .Z(n21525) );
  XNOR U22460 ( .A(n21526), .B(n21492), .Z(n21528) );
  XNOR U22461 ( .A(n21529), .B(n21530), .Z(n21492) );
  ANDN U22462 ( .B(n21531), .A(n21532), .Z(n21529) );
  XOR U22463 ( .A(n21530), .B(n21533), .Z(n21531) );
  XOR U22464 ( .A(n21526), .B(n21494), .Z(n21527) );
  XOR U22465 ( .A(n21534), .B(n21535), .Z(n21494) );
  AND U22466 ( .A(n962), .B(n21536), .Z(n21534) );
  XOR U22467 ( .A(n21537), .B(n21535), .Z(n21536) );
  XNOR U22468 ( .A(n21538), .B(n21539), .Z(n21526) );
  NAND U22469 ( .A(n21540), .B(n21541), .Z(n21539) );
  XOR U22470 ( .A(n21542), .B(n21518), .Z(n21541) );
  XOR U22471 ( .A(n21532), .B(n21533), .Z(n21518) );
  XOR U22472 ( .A(n21543), .B(n21544), .Z(n21533) );
  ANDN U22473 ( .B(n21545), .A(n21546), .Z(n21543) );
  XOR U22474 ( .A(n21544), .B(n21547), .Z(n21545) );
  XOR U22475 ( .A(n21548), .B(n21549), .Z(n21532) );
  XOR U22476 ( .A(n21550), .B(n21551), .Z(n21549) );
  ANDN U22477 ( .B(n21552), .A(n21553), .Z(n21550) );
  XOR U22478 ( .A(n21554), .B(n21551), .Z(n21552) );
  IV U22479 ( .A(n21530), .Z(n21548) );
  XOR U22480 ( .A(n21555), .B(n21556), .Z(n21530) );
  ANDN U22481 ( .B(n21557), .A(n21558), .Z(n21555) );
  XOR U22482 ( .A(n21556), .B(n21559), .Z(n21557) );
  IV U22483 ( .A(n21538), .Z(n21542) );
  XOR U22484 ( .A(n21538), .B(n21520), .Z(n21540) );
  XOR U22485 ( .A(n21560), .B(n21561), .Z(n21520) );
  AND U22486 ( .A(n962), .B(n21562), .Z(n21560) );
  XOR U22487 ( .A(n21563), .B(n21561), .Z(n21562) );
  NANDN U22488 ( .A(n21522), .B(n21524), .Z(n21538) );
  XOR U22489 ( .A(n21564), .B(n21565), .Z(n21524) );
  AND U22490 ( .A(n962), .B(n21566), .Z(n21564) );
  XOR U22491 ( .A(n21565), .B(n21567), .Z(n21566) );
  XOR U22492 ( .A(n21568), .B(n21569), .Z(n962) );
  AND U22493 ( .A(n21570), .B(n21571), .Z(n21568) );
  XNOR U22494 ( .A(n21569), .B(n21535), .Z(n21571) );
  XNOR U22495 ( .A(n21572), .B(n21573), .Z(n21535) );
  ANDN U22496 ( .B(n21574), .A(n21575), .Z(n21572) );
  XOR U22497 ( .A(n21573), .B(n21576), .Z(n21574) );
  XOR U22498 ( .A(n21569), .B(n21537), .Z(n21570) );
  XOR U22499 ( .A(n21577), .B(n21578), .Z(n21537) );
  AND U22500 ( .A(n966), .B(n21579), .Z(n21577) );
  XOR U22501 ( .A(n21580), .B(n21578), .Z(n21579) );
  XNOR U22502 ( .A(n21581), .B(n21582), .Z(n21569) );
  NAND U22503 ( .A(n21583), .B(n21584), .Z(n21582) );
  XOR U22504 ( .A(n21585), .B(n21561), .Z(n21584) );
  XOR U22505 ( .A(n21575), .B(n21576), .Z(n21561) );
  XOR U22506 ( .A(n21586), .B(n21587), .Z(n21576) );
  ANDN U22507 ( .B(n21588), .A(n21589), .Z(n21586) );
  XOR U22508 ( .A(n21587), .B(n21590), .Z(n21588) );
  XOR U22509 ( .A(n21591), .B(n21592), .Z(n21575) );
  XOR U22510 ( .A(n21593), .B(n21594), .Z(n21592) );
  ANDN U22511 ( .B(n21595), .A(n21596), .Z(n21593) );
  XOR U22512 ( .A(n21597), .B(n21594), .Z(n21595) );
  IV U22513 ( .A(n21573), .Z(n21591) );
  XOR U22514 ( .A(n21598), .B(n21599), .Z(n21573) );
  ANDN U22515 ( .B(n21600), .A(n21601), .Z(n21598) );
  XOR U22516 ( .A(n21599), .B(n21602), .Z(n21600) );
  IV U22517 ( .A(n21581), .Z(n21585) );
  XOR U22518 ( .A(n21581), .B(n21563), .Z(n21583) );
  XOR U22519 ( .A(n21603), .B(n21604), .Z(n21563) );
  AND U22520 ( .A(n966), .B(n21605), .Z(n21603) );
  XOR U22521 ( .A(n21606), .B(n21604), .Z(n21605) );
  NANDN U22522 ( .A(n21565), .B(n21567), .Z(n21581) );
  XOR U22523 ( .A(n21607), .B(n21608), .Z(n21567) );
  AND U22524 ( .A(n966), .B(n21609), .Z(n21607) );
  XOR U22525 ( .A(n21608), .B(n21610), .Z(n21609) );
  XOR U22526 ( .A(n21611), .B(n21612), .Z(n966) );
  AND U22527 ( .A(n21613), .B(n21614), .Z(n21611) );
  XNOR U22528 ( .A(n21612), .B(n21578), .Z(n21614) );
  XNOR U22529 ( .A(n21615), .B(n21616), .Z(n21578) );
  ANDN U22530 ( .B(n21617), .A(n21618), .Z(n21615) );
  XOR U22531 ( .A(n21616), .B(n21619), .Z(n21617) );
  XOR U22532 ( .A(n21612), .B(n21580), .Z(n21613) );
  XOR U22533 ( .A(n21620), .B(n21621), .Z(n21580) );
  AND U22534 ( .A(n970), .B(n21622), .Z(n21620) );
  XOR U22535 ( .A(n21623), .B(n21621), .Z(n21622) );
  XNOR U22536 ( .A(n21624), .B(n21625), .Z(n21612) );
  NAND U22537 ( .A(n21626), .B(n21627), .Z(n21625) );
  XOR U22538 ( .A(n21628), .B(n21604), .Z(n21627) );
  XOR U22539 ( .A(n21618), .B(n21619), .Z(n21604) );
  XOR U22540 ( .A(n21629), .B(n21630), .Z(n21619) );
  ANDN U22541 ( .B(n21631), .A(n21632), .Z(n21629) );
  XOR U22542 ( .A(n21630), .B(n21633), .Z(n21631) );
  XOR U22543 ( .A(n21634), .B(n21635), .Z(n21618) );
  XOR U22544 ( .A(n21636), .B(n21637), .Z(n21635) );
  ANDN U22545 ( .B(n21638), .A(n21639), .Z(n21636) );
  XOR U22546 ( .A(n21640), .B(n21637), .Z(n21638) );
  IV U22547 ( .A(n21616), .Z(n21634) );
  XOR U22548 ( .A(n21641), .B(n21642), .Z(n21616) );
  ANDN U22549 ( .B(n21643), .A(n21644), .Z(n21641) );
  XOR U22550 ( .A(n21642), .B(n21645), .Z(n21643) );
  IV U22551 ( .A(n21624), .Z(n21628) );
  XOR U22552 ( .A(n21624), .B(n21606), .Z(n21626) );
  XOR U22553 ( .A(n21646), .B(n21647), .Z(n21606) );
  AND U22554 ( .A(n970), .B(n21648), .Z(n21646) );
  XOR U22555 ( .A(n21649), .B(n21647), .Z(n21648) );
  NANDN U22556 ( .A(n21608), .B(n21610), .Z(n21624) );
  XOR U22557 ( .A(n21650), .B(n21651), .Z(n21610) );
  AND U22558 ( .A(n970), .B(n21652), .Z(n21650) );
  XOR U22559 ( .A(n21651), .B(n21653), .Z(n21652) );
  XOR U22560 ( .A(n21654), .B(n21655), .Z(n970) );
  AND U22561 ( .A(n21656), .B(n21657), .Z(n21654) );
  XNOR U22562 ( .A(n21655), .B(n21621), .Z(n21657) );
  XNOR U22563 ( .A(n21658), .B(n21659), .Z(n21621) );
  ANDN U22564 ( .B(n21660), .A(n21661), .Z(n21658) );
  XOR U22565 ( .A(n21659), .B(n21662), .Z(n21660) );
  XOR U22566 ( .A(n21655), .B(n21623), .Z(n21656) );
  XOR U22567 ( .A(n21663), .B(n21664), .Z(n21623) );
  AND U22568 ( .A(n974), .B(n21665), .Z(n21663) );
  XOR U22569 ( .A(n21666), .B(n21664), .Z(n21665) );
  XNOR U22570 ( .A(n21667), .B(n21668), .Z(n21655) );
  NAND U22571 ( .A(n21669), .B(n21670), .Z(n21668) );
  XOR U22572 ( .A(n21671), .B(n21647), .Z(n21670) );
  XOR U22573 ( .A(n21661), .B(n21662), .Z(n21647) );
  XOR U22574 ( .A(n21672), .B(n21673), .Z(n21662) );
  ANDN U22575 ( .B(n21674), .A(n21675), .Z(n21672) );
  XOR U22576 ( .A(n21673), .B(n21676), .Z(n21674) );
  XOR U22577 ( .A(n21677), .B(n21678), .Z(n21661) );
  XOR U22578 ( .A(n21679), .B(n21680), .Z(n21678) );
  ANDN U22579 ( .B(n21681), .A(n21682), .Z(n21679) );
  XOR U22580 ( .A(n21683), .B(n21680), .Z(n21681) );
  IV U22581 ( .A(n21659), .Z(n21677) );
  XOR U22582 ( .A(n21684), .B(n21685), .Z(n21659) );
  ANDN U22583 ( .B(n21686), .A(n21687), .Z(n21684) );
  XOR U22584 ( .A(n21685), .B(n21688), .Z(n21686) );
  IV U22585 ( .A(n21667), .Z(n21671) );
  XOR U22586 ( .A(n21667), .B(n21649), .Z(n21669) );
  XOR U22587 ( .A(n21689), .B(n21690), .Z(n21649) );
  AND U22588 ( .A(n974), .B(n21691), .Z(n21689) );
  XOR U22589 ( .A(n21692), .B(n21690), .Z(n21691) );
  NANDN U22590 ( .A(n21651), .B(n21653), .Z(n21667) );
  XOR U22591 ( .A(n21693), .B(n21694), .Z(n21653) );
  AND U22592 ( .A(n974), .B(n21695), .Z(n21693) );
  XOR U22593 ( .A(n21694), .B(n21696), .Z(n21695) );
  XOR U22594 ( .A(n21697), .B(n21698), .Z(n974) );
  AND U22595 ( .A(n21699), .B(n21700), .Z(n21697) );
  XNOR U22596 ( .A(n21698), .B(n21664), .Z(n21700) );
  XNOR U22597 ( .A(n21701), .B(n21702), .Z(n21664) );
  ANDN U22598 ( .B(n21703), .A(n21704), .Z(n21701) );
  XOR U22599 ( .A(n21702), .B(n21705), .Z(n21703) );
  XOR U22600 ( .A(n21698), .B(n21666), .Z(n21699) );
  XOR U22601 ( .A(n21706), .B(n21707), .Z(n21666) );
  AND U22602 ( .A(n978), .B(n21708), .Z(n21706) );
  XOR U22603 ( .A(n21709), .B(n21707), .Z(n21708) );
  XNOR U22604 ( .A(n21710), .B(n21711), .Z(n21698) );
  NAND U22605 ( .A(n21712), .B(n21713), .Z(n21711) );
  XOR U22606 ( .A(n21714), .B(n21690), .Z(n21713) );
  XOR U22607 ( .A(n21704), .B(n21705), .Z(n21690) );
  XOR U22608 ( .A(n21715), .B(n21716), .Z(n21705) );
  ANDN U22609 ( .B(n21717), .A(n21718), .Z(n21715) );
  XOR U22610 ( .A(n21716), .B(n21719), .Z(n21717) );
  XOR U22611 ( .A(n21720), .B(n21721), .Z(n21704) );
  XOR U22612 ( .A(n21722), .B(n21723), .Z(n21721) );
  ANDN U22613 ( .B(n21724), .A(n21725), .Z(n21722) );
  XOR U22614 ( .A(n21726), .B(n21723), .Z(n21724) );
  IV U22615 ( .A(n21702), .Z(n21720) );
  XOR U22616 ( .A(n21727), .B(n21728), .Z(n21702) );
  ANDN U22617 ( .B(n21729), .A(n21730), .Z(n21727) );
  XOR U22618 ( .A(n21728), .B(n21731), .Z(n21729) );
  IV U22619 ( .A(n21710), .Z(n21714) );
  XOR U22620 ( .A(n21710), .B(n21692), .Z(n21712) );
  XOR U22621 ( .A(n21732), .B(n21733), .Z(n21692) );
  AND U22622 ( .A(n978), .B(n21734), .Z(n21732) );
  XOR U22623 ( .A(n21735), .B(n21733), .Z(n21734) );
  NANDN U22624 ( .A(n21694), .B(n21696), .Z(n21710) );
  XOR U22625 ( .A(n21736), .B(n21737), .Z(n21696) );
  AND U22626 ( .A(n978), .B(n21738), .Z(n21736) );
  XOR U22627 ( .A(n21737), .B(n21739), .Z(n21738) );
  XOR U22628 ( .A(n21740), .B(n21741), .Z(n978) );
  AND U22629 ( .A(n21742), .B(n21743), .Z(n21740) );
  XNOR U22630 ( .A(n21741), .B(n21707), .Z(n21743) );
  XNOR U22631 ( .A(n21744), .B(n21745), .Z(n21707) );
  ANDN U22632 ( .B(n21746), .A(n21747), .Z(n21744) );
  XOR U22633 ( .A(n21745), .B(n21748), .Z(n21746) );
  XOR U22634 ( .A(n21741), .B(n21709), .Z(n21742) );
  XOR U22635 ( .A(n21749), .B(n21750), .Z(n21709) );
  AND U22636 ( .A(n982), .B(n21751), .Z(n21749) );
  XOR U22637 ( .A(n21752), .B(n21750), .Z(n21751) );
  XNOR U22638 ( .A(n21753), .B(n21754), .Z(n21741) );
  NAND U22639 ( .A(n21755), .B(n21756), .Z(n21754) );
  XOR U22640 ( .A(n21757), .B(n21733), .Z(n21756) );
  XOR U22641 ( .A(n21747), .B(n21748), .Z(n21733) );
  XOR U22642 ( .A(n21758), .B(n21759), .Z(n21748) );
  ANDN U22643 ( .B(n21760), .A(n21761), .Z(n21758) );
  XOR U22644 ( .A(n21759), .B(n21762), .Z(n21760) );
  XOR U22645 ( .A(n21763), .B(n21764), .Z(n21747) );
  XOR U22646 ( .A(n21765), .B(n21766), .Z(n21764) );
  ANDN U22647 ( .B(n21767), .A(n21768), .Z(n21765) );
  XOR U22648 ( .A(n21769), .B(n21766), .Z(n21767) );
  IV U22649 ( .A(n21745), .Z(n21763) );
  XOR U22650 ( .A(n21770), .B(n21771), .Z(n21745) );
  ANDN U22651 ( .B(n21772), .A(n21773), .Z(n21770) );
  XOR U22652 ( .A(n21771), .B(n21774), .Z(n21772) );
  IV U22653 ( .A(n21753), .Z(n21757) );
  XOR U22654 ( .A(n21753), .B(n21735), .Z(n21755) );
  XOR U22655 ( .A(n21775), .B(n21776), .Z(n21735) );
  AND U22656 ( .A(n982), .B(n21777), .Z(n21775) );
  XOR U22657 ( .A(n21778), .B(n21776), .Z(n21777) );
  NANDN U22658 ( .A(n21737), .B(n21739), .Z(n21753) );
  XOR U22659 ( .A(n21779), .B(n21780), .Z(n21739) );
  AND U22660 ( .A(n982), .B(n21781), .Z(n21779) );
  XOR U22661 ( .A(n21780), .B(n21782), .Z(n21781) );
  XOR U22662 ( .A(n21783), .B(n21784), .Z(n982) );
  AND U22663 ( .A(n21785), .B(n21786), .Z(n21783) );
  XNOR U22664 ( .A(n21784), .B(n21750), .Z(n21786) );
  XNOR U22665 ( .A(n21787), .B(n21788), .Z(n21750) );
  ANDN U22666 ( .B(n21789), .A(n21790), .Z(n21787) );
  XOR U22667 ( .A(n21788), .B(n21791), .Z(n21789) );
  XOR U22668 ( .A(n21784), .B(n21752), .Z(n21785) );
  XOR U22669 ( .A(n21792), .B(n21793), .Z(n21752) );
  AND U22670 ( .A(n986), .B(n21794), .Z(n21792) );
  XOR U22671 ( .A(n21795), .B(n21793), .Z(n21794) );
  XNOR U22672 ( .A(n21796), .B(n21797), .Z(n21784) );
  NAND U22673 ( .A(n21798), .B(n21799), .Z(n21797) );
  XOR U22674 ( .A(n21800), .B(n21776), .Z(n21799) );
  XOR U22675 ( .A(n21790), .B(n21791), .Z(n21776) );
  XOR U22676 ( .A(n21801), .B(n21802), .Z(n21791) );
  ANDN U22677 ( .B(n21803), .A(n21804), .Z(n21801) );
  XOR U22678 ( .A(n21802), .B(n21805), .Z(n21803) );
  XOR U22679 ( .A(n21806), .B(n21807), .Z(n21790) );
  XOR U22680 ( .A(n21808), .B(n21809), .Z(n21807) );
  ANDN U22681 ( .B(n21810), .A(n21811), .Z(n21808) );
  XOR U22682 ( .A(n21812), .B(n21809), .Z(n21810) );
  IV U22683 ( .A(n21788), .Z(n21806) );
  XOR U22684 ( .A(n21813), .B(n21814), .Z(n21788) );
  ANDN U22685 ( .B(n21815), .A(n21816), .Z(n21813) );
  XOR U22686 ( .A(n21814), .B(n21817), .Z(n21815) );
  IV U22687 ( .A(n21796), .Z(n21800) );
  XOR U22688 ( .A(n21796), .B(n21778), .Z(n21798) );
  XOR U22689 ( .A(n21818), .B(n21819), .Z(n21778) );
  AND U22690 ( .A(n986), .B(n21820), .Z(n21818) );
  XOR U22691 ( .A(n21821), .B(n21819), .Z(n21820) );
  NANDN U22692 ( .A(n21780), .B(n21782), .Z(n21796) );
  XOR U22693 ( .A(n21822), .B(n21823), .Z(n21782) );
  AND U22694 ( .A(n986), .B(n21824), .Z(n21822) );
  XOR U22695 ( .A(n21823), .B(n21825), .Z(n21824) );
  XOR U22696 ( .A(n21826), .B(n21827), .Z(n986) );
  AND U22697 ( .A(n21828), .B(n21829), .Z(n21826) );
  XNOR U22698 ( .A(n21827), .B(n21793), .Z(n21829) );
  XNOR U22699 ( .A(n21830), .B(n21831), .Z(n21793) );
  ANDN U22700 ( .B(n21832), .A(n21833), .Z(n21830) );
  XOR U22701 ( .A(n21831), .B(n21834), .Z(n21832) );
  XOR U22702 ( .A(n21827), .B(n21795), .Z(n21828) );
  XOR U22703 ( .A(n21835), .B(n21836), .Z(n21795) );
  AND U22704 ( .A(n990), .B(n21837), .Z(n21835) );
  XOR U22705 ( .A(n21838), .B(n21836), .Z(n21837) );
  XNOR U22706 ( .A(n21839), .B(n21840), .Z(n21827) );
  NAND U22707 ( .A(n21841), .B(n21842), .Z(n21840) );
  XOR U22708 ( .A(n21843), .B(n21819), .Z(n21842) );
  XOR U22709 ( .A(n21833), .B(n21834), .Z(n21819) );
  XOR U22710 ( .A(n21844), .B(n21845), .Z(n21834) );
  ANDN U22711 ( .B(n21846), .A(n21847), .Z(n21844) );
  XOR U22712 ( .A(n21845), .B(n21848), .Z(n21846) );
  XOR U22713 ( .A(n21849), .B(n21850), .Z(n21833) );
  XOR U22714 ( .A(n21851), .B(n21852), .Z(n21850) );
  ANDN U22715 ( .B(n21853), .A(n21854), .Z(n21851) );
  XOR U22716 ( .A(n21855), .B(n21852), .Z(n21853) );
  IV U22717 ( .A(n21831), .Z(n21849) );
  XOR U22718 ( .A(n21856), .B(n21857), .Z(n21831) );
  ANDN U22719 ( .B(n21858), .A(n21859), .Z(n21856) );
  XOR U22720 ( .A(n21857), .B(n21860), .Z(n21858) );
  IV U22721 ( .A(n21839), .Z(n21843) );
  XOR U22722 ( .A(n21839), .B(n21821), .Z(n21841) );
  XOR U22723 ( .A(n21861), .B(n21862), .Z(n21821) );
  AND U22724 ( .A(n990), .B(n21863), .Z(n21861) );
  XOR U22725 ( .A(n21864), .B(n21862), .Z(n21863) );
  NANDN U22726 ( .A(n21823), .B(n21825), .Z(n21839) );
  XOR U22727 ( .A(n21865), .B(n21866), .Z(n21825) );
  AND U22728 ( .A(n990), .B(n21867), .Z(n21865) );
  XOR U22729 ( .A(n21866), .B(n21868), .Z(n21867) );
  XOR U22730 ( .A(n21869), .B(n21870), .Z(n990) );
  AND U22731 ( .A(n21871), .B(n21872), .Z(n21869) );
  XNOR U22732 ( .A(n21870), .B(n21836), .Z(n21872) );
  XNOR U22733 ( .A(n21873), .B(n21874), .Z(n21836) );
  ANDN U22734 ( .B(n21875), .A(n21876), .Z(n21873) );
  XOR U22735 ( .A(n21874), .B(n21877), .Z(n21875) );
  XOR U22736 ( .A(n21870), .B(n21838), .Z(n21871) );
  XOR U22737 ( .A(n21878), .B(n21879), .Z(n21838) );
  AND U22738 ( .A(n994), .B(n21880), .Z(n21878) );
  XOR U22739 ( .A(n21881), .B(n21879), .Z(n21880) );
  XNOR U22740 ( .A(n21882), .B(n21883), .Z(n21870) );
  NAND U22741 ( .A(n21884), .B(n21885), .Z(n21883) );
  XOR U22742 ( .A(n21886), .B(n21862), .Z(n21885) );
  XOR U22743 ( .A(n21876), .B(n21877), .Z(n21862) );
  XOR U22744 ( .A(n21887), .B(n21888), .Z(n21877) );
  ANDN U22745 ( .B(n21889), .A(n21890), .Z(n21887) );
  XOR U22746 ( .A(n21888), .B(n21891), .Z(n21889) );
  XOR U22747 ( .A(n21892), .B(n21893), .Z(n21876) );
  XOR U22748 ( .A(n21894), .B(n21895), .Z(n21893) );
  ANDN U22749 ( .B(n21896), .A(n21897), .Z(n21894) );
  XOR U22750 ( .A(n21898), .B(n21895), .Z(n21896) );
  IV U22751 ( .A(n21874), .Z(n21892) );
  XOR U22752 ( .A(n21899), .B(n21900), .Z(n21874) );
  ANDN U22753 ( .B(n21901), .A(n21902), .Z(n21899) );
  XOR U22754 ( .A(n21900), .B(n21903), .Z(n21901) );
  IV U22755 ( .A(n21882), .Z(n21886) );
  XOR U22756 ( .A(n21882), .B(n21864), .Z(n21884) );
  XOR U22757 ( .A(n21904), .B(n21905), .Z(n21864) );
  AND U22758 ( .A(n994), .B(n21906), .Z(n21904) );
  XOR U22759 ( .A(n21907), .B(n21905), .Z(n21906) );
  NANDN U22760 ( .A(n21866), .B(n21868), .Z(n21882) );
  XOR U22761 ( .A(n21908), .B(n21909), .Z(n21868) );
  AND U22762 ( .A(n994), .B(n21910), .Z(n21908) );
  XOR U22763 ( .A(n21909), .B(n21911), .Z(n21910) );
  XOR U22764 ( .A(n21912), .B(n21913), .Z(n994) );
  AND U22765 ( .A(n21914), .B(n21915), .Z(n21912) );
  XNOR U22766 ( .A(n21913), .B(n21879), .Z(n21915) );
  XNOR U22767 ( .A(n21916), .B(n21917), .Z(n21879) );
  ANDN U22768 ( .B(n21918), .A(n21919), .Z(n21916) );
  XOR U22769 ( .A(n21917), .B(n21920), .Z(n21918) );
  XOR U22770 ( .A(n21913), .B(n21881), .Z(n21914) );
  XOR U22771 ( .A(n21921), .B(n21922), .Z(n21881) );
  AND U22772 ( .A(n998), .B(n21923), .Z(n21921) );
  XOR U22773 ( .A(n21924), .B(n21922), .Z(n21923) );
  XNOR U22774 ( .A(n21925), .B(n21926), .Z(n21913) );
  NAND U22775 ( .A(n21927), .B(n21928), .Z(n21926) );
  XOR U22776 ( .A(n21929), .B(n21905), .Z(n21928) );
  XOR U22777 ( .A(n21919), .B(n21920), .Z(n21905) );
  XOR U22778 ( .A(n21930), .B(n21931), .Z(n21920) );
  ANDN U22779 ( .B(n21932), .A(n21933), .Z(n21930) );
  XOR U22780 ( .A(n21931), .B(n21934), .Z(n21932) );
  XOR U22781 ( .A(n21935), .B(n21936), .Z(n21919) );
  XOR U22782 ( .A(n21937), .B(n21938), .Z(n21936) );
  ANDN U22783 ( .B(n21939), .A(n21940), .Z(n21937) );
  XOR U22784 ( .A(n21941), .B(n21938), .Z(n21939) );
  IV U22785 ( .A(n21917), .Z(n21935) );
  XOR U22786 ( .A(n21942), .B(n21943), .Z(n21917) );
  ANDN U22787 ( .B(n21944), .A(n21945), .Z(n21942) );
  XOR U22788 ( .A(n21943), .B(n21946), .Z(n21944) );
  IV U22789 ( .A(n21925), .Z(n21929) );
  XOR U22790 ( .A(n21925), .B(n21907), .Z(n21927) );
  XOR U22791 ( .A(n21947), .B(n21948), .Z(n21907) );
  AND U22792 ( .A(n998), .B(n21949), .Z(n21947) );
  XOR U22793 ( .A(n21950), .B(n21948), .Z(n21949) );
  NANDN U22794 ( .A(n21909), .B(n21911), .Z(n21925) );
  XOR U22795 ( .A(n21951), .B(n21952), .Z(n21911) );
  AND U22796 ( .A(n998), .B(n21953), .Z(n21951) );
  XOR U22797 ( .A(n21952), .B(n21954), .Z(n21953) );
  XOR U22798 ( .A(n21955), .B(n21956), .Z(n998) );
  AND U22799 ( .A(n21957), .B(n21958), .Z(n21955) );
  XNOR U22800 ( .A(n21956), .B(n21922), .Z(n21958) );
  XNOR U22801 ( .A(n21959), .B(n21960), .Z(n21922) );
  ANDN U22802 ( .B(n21961), .A(n21962), .Z(n21959) );
  XOR U22803 ( .A(n21960), .B(n21963), .Z(n21961) );
  XOR U22804 ( .A(n21956), .B(n21924), .Z(n21957) );
  XOR U22805 ( .A(n21964), .B(n21965), .Z(n21924) );
  AND U22806 ( .A(n1002), .B(n21966), .Z(n21964) );
  XOR U22807 ( .A(n21967), .B(n21965), .Z(n21966) );
  XNOR U22808 ( .A(n21968), .B(n21969), .Z(n21956) );
  NAND U22809 ( .A(n21970), .B(n21971), .Z(n21969) );
  XOR U22810 ( .A(n21972), .B(n21948), .Z(n21971) );
  XOR U22811 ( .A(n21962), .B(n21963), .Z(n21948) );
  XOR U22812 ( .A(n21973), .B(n21974), .Z(n21963) );
  ANDN U22813 ( .B(n21975), .A(n21976), .Z(n21973) );
  XOR U22814 ( .A(n21974), .B(n21977), .Z(n21975) );
  XOR U22815 ( .A(n21978), .B(n21979), .Z(n21962) );
  XOR U22816 ( .A(n21980), .B(n21981), .Z(n21979) );
  ANDN U22817 ( .B(n21982), .A(n21983), .Z(n21980) );
  XOR U22818 ( .A(n21984), .B(n21981), .Z(n21982) );
  IV U22819 ( .A(n21960), .Z(n21978) );
  XOR U22820 ( .A(n21985), .B(n21986), .Z(n21960) );
  ANDN U22821 ( .B(n21987), .A(n21988), .Z(n21985) );
  XOR U22822 ( .A(n21986), .B(n21989), .Z(n21987) );
  IV U22823 ( .A(n21968), .Z(n21972) );
  XOR U22824 ( .A(n21968), .B(n21950), .Z(n21970) );
  XOR U22825 ( .A(n21990), .B(n21991), .Z(n21950) );
  AND U22826 ( .A(n1002), .B(n21992), .Z(n21990) );
  XOR U22827 ( .A(n21993), .B(n21991), .Z(n21992) );
  NANDN U22828 ( .A(n21952), .B(n21954), .Z(n21968) );
  XOR U22829 ( .A(n21994), .B(n21995), .Z(n21954) );
  AND U22830 ( .A(n1002), .B(n21996), .Z(n21994) );
  XOR U22831 ( .A(n21995), .B(n21997), .Z(n21996) );
  XOR U22832 ( .A(n21998), .B(n21999), .Z(n1002) );
  AND U22833 ( .A(n22000), .B(n22001), .Z(n21998) );
  XNOR U22834 ( .A(n21999), .B(n21965), .Z(n22001) );
  XNOR U22835 ( .A(n22002), .B(n22003), .Z(n21965) );
  ANDN U22836 ( .B(n22004), .A(n22005), .Z(n22002) );
  XOR U22837 ( .A(n22003), .B(n22006), .Z(n22004) );
  XOR U22838 ( .A(n21999), .B(n21967), .Z(n22000) );
  XOR U22839 ( .A(n22007), .B(n22008), .Z(n21967) );
  AND U22840 ( .A(n1006), .B(n22009), .Z(n22007) );
  XOR U22841 ( .A(n22010), .B(n22008), .Z(n22009) );
  XNOR U22842 ( .A(n22011), .B(n22012), .Z(n21999) );
  NAND U22843 ( .A(n22013), .B(n22014), .Z(n22012) );
  XOR U22844 ( .A(n22015), .B(n21991), .Z(n22014) );
  XOR U22845 ( .A(n22005), .B(n22006), .Z(n21991) );
  XOR U22846 ( .A(n22016), .B(n22017), .Z(n22006) );
  ANDN U22847 ( .B(n22018), .A(n22019), .Z(n22016) );
  XOR U22848 ( .A(n22017), .B(n22020), .Z(n22018) );
  XOR U22849 ( .A(n22021), .B(n22022), .Z(n22005) );
  XOR U22850 ( .A(n22023), .B(n22024), .Z(n22022) );
  ANDN U22851 ( .B(n22025), .A(n22026), .Z(n22023) );
  XOR U22852 ( .A(n22027), .B(n22024), .Z(n22025) );
  IV U22853 ( .A(n22003), .Z(n22021) );
  XOR U22854 ( .A(n22028), .B(n22029), .Z(n22003) );
  ANDN U22855 ( .B(n22030), .A(n22031), .Z(n22028) );
  XOR U22856 ( .A(n22029), .B(n22032), .Z(n22030) );
  IV U22857 ( .A(n22011), .Z(n22015) );
  XOR U22858 ( .A(n22011), .B(n21993), .Z(n22013) );
  XOR U22859 ( .A(n22033), .B(n22034), .Z(n21993) );
  AND U22860 ( .A(n1006), .B(n22035), .Z(n22033) );
  XOR U22861 ( .A(n22036), .B(n22034), .Z(n22035) );
  NANDN U22862 ( .A(n21995), .B(n21997), .Z(n22011) );
  XOR U22863 ( .A(n22037), .B(n22038), .Z(n21997) );
  AND U22864 ( .A(n1006), .B(n22039), .Z(n22037) );
  XOR U22865 ( .A(n22038), .B(n22040), .Z(n22039) );
  XOR U22866 ( .A(n22041), .B(n22042), .Z(n1006) );
  AND U22867 ( .A(n22043), .B(n22044), .Z(n22041) );
  XNOR U22868 ( .A(n22042), .B(n22008), .Z(n22044) );
  XNOR U22869 ( .A(n22045), .B(n22046), .Z(n22008) );
  ANDN U22870 ( .B(n22047), .A(n22048), .Z(n22045) );
  XOR U22871 ( .A(n22046), .B(n22049), .Z(n22047) );
  XOR U22872 ( .A(n22042), .B(n22010), .Z(n22043) );
  XOR U22873 ( .A(n22050), .B(n22051), .Z(n22010) );
  AND U22874 ( .A(n1010), .B(n22052), .Z(n22050) );
  XOR U22875 ( .A(n22053), .B(n22051), .Z(n22052) );
  XNOR U22876 ( .A(n22054), .B(n22055), .Z(n22042) );
  NAND U22877 ( .A(n22056), .B(n22057), .Z(n22055) );
  XOR U22878 ( .A(n22058), .B(n22034), .Z(n22057) );
  XOR U22879 ( .A(n22048), .B(n22049), .Z(n22034) );
  XOR U22880 ( .A(n22059), .B(n22060), .Z(n22049) );
  ANDN U22881 ( .B(n22061), .A(n22062), .Z(n22059) );
  XOR U22882 ( .A(n22060), .B(n22063), .Z(n22061) );
  XOR U22883 ( .A(n22064), .B(n22065), .Z(n22048) );
  XOR U22884 ( .A(n22066), .B(n22067), .Z(n22065) );
  ANDN U22885 ( .B(n22068), .A(n22069), .Z(n22066) );
  XOR U22886 ( .A(n22070), .B(n22067), .Z(n22068) );
  IV U22887 ( .A(n22046), .Z(n22064) );
  XOR U22888 ( .A(n22071), .B(n22072), .Z(n22046) );
  ANDN U22889 ( .B(n22073), .A(n22074), .Z(n22071) );
  XOR U22890 ( .A(n22072), .B(n22075), .Z(n22073) );
  IV U22891 ( .A(n22054), .Z(n22058) );
  XOR U22892 ( .A(n22054), .B(n22036), .Z(n22056) );
  XOR U22893 ( .A(n22076), .B(n22077), .Z(n22036) );
  AND U22894 ( .A(n1010), .B(n22078), .Z(n22076) );
  XOR U22895 ( .A(n22079), .B(n22077), .Z(n22078) );
  NANDN U22896 ( .A(n22038), .B(n22040), .Z(n22054) );
  XOR U22897 ( .A(n22080), .B(n22081), .Z(n22040) );
  AND U22898 ( .A(n1010), .B(n22082), .Z(n22080) );
  XOR U22899 ( .A(n22081), .B(n22083), .Z(n22082) );
  XOR U22900 ( .A(n22084), .B(n22085), .Z(n1010) );
  AND U22901 ( .A(n22086), .B(n22087), .Z(n22084) );
  XNOR U22902 ( .A(n22085), .B(n22051), .Z(n22087) );
  XNOR U22903 ( .A(n22088), .B(n22089), .Z(n22051) );
  ANDN U22904 ( .B(n22090), .A(n22091), .Z(n22088) );
  XOR U22905 ( .A(n22089), .B(n22092), .Z(n22090) );
  XOR U22906 ( .A(n22085), .B(n22053), .Z(n22086) );
  XOR U22907 ( .A(n22093), .B(n22094), .Z(n22053) );
  AND U22908 ( .A(n1014), .B(n22095), .Z(n22093) );
  XOR U22909 ( .A(n22096), .B(n22094), .Z(n22095) );
  XNOR U22910 ( .A(n22097), .B(n22098), .Z(n22085) );
  NAND U22911 ( .A(n22099), .B(n22100), .Z(n22098) );
  XOR U22912 ( .A(n22101), .B(n22077), .Z(n22100) );
  XOR U22913 ( .A(n22091), .B(n22092), .Z(n22077) );
  XOR U22914 ( .A(n22102), .B(n22103), .Z(n22092) );
  ANDN U22915 ( .B(n22104), .A(n22105), .Z(n22102) );
  XOR U22916 ( .A(n22103), .B(n22106), .Z(n22104) );
  XOR U22917 ( .A(n22107), .B(n22108), .Z(n22091) );
  XOR U22918 ( .A(n22109), .B(n22110), .Z(n22108) );
  ANDN U22919 ( .B(n22111), .A(n22112), .Z(n22109) );
  XOR U22920 ( .A(n22113), .B(n22110), .Z(n22111) );
  IV U22921 ( .A(n22089), .Z(n22107) );
  XOR U22922 ( .A(n22114), .B(n22115), .Z(n22089) );
  ANDN U22923 ( .B(n22116), .A(n22117), .Z(n22114) );
  XOR U22924 ( .A(n22115), .B(n22118), .Z(n22116) );
  IV U22925 ( .A(n22097), .Z(n22101) );
  XOR U22926 ( .A(n22097), .B(n22079), .Z(n22099) );
  XOR U22927 ( .A(n22119), .B(n22120), .Z(n22079) );
  AND U22928 ( .A(n1014), .B(n22121), .Z(n22119) );
  XOR U22929 ( .A(n22122), .B(n22120), .Z(n22121) );
  NANDN U22930 ( .A(n22081), .B(n22083), .Z(n22097) );
  XOR U22931 ( .A(n22123), .B(n22124), .Z(n22083) );
  AND U22932 ( .A(n1014), .B(n22125), .Z(n22123) );
  XOR U22933 ( .A(n22124), .B(n22126), .Z(n22125) );
  XOR U22934 ( .A(n22127), .B(n22128), .Z(n1014) );
  AND U22935 ( .A(n22129), .B(n22130), .Z(n22127) );
  XNOR U22936 ( .A(n22128), .B(n22094), .Z(n22130) );
  XNOR U22937 ( .A(n22131), .B(n22132), .Z(n22094) );
  ANDN U22938 ( .B(n22133), .A(n22134), .Z(n22131) );
  XOR U22939 ( .A(n22132), .B(n22135), .Z(n22133) );
  XOR U22940 ( .A(n22128), .B(n22096), .Z(n22129) );
  XOR U22941 ( .A(n22136), .B(n22137), .Z(n22096) );
  AND U22942 ( .A(n1018), .B(n22138), .Z(n22136) );
  XOR U22943 ( .A(n22139), .B(n22137), .Z(n22138) );
  XNOR U22944 ( .A(n22140), .B(n22141), .Z(n22128) );
  NAND U22945 ( .A(n22142), .B(n22143), .Z(n22141) );
  XOR U22946 ( .A(n22144), .B(n22120), .Z(n22143) );
  XOR U22947 ( .A(n22134), .B(n22135), .Z(n22120) );
  XOR U22948 ( .A(n22145), .B(n22146), .Z(n22135) );
  ANDN U22949 ( .B(n22147), .A(n22148), .Z(n22145) );
  XOR U22950 ( .A(n22146), .B(n22149), .Z(n22147) );
  XOR U22951 ( .A(n22150), .B(n22151), .Z(n22134) );
  XOR U22952 ( .A(n22152), .B(n22153), .Z(n22151) );
  ANDN U22953 ( .B(n22154), .A(n22155), .Z(n22152) );
  XOR U22954 ( .A(n22156), .B(n22153), .Z(n22154) );
  IV U22955 ( .A(n22132), .Z(n22150) );
  XOR U22956 ( .A(n22157), .B(n22158), .Z(n22132) );
  ANDN U22957 ( .B(n22159), .A(n22160), .Z(n22157) );
  XOR U22958 ( .A(n22158), .B(n22161), .Z(n22159) );
  IV U22959 ( .A(n22140), .Z(n22144) );
  XOR U22960 ( .A(n22140), .B(n22122), .Z(n22142) );
  XOR U22961 ( .A(n22162), .B(n22163), .Z(n22122) );
  AND U22962 ( .A(n1018), .B(n22164), .Z(n22162) );
  XOR U22963 ( .A(n22165), .B(n22163), .Z(n22164) );
  NANDN U22964 ( .A(n22124), .B(n22126), .Z(n22140) );
  XOR U22965 ( .A(n22166), .B(n22167), .Z(n22126) );
  AND U22966 ( .A(n1018), .B(n22168), .Z(n22166) );
  XOR U22967 ( .A(n22167), .B(n22169), .Z(n22168) );
  XOR U22968 ( .A(n22170), .B(n22171), .Z(n1018) );
  AND U22969 ( .A(n22172), .B(n22173), .Z(n22170) );
  XNOR U22970 ( .A(n22171), .B(n22137), .Z(n22173) );
  XNOR U22971 ( .A(n22174), .B(n22175), .Z(n22137) );
  ANDN U22972 ( .B(n22176), .A(n22177), .Z(n22174) );
  XOR U22973 ( .A(n22175), .B(n22178), .Z(n22176) );
  XOR U22974 ( .A(n22171), .B(n22139), .Z(n22172) );
  XOR U22975 ( .A(n22179), .B(n22180), .Z(n22139) );
  AND U22976 ( .A(n1022), .B(n22181), .Z(n22179) );
  XOR U22977 ( .A(n22182), .B(n22180), .Z(n22181) );
  XNOR U22978 ( .A(n22183), .B(n22184), .Z(n22171) );
  NAND U22979 ( .A(n22185), .B(n22186), .Z(n22184) );
  XOR U22980 ( .A(n22187), .B(n22163), .Z(n22186) );
  XOR U22981 ( .A(n22177), .B(n22178), .Z(n22163) );
  XOR U22982 ( .A(n22188), .B(n22189), .Z(n22178) );
  ANDN U22983 ( .B(n22190), .A(n22191), .Z(n22188) );
  XOR U22984 ( .A(n22189), .B(n22192), .Z(n22190) );
  XOR U22985 ( .A(n22193), .B(n22194), .Z(n22177) );
  XOR U22986 ( .A(n22195), .B(n22196), .Z(n22194) );
  ANDN U22987 ( .B(n22197), .A(n22198), .Z(n22195) );
  XOR U22988 ( .A(n22199), .B(n22196), .Z(n22197) );
  IV U22989 ( .A(n22175), .Z(n22193) );
  XOR U22990 ( .A(n22200), .B(n22201), .Z(n22175) );
  ANDN U22991 ( .B(n22202), .A(n22203), .Z(n22200) );
  XOR U22992 ( .A(n22201), .B(n22204), .Z(n22202) );
  IV U22993 ( .A(n22183), .Z(n22187) );
  XOR U22994 ( .A(n22183), .B(n22165), .Z(n22185) );
  XOR U22995 ( .A(n22205), .B(n22206), .Z(n22165) );
  AND U22996 ( .A(n1022), .B(n22207), .Z(n22205) );
  XOR U22997 ( .A(n22208), .B(n22206), .Z(n22207) );
  NANDN U22998 ( .A(n22167), .B(n22169), .Z(n22183) );
  XOR U22999 ( .A(n22209), .B(n22210), .Z(n22169) );
  AND U23000 ( .A(n1022), .B(n22211), .Z(n22209) );
  XOR U23001 ( .A(n22210), .B(n22212), .Z(n22211) );
  XOR U23002 ( .A(n22213), .B(n22214), .Z(n1022) );
  AND U23003 ( .A(n22215), .B(n22216), .Z(n22213) );
  XNOR U23004 ( .A(n22214), .B(n22180), .Z(n22216) );
  XNOR U23005 ( .A(n22217), .B(n22218), .Z(n22180) );
  ANDN U23006 ( .B(n22219), .A(n22220), .Z(n22217) );
  XOR U23007 ( .A(n22218), .B(n22221), .Z(n22219) );
  XOR U23008 ( .A(n22214), .B(n22182), .Z(n22215) );
  XOR U23009 ( .A(n22222), .B(n22223), .Z(n22182) );
  AND U23010 ( .A(n1026), .B(n22224), .Z(n22222) );
  XOR U23011 ( .A(n22225), .B(n22223), .Z(n22224) );
  XNOR U23012 ( .A(n22226), .B(n22227), .Z(n22214) );
  NAND U23013 ( .A(n22228), .B(n22229), .Z(n22227) );
  XOR U23014 ( .A(n22230), .B(n22206), .Z(n22229) );
  XOR U23015 ( .A(n22220), .B(n22221), .Z(n22206) );
  XOR U23016 ( .A(n22231), .B(n22232), .Z(n22221) );
  ANDN U23017 ( .B(n22233), .A(n22234), .Z(n22231) );
  XOR U23018 ( .A(n22232), .B(n22235), .Z(n22233) );
  XOR U23019 ( .A(n22236), .B(n22237), .Z(n22220) );
  XOR U23020 ( .A(n22238), .B(n22239), .Z(n22237) );
  ANDN U23021 ( .B(n22240), .A(n22241), .Z(n22238) );
  XOR U23022 ( .A(n22242), .B(n22239), .Z(n22240) );
  IV U23023 ( .A(n22218), .Z(n22236) );
  XOR U23024 ( .A(n22243), .B(n22244), .Z(n22218) );
  ANDN U23025 ( .B(n22245), .A(n22246), .Z(n22243) );
  XOR U23026 ( .A(n22244), .B(n22247), .Z(n22245) );
  IV U23027 ( .A(n22226), .Z(n22230) );
  XOR U23028 ( .A(n22226), .B(n22208), .Z(n22228) );
  XOR U23029 ( .A(n22248), .B(n22249), .Z(n22208) );
  AND U23030 ( .A(n1026), .B(n22250), .Z(n22248) );
  XOR U23031 ( .A(n22251), .B(n22249), .Z(n22250) );
  NANDN U23032 ( .A(n22210), .B(n22212), .Z(n22226) );
  XOR U23033 ( .A(n22252), .B(n22253), .Z(n22212) );
  AND U23034 ( .A(n1026), .B(n22254), .Z(n22252) );
  XOR U23035 ( .A(n22253), .B(n22255), .Z(n22254) );
  XOR U23036 ( .A(n22256), .B(n22257), .Z(n1026) );
  AND U23037 ( .A(n22258), .B(n22259), .Z(n22256) );
  XNOR U23038 ( .A(n22257), .B(n22223), .Z(n22259) );
  XNOR U23039 ( .A(n22260), .B(n22261), .Z(n22223) );
  ANDN U23040 ( .B(n22262), .A(n22263), .Z(n22260) );
  XOR U23041 ( .A(n22261), .B(n22264), .Z(n22262) );
  XOR U23042 ( .A(n22257), .B(n22225), .Z(n22258) );
  XOR U23043 ( .A(n22265), .B(n22266), .Z(n22225) );
  AND U23044 ( .A(n1030), .B(n22267), .Z(n22265) );
  XOR U23045 ( .A(n22268), .B(n22266), .Z(n22267) );
  XNOR U23046 ( .A(n22269), .B(n22270), .Z(n22257) );
  NAND U23047 ( .A(n22271), .B(n22272), .Z(n22270) );
  XOR U23048 ( .A(n22273), .B(n22249), .Z(n22272) );
  XOR U23049 ( .A(n22263), .B(n22264), .Z(n22249) );
  XOR U23050 ( .A(n22274), .B(n22275), .Z(n22264) );
  ANDN U23051 ( .B(n22276), .A(n22277), .Z(n22274) );
  XOR U23052 ( .A(n22275), .B(n22278), .Z(n22276) );
  XOR U23053 ( .A(n22279), .B(n22280), .Z(n22263) );
  XOR U23054 ( .A(n22281), .B(n22282), .Z(n22280) );
  ANDN U23055 ( .B(n22283), .A(n22284), .Z(n22281) );
  XOR U23056 ( .A(n22285), .B(n22282), .Z(n22283) );
  IV U23057 ( .A(n22261), .Z(n22279) );
  XOR U23058 ( .A(n22286), .B(n22287), .Z(n22261) );
  ANDN U23059 ( .B(n22288), .A(n22289), .Z(n22286) );
  XOR U23060 ( .A(n22287), .B(n22290), .Z(n22288) );
  IV U23061 ( .A(n22269), .Z(n22273) );
  XOR U23062 ( .A(n22269), .B(n22251), .Z(n22271) );
  XOR U23063 ( .A(n22291), .B(n22292), .Z(n22251) );
  AND U23064 ( .A(n1030), .B(n22293), .Z(n22291) );
  XOR U23065 ( .A(n22294), .B(n22292), .Z(n22293) );
  NANDN U23066 ( .A(n22253), .B(n22255), .Z(n22269) );
  XOR U23067 ( .A(n22295), .B(n22296), .Z(n22255) );
  AND U23068 ( .A(n1030), .B(n22297), .Z(n22295) );
  XOR U23069 ( .A(n22296), .B(n22298), .Z(n22297) );
  XOR U23070 ( .A(n22299), .B(n22300), .Z(n1030) );
  AND U23071 ( .A(n22301), .B(n22302), .Z(n22299) );
  XNOR U23072 ( .A(n22300), .B(n22266), .Z(n22302) );
  XNOR U23073 ( .A(n22303), .B(n22304), .Z(n22266) );
  ANDN U23074 ( .B(n22305), .A(n22306), .Z(n22303) );
  XOR U23075 ( .A(n22304), .B(n22307), .Z(n22305) );
  XOR U23076 ( .A(n22300), .B(n22268), .Z(n22301) );
  XOR U23077 ( .A(n22308), .B(n22309), .Z(n22268) );
  AND U23078 ( .A(n1034), .B(n22310), .Z(n22308) );
  XOR U23079 ( .A(n22311), .B(n22309), .Z(n22310) );
  XNOR U23080 ( .A(n22312), .B(n22313), .Z(n22300) );
  NAND U23081 ( .A(n22314), .B(n22315), .Z(n22313) );
  XOR U23082 ( .A(n22316), .B(n22292), .Z(n22315) );
  XOR U23083 ( .A(n22306), .B(n22307), .Z(n22292) );
  XOR U23084 ( .A(n22317), .B(n22318), .Z(n22307) );
  ANDN U23085 ( .B(n22319), .A(n22320), .Z(n22317) );
  XOR U23086 ( .A(n22318), .B(n22321), .Z(n22319) );
  XOR U23087 ( .A(n22322), .B(n22323), .Z(n22306) );
  XOR U23088 ( .A(n22324), .B(n22325), .Z(n22323) );
  ANDN U23089 ( .B(n22326), .A(n22327), .Z(n22324) );
  XOR U23090 ( .A(n22328), .B(n22325), .Z(n22326) );
  IV U23091 ( .A(n22304), .Z(n22322) );
  XOR U23092 ( .A(n22329), .B(n22330), .Z(n22304) );
  ANDN U23093 ( .B(n22331), .A(n22332), .Z(n22329) );
  XOR U23094 ( .A(n22330), .B(n22333), .Z(n22331) );
  IV U23095 ( .A(n22312), .Z(n22316) );
  XOR U23096 ( .A(n22312), .B(n22294), .Z(n22314) );
  XOR U23097 ( .A(n22334), .B(n22335), .Z(n22294) );
  AND U23098 ( .A(n1034), .B(n22336), .Z(n22334) );
  XOR U23099 ( .A(n22337), .B(n22335), .Z(n22336) );
  NANDN U23100 ( .A(n22296), .B(n22298), .Z(n22312) );
  XOR U23101 ( .A(n22338), .B(n22339), .Z(n22298) );
  AND U23102 ( .A(n1034), .B(n22340), .Z(n22338) );
  XOR U23103 ( .A(n22339), .B(n22341), .Z(n22340) );
  XOR U23104 ( .A(n22342), .B(n22343), .Z(n1034) );
  AND U23105 ( .A(n22344), .B(n22345), .Z(n22342) );
  XNOR U23106 ( .A(n22343), .B(n22309), .Z(n22345) );
  XNOR U23107 ( .A(n22346), .B(n22347), .Z(n22309) );
  ANDN U23108 ( .B(n22348), .A(n22349), .Z(n22346) );
  XOR U23109 ( .A(n22347), .B(n22350), .Z(n22348) );
  XOR U23110 ( .A(n22343), .B(n22311), .Z(n22344) );
  XOR U23111 ( .A(n22351), .B(n22352), .Z(n22311) );
  AND U23112 ( .A(n1038), .B(n22353), .Z(n22351) );
  XOR U23113 ( .A(n22354), .B(n22352), .Z(n22353) );
  XNOR U23114 ( .A(n22355), .B(n22356), .Z(n22343) );
  NAND U23115 ( .A(n22357), .B(n22358), .Z(n22356) );
  XOR U23116 ( .A(n22359), .B(n22335), .Z(n22358) );
  XOR U23117 ( .A(n22349), .B(n22350), .Z(n22335) );
  XOR U23118 ( .A(n22360), .B(n22361), .Z(n22350) );
  ANDN U23119 ( .B(n22362), .A(n22363), .Z(n22360) );
  XOR U23120 ( .A(n22361), .B(n22364), .Z(n22362) );
  XOR U23121 ( .A(n22365), .B(n22366), .Z(n22349) );
  XOR U23122 ( .A(n22367), .B(n22368), .Z(n22366) );
  ANDN U23123 ( .B(n22369), .A(n22370), .Z(n22367) );
  XOR U23124 ( .A(n22371), .B(n22368), .Z(n22369) );
  IV U23125 ( .A(n22347), .Z(n22365) );
  XOR U23126 ( .A(n22372), .B(n22373), .Z(n22347) );
  ANDN U23127 ( .B(n22374), .A(n22375), .Z(n22372) );
  XOR U23128 ( .A(n22373), .B(n22376), .Z(n22374) );
  IV U23129 ( .A(n22355), .Z(n22359) );
  XOR U23130 ( .A(n22355), .B(n22337), .Z(n22357) );
  XOR U23131 ( .A(n22377), .B(n22378), .Z(n22337) );
  AND U23132 ( .A(n1038), .B(n22379), .Z(n22377) );
  XOR U23133 ( .A(n22380), .B(n22378), .Z(n22379) );
  NANDN U23134 ( .A(n22339), .B(n22341), .Z(n22355) );
  XOR U23135 ( .A(n22381), .B(n22382), .Z(n22341) );
  AND U23136 ( .A(n1038), .B(n22383), .Z(n22381) );
  XOR U23137 ( .A(n22382), .B(n22384), .Z(n22383) );
  XOR U23138 ( .A(n22385), .B(n22386), .Z(n1038) );
  AND U23139 ( .A(n22387), .B(n22388), .Z(n22385) );
  XNOR U23140 ( .A(n22386), .B(n22352), .Z(n22388) );
  XNOR U23141 ( .A(n22389), .B(n22390), .Z(n22352) );
  ANDN U23142 ( .B(n22391), .A(n22392), .Z(n22389) );
  XOR U23143 ( .A(n22390), .B(n22393), .Z(n22391) );
  XOR U23144 ( .A(n22386), .B(n22354), .Z(n22387) );
  XOR U23145 ( .A(n22394), .B(n22395), .Z(n22354) );
  AND U23146 ( .A(n1042), .B(n22396), .Z(n22394) );
  XOR U23147 ( .A(n22397), .B(n22395), .Z(n22396) );
  XNOR U23148 ( .A(n22398), .B(n22399), .Z(n22386) );
  NAND U23149 ( .A(n22400), .B(n22401), .Z(n22399) );
  XOR U23150 ( .A(n22402), .B(n22378), .Z(n22401) );
  XOR U23151 ( .A(n22392), .B(n22393), .Z(n22378) );
  XOR U23152 ( .A(n22403), .B(n22404), .Z(n22393) );
  ANDN U23153 ( .B(n22405), .A(n22406), .Z(n22403) );
  XOR U23154 ( .A(n22404), .B(n22407), .Z(n22405) );
  XOR U23155 ( .A(n22408), .B(n22409), .Z(n22392) );
  XOR U23156 ( .A(n22410), .B(n22411), .Z(n22409) );
  ANDN U23157 ( .B(n22412), .A(n22413), .Z(n22410) );
  XOR U23158 ( .A(n22414), .B(n22411), .Z(n22412) );
  IV U23159 ( .A(n22390), .Z(n22408) );
  XOR U23160 ( .A(n22415), .B(n22416), .Z(n22390) );
  ANDN U23161 ( .B(n22417), .A(n22418), .Z(n22415) );
  XOR U23162 ( .A(n22416), .B(n22419), .Z(n22417) );
  IV U23163 ( .A(n22398), .Z(n22402) );
  XOR U23164 ( .A(n22398), .B(n22380), .Z(n22400) );
  XOR U23165 ( .A(n22420), .B(n22421), .Z(n22380) );
  AND U23166 ( .A(n1042), .B(n22422), .Z(n22420) );
  XOR U23167 ( .A(n22423), .B(n22421), .Z(n22422) );
  NANDN U23168 ( .A(n22382), .B(n22384), .Z(n22398) );
  XOR U23169 ( .A(n22424), .B(n22425), .Z(n22384) );
  AND U23170 ( .A(n1042), .B(n22426), .Z(n22424) );
  XOR U23171 ( .A(n22425), .B(n22427), .Z(n22426) );
  XOR U23172 ( .A(n22428), .B(n22429), .Z(n1042) );
  AND U23173 ( .A(n22430), .B(n22431), .Z(n22428) );
  XNOR U23174 ( .A(n22429), .B(n22395), .Z(n22431) );
  XNOR U23175 ( .A(n22432), .B(n22433), .Z(n22395) );
  ANDN U23176 ( .B(n22434), .A(n22435), .Z(n22432) );
  XOR U23177 ( .A(n22433), .B(n22436), .Z(n22434) );
  XOR U23178 ( .A(n22429), .B(n22397), .Z(n22430) );
  XOR U23179 ( .A(n22437), .B(n22438), .Z(n22397) );
  AND U23180 ( .A(n1046), .B(n22439), .Z(n22437) );
  XOR U23181 ( .A(n22440), .B(n22438), .Z(n22439) );
  XNOR U23182 ( .A(n22441), .B(n22442), .Z(n22429) );
  NAND U23183 ( .A(n22443), .B(n22444), .Z(n22442) );
  XOR U23184 ( .A(n22445), .B(n22421), .Z(n22444) );
  XOR U23185 ( .A(n22435), .B(n22436), .Z(n22421) );
  XOR U23186 ( .A(n22446), .B(n22447), .Z(n22436) );
  ANDN U23187 ( .B(n22448), .A(n22449), .Z(n22446) );
  XOR U23188 ( .A(n22447), .B(n22450), .Z(n22448) );
  XOR U23189 ( .A(n22451), .B(n22452), .Z(n22435) );
  XOR U23190 ( .A(n22453), .B(n22454), .Z(n22452) );
  ANDN U23191 ( .B(n22455), .A(n22456), .Z(n22453) );
  XOR U23192 ( .A(n22457), .B(n22454), .Z(n22455) );
  IV U23193 ( .A(n22433), .Z(n22451) );
  XOR U23194 ( .A(n22458), .B(n22459), .Z(n22433) );
  ANDN U23195 ( .B(n22460), .A(n22461), .Z(n22458) );
  XOR U23196 ( .A(n22459), .B(n22462), .Z(n22460) );
  IV U23197 ( .A(n22441), .Z(n22445) );
  XOR U23198 ( .A(n22441), .B(n22423), .Z(n22443) );
  XOR U23199 ( .A(n22463), .B(n22464), .Z(n22423) );
  AND U23200 ( .A(n1046), .B(n22465), .Z(n22463) );
  XOR U23201 ( .A(n22466), .B(n22464), .Z(n22465) );
  NANDN U23202 ( .A(n22425), .B(n22427), .Z(n22441) );
  XOR U23203 ( .A(n22467), .B(n22468), .Z(n22427) );
  AND U23204 ( .A(n1046), .B(n22469), .Z(n22467) );
  XOR U23205 ( .A(n22468), .B(n22470), .Z(n22469) );
  XOR U23206 ( .A(n22471), .B(n22472), .Z(n1046) );
  AND U23207 ( .A(n22473), .B(n22474), .Z(n22471) );
  XNOR U23208 ( .A(n22472), .B(n22438), .Z(n22474) );
  XNOR U23209 ( .A(n22475), .B(n22476), .Z(n22438) );
  ANDN U23210 ( .B(n22477), .A(n22478), .Z(n22475) );
  XOR U23211 ( .A(n22476), .B(n22479), .Z(n22477) );
  XOR U23212 ( .A(n22472), .B(n22440), .Z(n22473) );
  XOR U23213 ( .A(n22480), .B(n22481), .Z(n22440) );
  AND U23214 ( .A(n1050), .B(n22482), .Z(n22480) );
  XOR U23215 ( .A(n22483), .B(n22481), .Z(n22482) );
  XNOR U23216 ( .A(n22484), .B(n22485), .Z(n22472) );
  NAND U23217 ( .A(n22486), .B(n22487), .Z(n22485) );
  XOR U23218 ( .A(n22488), .B(n22464), .Z(n22487) );
  XOR U23219 ( .A(n22478), .B(n22479), .Z(n22464) );
  XOR U23220 ( .A(n22489), .B(n22490), .Z(n22479) );
  ANDN U23221 ( .B(n22491), .A(n22492), .Z(n22489) );
  XOR U23222 ( .A(n22490), .B(n22493), .Z(n22491) );
  XOR U23223 ( .A(n22494), .B(n22495), .Z(n22478) );
  XOR U23224 ( .A(n22496), .B(n22497), .Z(n22495) );
  ANDN U23225 ( .B(n22498), .A(n22499), .Z(n22496) );
  XOR U23226 ( .A(n22500), .B(n22497), .Z(n22498) );
  IV U23227 ( .A(n22476), .Z(n22494) );
  XOR U23228 ( .A(n22501), .B(n22502), .Z(n22476) );
  ANDN U23229 ( .B(n22503), .A(n22504), .Z(n22501) );
  XOR U23230 ( .A(n22502), .B(n22505), .Z(n22503) );
  IV U23231 ( .A(n22484), .Z(n22488) );
  XOR U23232 ( .A(n22484), .B(n22466), .Z(n22486) );
  XOR U23233 ( .A(n22506), .B(n22507), .Z(n22466) );
  AND U23234 ( .A(n1050), .B(n22508), .Z(n22506) );
  XOR U23235 ( .A(n22509), .B(n22507), .Z(n22508) );
  NANDN U23236 ( .A(n22468), .B(n22470), .Z(n22484) );
  XOR U23237 ( .A(n22510), .B(n22511), .Z(n22470) );
  AND U23238 ( .A(n1050), .B(n22512), .Z(n22510) );
  XOR U23239 ( .A(n22511), .B(n22513), .Z(n22512) );
  XOR U23240 ( .A(n22514), .B(n22515), .Z(n1050) );
  AND U23241 ( .A(n22516), .B(n22517), .Z(n22514) );
  XNOR U23242 ( .A(n22515), .B(n22481), .Z(n22517) );
  XNOR U23243 ( .A(n22518), .B(n22519), .Z(n22481) );
  ANDN U23244 ( .B(n22520), .A(n22521), .Z(n22518) );
  XOR U23245 ( .A(n22519), .B(n22522), .Z(n22520) );
  XOR U23246 ( .A(n22515), .B(n22483), .Z(n22516) );
  XOR U23247 ( .A(n22523), .B(n22524), .Z(n22483) );
  AND U23248 ( .A(n1054), .B(n22525), .Z(n22523) );
  XOR U23249 ( .A(n22526), .B(n22524), .Z(n22525) );
  XNOR U23250 ( .A(n22527), .B(n22528), .Z(n22515) );
  NAND U23251 ( .A(n22529), .B(n22530), .Z(n22528) );
  XOR U23252 ( .A(n22531), .B(n22507), .Z(n22530) );
  XOR U23253 ( .A(n22521), .B(n22522), .Z(n22507) );
  XOR U23254 ( .A(n22532), .B(n22533), .Z(n22522) );
  ANDN U23255 ( .B(n22534), .A(n22535), .Z(n22532) );
  XOR U23256 ( .A(n22533), .B(n22536), .Z(n22534) );
  XOR U23257 ( .A(n22537), .B(n22538), .Z(n22521) );
  XOR U23258 ( .A(n22539), .B(n22540), .Z(n22538) );
  ANDN U23259 ( .B(n22541), .A(n22542), .Z(n22539) );
  XOR U23260 ( .A(n22543), .B(n22540), .Z(n22541) );
  IV U23261 ( .A(n22519), .Z(n22537) );
  XOR U23262 ( .A(n22544), .B(n22545), .Z(n22519) );
  ANDN U23263 ( .B(n22546), .A(n22547), .Z(n22544) );
  XOR U23264 ( .A(n22545), .B(n22548), .Z(n22546) );
  IV U23265 ( .A(n22527), .Z(n22531) );
  XOR U23266 ( .A(n22527), .B(n22509), .Z(n22529) );
  XOR U23267 ( .A(n22549), .B(n22550), .Z(n22509) );
  AND U23268 ( .A(n1054), .B(n22551), .Z(n22549) );
  XOR U23269 ( .A(n22552), .B(n22550), .Z(n22551) );
  NANDN U23270 ( .A(n22511), .B(n22513), .Z(n22527) );
  XOR U23271 ( .A(n22553), .B(n22554), .Z(n22513) );
  AND U23272 ( .A(n1054), .B(n22555), .Z(n22553) );
  XOR U23273 ( .A(n22554), .B(n22556), .Z(n22555) );
  XOR U23274 ( .A(n22557), .B(n22558), .Z(n1054) );
  AND U23275 ( .A(n22559), .B(n22560), .Z(n22557) );
  XNOR U23276 ( .A(n22558), .B(n22524), .Z(n22560) );
  XNOR U23277 ( .A(n22561), .B(n22562), .Z(n22524) );
  ANDN U23278 ( .B(n22563), .A(n22564), .Z(n22561) );
  XOR U23279 ( .A(n22562), .B(n22565), .Z(n22563) );
  XOR U23280 ( .A(n22558), .B(n22526), .Z(n22559) );
  XOR U23281 ( .A(n22566), .B(n22567), .Z(n22526) );
  AND U23282 ( .A(n1058), .B(n22568), .Z(n22566) );
  XOR U23283 ( .A(n22569), .B(n22567), .Z(n22568) );
  XNOR U23284 ( .A(n22570), .B(n22571), .Z(n22558) );
  NAND U23285 ( .A(n22572), .B(n22573), .Z(n22571) );
  XOR U23286 ( .A(n22574), .B(n22550), .Z(n22573) );
  XOR U23287 ( .A(n22564), .B(n22565), .Z(n22550) );
  XOR U23288 ( .A(n22575), .B(n22576), .Z(n22565) );
  ANDN U23289 ( .B(n22577), .A(n22578), .Z(n22575) );
  XOR U23290 ( .A(n22576), .B(n22579), .Z(n22577) );
  XOR U23291 ( .A(n22580), .B(n22581), .Z(n22564) );
  XOR U23292 ( .A(n22582), .B(n22583), .Z(n22581) );
  ANDN U23293 ( .B(n22584), .A(n22585), .Z(n22582) );
  XOR U23294 ( .A(n22586), .B(n22583), .Z(n22584) );
  IV U23295 ( .A(n22562), .Z(n22580) );
  XOR U23296 ( .A(n22587), .B(n22588), .Z(n22562) );
  ANDN U23297 ( .B(n22589), .A(n22590), .Z(n22587) );
  XOR U23298 ( .A(n22588), .B(n22591), .Z(n22589) );
  IV U23299 ( .A(n22570), .Z(n22574) );
  XOR U23300 ( .A(n22570), .B(n22552), .Z(n22572) );
  XOR U23301 ( .A(n22592), .B(n22593), .Z(n22552) );
  AND U23302 ( .A(n1058), .B(n22594), .Z(n22592) );
  XOR U23303 ( .A(n22595), .B(n22593), .Z(n22594) );
  NANDN U23304 ( .A(n22554), .B(n22556), .Z(n22570) );
  XOR U23305 ( .A(n22596), .B(n22597), .Z(n22556) );
  AND U23306 ( .A(n1058), .B(n22598), .Z(n22596) );
  XOR U23307 ( .A(n22597), .B(n22599), .Z(n22598) );
  XOR U23308 ( .A(n22600), .B(n22601), .Z(n1058) );
  AND U23309 ( .A(n22602), .B(n22603), .Z(n22600) );
  XNOR U23310 ( .A(n22601), .B(n22567), .Z(n22603) );
  XNOR U23311 ( .A(n22604), .B(n22605), .Z(n22567) );
  ANDN U23312 ( .B(n22606), .A(n22607), .Z(n22604) );
  XOR U23313 ( .A(n22605), .B(n22608), .Z(n22606) );
  XOR U23314 ( .A(n22601), .B(n22569), .Z(n22602) );
  XOR U23315 ( .A(n22609), .B(n22610), .Z(n22569) );
  AND U23316 ( .A(n1062), .B(n22611), .Z(n22609) );
  XOR U23317 ( .A(n22612), .B(n22610), .Z(n22611) );
  XNOR U23318 ( .A(n22613), .B(n22614), .Z(n22601) );
  NAND U23319 ( .A(n22615), .B(n22616), .Z(n22614) );
  XOR U23320 ( .A(n22617), .B(n22593), .Z(n22616) );
  XOR U23321 ( .A(n22607), .B(n22608), .Z(n22593) );
  XOR U23322 ( .A(n22618), .B(n22619), .Z(n22608) );
  ANDN U23323 ( .B(n22620), .A(n22621), .Z(n22618) );
  XOR U23324 ( .A(n22619), .B(n22622), .Z(n22620) );
  XOR U23325 ( .A(n22623), .B(n22624), .Z(n22607) );
  XOR U23326 ( .A(n22625), .B(n22626), .Z(n22624) );
  ANDN U23327 ( .B(n22627), .A(n22628), .Z(n22625) );
  XOR U23328 ( .A(n22629), .B(n22626), .Z(n22627) );
  IV U23329 ( .A(n22605), .Z(n22623) );
  XOR U23330 ( .A(n22630), .B(n22631), .Z(n22605) );
  ANDN U23331 ( .B(n22632), .A(n22633), .Z(n22630) );
  XOR U23332 ( .A(n22631), .B(n22634), .Z(n22632) );
  IV U23333 ( .A(n22613), .Z(n22617) );
  XOR U23334 ( .A(n22613), .B(n22595), .Z(n22615) );
  XOR U23335 ( .A(n22635), .B(n22636), .Z(n22595) );
  AND U23336 ( .A(n1062), .B(n22637), .Z(n22635) );
  XOR U23337 ( .A(n22638), .B(n22636), .Z(n22637) );
  NANDN U23338 ( .A(n22597), .B(n22599), .Z(n22613) );
  XOR U23339 ( .A(n22639), .B(n22640), .Z(n22599) );
  AND U23340 ( .A(n1062), .B(n22641), .Z(n22639) );
  XOR U23341 ( .A(n22640), .B(n22642), .Z(n22641) );
  XOR U23342 ( .A(n22643), .B(n22644), .Z(n1062) );
  AND U23343 ( .A(n22645), .B(n22646), .Z(n22643) );
  XNOR U23344 ( .A(n22644), .B(n22610), .Z(n22646) );
  XNOR U23345 ( .A(n22647), .B(n22648), .Z(n22610) );
  ANDN U23346 ( .B(n22649), .A(n22650), .Z(n22647) );
  XOR U23347 ( .A(n22648), .B(n22651), .Z(n22649) );
  XOR U23348 ( .A(n22644), .B(n22612), .Z(n22645) );
  XOR U23349 ( .A(n22652), .B(n22653), .Z(n22612) );
  AND U23350 ( .A(n1066), .B(n22654), .Z(n22652) );
  XOR U23351 ( .A(n22655), .B(n22653), .Z(n22654) );
  XNOR U23352 ( .A(n22656), .B(n22657), .Z(n22644) );
  NAND U23353 ( .A(n22658), .B(n22659), .Z(n22657) );
  XOR U23354 ( .A(n22660), .B(n22636), .Z(n22659) );
  XOR U23355 ( .A(n22650), .B(n22651), .Z(n22636) );
  XOR U23356 ( .A(n22661), .B(n22662), .Z(n22651) );
  ANDN U23357 ( .B(n22663), .A(n22664), .Z(n22661) );
  XOR U23358 ( .A(n22662), .B(n22665), .Z(n22663) );
  XOR U23359 ( .A(n22666), .B(n22667), .Z(n22650) );
  XOR U23360 ( .A(n22668), .B(n22669), .Z(n22667) );
  ANDN U23361 ( .B(n22670), .A(n22671), .Z(n22668) );
  XOR U23362 ( .A(n22672), .B(n22669), .Z(n22670) );
  IV U23363 ( .A(n22648), .Z(n22666) );
  XOR U23364 ( .A(n22673), .B(n22674), .Z(n22648) );
  ANDN U23365 ( .B(n22675), .A(n22676), .Z(n22673) );
  XOR U23366 ( .A(n22674), .B(n22677), .Z(n22675) );
  IV U23367 ( .A(n22656), .Z(n22660) );
  XOR U23368 ( .A(n22656), .B(n22638), .Z(n22658) );
  XOR U23369 ( .A(n22678), .B(n22679), .Z(n22638) );
  AND U23370 ( .A(n1066), .B(n22680), .Z(n22678) );
  XOR U23371 ( .A(n22681), .B(n22679), .Z(n22680) );
  NANDN U23372 ( .A(n22640), .B(n22642), .Z(n22656) );
  XOR U23373 ( .A(n22682), .B(n22683), .Z(n22642) );
  AND U23374 ( .A(n1066), .B(n22684), .Z(n22682) );
  XOR U23375 ( .A(n22683), .B(n22685), .Z(n22684) );
  XOR U23376 ( .A(n22686), .B(n22687), .Z(n1066) );
  AND U23377 ( .A(n22688), .B(n22689), .Z(n22686) );
  XNOR U23378 ( .A(n22687), .B(n22653), .Z(n22689) );
  XNOR U23379 ( .A(n22690), .B(n22691), .Z(n22653) );
  ANDN U23380 ( .B(n22692), .A(n22693), .Z(n22690) );
  XOR U23381 ( .A(n22691), .B(n22694), .Z(n22692) );
  XOR U23382 ( .A(n22687), .B(n22655), .Z(n22688) );
  XOR U23383 ( .A(n22695), .B(n22696), .Z(n22655) );
  AND U23384 ( .A(n1070), .B(n22697), .Z(n22695) );
  XOR U23385 ( .A(n22698), .B(n22696), .Z(n22697) );
  XNOR U23386 ( .A(n22699), .B(n22700), .Z(n22687) );
  NAND U23387 ( .A(n22701), .B(n22702), .Z(n22700) );
  XOR U23388 ( .A(n22703), .B(n22679), .Z(n22702) );
  XOR U23389 ( .A(n22693), .B(n22694), .Z(n22679) );
  XOR U23390 ( .A(n22704), .B(n22705), .Z(n22694) );
  ANDN U23391 ( .B(n22706), .A(n22707), .Z(n22704) );
  XOR U23392 ( .A(n22705), .B(n22708), .Z(n22706) );
  XOR U23393 ( .A(n22709), .B(n22710), .Z(n22693) );
  XOR U23394 ( .A(n22711), .B(n22712), .Z(n22710) );
  ANDN U23395 ( .B(n22713), .A(n22714), .Z(n22711) );
  XOR U23396 ( .A(n22715), .B(n22712), .Z(n22713) );
  IV U23397 ( .A(n22691), .Z(n22709) );
  XOR U23398 ( .A(n22716), .B(n22717), .Z(n22691) );
  ANDN U23399 ( .B(n22718), .A(n22719), .Z(n22716) );
  XOR U23400 ( .A(n22717), .B(n22720), .Z(n22718) );
  IV U23401 ( .A(n22699), .Z(n22703) );
  XOR U23402 ( .A(n22699), .B(n22681), .Z(n22701) );
  XOR U23403 ( .A(n22721), .B(n22722), .Z(n22681) );
  AND U23404 ( .A(n1070), .B(n22723), .Z(n22721) );
  XOR U23405 ( .A(n22724), .B(n22722), .Z(n22723) );
  NANDN U23406 ( .A(n22683), .B(n22685), .Z(n22699) );
  XOR U23407 ( .A(n22725), .B(n22726), .Z(n22685) );
  AND U23408 ( .A(n1070), .B(n22727), .Z(n22725) );
  XOR U23409 ( .A(n22726), .B(n22728), .Z(n22727) );
  XOR U23410 ( .A(n22729), .B(n22730), .Z(n1070) );
  AND U23411 ( .A(n22731), .B(n22732), .Z(n22729) );
  XNOR U23412 ( .A(n22730), .B(n22696), .Z(n22732) );
  XNOR U23413 ( .A(n22733), .B(n22734), .Z(n22696) );
  ANDN U23414 ( .B(n22735), .A(n22736), .Z(n22733) );
  XOR U23415 ( .A(n22734), .B(n22737), .Z(n22735) );
  XOR U23416 ( .A(n22730), .B(n22698), .Z(n22731) );
  XOR U23417 ( .A(n22738), .B(n22739), .Z(n22698) );
  AND U23418 ( .A(n1074), .B(n22740), .Z(n22738) );
  XOR U23419 ( .A(n22741), .B(n22739), .Z(n22740) );
  XNOR U23420 ( .A(n22742), .B(n22743), .Z(n22730) );
  NAND U23421 ( .A(n22744), .B(n22745), .Z(n22743) );
  XOR U23422 ( .A(n22746), .B(n22722), .Z(n22745) );
  XOR U23423 ( .A(n22736), .B(n22737), .Z(n22722) );
  XOR U23424 ( .A(n22747), .B(n22748), .Z(n22737) );
  ANDN U23425 ( .B(n22749), .A(n22750), .Z(n22747) );
  XOR U23426 ( .A(n22748), .B(n22751), .Z(n22749) );
  XOR U23427 ( .A(n22752), .B(n22753), .Z(n22736) );
  XOR U23428 ( .A(n22754), .B(n22755), .Z(n22753) );
  ANDN U23429 ( .B(n22756), .A(n22757), .Z(n22754) );
  XOR U23430 ( .A(n22758), .B(n22755), .Z(n22756) );
  IV U23431 ( .A(n22734), .Z(n22752) );
  XOR U23432 ( .A(n22759), .B(n22760), .Z(n22734) );
  ANDN U23433 ( .B(n22761), .A(n22762), .Z(n22759) );
  XOR U23434 ( .A(n22760), .B(n22763), .Z(n22761) );
  IV U23435 ( .A(n22742), .Z(n22746) );
  XOR U23436 ( .A(n22742), .B(n22724), .Z(n22744) );
  XOR U23437 ( .A(n22764), .B(n22765), .Z(n22724) );
  AND U23438 ( .A(n1074), .B(n22766), .Z(n22764) );
  XOR U23439 ( .A(n22767), .B(n22765), .Z(n22766) );
  NANDN U23440 ( .A(n22726), .B(n22728), .Z(n22742) );
  XOR U23441 ( .A(n22768), .B(n22769), .Z(n22728) );
  AND U23442 ( .A(n1074), .B(n22770), .Z(n22768) );
  XOR U23443 ( .A(n22769), .B(n22771), .Z(n22770) );
  XOR U23444 ( .A(n22772), .B(n22773), .Z(n1074) );
  AND U23445 ( .A(n22774), .B(n22775), .Z(n22772) );
  XNOR U23446 ( .A(n22773), .B(n22739), .Z(n22775) );
  XNOR U23447 ( .A(n22776), .B(n22777), .Z(n22739) );
  ANDN U23448 ( .B(n22778), .A(n22779), .Z(n22776) );
  XOR U23449 ( .A(n22777), .B(n22780), .Z(n22778) );
  XOR U23450 ( .A(n22773), .B(n22741), .Z(n22774) );
  XOR U23451 ( .A(n22781), .B(n22782), .Z(n22741) );
  AND U23452 ( .A(n1078), .B(n22783), .Z(n22781) );
  XOR U23453 ( .A(n22784), .B(n22782), .Z(n22783) );
  XNOR U23454 ( .A(n22785), .B(n22786), .Z(n22773) );
  NAND U23455 ( .A(n22787), .B(n22788), .Z(n22786) );
  XOR U23456 ( .A(n22789), .B(n22765), .Z(n22788) );
  XOR U23457 ( .A(n22779), .B(n22780), .Z(n22765) );
  XOR U23458 ( .A(n22790), .B(n22791), .Z(n22780) );
  ANDN U23459 ( .B(n22792), .A(n22793), .Z(n22790) );
  XOR U23460 ( .A(n22791), .B(n22794), .Z(n22792) );
  XOR U23461 ( .A(n22795), .B(n22796), .Z(n22779) );
  XOR U23462 ( .A(n22797), .B(n22798), .Z(n22796) );
  ANDN U23463 ( .B(n22799), .A(n22800), .Z(n22797) );
  XOR U23464 ( .A(n22801), .B(n22798), .Z(n22799) );
  IV U23465 ( .A(n22777), .Z(n22795) );
  XOR U23466 ( .A(n22802), .B(n22803), .Z(n22777) );
  ANDN U23467 ( .B(n22804), .A(n22805), .Z(n22802) );
  XOR U23468 ( .A(n22803), .B(n22806), .Z(n22804) );
  IV U23469 ( .A(n22785), .Z(n22789) );
  XOR U23470 ( .A(n22785), .B(n22767), .Z(n22787) );
  XOR U23471 ( .A(n22807), .B(n22808), .Z(n22767) );
  AND U23472 ( .A(n1078), .B(n22809), .Z(n22807) );
  XOR U23473 ( .A(n22810), .B(n22808), .Z(n22809) );
  NANDN U23474 ( .A(n22769), .B(n22771), .Z(n22785) );
  XOR U23475 ( .A(n22811), .B(n22812), .Z(n22771) );
  AND U23476 ( .A(n1078), .B(n22813), .Z(n22811) );
  XOR U23477 ( .A(n22812), .B(n22814), .Z(n22813) );
  XOR U23478 ( .A(n22815), .B(n22816), .Z(n1078) );
  AND U23479 ( .A(n22817), .B(n22818), .Z(n22815) );
  XNOR U23480 ( .A(n22816), .B(n22782), .Z(n22818) );
  XNOR U23481 ( .A(n22819), .B(n22820), .Z(n22782) );
  ANDN U23482 ( .B(n22821), .A(n22822), .Z(n22819) );
  XOR U23483 ( .A(n22820), .B(n22823), .Z(n22821) );
  XOR U23484 ( .A(n22816), .B(n22784), .Z(n22817) );
  XOR U23485 ( .A(n22824), .B(n22825), .Z(n22784) );
  AND U23486 ( .A(n1082), .B(n22826), .Z(n22824) );
  XOR U23487 ( .A(n22827), .B(n22825), .Z(n22826) );
  XNOR U23488 ( .A(n22828), .B(n22829), .Z(n22816) );
  NAND U23489 ( .A(n22830), .B(n22831), .Z(n22829) );
  XOR U23490 ( .A(n22832), .B(n22808), .Z(n22831) );
  XOR U23491 ( .A(n22822), .B(n22823), .Z(n22808) );
  XOR U23492 ( .A(n22833), .B(n22834), .Z(n22823) );
  ANDN U23493 ( .B(n22835), .A(n22836), .Z(n22833) );
  XOR U23494 ( .A(n22834), .B(n22837), .Z(n22835) );
  XOR U23495 ( .A(n22838), .B(n22839), .Z(n22822) );
  XOR U23496 ( .A(n22840), .B(n22841), .Z(n22839) );
  ANDN U23497 ( .B(n22842), .A(n22843), .Z(n22840) );
  XOR U23498 ( .A(n22844), .B(n22841), .Z(n22842) );
  IV U23499 ( .A(n22820), .Z(n22838) );
  XOR U23500 ( .A(n22845), .B(n22846), .Z(n22820) );
  ANDN U23501 ( .B(n22847), .A(n22848), .Z(n22845) );
  XOR U23502 ( .A(n22846), .B(n22849), .Z(n22847) );
  IV U23503 ( .A(n22828), .Z(n22832) );
  XOR U23504 ( .A(n22828), .B(n22810), .Z(n22830) );
  XOR U23505 ( .A(n22850), .B(n22851), .Z(n22810) );
  AND U23506 ( .A(n1082), .B(n22852), .Z(n22850) );
  XOR U23507 ( .A(n22853), .B(n22851), .Z(n22852) );
  NANDN U23508 ( .A(n22812), .B(n22814), .Z(n22828) );
  XOR U23509 ( .A(n22854), .B(n22855), .Z(n22814) );
  AND U23510 ( .A(n1082), .B(n22856), .Z(n22854) );
  XOR U23511 ( .A(n22855), .B(n22857), .Z(n22856) );
  XOR U23512 ( .A(n22858), .B(n22859), .Z(n1082) );
  AND U23513 ( .A(n22860), .B(n22861), .Z(n22858) );
  XNOR U23514 ( .A(n22859), .B(n22825), .Z(n22861) );
  XNOR U23515 ( .A(n22862), .B(n22863), .Z(n22825) );
  ANDN U23516 ( .B(n22864), .A(n22865), .Z(n22862) );
  XOR U23517 ( .A(n22863), .B(n22866), .Z(n22864) );
  XOR U23518 ( .A(n22859), .B(n22827), .Z(n22860) );
  XOR U23519 ( .A(n22867), .B(n22868), .Z(n22827) );
  AND U23520 ( .A(n1086), .B(n22869), .Z(n22867) );
  XOR U23521 ( .A(n22870), .B(n22868), .Z(n22869) );
  XNOR U23522 ( .A(n22871), .B(n22872), .Z(n22859) );
  NAND U23523 ( .A(n22873), .B(n22874), .Z(n22872) );
  XOR U23524 ( .A(n22875), .B(n22851), .Z(n22874) );
  XOR U23525 ( .A(n22865), .B(n22866), .Z(n22851) );
  XOR U23526 ( .A(n22876), .B(n22877), .Z(n22866) );
  ANDN U23527 ( .B(n22878), .A(n22879), .Z(n22876) );
  XOR U23528 ( .A(n22877), .B(n22880), .Z(n22878) );
  XOR U23529 ( .A(n22881), .B(n22882), .Z(n22865) );
  XOR U23530 ( .A(n22883), .B(n22884), .Z(n22882) );
  ANDN U23531 ( .B(n22885), .A(n22886), .Z(n22883) );
  XOR U23532 ( .A(n22887), .B(n22884), .Z(n22885) );
  IV U23533 ( .A(n22863), .Z(n22881) );
  XOR U23534 ( .A(n22888), .B(n22889), .Z(n22863) );
  ANDN U23535 ( .B(n22890), .A(n22891), .Z(n22888) );
  XOR U23536 ( .A(n22889), .B(n22892), .Z(n22890) );
  IV U23537 ( .A(n22871), .Z(n22875) );
  XOR U23538 ( .A(n22871), .B(n22853), .Z(n22873) );
  XOR U23539 ( .A(n22893), .B(n22894), .Z(n22853) );
  AND U23540 ( .A(n1086), .B(n22895), .Z(n22893) );
  XOR U23541 ( .A(n22896), .B(n22894), .Z(n22895) );
  NANDN U23542 ( .A(n22855), .B(n22857), .Z(n22871) );
  XOR U23543 ( .A(n22897), .B(n22898), .Z(n22857) );
  AND U23544 ( .A(n1086), .B(n22899), .Z(n22897) );
  XOR U23545 ( .A(n22898), .B(n22900), .Z(n22899) );
  XOR U23546 ( .A(n22901), .B(n22902), .Z(n1086) );
  AND U23547 ( .A(n22903), .B(n22904), .Z(n22901) );
  XNOR U23548 ( .A(n22902), .B(n22868), .Z(n22904) );
  XNOR U23549 ( .A(n22905), .B(n22906), .Z(n22868) );
  ANDN U23550 ( .B(n22907), .A(n22908), .Z(n22905) );
  XOR U23551 ( .A(n22906), .B(n22909), .Z(n22907) );
  XOR U23552 ( .A(n22902), .B(n22870), .Z(n22903) );
  XOR U23553 ( .A(n22910), .B(n22911), .Z(n22870) );
  AND U23554 ( .A(n1090), .B(n22912), .Z(n22910) );
  XOR U23555 ( .A(n22913), .B(n22911), .Z(n22912) );
  XNOR U23556 ( .A(n22914), .B(n22915), .Z(n22902) );
  NAND U23557 ( .A(n22916), .B(n22917), .Z(n22915) );
  XOR U23558 ( .A(n22918), .B(n22894), .Z(n22917) );
  XOR U23559 ( .A(n22908), .B(n22909), .Z(n22894) );
  XOR U23560 ( .A(n22919), .B(n22920), .Z(n22909) );
  ANDN U23561 ( .B(n22921), .A(n22922), .Z(n22919) );
  XOR U23562 ( .A(n22920), .B(n22923), .Z(n22921) );
  XOR U23563 ( .A(n22924), .B(n22925), .Z(n22908) );
  XOR U23564 ( .A(n22926), .B(n22927), .Z(n22925) );
  ANDN U23565 ( .B(n22928), .A(n22929), .Z(n22926) );
  XOR U23566 ( .A(n22930), .B(n22927), .Z(n22928) );
  IV U23567 ( .A(n22906), .Z(n22924) );
  XOR U23568 ( .A(n22931), .B(n22932), .Z(n22906) );
  ANDN U23569 ( .B(n22933), .A(n22934), .Z(n22931) );
  XOR U23570 ( .A(n22932), .B(n22935), .Z(n22933) );
  IV U23571 ( .A(n22914), .Z(n22918) );
  XOR U23572 ( .A(n22914), .B(n22896), .Z(n22916) );
  XOR U23573 ( .A(n22936), .B(n22937), .Z(n22896) );
  AND U23574 ( .A(n1090), .B(n22938), .Z(n22936) );
  XOR U23575 ( .A(n22939), .B(n22937), .Z(n22938) );
  NANDN U23576 ( .A(n22898), .B(n22900), .Z(n22914) );
  XOR U23577 ( .A(n22940), .B(n22941), .Z(n22900) );
  AND U23578 ( .A(n1090), .B(n22942), .Z(n22940) );
  XOR U23579 ( .A(n22941), .B(n22943), .Z(n22942) );
  XOR U23580 ( .A(n22944), .B(n22945), .Z(n1090) );
  AND U23581 ( .A(n22946), .B(n22947), .Z(n22944) );
  XNOR U23582 ( .A(n22945), .B(n22911), .Z(n22947) );
  XNOR U23583 ( .A(n22948), .B(n22949), .Z(n22911) );
  ANDN U23584 ( .B(n22950), .A(n22951), .Z(n22948) );
  XOR U23585 ( .A(n22949), .B(n22952), .Z(n22950) );
  XOR U23586 ( .A(n22945), .B(n22913), .Z(n22946) );
  XOR U23587 ( .A(n22953), .B(n22954), .Z(n22913) );
  AND U23588 ( .A(n1094), .B(n22955), .Z(n22953) );
  XOR U23589 ( .A(n22956), .B(n22954), .Z(n22955) );
  XNOR U23590 ( .A(n22957), .B(n22958), .Z(n22945) );
  NAND U23591 ( .A(n22959), .B(n22960), .Z(n22958) );
  XOR U23592 ( .A(n22961), .B(n22937), .Z(n22960) );
  XOR U23593 ( .A(n22951), .B(n22952), .Z(n22937) );
  XOR U23594 ( .A(n22962), .B(n22963), .Z(n22952) );
  ANDN U23595 ( .B(n22964), .A(n22965), .Z(n22962) );
  XOR U23596 ( .A(n22963), .B(n22966), .Z(n22964) );
  XOR U23597 ( .A(n22967), .B(n22968), .Z(n22951) );
  XOR U23598 ( .A(n22969), .B(n22970), .Z(n22968) );
  ANDN U23599 ( .B(n22971), .A(n22972), .Z(n22969) );
  XOR U23600 ( .A(n22973), .B(n22970), .Z(n22971) );
  IV U23601 ( .A(n22949), .Z(n22967) );
  XOR U23602 ( .A(n22974), .B(n22975), .Z(n22949) );
  ANDN U23603 ( .B(n22976), .A(n22977), .Z(n22974) );
  XOR U23604 ( .A(n22975), .B(n22978), .Z(n22976) );
  IV U23605 ( .A(n22957), .Z(n22961) );
  XOR U23606 ( .A(n22957), .B(n22939), .Z(n22959) );
  XOR U23607 ( .A(n22979), .B(n22980), .Z(n22939) );
  AND U23608 ( .A(n1094), .B(n22981), .Z(n22979) );
  XOR U23609 ( .A(n22982), .B(n22980), .Z(n22981) );
  NANDN U23610 ( .A(n22941), .B(n22943), .Z(n22957) );
  XOR U23611 ( .A(n22983), .B(n22984), .Z(n22943) );
  AND U23612 ( .A(n1094), .B(n22985), .Z(n22983) );
  XOR U23613 ( .A(n22984), .B(n22986), .Z(n22985) );
  XOR U23614 ( .A(n22987), .B(n22988), .Z(n1094) );
  AND U23615 ( .A(n22989), .B(n22990), .Z(n22987) );
  XNOR U23616 ( .A(n22988), .B(n22954), .Z(n22990) );
  XNOR U23617 ( .A(n22991), .B(n22992), .Z(n22954) );
  ANDN U23618 ( .B(n22993), .A(n22994), .Z(n22991) );
  XOR U23619 ( .A(n22992), .B(n22995), .Z(n22993) );
  XOR U23620 ( .A(n22988), .B(n22956), .Z(n22989) );
  XOR U23621 ( .A(n22996), .B(n22997), .Z(n22956) );
  AND U23622 ( .A(n1098), .B(n22998), .Z(n22996) );
  XOR U23623 ( .A(n22999), .B(n22997), .Z(n22998) );
  XNOR U23624 ( .A(n23000), .B(n23001), .Z(n22988) );
  NAND U23625 ( .A(n23002), .B(n23003), .Z(n23001) );
  XOR U23626 ( .A(n23004), .B(n22980), .Z(n23003) );
  XOR U23627 ( .A(n22994), .B(n22995), .Z(n22980) );
  XOR U23628 ( .A(n23005), .B(n23006), .Z(n22995) );
  ANDN U23629 ( .B(n23007), .A(n23008), .Z(n23005) );
  XOR U23630 ( .A(n23006), .B(n23009), .Z(n23007) );
  XOR U23631 ( .A(n23010), .B(n23011), .Z(n22994) );
  XOR U23632 ( .A(n23012), .B(n23013), .Z(n23011) );
  ANDN U23633 ( .B(n23014), .A(n23015), .Z(n23012) );
  XOR U23634 ( .A(n23016), .B(n23013), .Z(n23014) );
  IV U23635 ( .A(n22992), .Z(n23010) );
  XOR U23636 ( .A(n23017), .B(n23018), .Z(n22992) );
  ANDN U23637 ( .B(n23019), .A(n23020), .Z(n23017) );
  XOR U23638 ( .A(n23018), .B(n23021), .Z(n23019) );
  IV U23639 ( .A(n23000), .Z(n23004) );
  XOR U23640 ( .A(n23000), .B(n22982), .Z(n23002) );
  XOR U23641 ( .A(n23022), .B(n23023), .Z(n22982) );
  AND U23642 ( .A(n1098), .B(n23024), .Z(n23022) );
  XOR U23643 ( .A(n23025), .B(n23023), .Z(n23024) );
  NANDN U23644 ( .A(n22984), .B(n22986), .Z(n23000) );
  XOR U23645 ( .A(n23026), .B(n23027), .Z(n22986) );
  AND U23646 ( .A(n1098), .B(n23028), .Z(n23026) );
  XOR U23647 ( .A(n23027), .B(n23029), .Z(n23028) );
  XOR U23648 ( .A(n23030), .B(n23031), .Z(n1098) );
  AND U23649 ( .A(n23032), .B(n23033), .Z(n23030) );
  XNOR U23650 ( .A(n23031), .B(n22997), .Z(n23033) );
  XNOR U23651 ( .A(n23034), .B(n23035), .Z(n22997) );
  ANDN U23652 ( .B(n23036), .A(n23037), .Z(n23034) );
  XOR U23653 ( .A(n23035), .B(n23038), .Z(n23036) );
  XOR U23654 ( .A(n23031), .B(n22999), .Z(n23032) );
  XOR U23655 ( .A(n23039), .B(n23040), .Z(n22999) );
  AND U23656 ( .A(n1102), .B(n23041), .Z(n23039) );
  XOR U23657 ( .A(n23042), .B(n23040), .Z(n23041) );
  XNOR U23658 ( .A(n23043), .B(n23044), .Z(n23031) );
  NAND U23659 ( .A(n23045), .B(n23046), .Z(n23044) );
  XOR U23660 ( .A(n23047), .B(n23023), .Z(n23046) );
  XOR U23661 ( .A(n23037), .B(n23038), .Z(n23023) );
  XOR U23662 ( .A(n23048), .B(n23049), .Z(n23038) );
  ANDN U23663 ( .B(n23050), .A(n23051), .Z(n23048) );
  XOR U23664 ( .A(n23049), .B(n23052), .Z(n23050) );
  XOR U23665 ( .A(n23053), .B(n23054), .Z(n23037) );
  XOR U23666 ( .A(n23055), .B(n23056), .Z(n23054) );
  ANDN U23667 ( .B(n23057), .A(n23058), .Z(n23055) );
  XOR U23668 ( .A(n23059), .B(n23056), .Z(n23057) );
  IV U23669 ( .A(n23035), .Z(n23053) );
  XOR U23670 ( .A(n23060), .B(n23061), .Z(n23035) );
  ANDN U23671 ( .B(n23062), .A(n23063), .Z(n23060) );
  XOR U23672 ( .A(n23061), .B(n23064), .Z(n23062) );
  IV U23673 ( .A(n23043), .Z(n23047) );
  XOR U23674 ( .A(n23043), .B(n23025), .Z(n23045) );
  XOR U23675 ( .A(n23065), .B(n23066), .Z(n23025) );
  AND U23676 ( .A(n1102), .B(n23067), .Z(n23065) );
  XOR U23677 ( .A(n23068), .B(n23066), .Z(n23067) );
  NANDN U23678 ( .A(n23027), .B(n23029), .Z(n23043) );
  XOR U23679 ( .A(n23069), .B(n23070), .Z(n23029) );
  AND U23680 ( .A(n1102), .B(n23071), .Z(n23069) );
  XOR U23681 ( .A(n23070), .B(n23072), .Z(n23071) );
  XOR U23682 ( .A(n23073), .B(n23074), .Z(n1102) );
  AND U23683 ( .A(n23075), .B(n23076), .Z(n23073) );
  XNOR U23684 ( .A(n23074), .B(n23040), .Z(n23076) );
  XNOR U23685 ( .A(n23077), .B(n23078), .Z(n23040) );
  ANDN U23686 ( .B(n23079), .A(n23080), .Z(n23077) );
  XOR U23687 ( .A(n23078), .B(n23081), .Z(n23079) );
  XOR U23688 ( .A(n23074), .B(n23042), .Z(n23075) );
  XOR U23689 ( .A(n23082), .B(n23083), .Z(n23042) );
  AND U23690 ( .A(n1106), .B(n23084), .Z(n23082) );
  XOR U23691 ( .A(n23085), .B(n23083), .Z(n23084) );
  XNOR U23692 ( .A(n23086), .B(n23087), .Z(n23074) );
  NAND U23693 ( .A(n23088), .B(n23089), .Z(n23087) );
  XOR U23694 ( .A(n23090), .B(n23066), .Z(n23089) );
  XOR U23695 ( .A(n23080), .B(n23081), .Z(n23066) );
  XOR U23696 ( .A(n23091), .B(n23092), .Z(n23081) );
  ANDN U23697 ( .B(n23093), .A(n23094), .Z(n23091) );
  XOR U23698 ( .A(n23092), .B(n23095), .Z(n23093) );
  XOR U23699 ( .A(n23096), .B(n23097), .Z(n23080) );
  XOR U23700 ( .A(n23098), .B(n23099), .Z(n23097) );
  ANDN U23701 ( .B(n23100), .A(n23101), .Z(n23098) );
  XOR U23702 ( .A(n23102), .B(n23099), .Z(n23100) );
  IV U23703 ( .A(n23078), .Z(n23096) );
  XOR U23704 ( .A(n23103), .B(n23104), .Z(n23078) );
  ANDN U23705 ( .B(n23105), .A(n23106), .Z(n23103) );
  XOR U23706 ( .A(n23104), .B(n23107), .Z(n23105) );
  IV U23707 ( .A(n23086), .Z(n23090) );
  XOR U23708 ( .A(n23086), .B(n23068), .Z(n23088) );
  XOR U23709 ( .A(n23108), .B(n23109), .Z(n23068) );
  AND U23710 ( .A(n1106), .B(n23110), .Z(n23108) );
  XOR U23711 ( .A(n23111), .B(n23109), .Z(n23110) );
  NANDN U23712 ( .A(n23070), .B(n23072), .Z(n23086) );
  XOR U23713 ( .A(n23112), .B(n23113), .Z(n23072) );
  AND U23714 ( .A(n1106), .B(n23114), .Z(n23112) );
  XOR U23715 ( .A(n23113), .B(n23115), .Z(n23114) );
  XOR U23716 ( .A(n23116), .B(n23117), .Z(n1106) );
  AND U23717 ( .A(n23118), .B(n23119), .Z(n23116) );
  XNOR U23718 ( .A(n23117), .B(n23083), .Z(n23119) );
  XNOR U23719 ( .A(n23120), .B(n23121), .Z(n23083) );
  ANDN U23720 ( .B(n23122), .A(n23123), .Z(n23120) );
  XOR U23721 ( .A(n23121), .B(n23124), .Z(n23122) );
  XOR U23722 ( .A(n23117), .B(n23085), .Z(n23118) );
  XOR U23723 ( .A(n23125), .B(n23126), .Z(n23085) );
  AND U23724 ( .A(n1110), .B(n23127), .Z(n23125) );
  XOR U23725 ( .A(n23128), .B(n23126), .Z(n23127) );
  XNOR U23726 ( .A(n23129), .B(n23130), .Z(n23117) );
  NAND U23727 ( .A(n23131), .B(n23132), .Z(n23130) );
  XOR U23728 ( .A(n23133), .B(n23109), .Z(n23132) );
  XOR U23729 ( .A(n23123), .B(n23124), .Z(n23109) );
  XOR U23730 ( .A(n23134), .B(n23135), .Z(n23124) );
  ANDN U23731 ( .B(n23136), .A(n23137), .Z(n23134) );
  XOR U23732 ( .A(n23135), .B(n23138), .Z(n23136) );
  XOR U23733 ( .A(n23139), .B(n23140), .Z(n23123) );
  XOR U23734 ( .A(n23141), .B(n23142), .Z(n23140) );
  ANDN U23735 ( .B(n23143), .A(n23144), .Z(n23141) );
  XOR U23736 ( .A(n23145), .B(n23142), .Z(n23143) );
  IV U23737 ( .A(n23121), .Z(n23139) );
  XOR U23738 ( .A(n23146), .B(n23147), .Z(n23121) );
  ANDN U23739 ( .B(n23148), .A(n23149), .Z(n23146) );
  XOR U23740 ( .A(n23147), .B(n23150), .Z(n23148) );
  IV U23741 ( .A(n23129), .Z(n23133) );
  XOR U23742 ( .A(n23129), .B(n23111), .Z(n23131) );
  XOR U23743 ( .A(n23151), .B(n23152), .Z(n23111) );
  AND U23744 ( .A(n1110), .B(n23153), .Z(n23151) );
  XOR U23745 ( .A(n23154), .B(n23152), .Z(n23153) );
  NANDN U23746 ( .A(n23113), .B(n23115), .Z(n23129) );
  XOR U23747 ( .A(n23155), .B(n23156), .Z(n23115) );
  AND U23748 ( .A(n1110), .B(n23157), .Z(n23155) );
  XOR U23749 ( .A(n23156), .B(n23158), .Z(n23157) );
  XOR U23750 ( .A(n23159), .B(n23160), .Z(n1110) );
  AND U23751 ( .A(n23161), .B(n23162), .Z(n23159) );
  XNOR U23752 ( .A(n23160), .B(n23126), .Z(n23162) );
  XNOR U23753 ( .A(n23163), .B(n23164), .Z(n23126) );
  ANDN U23754 ( .B(n23165), .A(n23166), .Z(n23163) );
  XOR U23755 ( .A(n23164), .B(n23167), .Z(n23165) );
  XOR U23756 ( .A(n23160), .B(n23128), .Z(n23161) );
  XOR U23757 ( .A(n23168), .B(n23169), .Z(n23128) );
  AND U23758 ( .A(n1114), .B(n23170), .Z(n23168) );
  XOR U23759 ( .A(n23171), .B(n23169), .Z(n23170) );
  XNOR U23760 ( .A(n23172), .B(n23173), .Z(n23160) );
  NAND U23761 ( .A(n23174), .B(n23175), .Z(n23173) );
  XOR U23762 ( .A(n23176), .B(n23152), .Z(n23175) );
  XOR U23763 ( .A(n23166), .B(n23167), .Z(n23152) );
  XOR U23764 ( .A(n23177), .B(n23178), .Z(n23167) );
  ANDN U23765 ( .B(n23179), .A(n23180), .Z(n23177) );
  XOR U23766 ( .A(n23178), .B(n23181), .Z(n23179) );
  XOR U23767 ( .A(n23182), .B(n23183), .Z(n23166) );
  XOR U23768 ( .A(n23184), .B(n23185), .Z(n23183) );
  ANDN U23769 ( .B(n23186), .A(n23187), .Z(n23184) );
  XOR U23770 ( .A(n23188), .B(n23185), .Z(n23186) );
  IV U23771 ( .A(n23164), .Z(n23182) );
  XOR U23772 ( .A(n23189), .B(n23190), .Z(n23164) );
  ANDN U23773 ( .B(n23191), .A(n23192), .Z(n23189) );
  XOR U23774 ( .A(n23190), .B(n23193), .Z(n23191) );
  IV U23775 ( .A(n23172), .Z(n23176) );
  XOR U23776 ( .A(n23172), .B(n23154), .Z(n23174) );
  XOR U23777 ( .A(n23194), .B(n23195), .Z(n23154) );
  AND U23778 ( .A(n1114), .B(n23196), .Z(n23194) );
  XOR U23779 ( .A(n23197), .B(n23195), .Z(n23196) );
  NANDN U23780 ( .A(n23156), .B(n23158), .Z(n23172) );
  XOR U23781 ( .A(n23198), .B(n23199), .Z(n23158) );
  AND U23782 ( .A(n1114), .B(n23200), .Z(n23198) );
  XOR U23783 ( .A(n23199), .B(n23201), .Z(n23200) );
  XOR U23784 ( .A(n23202), .B(n23203), .Z(n1114) );
  AND U23785 ( .A(n23204), .B(n23205), .Z(n23202) );
  XNOR U23786 ( .A(n23203), .B(n23169), .Z(n23205) );
  XNOR U23787 ( .A(n23206), .B(n23207), .Z(n23169) );
  ANDN U23788 ( .B(n23208), .A(n23209), .Z(n23206) );
  XOR U23789 ( .A(n23207), .B(n23210), .Z(n23208) );
  XOR U23790 ( .A(n23203), .B(n23171), .Z(n23204) );
  XOR U23791 ( .A(n23211), .B(n23212), .Z(n23171) );
  AND U23792 ( .A(n1118), .B(n23213), .Z(n23211) );
  XOR U23793 ( .A(n23214), .B(n23212), .Z(n23213) );
  XNOR U23794 ( .A(n23215), .B(n23216), .Z(n23203) );
  NAND U23795 ( .A(n23217), .B(n23218), .Z(n23216) );
  XOR U23796 ( .A(n23219), .B(n23195), .Z(n23218) );
  XOR U23797 ( .A(n23209), .B(n23210), .Z(n23195) );
  XOR U23798 ( .A(n23220), .B(n23221), .Z(n23210) );
  ANDN U23799 ( .B(n23222), .A(n23223), .Z(n23220) );
  XOR U23800 ( .A(n23221), .B(n23224), .Z(n23222) );
  XOR U23801 ( .A(n23225), .B(n23226), .Z(n23209) );
  XOR U23802 ( .A(n23227), .B(n23228), .Z(n23226) );
  ANDN U23803 ( .B(n23229), .A(n23230), .Z(n23227) );
  XOR U23804 ( .A(n23231), .B(n23228), .Z(n23229) );
  IV U23805 ( .A(n23207), .Z(n23225) );
  XOR U23806 ( .A(n23232), .B(n23233), .Z(n23207) );
  ANDN U23807 ( .B(n23234), .A(n23235), .Z(n23232) );
  XOR U23808 ( .A(n23233), .B(n23236), .Z(n23234) );
  IV U23809 ( .A(n23215), .Z(n23219) );
  XOR U23810 ( .A(n23215), .B(n23197), .Z(n23217) );
  XOR U23811 ( .A(n23237), .B(n23238), .Z(n23197) );
  AND U23812 ( .A(n1118), .B(n23239), .Z(n23237) );
  XOR U23813 ( .A(n23240), .B(n23238), .Z(n23239) );
  NANDN U23814 ( .A(n23199), .B(n23201), .Z(n23215) );
  XOR U23815 ( .A(n23241), .B(n23242), .Z(n23201) );
  AND U23816 ( .A(n1118), .B(n23243), .Z(n23241) );
  XOR U23817 ( .A(n23242), .B(n23244), .Z(n23243) );
  XOR U23818 ( .A(n23245), .B(n23246), .Z(n1118) );
  AND U23819 ( .A(n23247), .B(n23248), .Z(n23245) );
  XNOR U23820 ( .A(n23246), .B(n23212), .Z(n23248) );
  XNOR U23821 ( .A(n23249), .B(n23250), .Z(n23212) );
  ANDN U23822 ( .B(n23251), .A(n23252), .Z(n23249) );
  XOR U23823 ( .A(n23250), .B(n23253), .Z(n23251) );
  XOR U23824 ( .A(n23246), .B(n23214), .Z(n23247) );
  XOR U23825 ( .A(n23254), .B(n23255), .Z(n23214) );
  AND U23826 ( .A(n1122), .B(n23256), .Z(n23254) );
  XOR U23827 ( .A(n23257), .B(n23255), .Z(n23256) );
  XNOR U23828 ( .A(n23258), .B(n23259), .Z(n23246) );
  NAND U23829 ( .A(n23260), .B(n23261), .Z(n23259) );
  XOR U23830 ( .A(n23262), .B(n23238), .Z(n23261) );
  XOR U23831 ( .A(n23252), .B(n23253), .Z(n23238) );
  XOR U23832 ( .A(n23263), .B(n23264), .Z(n23253) );
  ANDN U23833 ( .B(n23265), .A(n23266), .Z(n23263) );
  XOR U23834 ( .A(n23264), .B(n23267), .Z(n23265) );
  XOR U23835 ( .A(n23268), .B(n23269), .Z(n23252) );
  XOR U23836 ( .A(n23270), .B(n23271), .Z(n23269) );
  ANDN U23837 ( .B(n23272), .A(n23273), .Z(n23270) );
  XOR U23838 ( .A(n23274), .B(n23271), .Z(n23272) );
  IV U23839 ( .A(n23250), .Z(n23268) );
  XOR U23840 ( .A(n23275), .B(n23276), .Z(n23250) );
  ANDN U23841 ( .B(n23277), .A(n23278), .Z(n23275) );
  XOR U23842 ( .A(n23276), .B(n23279), .Z(n23277) );
  IV U23843 ( .A(n23258), .Z(n23262) );
  XOR U23844 ( .A(n23258), .B(n23240), .Z(n23260) );
  XOR U23845 ( .A(n23280), .B(n23281), .Z(n23240) );
  AND U23846 ( .A(n1122), .B(n23282), .Z(n23280) );
  XOR U23847 ( .A(n23283), .B(n23281), .Z(n23282) );
  NANDN U23848 ( .A(n23242), .B(n23244), .Z(n23258) );
  XOR U23849 ( .A(n23284), .B(n23285), .Z(n23244) );
  AND U23850 ( .A(n1122), .B(n23286), .Z(n23284) );
  XOR U23851 ( .A(n23285), .B(n23287), .Z(n23286) );
  XOR U23852 ( .A(n23288), .B(n23289), .Z(n1122) );
  AND U23853 ( .A(n23290), .B(n23291), .Z(n23288) );
  XNOR U23854 ( .A(n23289), .B(n23255), .Z(n23291) );
  XNOR U23855 ( .A(n23292), .B(n23293), .Z(n23255) );
  ANDN U23856 ( .B(n23294), .A(n23295), .Z(n23292) );
  XOR U23857 ( .A(n23293), .B(n23296), .Z(n23294) );
  XOR U23858 ( .A(n23289), .B(n23257), .Z(n23290) );
  XOR U23859 ( .A(n23297), .B(n23298), .Z(n23257) );
  AND U23860 ( .A(n1126), .B(n23299), .Z(n23297) );
  XOR U23861 ( .A(n23300), .B(n23298), .Z(n23299) );
  XNOR U23862 ( .A(n23301), .B(n23302), .Z(n23289) );
  NAND U23863 ( .A(n23303), .B(n23304), .Z(n23302) );
  XOR U23864 ( .A(n23305), .B(n23281), .Z(n23304) );
  XOR U23865 ( .A(n23295), .B(n23296), .Z(n23281) );
  XOR U23866 ( .A(n23306), .B(n23307), .Z(n23296) );
  ANDN U23867 ( .B(n23308), .A(n23309), .Z(n23306) );
  XOR U23868 ( .A(n23307), .B(n23310), .Z(n23308) );
  XOR U23869 ( .A(n23311), .B(n23312), .Z(n23295) );
  XOR U23870 ( .A(n23313), .B(n23314), .Z(n23312) );
  ANDN U23871 ( .B(n23315), .A(n23316), .Z(n23313) );
  XOR U23872 ( .A(n23317), .B(n23314), .Z(n23315) );
  IV U23873 ( .A(n23293), .Z(n23311) );
  XOR U23874 ( .A(n23318), .B(n23319), .Z(n23293) );
  ANDN U23875 ( .B(n23320), .A(n23321), .Z(n23318) );
  XOR U23876 ( .A(n23319), .B(n23322), .Z(n23320) );
  IV U23877 ( .A(n23301), .Z(n23305) );
  XOR U23878 ( .A(n23301), .B(n23283), .Z(n23303) );
  XOR U23879 ( .A(n23323), .B(n23324), .Z(n23283) );
  AND U23880 ( .A(n1126), .B(n23325), .Z(n23323) );
  XOR U23881 ( .A(n23326), .B(n23324), .Z(n23325) );
  NANDN U23882 ( .A(n23285), .B(n23287), .Z(n23301) );
  XOR U23883 ( .A(n23327), .B(n23328), .Z(n23287) );
  AND U23884 ( .A(n1126), .B(n23329), .Z(n23327) );
  XOR U23885 ( .A(n23328), .B(n23330), .Z(n23329) );
  XOR U23886 ( .A(n23331), .B(n23332), .Z(n1126) );
  AND U23887 ( .A(n23333), .B(n23334), .Z(n23331) );
  XNOR U23888 ( .A(n23332), .B(n23298), .Z(n23334) );
  XNOR U23889 ( .A(n23335), .B(n23336), .Z(n23298) );
  ANDN U23890 ( .B(n23337), .A(n23338), .Z(n23335) );
  XOR U23891 ( .A(n23336), .B(n23339), .Z(n23337) );
  XOR U23892 ( .A(n23332), .B(n23300), .Z(n23333) );
  XOR U23893 ( .A(n23340), .B(n23341), .Z(n23300) );
  AND U23894 ( .A(n1130), .B(n23342), .Z(n23340) );
  XOR U23895 ( .A(n23343), .B(n23341), .Z(n23342) );
  XNOR U23896 ( .A(n23344), .B(n23345), .Z(n23332) );
  NAND U23897 ( .A(n23346), .B(n23347), .Z(n23345) );
  XOR U23898 ( .A(n23348), .B(n23324), .Z(n23347) );
  XOR U23899 ( .A(n23338), .B(n23339), .Z(n23324) );
  XOR U23900 ( .A(n23349), .B(n23350), .Z(n23339) );
  ANDN U23901 ( .B(n23351), .A(n23352), .Z(n23349) );
  XOR U23902 ( .A(n23350), .B(n23353), .Z(n23351) );
  XOR U23903 ( .A(n23354), .B(n23355), .Z(n23338) );
  XOR U23904 ( .A(n23356), .B(n23357), .Z(n23355) );
  ANDN U23905 ( .B(n23358), .A(n23359), .Z(n23356) );
  XOR U23906 ( .A(n23360), .B(n23357), .Z(n23358) );
  IV U23907 ( .A(n23336), .Z(n23354) );
  XOR U23908 ( .A(n23361), .B(n23362), .Z(n23336) );
  ANDN U23909 ( .B(n23363), .A(n23364), .Z(n23361) );
  XOR U23910 ( .A(n23362), .B(n23365), .Z(n23363) );
  IV U23911 ( .A(n23344), .Z(n23348) );
  XOR U23912 ( .A(n23344), .B(n23326), .Z(n23346) );
  XOR U23913 ( .A(n23366), .B(n23367), .Z(n23326) );
  AND U23914 ( .A(n1130), .B(n23368), .Z(n23366) );
  XOR U23915 ( .A(n23369), .B(n23367), .Z(n23368) );
  NANDN U23916 ( .A(n23328), .B(n23330), .Z(n23344) );
  XOR U23917 ( .A(n23370), .B(n23371), .Z(n23330) );
  AND U23918 ( .A(n1130), .B(n23372), .Z(n23370) );
  XOR U23919 ( .A(n23371), .B(n23373), .Z(n23372) );
  XOR U23920 ( .A(n23374), .B(n23375), .Z(n1130) );
  AND U23921 ( .A(n23376), .B(n23377), .Z(n23374) );
  XNOR U23922 ( .A(n23375), .B(n23341), .Z(n23377) );
  XNOR U23923 ( .A(n23378), .B(n23379), .Z(n23341) );
  ANDN U23924 ( .B(n23380), .A(n23381), .Z(n23378) );
  XOR U23925 ( .A(n23379), .B(n23382), .Z(n23380) );
  XOR U23926 ( .A(n23375), .B(n23343), .Z(n23376) );
  XOR U23927 ( .A(n23383), .B(n23384), .Z(n23343) );
  AND U23928 ( .A(n1134), .B(n23385), .Z(n23383) );
  XOR U23929 ( .A(n23386), .B(n23384), .Z(n23385) );
  XNOR U23930 ( .A(n23387), .B(n23388), .Z(n23375) );
  NAND U23931 ( .A(n23389), .B(n23390), .Z(n23388) );
  XOR U23932 ( .A(n23391), .B(n23367), .Z(n23390) );
  XOR U23933 ( .A(n23381), .B(n23382), .Z(n23367) );
  XOR U23934 ( .A(n23392), .B(n23393), .Z(n23382) );
  ANDN U23935 ( .B(n23394), .A(n23395), .Z(n23392) );
  XOR U23936 ( .A(n23393), .B(n23396), .Z(n23394) );
  XOR U23937 ( .A(n23397), .B(n23398), .Z(n23381) );
  XOR U23938 ( .A(n23399), .B(n23400), .Z(n23398) );
  ANDN U23939 ( .B(n23401), .A(n23402), .Z(n23399) );
  XOR U23940 ( .A(n23403), .B(n23400), .Z(n23401) );
  IV U23941 ( .A(n23379), .Z(n23397) );
  XOR U23942 ( .A(n23404), .B(n23405), .Z(n23379) );
  ANDN U23943 ( .B(n23406), .A(n23407), .Z(n23404) );
  XOR U23944 ( .A(n23405), .B(n23408), .Z(n23406) );
  IV U23945 ( .A(n23387), .Z(n23391) );
  XOR U23946 ( .A(n23387), .B(n23369), .Z(n23389) );
  XOR U23947 ( .A(n23409), .B(n23410), .Z(n23369) );
  AND U23948 ( .A(n1134), .B(n23411), .Z(n23409) );
  XOR U23949 ( .A(n23412), .B(n23410), .Z(n23411) );
  NANDN U23950 ( .A(n23371), .B(n23373), .Z(n23387) );
  XOR U23951 ( .A(n23413), .B(n23414), .Z(n23373) );
  AND U23952 ( .A(n1134), .B(n23415), .Z(n23413) );
  XOR U23953 ( .A(n23414), .B(n23416), .Z(n23415) );
  XOR U23954 ( .A(n23417), .B(n23418), .Z(n1134) );
  AND U23955 ( .A(n23419), .B(n23420), .Z(n23417) );
  XNOR U23956 ( .A(n23418), .B(n23384), .Z(n23420) );
  XNOR U23957 ( .A(n23421), .B(n23422), .Z(n23384) );
  ANDN U23958 ( .B(n23423), .A(n23424), .Z(n23421) );
  XOR U23959 ( .A(n23422), .B(n23425), .Z(n23423) );
  XOR U23960 ( .A(n23418), .B(n23386), .Z(n23419) );
  XOR U23961 ( .A(n23426), .B(n23427), .Z(n23386) );
  AND U23962 ( .A(n1138), .B(n23428), .Z(n23426) );
  XOR U23963 ( .A(n23429), .B(n23427), .Z(n23428) );
  XNOR U23964 ( .A(n23430), .B(n23431), .Z(n23418) );
  NAND U23965 ( .A(n23432), .B(n23433), .Z(n23431) );
  XOR U23966 ( .A(n23434), .B(n23410), .Z(n23433) );
  XOR U23967 ( .A(n23424), .B(n23425), .Z(n23410) );
  XOR U23968 ( .A(n23435), .B(n23436), .Z(n23425) );
  ANDN U23969 ( .B(n23437), .A(n23438), .Z(n23435) );
  XOR U23970 ( .A(n23436), .B(n23439), .Z(n23437) );
  XOR U23971 ( .A(n23440), .B(n23441), .Z(n23424) );
  XOR U23972 ( .A(n23442), .B(n23443), .Z(n23441) );
  ANDN U23973 ( .B(n23444), .A(n23445), .Z(n23442) );
  XOR U23974 ( .A(n23446), .B(n23443), .Z(n23444) );
  IV U23975 ( .A(n23422), .Z(n23440) );
  XOR U23976 ( .A(n23447), .B(n23448), .Z(n23422) );
  ANDN U23977 ( .B(n23449), .A(n23450), .Z(n23447) );
  XOR U23978 ( .A(n23448), .B(n23451), .Z(n23449) );
  IV U23979 ( .A(n23430), .Z(n23434) );
  XOR U23980 ( .A(n23430), .B(n23412), .Z(n23432) );
  XOR U23981 ( .A(n23452), .B(n23453), .Z(n23412) );
  AND U23982 ( .A(n1138), .B(n23454), .Z(n23452) );
  XOR U23983 ( .A(n23455), .B(n23453), .Z(n23454) );
  NANDN U23984 ( .A(n23414), .B(n23416), .Z(n23430) );
  XOR U23985 ( .A(n23456), .B(n23457), .Z(n23416) );
  AND U23986 ( .A(n1138), .B(n23458), .Z(n23456) );
  XOR U23987 ( .A(n23457), .B(n23459), .Z(n23458) );
  XOR U23988 ( .A(n23460), .B(n23461), .Z(n1138) );
  AND U23989 ( .A(n23462), .B(n23463), .Z(n23460) );
  XNOR U23990 ( .A(n23461), .B(n23427), .Z(n23463) );
  XNOR U23991 ( .A(n23464), .B(n23465), .Z(n23427) );
  ANDN U23992 ( .B(n23466), .A(n23467), .Z(n23464) );
  XOR U23993 ( .A(n23465), .B(n23468), .Z(n23466) );
  XOR U23994 ( .A(n23461), .B(n23429), .Z(n23462) );
  XOR U23995 ( .A(n23469), .B(n23470), .Z(n23429) );
  AND U23996 ( .A(n1142), .B(n23471), .Z(n23469) );
  XOR U23997 ( .A(n23472), .B(n23470), .Z(n23471) );
  XNOR U23998 ( .A(n23473), .B(n23474), .Z(n23461) );
  NAND U23999 ( .A(n23475), .B(n23476), .Z(n23474) );
  XOR U24000 ( .A(n23477), .B(n23453), .Z(n23476) );
  XOR U24001 ( .A(n23467), .B(n23468), .Z(n23453) );
  XOR U24002 ( .A(n23478), .B(n23479), .Z(n23468) );
  ANDN U24003 ( .B(n23480), .A(n23481), .Z(n23478) );
  XOR U24004 ( .A(n23479), .B(n23482), .Z(n23480) );
  XOR U24005 ( .A(n23483), .B(n23484), .Z(n23467) );
  XOR U24006 ( .A(n23485), .B(n23486), .Z(n23484) );
  ANDN U24007 ( .B(n23487), .A(n23488), .Z(n23485) );
  XOR U24008 ( .A(n23489), .B(n23486), .Z(n23487) );
  IV U24009 ( .A(n23465), .Z(n23483) );
  XOR U24010 ( .A(n23490), .B(n23491), .Z(n23465) );
  ANDN U24011 ( .B(n23492), .A(n23493), .Z(n23490) );
  XOR U24012 ( .A(n23491), .B(n23494), .Z(n23492) );
  IV U24013 ( .A(n23473), .Z(n23477) );
  XOR U24014 ( .A(n23473), .B(n23455), .Z(n23475) );
  XOR U24015 ( .A(n23495), .B(n23496), .Z(n23455) );
  AND U24016 ( .A(n1142), .B(n23497), .Z(n23495) );
  XOR U24017 ( .A(n23498), .B(n23496), .Z(n23497) );
  NANDN U24018 ( .A(n23457), .B(n23459), .Z(n23473) );
  XOR U24019 ( .A(n23499), .B(n23500), .Z(n23459) );
  AND U24020 ( .A(n1142), .B(n23501), .Z(n23499) );
  XOR U24021 ( .A(n23500), .B(n23502), .Z(n23501) );
  XOR U24022 ( .A(n23503), .B(n23504), .Z(n1142) );
  AND U24023 ( .A(n23505), .B(n23506), .Z(n23503) );
  XNOR U24024 ( .A(n23504), .B(n23470), .Z(n23506) );
  XNOR U24025 ( .A(n23507), .B(n23508), .Z(n23470) );
  ANDN U24026 ( .B(n23509), .A(n23510), .Z(n23507) );
  XOR U24027 ( .A(n23508), .B(n23511), .Z(n23509) );
  XOR U24028 ( .A(n23504), .B(n23472), .Z(n23505) );
  XOR U24029 ( .A(n23512), .B(n23513), .Z(n23472) );
  AND U24030 ( .A(n1146), .B(n23514), .Z(n23512) );
  XOR U24031 ( .A(n23515), .B(n23513), .Z(n23514) );
  XNOR U24032 ( .A(n23516), .B(n23517), .Z(n23504) );
  NAND U24033 ( .A(n23518), .B(n23519), .Z(n23517) );
  XOR U24034 ( .A(n23520), .B(n23496), .Z(n23519) );
  XOR U24035 ( .A(n23510), .B(n23511), .Z(n23496) );
  XOR U24036 ( .A(n23521), .B(n23522), .Z(n23511) );
  ANDN U24037 ( .B(n23523), .A(n23524), .Z(n23521) );
  XOR U24038 ( .A(n23522), .B(n23525), .Z(n23523) );
  XOR U24039 ( .A(n23526), .B(n23527), .Z(n23510) );
  XOR U24040 ( .A(n23528), .B(n23529), .Z(n23527) );
  ANDN U24041 ( .B(n23530), .A(n23531), .Z(n23528) );
  XOR U24042 ( .A(n23532), .B(n23529), .Z(n23530) );
  IV U24043 ( .A(n23508), .Z(n23526) );
  XOR U24044 ( .A(n23533), .B(n23534), .Z(n23508) );
  ANDN U24045 ( .B(n23535), .A(n23536), .Z(n23533) );
  XOR U24046 ( .A(n23534), .B(n23537), .Z(n23535) );
  IV U24047 ( .A(n23516), .Z(n23520) );
  XOR U24048 ( .A(n23516), .B(n23498), .Z(n23518) );
  XOR U24049 ( .A(n23538), .B(n23539), .Z(n23498) );
  AND U24050 ( .A(n1146), .B(n23540), .Z(n23538) );
  XOR U24051 ( .A(n23541), .B(n23539), .Z(n23540) );
  NANDN U24052 ( .A(n23500), .B(n23502), .Z(n23516) );
  XOR U24053 ( .A(n23542), .B(n23543), .Z(n23502) );
  AND U24054 ( .A(n1146), .B(n23544), .Z(n23542) );
  XOR U24055 ( .A(n23543), .B(n23545), .Z(n23544) );
  XOR U24056 ( .A(n23546), .B(n23547), .Z(n1146) );
  AND U24057 ( .A(n23548), .B(n23549), .Z(n23546) );
  XNOR U24058 ( .A(n23547), .B(n23513), .Z(n23549) );
  XNOR U24059 ( .A(n23550), .B(n23551), .Z(n23513) );
  ANDN U24060 ( .B(n23552), .A(n23553), .Z(n23550) );
  XOR U24061 ( .A(n23551), .B(n23554), .Z(n23552) );
  XOR U24062 ( .A(n23547), .B(n23515), .Z(n23548) );
  XOR U24063 ( .A(n23555), .B(n23556), .Z(n23515) );
  AND U24064 ( .A(n1150), .B(n23557), .Z(n23555) );
  XOR U24065 ( .A(n23558), .B(n23556), .Z(n23557) );
  XNOR U24066 ( .A(n23559), .B(n23560), .Z(n23547) );
  NAND U24067 ( .A(n23561), .B(n23562), .Z(n23560) );
  XOR U24068 ( .A(n23563), .B(n23539), .Z(n23562) );
  XOR U24069 ( .A(n23553), .B(n23554), .Z(n23539) );
  XOR U24070 ( .A(n23564), .B(n23565), .Z(n23554) );
  ANDN U24071 ( .B(n23566), .A(n23567), .Z(n23564) );
  XOR U24072 ( .A(n23565), .B(n23568), .Z(n23566) );
  XOR U24073 ( .A(n23569), .B(n23570), .Z(n23553) );
  XOR U24074 ( .A(n23571), .B(n23572), .Z(n23570) );
  ANDN U24075 ( .B(n23573), .A(n23574), .Z(n23571) );
  XOR U24076 ( .A(n23575), .B(n23572), .Z(n23573) );
  IV U24077 ( .A(n23551), .Z(n23569) );
  XOR U24078 ( .A(n23576), .B(n23577), .Z(n23551) );
  ANDN U24079 ( .B(n23578), .A(n23579), .Z(n23576) );
  XOR U24080 ( .A(n23577), .B(n23580), .Z(n23578) );
  IV U24081 ( .A(n23559), .Z(n23563) );
  XOR U24082 ( .A(n23559), .B(n23541), .Z(n23561) );
  XOR U24083 ( .A(n23581), .B(n23582), .Z(n23541) );
  AND U24084 ( .A(n1150), .B(n23583), .Z(n23581) );
  XOR U24085 ( .A(n23584), .B(n23582), .Z(n23583) );
  NANDN U24086 ( .A(n23543), .B(n23545), .Z(n23559) );
  XOR U24087 ( .A(n23585), .B(n23586), .Z(n23545) );
  AND U24088 ( .A(n1150), .B(n23587), .Z(n23585) );
  XOR U24089 ( .A(n23586), .B(n23588), .Z(n23587) );
  XOR U24090 ( .A(n23589), .B(n23590), .Z(n1150) );
  AND U24091 ( .A(n23591), .B(n23592), .Z(n23589) );
  XNOR U24092 ( .A(n23590), .B(n23556), .Z(n23592) );
  XNOR U24093 ( .A(n23593), .B(n23594), .Z(n23556) );
  ANDN U24094 ( .B(n23595), .A(n23596), .Z(n23593) );
  XOR U24095 ( .A(n23594), .B(n23597), .Z(n23595) );
  XOR U24096 ( .A(n23590), .B(n23558), .Z(n23591) );
  XOR U24097 ( .A(n23598), .B(n23599), .Z(n23558) );
  AND U24098 ( .A(n1154), .B(n23600), .Z(n23598) );
  XOR U24099 ( .A(n23601), .B(n23599), .Z(n23600) );
  XNOR U24100 ( .A(n23602), .B(n23603), .Z(n23590) );
  NAND U24101 ( .A(n23604), .B(n23605), .Z(n23603) );
  XOR U24102 ( .A(n23606), .B(n23582), .Z(n23605) );
  XOR U24103 ( .A(n23596), .B(n23597), .Z(n23582) );
  XOR U24104 ( .A(n23607), .B(n23608), .Z(n23597) );
  ANDN U24105 ( .B(n23609), .A(n23610), .Z(n23607) );
  XOR U24106 ( .A(n23608), .B(n23611), .Z(n23609) );
  XOR U24107 ( .A(n23612), .B(n23613), .Z(n23596) );
  XOR U24108 ( .A(n23614), .B(n23615), .Z(n23613) );
  ANDN U24109 ( .B(n23616), .A(n23617), .Z(n23614) );
  XOR U24110 ( .A(n23618), .B(n23615), .Z(n23616) );
  IV U24111 ( .A(n23594), .Z(n23612) );
  XOR U24112 ( .A(n23619), .B(n23620), .Z(n23594) );
  ANDN U24113 ( .B(n23621), .A(n23622), .Z(n23619) );
  XOR U24114 ( .A(n23620), .B(n23623), .Z(n23621) );
  IV U24115 ( .A(n23602), .Z(n23606) );
  XOR U24116 ( .A(n23602), .B(n23584), .Z(n23604) );
  XOR U24117 ( .A(n23624), .B(n23625), .Z(n23584) );
  AND U24118 ( .A(n1154), .B(n23626), .Z(n23624) );
  XOR U24119 ( .A(n23627), .B(n23625), .Z(n23626) );
  NANDN U24120 ( .A(n23586), .B(n23588), .Z(n23602) );
  XOR U24121 ( .A(n23628), .B(n23629), .Z(n23588) );
  AND U24122 ( .A(n1154), .B(n23630), .Z(n23628) );
  XOR U24123 ( .A(n23629), .B(n23631), .Z(n23630) );
  XOR U24124 ( .A(n23632), .B(n23633), .Z(n1154) );
  AND U24125 ( .A(n23634), .B(n23635), .Z(n23632) );
  XNOR U24126 ( .A(n23633), .B(n23599), .Z(n23635) );
  XNOR U24127 ( .A(n23636), .B(n23637), .Z(n23599) );
  ANDN U24128 ( .B(n23638), .A(n23639), .Z(n23636) );
  XOR U24129 ( .A(n23637), .B(n23640), .Z(n23638) );
  XOR U24130 ( .A(n23633), .B(n23601), .Z(n23634) );
  XOR U24131 ( .A(n23641), .B(n23642), .Z(n23601) );
  AND U24132 ( .A(n1158), .B(n23643), .Z(n23641) );
  XOR U24133 ( .A(n23644), .B(n23642), .Z(n23643) );
  XNOR U24134 ( .A(n23645), .B(n23646), .Z(n23633) );
  NAND U24135 ( .A(n23647), .B(n23648), .Z(n23646) );
  XOR U24136 ( .A(n23649), .B(n23625), .Z(n23648) );
  XOR U24137 ( .A(n23639), .B(n23640), .Z(n23625) );
  XOR U24138 ( .A(n23650), .B(n23651), .Z(n23640) );
  ANDN U24139 ( .B(n23652), .A(n23653), .Z(n23650) );
  XOR U24140 ( .A(n23651), .B(n23654), .Z(n23652) );
  XOR U24141 ( .A(n23655), .B(n23656), .Z(n23639) );
  XOR U24142 ( .A(n23657), .B(n23658), .Z(n23656) );
  ANDN U24143 ( .B(n23659), .A(n23660), .Z(n23657) );
  XOR U24144 ( .A(n23661), .B(n23658), .Z(n23659) );
  IV U24145 ( .A(n23637), .Z(n23655) );
  XOR U24146 ( .A(n23662), .B(n23663), .Z(n23637) );
  ANDN U24147 ( .B(n23664), .A(n23665), .Z(n23662) );
  XOR U24148 ( .A(n23663), .B(n23666), .Z(n23664) );
  IV U24149 ( .A(n23645), .Z(n23649) );
  XOR U24150 ( .A(n23645), .B(n23627), .Z(n23647) );
  XOR U24151 ( .A(n23667), .B(n23668), .Z(n23627) );
  AND U24152 ( .A(n1158), .B(n23669), .Z(n23667) );
  XOR U24153 ( .A(n23670), .B(n23668), .Z(n23669) );
  NANDN U24154 ( .A(n23629), .B(n23631), .Z(n23645) );
  XOR U24155 ( .A(n23671), .B(n23672), .Z(n23631) );
  AND U24156 ( .A(n1158), .B(n23673), .Z(n23671) );
  XOR U24157 ( .A(n23672), .B(n23674), .Z(n23673) );
  XOR U24158 ( .A(n23675), .B(n23676), .Z(n1158) );
  AND U24159 ( .A(n23677), .B(n23678), .Z(n23675) );
  XNOR U24160 ( .A(n23676), .B(n23642), .Z(n23678) );
  XNOR U24161 ( .A(n23679), .B(n23680), .Z(n23642) );
  ANDN U24162 ( .B(n23681), .A(n23682), .Z(n23679) );
  XOR U24163 ( .A(n23680), .B(n23683), .Z(n23681) );
  XOR U24164 ( .A(n23676), .B(n23644), .Z(n23677) );
  XOR U24165 ( .A(n23684), .B(n23685), .Z(n23644) );
  AND U24166 ( .A(n1162), .B(n23686), .Z(n23684) );
  XOR U24167 ( .A(n23687), .B(n23685), .Z(n23686) );
  XNOR U24168 ( .A(n23688), .B(n23689), .Z(n23676) );
  NAND U24169 ( .A(n23690), .B(n23691), .Z(n23689) );
  XOR U24170 ( .A(n23692), .B(n23668), .Z(n23691) );
  XOR U24171 ( .A(n23682), .B(n23683), .Z(n23668) );
  XOR U24172 ( .A(n23693), .B(n23694), .Z(n23683) );
  ANDN U24173 ( .B(n23695), .A(n23696), .Z(n23693) );
  XOR U24174 ( .A(n23694), .B(n23697), .Z(n23695) );
  XOR U24175 ( .A(n23698), .B(n23699), .Z(n23682) );
  XOR U24176 ( .A(n23700), .B(n23701), .Z(n23699) );
  ANDN U24177 ( .B(n23702), .A(n23703), .Z(n23700) );
  XOR U24178 ( .A(n23704), .B(n23701), .Z(n23702) );
  IV U24179 ( .A(n23680), .Z(n23698) );
  XOR U24180 ( .A(n23705), .B(n23706), .Z(n23680) );
  ANDN U24181 ( .B(n23707), .A(n23708), .Z(n23705) );
  XOR U24182 ( .A(n23706), .B(n23709), .Z(n23707) );
  IV U24183 ( .A(n23688), .Z(n23692) );
  XOR U24184 ( .A(n23688), .B(n23670), .Z(n23690) );
  XOR U24185 ( .A(n23710), .B(n23711), .Z(n23670) );
  AND U24186 ( .A(n1162), .B(n23712), .Z(n23710) );
  XOR U24187 ( .A(n23713), .B(n23711), .Z(n23712) );
  NANDN U24188 ( .A(n23672), .B(n23674), .Z(n23688) );
  XOR U24189 ( .A(n23714), .B(n23715), .Z(n23674) );
  AND U24190 ( .A(n1162), .B(n23716), .Z(n23714) );
  XOR U24191 ( .A(n23715), .B(n23717), .Z(n23716) );
  XOR U24192 ( .A(n23718), .B(n23719), .Z(n1162) );
  AND U24193 ( .A(n23720), .B(n23721), .Z(n23718) );
  XNOR U24194 ( .A(n23719), .B(n23685), .Z(n23721) );
  XNOR U24195 ( .A(n23722), .B(n23723), .Z(n23685) );
  ANDN U24196 ( .B(n23724), .A(n23725), .Z(n23722) );
  XOR U24197 ( .A(n23723), .B(n23726), .Z(n23724) );
  XOR U24198 ( .A(n23719), .B(n23687), .Z(n23720) );
  XOR U24199 ( .A(n23727), .B(n23728), .Z(n23687) );
  AND U24200 ( .A(n1166), .B(n23729), .Z(n23727) );
  XOR U24201 ( .A(n23730), .B(n23728), .Z(n23729) );
  XNOR U24202 ( .A(n23731), .B(n23732), .Z(n23719) );
  NAND U24203 ( .A(n23733), .B(n23734), .Z(n23732) );
  XOR U24204 ( .A(n23735), .B(n23711), .Z(n23734) );
  XOR U24205 ( .A(n23725), .B(n23726), .Z(n23711) );
  XOR U24206 ( .A(n23736), .B(n23737), .Z(n23726) );
  ANDN U24207 ( .B(n23738), .A(n23739), .Z(n23736) );
  XOR U24208 ( .A(n23737), .B(n23740), .Z(n23738) );
  XOR U24209 ( .A(n23741), .B(n23742), .Z(n23725) );
  XOR U24210 ( .A(n23743), .B(n23744), .Z(n23742) );
  ANDN U24211 ( .B(n23745), .A(n23746), .Z(n23743) );
  XOR U24212 ( .A(n23747), .B(n23744), .Z(n23745) );
  IV U24213 ( .A(n23723), .Z(n23741) );
  XOR U24214 ( .A(n23748), .B(n23749), .Z(n23723) );
  ANDN U24215 ( .B(n23750), .A(n23751), .Z(n23748) );
  XOR U24216 ( .A(n23749), .B(n23752), .Z(n23750) );
  IV U24217 ( .A(n23731), .Z(n23735) );
  XOR U24218 ( .A(n23731), .B(n23713), .Z(n23733) );
  XOR U24219 ( .A(n23753), .B(n23754), .Z(n23713) );
  AND U24220 ( .A(n1166), .B(n23755), .Z(n23753) );
  XOR U24221 ( .A(n23756), .B(n23754), .Z(n23755) );
  NANDN U24222 ( .A(n23715), .B(n23717), .Z(n23731) );
  XOR U24223 ( .A(n23757), .B(n23758), .Z(n23717) );
  AND U24224 ( .A(n1166), .B(n23759), .Z(n23757) );
  XOR U24225 ( .A(n23758), .B(n23760), .Z(n23759) );
  XOR U24226 ( .A(n23761), .B(n23762), .Z(n1166) );
  AND U24227 ( .A(n23763), .B(n23764), .Z(n23761) );
  XNOR U24228 ( .A(n23762), .B(n23728), .Z(n23764) );
  XNOR U24229 ( .A(n23765), .B(n23766), .Z(n23728) );
  ANDN U24230 ( .B(n23767), .A(n23768), .Z(n23765) );
  XOR U24231 ( .A(n23766), .B(n23769), .Z(n23767) );
  XOR U24232 ( .A(n23762), .B(n23730), .Z(n23763) );
  XOR U24233 ( .A(n23770), .B(n23771), .Z(n23730) );
  AND U24234 ( .A(n1170), .B(n23772), .Z(n23770) );
  XOR U24235 ( .A(n23773), .B(n23771), .Z(n23772) );
  XNOR U24236 ( .A(n23774), .B(n23775), .Z(n23762) );
  NAND U24237 ( .A(n23776), .B(n23777), .Z(n23775) );
  XOR U24238 ( .A(n23778), .B(n23754), .Z(n23777) );
  XOR U24239 ( .A(n23768), .B(n23769), .Z(n23754) );
  XOR U24240 ( .A(n23779), .B(n23780), .Z(n23769) );
  ANDN U24241 ( .B(n23781), .A(n23782), .Z(n23779) );
  XOR U24242 ( .A(n23780), .B(n23783), .Z(n23781) );
  XOR U24243 ( .A(n23784), .B(n23785), .Z(n23768) );
  XOR U24244 ( .A(n23786), .B(n23787), .Z(n23785) );
  ANDN U24245 ( .B(n23788), .A(n23789), .Z(n23786) );
  XOR U24246 ( .A(n23790), .B(n23787), .Z(n23788) );
  IV U24247 ( .A(n23766), .Z(n23784) );
  XOR U24248 ( .A(n23791), .B(n23792), .Z(n23766) );
  ANDN U24249 ( .B(n23793), .A(n23794), .Z(n23791) );
  XOR U24250 ( .A(n23792), .B(n23795), .Z(n23793) );
  IV U24251 ( .A(n23774), .Z(n23778) );
  XOR U24252 ( .A(n23774), .B(n23756), .Z(n23776) );
  XOR U24253 ( .A(n23796), .B(n23797), .Z(n23756) );
  AND U24254 ( .A(n1170), .B(n23798), .Z(n23796) );
  XOR U24255 ( .A(n23799), .B(n23797), .Z(n23798) );
  NANDN U24256 ( .A(n23758), .B(n23760), .Z(n23774) );
  XOR U24257 ( .A(n23800), .B(n23801), .Z(n23760) );
  AND U24258 ( .A(n1170), .B(n23802), .Z(n23800) );
  XOR U24259 ( .A(n23801), .B(n23803), .Z(n23802) );
  XOR U24260 ( .A(n23804), .B(n23805), .Z(n1170) );
  AND U24261 ( .A(n23806), .B(n23807), .Z(n23804) );
  XNOR U24262 ( .A(n23805), .B(n23771), .Z(n23807) );
  XNOR U24263 ( .A(n23808), .B(n23809), .Z(n23771) );
  ANDN U24264 ( .B(n23810), .A(n23811), .Z(n23808) );
  XOR U24265 ( .A(n23809), .B(n23812), .Z(n23810) );
  XOR U24266 ( .A(n23805), .B(n23773), .Z(n23806) );
  XOR U24267 ( .A(n23813), .B(n23814), .Z(n23773) );
  AND U24268 ( .A(n1174), .B(n23815), .Z(n23813) );
  XOR U24269 ( .A(n23816), .B(n23814), .Z(n23815) );
  XNOR U24270 ( .A(n23817), .B(n23818), .Z(n23805) );
  NAND U24271 ( .A(n23819), .B(n23820), .Z(n23818) );
  XOR U24272 ( .A(n23821), .B(n23797), .Z(n23820) );
  XOR U24273 ( .A(n23811), .B(n23812), .Z(n23797) );
  XOR U24274 ( .A(n23822), .B(n23823), .Z(n23812) );
  ANDN U24275 ( .B(n23824), .A(n23825), .Z(n23822) );
  XOR U24276 ( .A(n23823), .B(n23826), .Z(n23824) );
  XOR U24277 ( .A(n23827), .B(n23828), .Z(n23811) );
  XOR U24278 ( .A(n23829), .B(n23830), .Z(n23828) );
  ANDN U24279 ( .B(n23831), .A(n23832), .Z(n23829) );
  XOR U24280 ( .A(n23833), .B(n23830), .Z(n23831) );
  IV U24281 ( .A(n23809), .Z(n23827) );
  XOR U24282 ( .A(n23834), .B(n23835), .Z(n23809) );
  ANDN U24283 ( .B(n23836), .A(n23837), .Z(n23834) );
  XOR U24284 ( .A(n23835), .B(n23838), .Z(n23836) );
  IV U24285 ( .A(n23817), .Z(n23821) );
  XOR U24286 ( .A(n23817), .B(n23799), .Z(n23819) );
  XOR U24287 ( .A(n23839), .B(n23840), .Z(n23799) );
  AND U24288 ( .A(n1174), .B(n23841), .Z(n23839) );
  XOR U24289 ( .A(n23842), .B(n23840), .Z(n23841) );
  NANDN U24290 ( .A(n23801), .B(n23803), .Z(n23817) );
  XOR U24291 ( .A(n23843), .B(n23844), .Z(n23803) );
  AND U24292 ( .A(n1174), .B(n23845), .Z(n23843) );
  XOR U24293 ( .A(n23844), .B(n23846), .Z(n23845) );
  XOR U24294 ( .A(n23847), .B(n23848), .Z(n1174) );
  AND U24295 ( .A(n23849), .B(n23850), .Z(n23847) );
  XNOR U24296 ( .A(n23848), .B(n23814), .Z(n23850) );
  XNOR U24297 ( .A(n23851), .B(n23852), .Z(n23814) );
  ANDN U24298 ( .B(n23853), .A(n23854), .Z(n23851) );
  XOR U24299 ( .A(n23852), .B(n23855), .Z(n23853) );
  XOR U24300 ( .A(n23848), .B(n23816), .Z(n23849) );
  XOR U24301 ( .A(n23856), .B(n23857), .Z(n23816) );
  AND U24302 ( .A(n1178), .B(n23858), .Z(n23856) );
  XOR U24303 ( .A(n23859), .B(n23857), .Z(n23858) );
  XNOR U24304 ( .A(n23860), .B(n23861), .Z(n23848) );
  NAND U24305 ( .A(n23862), .B(n23863), .Z(n23861) );
  XOR U24306 ( .A(n23864), .B(n23840), .Z(n23863) );
  XOR U24307 ( .A(n23854), .B(n23855), .Z(n23840) );
  XOR U24308 ( .A(n23865), .B(n23866), .Z(n23855) );
  ANDN U24309 ( .B(n23867), .A(n23868), .Z(n23865) );
  XOR U24310 ( .A(n23866), .B(n23869), .Z(n23867) );
  XOR U24311 ( .A(n23870), .B(n23871), .Z(n23854) );
  XOR U24312 ( .A(n23872), .B(n23873), .Z(n23871) );
  ANDN U24313 ( .B(n23874), .A(n23875), .Z(n23872) );
  XOR U24314 ( .A(n23876), .B(n23873), .Z(n23874) );
  IV U24315 ( .A(n23852), .Z(n23870) );
  XOR U24316 ( .A(n23877), .B(n23878), .Z(n23852) );
  ANDN U24317 ( .B(n23879), .A(n23880), .Z(n23877) );
  XOR U24318 ( .A(n23878), .B(n23881), .Z(n23879) );
  IV U24319 ( .A(n23860), .Z(n23864) );
  XOR U24320 ( .A(n23860), .B(n23842), .Z(n23862) );
  XOR U24321 ( .A(n23882), .B(n23883), .Z(n23842) );
  AND U24322 ( .A(n1178), .B(n23884), .Z(n23882) );
  XOR U24323 ( .A(n23885), .B(n23883), .Z(n23884) );
  NANDN U24324 ( .A(n23844), .B(n23846), .Z(n23860) );
  XOR U24325 ( .A(n23886), .B(n23887), .Z(n23846) );
  AND U24326 ( .A(n1178), .B(n23888), .Z(n23886) );
  XOR U24327 ( .A(n23887), .B(n23889), .Z(n23888) );
  XOR U24328 ( .A(n23890), .B(n23891), .Z(n1178) );
  AND U24329 ( .A(n23892), .B(n23893), .Z(n23890) );
  XNOR U24330 ( .A(n23891), .B(n23857), .Z(n23893) );
  XNOR U24331 ( .A(n23894), .B(n23895), .Z(n23857) );
  ANDN U24332 ( .B(n23896), .A(n23897), .Z(n23894) );
  XOR U24333 ( .A(n23895), .B(n23898), .Z(n23896) );
  XOR U24334 ( .A(n23891), .B(n23859), .Z(n23892) );
  XOR U24335 ( .A(n23899), .B(n23900), .Z(n23859) );
  AND U24336 ( .A(n1182), .B(n23901), .Z(n23899) );
  XOR U24337 ( .A(n23902), .B(n23900), .Z(n23901) );
  XNOR U24338 ( .A(n23903), .B(n23904), .Z(n23891) );
  NAND U24339 ( .A(n23905), .B(n23906), .Z(n23904) );
  XOR U24340 ( .A(n23907), .B(n23883), .Z(n23906) );
  XOR U24341 ( .A(n23897), .B(n23898), .Z(n23883) );
  XOR U24342 ( .A(n23908), .B(n23909), .Z(n23898) );
  ANDN U24343 ( .B(n23910), .A(n23911), .Z(n23908) );
  XOR U24344 ( .A(n23909), .B(n23912), .Z(n23910) );
  XOR U24345 ( .A(n23913), .B(n23914), .Z(n23897) );
  XOR U24346 ( .A(n23915), .B(n23916), .Z(n23914) );
  ANDN U24347 ( .B(n23917), .A(n23918), .Z(n23915) );
  XOR U24348 ( .A(n23919), .B(n23916), .Z(n23917) );
  IV U24349 ( .A(n23895), .Z(n23913) );
  XOR U24350 ( .A(n23920), .B(n23921), .Z(n23895) );
  ANDN U24351 ( .B(n23922), .A(n23923), .Z(n23920) );
  XOR U24352 ( .A(n23921), .B(n23924), .Z(n23922) );
  IV U24353 ( .A(n23903), .Z(n23907) );
  XOR U24354 ( .A(n23903), .B(n23885), .Z(n23905) );
  XOR U24355 ( .A(n23925), .B(n23926), .Z(n23885) );
  AND U24356 ( .A(n1182), .B(n23927), .Z(n23925) );
  XOR U24357 ( .A(n23928), .B(n23926), .Z(n23927) );
  NANDN U24358 ( .A(n23887), .B(n23889), .Z(n23903) );
  XOR U24359 ( .A(n23929), .B(n23930), .Z(n23889) );
  AND U24360 ( .A(n1182), .B(n23931), .Z(n23929) );
  XOR U24361 ( .A(n23930), .B(n23932), .Z(n23931) );
  XOR U24362 ( .A(n23933), .B(n23934), .Z(n1182) );
  AND U24363 ( .A(n23935), .B(n23936), .Z(n23933) );
  XNOR U24364 ( .A(n23934), .B(n23900), .Z(n23936) );
  XNOR U24365 ( .A(n23937), .B(n23938), .Z(n23900) );
  ANDN U24366 ( .B(n23939), .A(n23940), .Z(n23937) );
  XOR U24367 ( .A(n23938), .B(n23941), .Z(n23939) );
  XOR U24368 ( .A(n23934), .B(n23902), .Z(n23935) );
  XOR U24369 ( .A(n23942), .B(n23943), .Z(n23902) );
  AND U24370 ( .A(n1186), .B(n23944), .Z(n23942) );
  XOR U24371 ( .A(n23945), .B(n23943), .Z(n23944) );
  XNOR U24372 ( .A(n23946), .B(n23947), .Z(n23934) );
  NAND U24373 ( .A(n23948), .B(n23949), .Z(n23947) );
  XOR U24374 ( .A(n23950), .B(n23926), .Z(n23949) );
  XOR U24375 ( .A(n23940), .B(n23941), .Z(n23926) );
  XOR U24376 ( .A(n23951), .B(n23952), .Z(n23941) );
  ANDN U24377 ( .B(n23953), .A(n23954), .Z(n23951) );
  XOR U24378 ( .A(n23952), .B(n23955), .Z(n23953) );
  XOR U24379 ( .A(n23956), .B(n23957), .Z(n23940) );
  XOR U24380 ( .A(n23958), .B(n23959), .Z(n23957) );
  ANDN U24381 ( .B(n23960), .A(n23961), .Z(n23958) );
  XOR U24382 ( .A(n23962), .B(n23959), .Z(n23960) );
  IV U24383 ( .A(n23938), .Z(n23956) );
  XOR U24384 ( .A(n23963), .B(n23964), .Z(n23938) );
  ANDN U24385 ( .B(n23965), .A(n23966), .Z(n23963) );
  XOR U24386 ( .A(n23964), .B(n23967), .Z(n23965) );
  IV U24387 ( .A(n23946), .Z(n23950) );
  XOR U24388 ( .A(n23946), .B(n23928), .Z(n23948) );
  XOR U24389 ( .A(n23968), .B(n23969), .Z(n23928) );
  AND U24390 ( .A(n1186), .B(n23970), .Z(n23968) );
  XOR U24391 ( .A(n23971), .B(n23969), .Z(n23970) );
  NANDN U24392 ( .A(n23930), .B(n23932), .Z(n23946) );
  XOR U24393 ( .A(n23972), .B(n23973), .Z(n23932) );
  AND U24394 ( .A(n1186), .B(n23974), .Z(n23972) );
  XOR U24395 ( .A(n23973), .B(n23975), .Z(n23974) );
  XOR U24396 ( .A(n23976), .B(n23977), .Z(n1186) );
  AND U24397 ( .A(n23978), .B(n23979), .Z(n23976) );
  XNOR U24398 ( .A(n23977), .B(n23943), .Z(n23979) );
  XNOR U24399 ( .A(n23980), .B(n23981), .Z(n23943) );
  ANDN U24400 ( .B(n23982), .A(n23983), .Z(n23980) );
  XOR U24401 ( .A(n23981), .B(n23984), .Z(n23982) );
  XOR U24402 ( .A(n23977), .B(n23945), .Z(n23978) );
  XOR U24403 ( .A(n23985), .B(n23986), .Z(n23945) );
  AND U24404 ( .A(n1190), .B(n23987), .Z(n23985) );
  XOR U24405 ( .A(n23988), .B(n23986), .Z(n23987) );
  XNOR U24406 ( .A(n23989), .B(n23990), .Z(n23977) );
  NAND U24407 ( .A(n23991), .B(n23992), .Z(n23990) );
  XOR U24408 ( .A(n23993), .B(n23969), .Z(n23992) );
  XOR U24409 ( .A(n23983), .B(n23984), .Z(n23969) );
  XOR U24410 ( .A(n23994), .B(n23995), .Z(n23984) );
  ANDN U24411 ( .B(n23996), .A(n23997), .Z(n23994) );
  XOR U24412 ( .A(n23995), .B(n23998), .Z(n23996) );
  XOR U24413 ( .A(n23999), .B(n24000), .Z(n23983) );
  XOR U24414 ( .A(n24001), .B(n24002), .Z(n24000) );
  ANDN U24415 ( .B(n24003), .A(n24004), .Z(n24001) );
  XOR U24416 ( .A(n24005), .B(n24002), .Z(n24003) );
  IV U24417 ( .A(n23981), .Z(n23999) );
  XOR U24418 ( .A(n24006), .B(n24007), .Z(n23981) );
  ANDN U24419 ( .B(n24008), .A(n24009), .Z(n24006) );
  XOR U24420 ( .A(n24007), .B(n24010), .Z(n24008) );
  IV U24421 ( .A(n23989), .Z(n23993) );
  XOR U24422 ( .A(n23989), .B(n23971), .Z(n23991) );
  XOR U24423 ( .A(n24011), .B(n24012), .Z(n23971) );
  AND U24424 ( .A(n1190), .B(n24013), .Z(n24011) );
  XOR U24425 ( .A(n24014), .B(n24012), .Z(n24013) );
  NANDN U24426 ( .A(n23973), .B(n23975), .Z(n23989) );
  XOR U24427 ( .A(n24015), .B(n24016), .Z(n23975) );
  AND U24428 ( .A(n1190), .B(n24017), .Z(n24015) );
  XOR U24429 ( .A(n24016), .B(n24018), .Z(n24017) );
  XOR U24430 ( .A(n24019), .B(n24020), .Z(n1190) );
  AND U24431 ( .A(n24021), .B(n24022), .Z(n24019) );
  XNOR U24432 ( .A(n24020), .B(n23986), .Z(n24022) );
  XNOR U24433 ( .A(n24023), .B(n24024), .Z(n23986) );
  ANDN U24434 ( .B(n24025), .A(n24026), .Z(n24023) );
  XOR U24435 ( .A(n24024), .B(n24027), .Z(n24025) );
  XOR U24436 ( .A(n24020), .B(n23988), .Z(n24021) );
  XOR U24437 ( .A(n24028), .B(n24029), .Z(n23988) );
  AND U24438 ( .A(n1194), .B(n24030), .Z(n24028) );
  XOR U24439 ( .A(n24031), .B(n24029), .Z(n24030) );
  XNOR U24440 ( .A(n24032), .B(n24033), .Z(n24020) );
  NAND U24441 ( .A(n24034), .B(n24035), .Z(n24033) );
  XOR U24442 ( .A(n24036), .B(n24012), .Z(n24035) );
  XOR U24443 ( .A(n24026), .B(n24027), .Z(n24012) );
  XOR U24444 ( .A(n24037), .B(n24038), .Z(n24027) );
  ANDN U24445 ( .B(n24039), .A(n24040), .Z(n24037) );
  XOR U24446 ( .A(n24038), .B(n24041), .Z(n24039) );
  XOR U24447 ( .A(n24042), .B(n24043), .Z(n24026) );
  XOR U24448 ( .A(n24044), .B(n24045), .Z(n24043) );
  ANDN U24449 ( .B(n24046), .A(n24047), .Z(n24044) );
  XOR U24450 ( .A(n24048), .B(n24045), .Z(n24046) );
  IV U24451 ( .A(n24024), .Z(n24042) );
  XOR U24452 ( .A(n24049), .B(n24050), .Z(n24024) );
  ANDN U24453 ( .B(n24051), .A(n24052), .Z(n24049) );
  XOR U24454 ( .A(n24050), .B(n24053), .Z(n24051) );
  IV U24455 ( .A(n24032), .Z(n24036) );
  XOR U24456 ( .A(n24032), .B(n24014), .Z(n24034) );
  XOR U24457 ( .A(n24054), .B(n24055), .Z(n24014) );
  AND U24458 ( .A(n1194), .B(n24056), .Z(n24054) );
  XOR U24459 ( .A(n24057), .B(n24055), .Z(n24056) );
  NANDN U24460 ( .A(n24016), .B(n24018), .Z(n24032) );
  XOR U24461 ( .A(n24058), .B(n24059), .Z(n24018) );
  AND U24462 ( .A(n1194), .B(n24060), .Z(n24058) );
  XOR U24463 ( .A(n24059), .B(n24061), .Z(n24060) );
  XOR U24464 ( .A(n24062), .B(n24063), .Z(n1194) );
  AND U24465 ( .A(n24064), .B(n24065), .Z(n24062) );
  XNOR U24466 ( .A(n24063), .B(n24029), .Z(n24065) );
  XNOR U24467 ( .A(n24066), .B(n24067), .Z(n24029) );
  ANDN U24468 ( .B(n24068), .A(n24069), .Z(n24066) );
  XOR U24469 ( .A(n24067), .B(n24070), .Z(n24068) );
  XOR U24470 ( .A(n24063), .B(n24031), .Z(n24064) );
  XOR U24471 ( .A(n24071), .B(n24072), .Z(n24031) );
  AND U24472 ( .A(n1198), .B(n24073), .Z(n24071) );
  XOR U24473 ( .A(n24074), .B(n24072), .Z(n24073) );
  XNOR U24474 ( .A(n24075), .B(n24076), .Z(n24063) );
  NAND U24475 ( .A(n24077), .B(n24078), .Z(n24076) );
  XOR U24476 ( .A(n24079), .B(n24055), .Z(n24078) );
  XOR U24477 ( .A(n24069), .B(n24070), .Z(n24055) );
  XOR U24478 ( .A(n24080), .B(n24081), .Z(n24070) );
  ANDN U24479 ( .B(n24082), .A(n24083), .Z(n24080) );
  XOR U24480 ( .A(n24081), .B(n24084), .Z(n24082) );
  XOR U24481 ( .A(n24085), .B(n24086), .Z(n24069) );
  XOR U24482 ( .A(n24087), .B(n24088), .Z(n24086) );
  ANDN U24483 ( .B(n24089), .A(n24090), .Z(n24087) );
  XOR U24484 ( .A(n24091), .B(n24088), .Z(n24089) );
  IV U24485 ( .A(n24067), .Z(n24085) );
  XOR U24486 ( .A(n24092), .B(n24093), .Z(n24067) );
  ANDN U24487 ( .B(n24094), .A(n24095), .Z(n24092) );
  XOR U24488 ( .A(n24093), .B(n24096), .Z(n24094) );
  IV U24489 ( .A(n24075), .Z(n24079) );
  XOR U24490 ( .A(n24075), .B(n24057), .Z(n24077) );
  XOR U24491 ( .A(n24097), .B(n24098), .Z(n24057) );
  AND U24492 ( .A(n1198), .B(n24099), .Z(n24097) );
  XOR U24493 ( .A(n24100), .B(n24098), .Z(n24099) );
  NANDN U24494 ( .A(n24059), .B(n24061), .Z(n24075) );
  XOR U24495 ( .A(n24101), .B(n24102), .Z(n24061) );
  AND U24496 ( .A(n1198), .B(n24103), .Z(n24101) );
  XOR U24497 ( .A(n24102), .B(n24104), .Z(n24103) );
  XOR U24498 ( .A(n24105), .B(n24106), .Z(n1198) );
  AND U24499 ( .A(n24107), .B(n24108), .Z(n24105) );
  XNOR U24500 ( .A(n24106), .B(n24072), .Z(n24108) );
  XNOR U24501 ( .A(n24109), .B(n24110), .Z(n24072) );
  ANDN U24502 ( .B(n24111), .A(n24112), .Z(n24109) );
  XOR U24503 ( .A(n24110), .B(n24113), .Z(n24111) );
  XOR U24504 ( .A(n24106), .B(n24074), .Z(n24107) );
  XOR U24505 ( .A(n24114), .B(n24115), .Z(n24074) );
  AND U24506 ( .A(n1202), .B(n24116), .Z(n24114) );
  XOR U24507 ( .A(n24117), .B(n24115), .Z(n24116) );
  XNOR U24508 ( .A(n24118), .B(n24119), .Z(n24106) );
  NAND U24509 ( .A(n24120), .B(n24121), .Z(n24119) );
  XOR U24510 ( .A(n24122), .B(n24098), .Z(n24121) );
  XOR U24511 ( .A(n24112), .B(n24113), .Z(n24098) );
  XOR U24512 ( .A(n24123), .B(n24124), .Z(n24113) );
  ANDN U24513 ( .B(n24125), .A(n24126), .Z(n24123) );
  XOR U24514 ( .A(n24124), .B(n24127), .Z(n24125) );
  XOR U24515 ( .A(n24128), .B(n24129), .Z(n24112) );
  XOR U24516 ( .A(n24130), .B(n24131), .Z(n24129) );
  ANDN U24517 ( .B(n24132), .A(n24133), .Z(n24130) );
  XOR U24518 ( .A(n24134), .B(n24131), .Z(n24132) );
  IV U24519 ( .A(n24110), .Z(n24128) );
  XOR U24520 ( .A(n24135), .B(n24136), .Z(n24110) );
  ANDN U24521 ( .B(n24137), .A(n24138), .Z(n24135) );
  XOR U24522 ( .A(n24136), .B(n24139), .Z(n24137) );
  IV U24523 ( .A(n24118), .Z(n24122) );
  XOR U24524 ( .A(n24118), .B(n24100), .Z(n24120) );
  XOR U24525 ( .A(n24140), .B(n24141), .Z(n24100) );
  AND U24526 ( .A(n1202), .B(n24142), .Z(n24140) );
  XOR U24527 ( .A(n24143), .B(n24141), .Z(n24142) );
  NANDN U24528 ( .A(n24102), .B(n24104), .Z(n24118) );
  XOR U24529 ( .A(n24144), .B(n24145), .Z(n24104) );
  AND U24530 ( .A(n1202), .B(n24146), .Z(n24144) );
  XOR U24531 ( .A(n24145), .B(n24147), .Z(n24146) );
  XOR U24532 ( .A(n24148), .B(n24149), .Z(n1202) );
  AND U24533 ( .A(n24150), .B(n24151), .Z(n24148) );
  XNOR U24534 ( .A(n24149), .B(n24115), .Z(n24151) );
  XNOR U24535 ( .A(n24152), .B(n24153), .Z(n24115) );
  ANDN U24536 ( .B(n24154), .A(n24155), .Z(n24152) );
  XOR U24537 ( .A(n24153), .B(n24156), .Z(n24154) );
  XOR U24538 ( .A(n24149), .B(n24117), .Z(n24150) );
  XOR U24539 ( .A(n24157), .B(n24158), .Z(n24117) );
  AND U24540 ( .A(n1206), .B(n24159), .Z(n24157) );
  XOR U24541 ( .A(n24160), .B(n24158), .Z(n24159) );
  XNOR U24542 ( .A(n24161), .B(n24162), .Z(n24149) );
  NAND U24543 ( .A(n24163), .B(n24164), .Z(n24162) );
  XOR U24544 ( .A(n24165), .B(n24141), .Z(n24164) );
  XOR U24545 ( .A(n24155), .B(n24156), .Z(n24141) );
  XOR U24546 ( .A(n24166), .B(n24167), .Z(n24156) );
  ANDN U24547 ( .B(n24168), .A(n24169), .Z(n24166) );
  XOR U24548 ( .A(n24167), .B(n24170), .Z(n24168) );
  XOR U24549 ( .A(n24171), .B(n24172), .Z(n24155) );
  XOR U24550 ( .A(n24173), .B(n24174), .Z(n24172) );
  ANDN U24551 ( .B(n24175), .A(n24176), .Z(n24173) );
  XOR U24552 ( .A(n24177), .B(n24174), .Z(n24175) );
  IV U24553 ( .A(n24153), .Z(n24171) );
  XOR U24554 ( .A(n24178), .B(n24179), .Z(n24153) );
  ANDN U24555 ( .B(n24180), .A(n24181), .Z(n24178) );
  XOR U24556 ( .A(n24179), .B(n24182), .Z(n24180) );
  IV U24557 ( .A(n24161), .Z(n24165) );
  XOR U24558 ( .A(n24161), .B(n24143), .Z(n24163) );
  XOR U24559 ( .A(n24183), .B(n24184), .Z(n24143) );
  AND U24560 ( .A(n1206), .B(n24185), .Z(n24183) );
  XOR U24561 ( .A(n24186), .B(n24184), .Z(n24185) );
  NANDN U24562 ( .A(n24145), .B(n24147), .Z(n24161) );
  XOR U24563 ( .A(n24187), .B(n24188), .Z(n24147) );
  AND U24564 ( .A(n1206), .B(n24189), .Z(n24187) );
  XOR U24565 ( .A(n24188), .B(n24190), .Z(n24189) );
  XOR U24566 ( .A(n24191), .B(n24192), .Z(n1206) );
  AND U24567 ( .A(n24193), .B(n24194), .Z(n24191) );
  XNOR U24568 ( .A(n24192), .B(n24158), .Z(n24194) );
  XNOR U24569 ( .A(n24195), .B(n24196), .Z(n24158) );
  ANDN U24570 ( .B(n24197), .A(n24198), .Z(n24195) );
  XOR U24571 ( .A(n24196), .B(n24199), .Z(n24197) );
  XOR U24572 ( .A(n24192), .B(n24160), .Z(n24193) );
  XOR U24573 ( .A(n24200), .B(n24201), .Z(n24160) );
  AND U24574 ( .A(n1210), .B(n24202), .Z(n24200) );
  XOR U24575 ( .A(n24203), .B(n24201), .Z(n24202) );
  XNOR U24576 ( .A(n24204), .B(n24205), .Z(n24192) );
  NAND U24577 ( .A(n24206), .B(n24207), .Z(n24205) );
  XOR U24578 ( .A(n24208), .B(n24184), .Z(n24207) );
  XOR U24579 ( .A(n24198), .B(n24199), .Z(n24184) );
  XOR U24580 ( .A(n24209), .B(n24210), .Z(n24199) );
  ANDN U24581 ( .B(n24211), .A(n24212), .Z(n24209) );
  XOR U24582 ( .A(n24210), .B(n24213), .Z(n24211) );
  XOR U24583 ( .A(n24214), .B(n24215), .Z(n24198) );
  XOR U24584 ( .A(n24216), .B(n24217), .Z(n24215) );
  ANDN U24585 ( .B(n24218), .A(n24219), .Z(n24216) );
  XOR U24586 ( .A(n24220), .B(n24217), .Z(n24218) );
  IV U24587 ( .A(n24196), .Z(n24214) );
  XOR U24588 ( .A(n24221), .B(n24222), .Z(n24196) );
  ANDN U24589 ( .B(n24223), .A(n24224), .Z(n24221) );
  XOR U24590 ( .A(n24222), .B(n24225), .Z(n24223) );
  IV U24591 ( .A(n24204), .Z(n24208) );
  XOR U24592 ( .A(n24204), .B(n24186), .Z(n24206) );
  XOR U24593 ( .A(n24226), .B(n24227), .Z(n24186) );
  AND U24594 ( .A(n1210), .B(n24228), .Z(n24226) );
  XOR U24595 ( .A(n24229), .B(n24227), .Z(n24228) );
  NANDN U24596 ( .A(n24188), .B(n24190), .Z(n24204) );
  XOR U24597 ( .A(n24230), .B(n24231), .Z(n24190) );
  AND U24598 ( .A(n1210), .B(n24232), .Z(n24230) );
  XOR U24599 ( .A(n24231), .B(n24233), .Z(n24232) );
  XOR U24600 ( .A(n24234), .B(n24235), .Z(n1210) );
  AND U24601 ( .A(n24236), .B(n24237), .Z(n24234) );
  XNOR U24602 ( .A(n24235), .B(n24201), .Z(n24237) );
  XNOR U24603 ( .A(n24238), .B(n24239), .Z(n24201) );
  ANDN U24604 ( .B(n24240), .A(n24241), .Z(n24238) );
  XOR U24605 ( .A(n24239), .B(n24242), .Z(n24240) );
  XOR U24606 ( .A(n24235), .B(n24203), .Z(n24236) );
  XOR U24607 ( .A(n24243), .B(n24244), .Z(n24203) );
  AND U24608 ( .A(n1214), .B(n24245), .Z(n24243) );
  XOR U24609 ( .A(n24246), .B(n24244), .Z(n24245) );
  XNOR U24610 ( .A(n24247), .B(n24248), .Z(n24235) );
  NAND U24611 ( .A(n24249), .B(n24250), .Z(n24248) );
  XOR U24612 ( .A(n24251), .B(n24227), .Z(n24250) );
  XOR U24613 ( .A(n24241), .B(n24242), .Z(n24227) );
  XOR U24614 ( .A(n24252), .B(n24253), .Z(n24242) );
  ANDN U24615 ( .B(n24254), .A(n24255), .Z(n24252) );
  XOR U24616 ( .A(n24253), .B(n24256), .Z(n24254) );
  XOR U24617 ( .A(n24257), .B(n24258), .Z(n24241) );
  XOR U24618 ( .A(n24259), .B(n24260), .Z(n24258) );
  ANDN U24619 ( .B(n24261), .A(n24262), .Z(n24259) );
  XOR U24620 ( .A(n24263), .B(n24260), .Z(n24261) );
  IV U24621 ( .A(n24239), .Z(n24257) );
  XOR U24622 ( .A(n24264), .B(n24265), .Z(n24239) );
  ANDN U24623 ( .B(n24266), .A(n24267), .Z(n24264) );
  XOR U24624 ( .A(n24265), .B(n24268), .Z(n24266) );
  IV U24625 ( .A(n24247), .Z(n24251) );
  XOR U24626 ( .A(n24247), .B(n24229), .Z(n24249) );
  XOR U24627 ( .A(n24269), .B(n24270), .Z(n24229) );
  AND U24628 ( .A(n1214), .B(n24271), .Z(n24269) );
  XOR U24629 ( .A(n24272), .B(n24270), .Z(n24271) );
  NANDN U24630 ( .A(n24231), .B(n24233), .Z(n24247) );
  XOR U24631 ( .A(n24273), .B(n24274), .Z(n24233) );
  AND U24632 ( .A(n1214), .B(n24275), .Z(n24273) );
  XOR U24633 ( .A(n24274), .B(n24276), .Z(n24275) );
  XOR U24634 ( .A(n24277), .B(n24278), .Z(n1214) );
  AND U24635 ( .A(n24279), .B(n24280), .Z(n24277) );
  XNOR U24636 ( .A(n24278), .B(n24244), .Z(n24280) );
  XNOR U24637 ( .A(n24281), .B(n24282), .Z(n24244) );
  ANDN U24638 ( .B(n24283), .A(n24284), .Z(n24281) );
  XOR U24639 ( .A(n24282), .B(n24285), .Z(n24283) );
  XOR U24640 ( .A(n24278), .B(n24246), .Z(n24279) );
  XOR U24641 ( .A(n24286), .B(n24287), .Z(n24246) );
  AND U24642 ( .A(n1218), .B(n24288), .Z(n24286) );
  XOR U24643 ( .A(n24289), .B(n24287), .Z(n24288) );
  XNOR U24644 ( .A(n24290), .B(n24291), .Z(n24278) );
  NAND U24645 ( .A(n24292), .B(n24293), .Z(n24291) );
  XOR U24646 ( .A(n24294), .B(n24270), .Z(n24293) );
  XOR U24647 ( .A(n24284), .B(n24285), .Z(n24270) );
  XOR U24648 ( .A(n24295), .B(n24296), .Z(n24285) );
  ANDN U24649 ( .B(n24297), .A(n24298), .Z(n24295) );
  XOR U24650 ( .A(n24296), .B(n24299), .Z(n24297) );
  XOR U24651 ( .A(n24300), .B(n24301), .Z(n24284) );
  XOR U24652 ( .A(n24302), .B(n24303), .Z(n24301) );
  ANDN U24653 ( .B(n24304), .A(n24305), .Z(n24302) );
  XOR U24654 ( .A(n24306), .B(n24303), .Z(n24304) );
  IV U24655 ( .A(n24282), .Z(n24300) );
  XOR U24656 ( .A(n24307), .B(n24308), .Z(n24282) );
  ANDN U24657 ( .B(n24309), .A(n24310), .Z(n24307) );
  XOR U24658 ( .A(n24308), .B(n24311), .Z(n24309) );
  IV U24659 ( .A(n24290), .Z(n24294) );
  XOR U24660 ( .A(n24290), .B(n24272), .Z(n24292) );
  XOR U24661 ( .A(n24312), .B(n24313), .Z(n24272) );
  AND U24662 ( .A(n1218), .B(n24314), .Z(n24312) );
  XOR U24663 ( .A(n24315), .B(n24313), .Z(n24314) );
  NANDN U24664 ( .A(n24274), .B(n24276), .Z(n24290) );
  XOR U24665 ( .A(n24316), .B(n24317), .Z(n24276) );
  AND U24666 ( .A(n1218), .B(n24318), .Z(n24316) );
  XOR U24667 ( .A(n24317), .B(n24319), .Z(n24318) );
  XOR U24668 ( .A(n24320), .B(n24321), .Z(n1218) );
  AND U24669 ( .A(n24322), .B(n24323), .Z(n24320) );
  XNOR U24670 ( .A(n24321), .B(n24287), .Z(n24323) );
  XNOR U24671 ( .A(n24324), .B(n24325), .Z(n24287) );
  ANDN U24672 ( .B(n24326), .A(n24327), .Z(n24324) );
  XOR U24673 ( .A(n24325), .B(n24328), .Z(n24326) );
  XOR U24674 ( .A(n24321), .B(n24289), .Z(n24322) );
  XOR U24675 ( .A(n24329), .B(n24330), .Z(n24289) );
  AND U24676 ( .A(n1222), .B(n24331), .Z(n24329) );
  XOR U24677 ( .A(n24332), .B(n24330), .Z(n24331) );
  XNOR U24678 ( .A(n24333), .B(n24334), .Z(n24321) );
  NAND U24679 ( .A(n24335), .B(n24336), .Z(n24334) );
  XOR U24680 ( .A(n24337), .B(n24313), .Z(n24336) );
  XOR U24681 ( .A(n24327), .B(n24328), .Z(n24313) );
  XOR U24682 ( .A(n24338), .B(n24339), .Z(n24328) );
  ANDN U24683 ( .B(n24340), .A(n24341), .Z(n24338) );
  XOR U24684 ( .A(n24339), .B(n24342), .Z(n24340) );
  XOR U24685 ( .A(n24343), .B(n24344), .Z(n24327) );
  XOR U24686 ( .A(n24345), .B(n24346), .Z(n24344) );
  ANDN U24687 ( .B(n24347), .A(n24348), .Z(n24345) );
  XOR U24688 ( .A(n24349), .B(n24346), .Z(n24347) );
  IV U24689 ( .A(n24325), .Z(n24343) );
  XOR U24690 ( .A(n24350), .B(n24351), .Z(n24325) );
  ANDN U24691 ( .B(n24352), .A(n24353), .Z(n24350) );
  XOR U24692 ( .A(n24351), .B(n24354), .Z(n24352) );
  IV U24693 ( .A(n24333), .Z(n24337) );
  XOR U24694 ( .A(n24333), .B(n24315), .Z(n24335) );
  XOR U24695 ( .A(n24355), .B(n24356), .Z(n24315) );
  AND U24696 ( .A(n1222), .B(n24357), .Z(n24355) );
  XOR U24697 ( .A(n24358), .B(n24356), .Z(n24357) );
  NANDN U24698 ( .A(n24317), .B(n24319), .Z(n24333) );
  XOR U24699 ( .A(n24359), .B(n24360), .Z(n24319) );
  AND U24700 ( .A(n1222), .B(n24361), .Z(n24359) );
  XOR U24701 ( .A(n24360), .B(n24362), .Z(n24361) );
  XOR U24702 ( .A(n24363), .B(n24364), .Z(n1222) );
  AND U24703 ( .A(n24365), .B(n24366), .Z(n24363) );
  XNOR U24704 ( .A(n24364), .B(n24330), .Z(n24366) );
  XNOR U24705 ( .A(n24367), .B(n24368), .Z(n24330) );
  ANDN U24706 ( .B(n24369), .A(n24370), .Z(n24367) );
  XOR U24707 ( .A(n24368), .B(n24371), .Z(n24369) );
  XOR U24708 ( .A(n24364), .B(n24332), .Z(n24365) );
  XOR U24709 ( .A(n24372), .B(n24373), .Z(n24332) );
  AND U24710 ( .A(n1226), .B(n24374), .Z(n24372) );
  XOR U24711 ( .A(n24375), .B(n24373), .Z(n24374) );
  XNOR U24712 ( .A(n24376), .B(n24377), .Z(n24364) );
  NAND U24713 ( .A(n24378), .B(n24379), .Z(n24377) );
  XOR U24714 ( .A(n24380), .B(n24356), .Z(n24379) );
  XOR U24715 ( .A(n24370), .B(n24371), .Z(n24356) );
  XOR U24716 ( .A(n24381), .B(n24382), .Z(n24371) );
  ANDN U24717 ( .B(n24383), .A(n24384), .Z(n24381) );
  XOR U24718 ( .A(n24382), .B(n24385), .Z(n24383) );
  XOR U24719 ( .A(n24386), .B(n24387), .Z(n24370) );
  XOR U24720 ( .A(n24388), .B(n24389), .Z(n24387) );
  ANDN U24721 ( .B(n24390), .A(n24391), .Z(n24388) );
  XOR U24722 ( .A(n24392), .B(n24389), .Z(n24390) );
  IV U24723 ( .A(n24368), .Z(n24386) );
  XOR U24724 ( .A(n24393), .B(n24394), .Z(n24368) );
  ANDN U24725 ( .B(n24395), .A(n24396), .Z(n24393) );
  XOR U24726 ( .A(n24394), .B(n24397), .Z(n24395) );
  IV U24727 ( .A(n24376), .Z(n24380) );
  XOR U24728 ( .A(n24376), .B(n24358), .Z(n24378) );
  XOR U24729 ( .A(n24398), .B(n24399), .Z(n24358) );
  AND U24730 ( .A(n1226), .B(n24400), .Z(n24398) );
  XOR U24731 ( .A(n24401), .B(n24399), .Z(n24400) );
  NANDN U24732 ( .A(n24360), .B(n24362), .Z(n24376) );
  XOR U24733 ( .A(n24402), .B(n24403), .Z(n24362) );
  AND U24734 ( .A(n1226), .B(n24404), .Z(n24402) );
  XOR U24735 ( .A(n24403), .B(n24405), .Z(n24404) );
  XOR U24736 ( .A(n24406), .B(n24407), .Z(n1226) );
  AND U24737 ( .A(n24408), .B(n24409), .Z(n24406) );
  XNOR U24738 ( .A(n24407), .B(n24373), .Z(n24409) );
  XNOR U24739 ( .A(n24410), .B(n24411), .Z(n24373) );
  ANDN U24740 ( .B(n24412), .A(n24413), .Z(n24410) );
  XOR U24741 ( .A(n24411), .B(n24414), .Z(n24412) );
  XOR U24742 ( .A(n24407), .B(n24375), .Z(n24408) );
  XOR U24743 ( .A(n24415), .B(n24416), .Z(n24375) );
  AND U24744 ( .A(n1230), .B(n24417), .Z(n24415) );
  XOR U24745 ( .A(n24418), .B(n24416), .Z(n24417) );
  XNOR U24746 ( .A(n24419), .B(n24420), .Z(n24407) );
  NAND U24747 ( .A(n24421), .B(n24422), .Z(n24420) );
  XOR U24748 ( .A(n24423), .B(n24399), .Z(n24422) );
  XOR U24749 ( .A(n24413), .B(n24414), .Z(n24399) );
  XOR U24750 ( .A(n24424), .B(n24425), .Z(n24414) );
  ANDN U24751 ( .B(n24426), .A(n24427), .Z(n24424) );
  XOR U24752 ( .A(n24425), .B(n24428), .Z(n24426) );
  XOR U24753 ( .A(n24429), .B(n24430), .Z(n24413) );
  XOR U24754 ( .A(n24431), .B(n24432), .Z(n24430) );
  ANDN U24755 ( .B(n24433), .A(n24434), .Z(n24431) );
  XOR U24756 ( .A(n24435), .B(n24432), .Z(n24433) );
  IV U24757 ( .A(n24411), .Z(n24429) );
  XOR U24758 ( .A(n24436), .B(n24437), .Z(n24411) );
  ANDN U24759 ( .B(n24438), .A(n24439), .Z(n24436) );
  XOR U24760 ( .A(n24437), .B(n24440), .Z(n24438) );
  IV U24761 ( .A(n24419), .Z(n24423) );
  XOR U24762 ( .A(n24419), .B(n24401), .Z(n24421) );
  XOR U24763 ( .A(n24441), .B(n24442), .Z(n24401) );
  AND U24764 ( .A(n1230), .B(n24443), .Z(n24441) );
  XOR U24765 ( .A(n24444), .B(n24442), .Z(n24443) );
  NANDN U24766 ( .A(n24403), .B(n24405), .Z(n24419) );
  XOR U24767 ( .A(n24445), .B(n24446), .Z(n24405) );
  AND U24768 ( .A(n1230), .B(n24447), .Z(n24445) );
  XOR U24769 ( .A(n24446), .B(n24448), .Z(n24447) );
  XOR U24770 ( .A(n24449), .B(n24450), .Z(n1230) );
  AND U24771 ( .A(n24451), .B(n24452), .Z(n24449) );
  XNOR U24772 ( .A(n24450), .B(n24416), .Z(n24452) );
  XNOR U24773 ( .A(n24453), .B(n24454), .Z(n24416) );
  ANDN U24774 ( .B(n24455), .A(n24456), .Z(n24453) );
  XOR U24775 ( .A(n24454), .B(n24457), .Z(n24455) );
  XOR U24776 ( .A(n24450), .B(n24418), .Z(n24451) );
  XOR U24777 ( .A(n24458), .B(n24459), .Z(n24418) );
  AND U24778 ( .A(n1234), .B(n24460), .Z(n24458) );
  XOR U24779 ( .A(n24461), .B(n24459), .Z(n24460) );
  XNOR U24780 ( .A(n24462), .B(n24463), .Z(n24450) );
  NAND U24781 ( .A(n24464), .B(n24465), .Z(n24463) );
  XOR U24782 ( .A(n24466), .B(n24442), .Z(n24465) );
  XOR U24783 ( .A(n24456), .B(n24457), .Z(n24442) );
  XOR U24784 ( .A(n24467), .B(n24468), .Z(n24457) );
  ANDN U24785 ( .B(n24469), .A(n24470), .Z(n24467) );
  XOR U24786 ( .A(n24468), .B(n24471), .Z(n24469) );
  XOR U24787 ( .A(n24472), .B(n24473), .Z(n24456) );
  XOR U24788 ( .A(n24474), .B(n24475), .Z(n24473) );
  ANDN U24789 ( .B(n24476), .A(n24477), .Z(n24474) );
  XOR U24790 ( .A(n24478), .B(n24475), .Z(n24476) );
  IV U24791 ( .A(n24454), .Z(n24472) );
  XOR U24792 ( .A(n24479), .B(n24480), .Z(n24454) );
  ANDN U24793 ( .B(n24481), .A(n24482), .Z(n24479) );
  XOR U24794 ( .A(n24480), .B(n24483), .Z(n24481) );
  IV U24795 ( .A(n24462), .Z(n24466) );
  XOR U24796 ( .A(n24462), .B(n24444), .Z(n24464) );
  XOR U24797 ( .A(n24484), .B(n24485), .Z(n24444) );
  AND U24798 ( .A(n1234), .B(n24486), .Z(n24484) );
  XOR U24799 ( .A(n24487), .B(n24485), .Z(n24486) );
  NANDN U24800 ( .A(n24446), .B(n24448), .Z(n24462) );
  XOR U24801 ( .A(n24488), .B(n24489), .Z(n24448) );
  AND U24802 ( .A(n1234), .B(n24490), .Z(n24488) );
  XOR U24803 ( .A(n24489), .B(n24491), .Z(n24490) );
  XOR U24804 ( .A(n24492), .B(n24493), .Z(n1234) );
  AND U24805 ( .A(n24494), .B(n24495), .Z(n24492) );
  XNOR U24806 ( .A(n24493), .B(n24459), .Z(n24495) );
  XNOR U24807 ( .A(n24496), .B(n24497), .Z(n24459) );
  ANDN U24808 ( .B(n24498), .A(n24499), .Z(n24496) );
  XOR U24809 ( .A(n24497), .B(n24500), .Z(n24498) );
  XOR U24810 ( .A(n24493), .B(n24461), .Z(n24494) );
  XOR U24811 ( .A(n24501), .B(n24502), .Z(n24461) );
  AND U24812 ( .A(n1238), .B(n24503), .Z(n24501) );
  XOR U24813 ( .A(n24504), .B(n24502), .Z(n24503) );
  XNOR U24814 ( .A(n24505), .B(n24506), .Z(n24493) );
  NAND U24815 ( .A(n24507), .B(n24508), .Z(n24506) );
  XOR U24816 ( .A(n24509), .B(n24485), .Z(n24508) );
  XOR U24817 ( .A(n24499), .B(n24500), .Z(n24485) );
  XOR U24818 ( .A(n24510), .B(n24511), .Z(n24500) );
  ANDN U24819 ( .B(n24512), .A(n24513), .Z(n24510) );
  XOR U24820 ( .A(n24511), .B(n24514), .Z(n24512) );
  XOR U24821 ( .A(n24515), .B(n24516), .Z(n24499) );
  XOR U24822 ( .A(n24517), .B(n24518), .Z(n24516) );
  ANDN U24823 ( .B(n24519), .A(n24520), .Z(n24517) );
  XOR U24824 ( .A(n24521), .B(n24518), .Z(n24519) );
  IV U24825 ( .A(n24497), .Z(n24515) );
  XOR U24826 ( .A(n24522), .B(n24523), .Z(n24497) );
  ANDN U24827 ( .B(n24524), .A(n24525), .Z(n24522) );
  XOR U24828 ( .A(n24523), .B(n24526), .Z(n24524) );
  IV U24829 ( .A(n24505), .Z(n24509) );
  XOR U24830 ( .A(n24505), .B(n24487), .Z(n24507) );
  XOR U24831 ( .A(n24527), .B(n24528), .Z(n24487) );
  AND U24832 ( .A(n1238), .B(n24529), .Z(n24527) );
  XOR U24833 ( .A(n24530), .B(n24528), .Z(n24529) );
  NANDN U24834 ( .A(n24489), .B(n24491), .Z(n24505) );
  XOR U24835 ( .A(n24531), .B(n24532), .Z(n24491) );
  AND U24836 ( .A(n1238), .B(n24533), .Z(n24531) );
  XOR U24837 ( .A(n24532), .B(n24534), .Z(n24533) );
  XOR U24838 ( .A(n24535), .B(n24536), .Z(n1238) );
  AND U24839 ( .A(n24537), .B(n24538), .Z(n24535) );
  XNOR U24840 ( .A(n24536), .B(n24502), .Z(n24538) );
  XNOR U24841 ( .A(n24539), .B(n24540), .Z(n24502) );
  ANDN U24842 ( .B(n24541), .A(n24542), .Z(n24539) );
  XOR U24843 ( .A(n24540), .B(n24543), .Z(n24541) );
  XOR U24844 ( .A(n24536), .B(n24504), .Z(n24537) );
  XOR U24845 ( .A(n24544), .B(n24545), .Z(n24504) );
  AND U24846 ( .A(n1242), .B(n24546), .Z(n24544) );
  XOR U24847 ( .A(n24547), .B(n24545), .Z(n24546) );
  XNOR U24848 ( .A(n24548), .B(n24549), .Z(n24536) );
  NAND U24849 ( .A(n24550), .B(n24551), .Z(n24549) );
  XOR U24850 ( .A(n24552), .B(n24528), .Z(n24551) );
  XOR U24851 ( .A(n24542), .B(n24543), .Z(n24528) );
  XOR U24852 ( .A(n24553), .B(n24554), .Z(n24543) );
  ANDN U24853 ( .B(n24555), .A(n24556), .Z(n24553) );
  XOR U24854 ( .A(n24554), .B(n24557), .Z(n24555) );
  XOR U24855 ( .A(n24558), .B(n24559), .Z(n24542) );
  XOR U24856 ( .A(n24560), .B(n24561), .Z(n24559) );
  ANDN U24857 ( .B(n24562), .A(n24563), .Z(n24560) );
  XOR U24858 ( .A(n24564), .B(n24561), .Z(n24562) );
  IV U24859 ( .A(n24540), .Z(n24558) );
  XOR U24860 ( .A(n24565), .B(n24566), .Z(n24540) );
  ANDN U24861 ( .B(n24567), .A(n24568), .Z(n24565) );
  XOR U24862 ( .A(n24566), .B(n24569), .Z(n24567) );
  IV U24863 ( .A(n24548), .Z(n24552) );
  XOR U24864 ( .A(n24548), .B(n24530), .Z(n24550) );
  XOR U24865 ( .A(n24570), .B(n24571), .Z(n24530) );
  AND U24866 ( .A(n1242), .B(n24572), .Z(n24570) );
  XOR U24867 ( .A(n24573), .B(n24571), .Z(n24572) );
  NANDN U24868 ( .A(n24532), .B(n24534), .Z(n24548) );
  XOR U24869 ( .A(n24574), .B(n24575), .Z(n24534) );
  AND U24870 ( .A(n1242), .B(n24576), .Z(n24574) );
  XOR U24871 ( .A(n24575), .B(n24577), .Z(n24576) );
  XOR U24872 ( .A(n24578), .B(n24579), .Z(n1242) );
  AND U24873 ( .A(n24580), .B(n24581), .Z(n24578) );
  XNOR U24874 ( .A(n24579), .B(n24545), .Z(n24581) );
  XNOR U24875 ( .A(n24582), .B(n24583), .Z(n24545) );
  ANDN U24876 ( .B(n24584), .A(n24585), .Z(n24582) );
  XOR U24877 ( .A(n24583), .B(n24586), .Z(n24584) );
  XOR U24878 ( .A(n24579), .B(n24547), .Z(n24580) );
  XOR U24879 ( .A(n24587), .B(n24588), .Z(n24547) );
  AND U24880 ( .A(n1246), .B(n24589), .Z(n24587) );
  XOR U24881 ( .A(n24590), .B(n24588), .Z(n24589) );
  XNOR U24882 ( .A(n24591), .B(n24592), .Z(n24579) );
  NAND U24883 ( .A(n24593), .B(n24594), .Z(n24592) );
  XOR U24884 ( .A(n24595), .B(n24571), .Z(n24594) );
  XOR U24885 ( .A(n24585), .B(n24586), .Z(n24571) );
  XOR U24886 ( .A(n24596), .B(n24597), .Z(n24586) );
  ANDN U24887 ( .B(n24598), .A(n24599), .Z(n24596) );
  XOR U24888 ( .A(n24597), .B(n24600), .Z(n24598) );
  XOR U24889 ( .A(n24601), .B(n24602), .Z(n24585) );
  XOR U24890 ( .A(n24603), .B(n24604), .Z(n24602) );
  ANDN U24891 ( .B(n24605), .A(n24606), .Z(n24603) );
  XOR U24892 ( .A(n24607), .B(n24604), .Z(n24605) );
  IV U24893 ( .A(n24583), .Z(n24601) );
  XOR U24894 ( .A(n24608), .B(n24609), .Z(n24583) );
  ANDN U24895 ( .B(n24610), .A(n24611), .Z(n24608) );
  XOR U24896 ( .A(n24609), .B(n24612), .Z(n24610) );
  IV U24897 ( .A(n24591), .Z(n24595) );
  XOR U24898 ( .A(n24591), .B(n24573), .Z(n24593) );
  XOR U24899 ( .A(n24613), .B(n24614), .Z(n24573) );
  AND U24900 ( .A(n1246), .B(n24615), .Z(n24613) );
  XOR U24901 ( .A(n24616), .B(n24614), .Z(n24615) );
  NANDN U24902 ( .A(n24575), .B(n24577), .Z(n24591) );
  XOR U24903 ( .A(n24617), .B(n24618), .Z(n24577) );
  AND U24904 ( .A(n1246), .B(n24619), .Z(n24617) );
  XOR U24905 ( .A(n24618), .B(n24620), .Z(n24619) );
  XOR U24906 ( .A(n24621), .B(n24622), .Z(n1246) );
  AND U24907 ( .A(n24623), .B(n24624), .Z(n24621) );
  XNOR U24908 ( .A(n24622), .B(n24588), .Z(n24624) );
  XNOR U24909 ( .A(n24625), .B(n24626), .Z(n24588) );
  ANDN U24910 ( .B(n24627), .A(n24628), .Z(n24625) );
  XOR U24911 ( .A(n24626), .B(n24629), .Z(n24627) );
  XOR U24912 ( .A(n24622), .B(n24590), .Z(n24623) );
  XOR U24913 ( .A(n24630), .B(n24631), .Z(n24590) );
  AND U24914 ( .A(n1250), .B(n24632), .Z(n24630) );
  XOR U24915 ( .A(n24633), .B(n24631), .Z(n24632) );
  XNOR U24916 ( .A(n24634), .B(n24635), .Z(n24622) );
  NAND U24917 ( .A(n24636), .B(n24637), .Z(n24635) );
  XOR U24918 ( .A(n24638), .B(n24614), .Z(n24637) );
  XOR U24919 ( .A(n24628), .B(n24629), .Z(n24614) );
  XOR U24920 ( .A(n24639), .B(n24640), .Z(n24629) );
  ANDN U24921 ( .B(n24641), .A(n24642), .Z(n24639) );
  XOR U24922 ( .A(n24640), .B(n24643), .Z(n24641) );
  XOR U24923 ( .A(n24644), .B(n24645), .Z(n24628) );
  XOR U24924 ( .A(n24646), .B(n24647), .Z(n24645) );
  ANDN U24925 ( .B(n24648), .A(n24649), .Z(n24646) );
  XOR U24926 ( .A(n24650), .B(n24647), .Z(n24648) );
  IV U24927 ( .A(n24626), .Z(n24644) );
  XOR U24928 ( .A(n24651), .B(n24652), .Z(n24626) );
  ANDN U24929 ( .B(n24653), .A(n24654), .Z(n24651) );
  XOR U24930 ( .A(n24652), .B(n24655), .Z(n24653) );
  IV U24931 ( .A(n24634), .Z(n24638) );
  XOR U24932 ( .A(n24634), .B(n24616), .Z(n24636) );
  XOR U24933 ( .A(n24656), .B(n24657), .Z(n24616) );
  AND U24934 ( .A(n1250), .B(n24658), .Z(n24656) );
  XOR U24935 ( .A(n24659), .B(n24657), .Z(n24658) );
  NANDN U24936 ( .A(n24618), .B(n24620), .Z(n24634) );
  XOR U24937 ( .A(n24660), .B(n24661), .Z(n24620) );
  AND U24938 ( .A(n1250), .B(n24662), .Z(n24660) );
  XOR U24939 ( .A(n24661), .B(n24663), .Z(n24662) );
  XOR U24940 ( .A(n24664), .B(n24665), .Z(n1250) );
  AND U24941 ( .A(n24666), .B(n24667), .Z(n24664) );
  XNOR U24942 ( .A(n24665), .B(n24631), .Z(n24667) );
  XNOR U24943 ( .A(n24668), .B(n24669), .Z(n24631) );
  ANDN U24944 ( .B(n24670), .A(n24671), .Z(n24668) );
  XOR U24945 ( .A(n24669), .B(n24672), .Z(n24670) );
  XOR U24946 ( .A(n24665), .B(n24633), .Z(n24666) );
  XOR U24947 ( .A(n24673), .B(n24674), .Z(n24633) );
  AND U24948 ( .A(n1254), .B(n24675), .Z(n24673) );
  XOR U24949 ( .A(n24676), .B(n24674), .Z(n24675) );
  XNOR U24950 ( .A(n24677), .B(n24678), .Z(n24665) );
  NAND U24951 ( .A(n24679), .B(n24680), .Z(n24678) );
  XOR U24952 ( .A(n24681), .B(n24657), .Z(n24680) );
  XOR U24953 ( .A(n24671), .B(n24672), .Z(n24657) );
  XOR U24954 ( .A(n24682), .B(n24683), .Z(n24672) );
  ANDN U24955 ( .B(n24684), .A(n24685), .Z(n24682) );
  XOR U24956 ( .A(n24683), .B(n24686), .Z(n24684) );
  XOR U24957 ( .A(n24687), .B(n24688), .Z(n24671) );
  XOR U24958 ( .A(n24689), .B(n24690), .Z(n24688) );
  ANDN U24959 ( .B(n24691), .A(n24692), .Z(n24689) );
  XOR U24960 ( .A(n24693), .B(n24690), .Z(n24691) );
  IV U24961 ( .A(n24669), .Z(n24687) );
  XOR U24962 ( .A(n24694), .B(n24695), .Z(n24669) );
  ANDN U24963 ( .B(n24696), .A(n24697), .Z(n24694) );
  XOR U24964 ( .A(n24695), .B(n24698), .Z(n24696) );
  IV U24965 ( .A(n24677), .Z(n24681) );
  XOR U24966 ( .A(n24677), .B(n24659), .Z(n24679) );
  XOR U24967 ( .A(n24699), .B(n24700), .Z(n24659) );
  AND U24968 ( .A(n1254), .B(n24701), .Z(n24699) );
  XOR U24969 ( .A(n24702), .B(n24700), .Z(n24701) );
  NANDN U24970 ( .A(n24661), .B(n24663), .Z(n24677) );
  XOR U24971 ( .A(n24703), .B(n24704), .Z(n24663) );
  AND U24972 ( .A(n1254), .B(n24705), .Z(n24703) );
  XOR U24973 ( .A(n24704), .B(n24706), .Z(n24705) );
  XOR U24974 ( .A(n24707), .B(n24708), .Z(n1254) );
  AND U24975 ( .A(n24709), .B(n24710), .Z(n24707) );
  XNOR U24976 ( .A(n24708), .B(n24674), .Z(n24710) );
  XNOR U24977 ( .A(n24711), .B(n24712), .Z(n24674) );
  ANDN U24978 ( .B(n24713), .A(n24714), .Z(n24711) );
  XOR U24979 ( .A(n24712), .B(n24715), .Z(n24713) );
  XOR U24980 ( .A(n24708), .B(n24676), .Z(n24709) );
  XOR U24981 ( .A(n24716), .B(n24717), .Z(n24676) );
  AND U24982 ( .A(n1258), .B(n24718), .Z(n24716) );
  XOR U24983 ( .A(n24719), .B(n24717), .Z(n24718) );
  XNOR U24984 ( .A(n24720), .B(n24721), .Z(n24708) );
  NAND U24985 ( .A(n24722), .B(n24723), .Z(n24721) );
  XOR U24986 ( .A(n24724), .B(n24700), .Z(n24723) );
  XOR U24987 ( .A(n24714), .B(n24715), .Z(n24700) );
  XOR U24988 ( .A(n24725), .B(n24726), .Z(n24715) );
  ANDN U24989 ( .B(n24727), .A(n24728), .Z(n24725) );
  XOR U24990 ( .A(n24726), .B(n24729), .Z(n24727) );
  XOR U24991 ( .A(n24730), .B(n24731), .Z(n24714) );
  XOR U24992 ( .A(n24732), .B(n24733), .Z(n24731) );
  ANDN U24993 ( .B(n24734), .A(n24735), .Z(n24732) );
  XOR U24994 ( .A(n24736), .B(n24733), .Z(n24734) );
  IV U24995 ( .A(n24712), .Z(n24730) );
  XOR U24996 ( .A(n24737), .B(n24738), .Z(n24712) );
  ANDN U24997 ( .B(n24739), .A(n24740), .Z(n24737) );
  XOR U24998 ( .A(n24738), .B(n24741), .Z(n24739) );
  IV U24999 ( .A(n24720), .Z(n24724) );
  XOR U25000 ( .A(n24720), .B(n24702), .Z(n24722) );
  XOR U25001 ( .A(n24742), .B(n24743), .Z(n24702) );
  AND U25002 ( .A(n1258), .B(n24744), .Z(n24742) );
  XOR U25003 ( .A(n24745), .B(n24743), .Z(n24744) );
  NANDN U25004 ( .A(n24704), .B(n24706), .Z(n24720) );
  XOR U25005 ( .A(n24746), .B(n24747), .Z(n24706) );
  AND U25006 ( .A(n1258), .B(n24748), .Z(n24746) );
  XOR U25007 ( .A(n24747), .B(n24749), .Z(n24748) );
  XOR U25008 ( .A(n24750), .B(n24751), .Z(n1258) );
  AND U25009 ( .A(n24752), .B(n24753), .Z(n24750) );
  XNOR U25010 ( .A(n24751), .B(n24717), .Z(n24753) );
  XNOR U25011 ( .A(n24754), .B(n24755), .Z(n24717) );
  ANDN U25012 ( .B(n24756), .A(n24757), .Z(n24754) );
  XOR U25013 ( .A(n24755), .B(n24758), .Z(n24756) );
  XOR U25014 ( .A(n24751), .B(n24719), .Z(n24752) );
  XOR U25015 ( .A(n24759), .B(n24760), .Z(n24719) );
  AND U25016 ( .A(n1262), .B(n24761), .Z(n24759) );
  XOR U25017 ( .A(n24762), .B(n24760), .Z(n24761) );
  XNOR U25018 ( .A(n24763), .B(n24764), .Z(n24751) );
  NAND U25019 ( .A(n24765), .B(n24766), .Z(n24764) );
  XOR U25020 ( .A(n24767), .B(n24743), .Z(n24766) );
  XOR U25021 ( .A(n24757), .B(n24758), .Z(n24743) );
  XOR U25022 ( .A(n24768), .B(n24769), .Z(n24758) );
  ANDN U25023 ( .B(n24770), .A(n24771), .Z(n24768) );
  XOR U25024 ( .A(n24769), .B(n24772), .Z(n24770) );
  XOR U25025 ( .A(n24773), .B(n24774), .Z(n24757) );
  XOR U25026 ( .A(n24775), .B(n24776), .Z(n24774) );
  ANDN U25027 ( .B(n24777), .A(n24778), .Z(n24775) );
  XOR U25028 ( .A(n24779), .B(n24776), .Z(n24777) );
  IV U25029 ( .A(n24755), .Z(n24773) );
  XOR U25030 ( .A(n24780), .B(n24781), .Z(n24755) );
  ANDN U25031 ( .B(n24782), .A(n24783), .Z(n24780) );
  XOR U25032 ( .A(n24781), .B(n24784), .Z(n24782) );
  IV U25033 ( .A(n24763), .Z(n24767) );
  XOR U25034 ( .A(n24763), .B(n24745), .Z(n24765) );
  XOR U25035 ( .A(n24785), .B(n24786), .Z(n24745) );
  AND U25036 ( .A(n1262), .B(n24787), .Z(n24785) );
  XOR U25037 ( .A(n24788), .B(n24786), .Z(n24787) );
  NANDN U25038 ( .A(n24747), .B(n24749), .Z(n24763) );
  XOR U25039 ( .A(n24789), .B(n24790), .Z(n24749) );
  AND U25040 ( .A(n1262), .B(n24791), .Z(n24789) );
  XOR U25041 ( .A(n24790), .B(n24792), .Z(n24791) );
  XOR U25042 ( .A(n24793), .B(n24794), .Z(n1262) );
  AND U25043 ( .A(n24795), .B(n24796), .Z(n24793) );
  XNOR U25044 ( .A(n24794), .B(n24760), .Z(n24796) );
  XNOR U25045 ( .A(n24797), .B(n24798), .Z(n24760) );
  ANDN U25046 ( .B(n24799), .A(n24800), .Z(n24797) );
  XOR U25047 ( .A(n24798), .B(n24801), .Z(n24799) );
  XOR U25048 ( .A(n24794), .B(n24762), .Z(n24795) );
  XOR U25049 ( .A(n24802), .B(n24803), .Z(n24762) );
  AND U25050 ( .A(n1266), .B(n24804), .Z(n24802) );
  XOR U25051 ( .A(n24805), .B(n24803), .Z(n24804) );
  XNOR U25052 ( .A(n24806), .B(n24807), .Z(n24794) );
  NAND U25053 ( .A(n24808), .B(n24809), .Z(n24807) );
  XOR U25054 ( .A(n24810), .B(n24786), .Z(n24809) );
  XOR U25055 ( .A(n24800), .B(n24801), .Z(n24786) );
  XOR U25056 ( .A(n24811), .B(n24812), .Z(n24801) );
  ANDN U25057 ( .B(n24813), .A(n24814), .Z(n24811) );
  XOR U25058 ( .A(n24812), .B(n24815), .Z(n24813) );
  XOR U25059 ( .A(n24816), .B(n24817), .Z(n24800) );
  XOR U25060 ( .A(n24818), .B(n24819), .Z(n24817) );
  ANDN U25061 ( .B(n24820), .A(n24821), .Z(n24818) );
  XOR U25062 ( .A(n24822), .B(n24819), .Z(n24820) );
  IV U25063 ( .A(n24798), .Z(n24816) );
  XOR U25064 ( .A(n24823), .B(n24824), .Z(n24798) );
  ANDN U25065 ( .B(n24825), .A(n24826), .Z(n24823) );
  XOR U25066 ( .A(n24824), .B(n24827), .Z(n24825) );
  IV U25067 ( .A(n24806), .Z(n24810) );
  XOR U25068 ( .A(n24806), .B(n24788), .Z(n24808) );
  XOR U25069 ( .A(n24828), .B(n24829), .Z(n24788) );
  AND U25070 ( .A(n1266), .B(n24830), .Z(n24828) );
  XOR U25071 ( .A(n24831), .B(n24829), .Z(n24830) );
  NANDN U25072 ( .A(n24790), .B(n24792), .Z(n24806) );
  XOR U25073 ( .A(n24832), .B(n24833), .Z(n24792) );
  AND U25074 ( .A(n1266), .B(n24834), .Z(n24832) );
  XOR U25075 ( .A(n24833), .B(n24835), .Z(n24834) );
  XOR U25076 ( .A(n24836), .B(n24837), .Z(n1266) );
  AND U25077 ( .A(n24838), .B(n24839), .Z(n24836) );
  XNOR U25078 ( .A(n24837), .B(n24803), .Z(n24839) );
  XNOR U25079 ( .A(n24840), .B(n24841), .Z(n24803) );
  ANDN U25080 ( .B(n24842), .A(n24843), .Z(n24840) );
  XOR U25081 ( .A(n24841), .B(n24844), .Z(n24842) );
  XOR U25082 ( .A(n24837), .B(n24805), .Z(n24838) );
  XOR U25083 ( .A(n24845), .B(n24846), .Z(n24805) );
  AND U25084 ( .A(n1270), .B(n24847), .Z(n24845) );
  XOR U25085 ( .A(n24848), .B(n24846), .Z(n24847) );
  XNOR U25086 ( .A(n24849), .B(n24850), .Z(n24837) );
  NAND U25087 ( .A(n24851), .B(n24852), .Z(n24850) );
  XOR U25088 ( .A(n24853), .B(n24829), .Z(n24852) );
  XOR U25089 ( .A(n24843), .B(n24844), .Z(n24829) );
  XOR U25090 ( .A(n24854), .B(n24855), .Z(n24844) );
  ANDN U25091 ( .B(n24856), .A(n24857), .Z(n24854) );
  XOR U25092 ( .A(n24855), .B(n24858), .Z(n24856) );
  XOR U25093 ( .A(n24859), .B(n24860), .Z(n24843) );
  XOR U25094 ( .A(n24861), .B(n24862), .Z(n24860) );
  ANDN U25095 ( .B(n24863), .A(n24864), .Z(n24861) );
  XOR U25096 ( .A(n24865), .B(n24862), .Z(n24863) );
  IV U25097 ( .A(n24841), .Z(n24859) );
  XOR U25098 ( .A(n24866), .B(n24867), .Z(n24841) );
  ANDN U25099 ( .B(n24868), .A(n24869), .Z(n24866) );
  XOR U25100 ( .A(n24867), .B(n24870), .Z(n24868) );
  IV U25101 ( .A(n24849), .Z(n24853) );
  XOR U25102 ( .A(n24849), .B(n24831), .Z(n24851) );
  XOR U25103 ( .A(n24871), .B(n24872), .Z(n24831) );
  AND U25104 ( .A(n1270), .B(n24873), .Z(n24871) );
  XOR U25105 ( .A(n24874), .B(n24872), .Z(n24873) );
  NANDN U25106 ( .A(n24833), .B(n24835), .Z(n24849) );
  XOR U25107 ( .A(n24875), .B(n24876), .Z(n24835) );
  AND U25108 ( .A(n1270), .B(n24877), .Z(n24875) );
  XOR U25109 ( .A(n24876), .B(n24878), .Z(n24877) );
  XOR U25110 ( .A(n24879), .B(n24880), .Z(n1270) );
  AND U25111 ( .A(n24881), .B(n24882), .Z(n24879) );
  XNOR U25112 ( .A(n24880), .B(n24846), .Z(n24882) );
  XNOR U25113 ( .A(n24883), .B(n24884), .Z(n24846) );
  ANDN U25114 ( .B(n24885), .A(n24886), .Z(n24883) );
  XOR U25115 ( .A(n24884), .B(n24887), .Z(n24885) );
  XOR U25116 ( .A(n24880), .B(n24848), .Z(n24881) );
  XOR U25117 ( .A(n24888), .B(n24889), .Z(n24848) );
  AND U25118 ( .A(n1274), .B(n24890), .Z(n24888) );
  XOR U25119 ( .A(n24891), .B(n24889), .Z(n24890) );
  XNOR U25120 ( .A(n24892), .B(n24893), .Z(n24880) );
  NAND U25121 ( .A(n24894), .B(n24895), .Z(n24893) );
  XOR U25122 ( .A(n24896), .B(n24872), .Z(n24895) );
  XOR U25123 ( .A(n24886), .B(n24887), .Z(n24872) );
  XOR U25124 ( .A(n24897), .B(n24898), .Z(n24887) );
  ANDN U25125 ( .B(n24899), .A(n24900), .Z(n24897) );
  XOR U25126 ( .A(n24898), .B(n24901), .Z(n24899) );
  XOR U25127 ( .A(n24902), .B(n24903), .Z(n24886) );
  XOR U25128 ( .A(n24904), .B(n24905), .Z(n24903) );
  ANDN U25129 ( .B(n24906), .A(n24907), .Z(n24904) );
  XOR U25130 ( .A(n24908), .B(n24905), .Z(n24906) );
  IV U25131 ( .A(n24884), .Z(n24902) );
  XOR U25132 ( .A(n24909), .B(n24910), .Z(n24884) );
  ANDN U25133 ( .B(n24911), .A(n24912), .Z(n24909) );
  XOR U25134 ( .A(n24910), .B(n24913), .Z(n24911) );
  IV U25135 ( .A(n24892), .Z(n24896) );
  XOR U25136 ( .A(n24892), .B(n24874), .Z(n24894) );
  XOR U25137 ( .A(n24914), .B(n24915), .Z(n24874) );
  AND U25138 ( .A(n1274), .B(n24916), .Z(n24914) );
  XOR U25139 ( .A(n24917), .B(n24915), .Z(n24916) );
  NANDN U25140 ( .A(n24876), .B(n24878), .Z(n24892) );
  XOR U25141 ( .A(n24918), .B(n24919), .Z(n24878) );
  AND U25142 ( .A(n1274), .B(n24920), .Z(n24918) );
  XOR U25143 ( .A(n24919), .B(n24921), .Z(n24920) );
  XOR U25144 ( .A(n24922), .B(n24923), .Z(n1274) );
  AND U25145 ( .A(n24924), .B(n24925), .Z(n24922) );
  XNOR U25146 ( .A(n24923), .B(n24889), .Z(n24925) );
  XNOR U25147 ( .A(n24926), .B(n24927), .Z(n24889) );
  ANDN U25148 ( .B(n24928), .A(n24929), .Z(n24926) );
  XOR U25149 ( .A(n24927), .B(n24930), .Z(n24928) );
  XOR U25150 ( .A(n24923), .B(n24891), .Z(n24924) );
  XOR U25151 ( .A(n24931), .B(n24932), .Z(n24891) );
  AND U25152 ( .A(n1278), .B(n24933), .Z(n24931) );
  XOR U25153 ( .A(n24934), .B(n24932), .Z(n24933) );
  XNOR U25154 ( .A(n24935), .B(n24936), .Z(n24923) );
  NAND U25155 ( .A(n24937), .B(n24938), .Z(n24936) );
  XOR U25156 ( .A(n24939), .B(n24915), .Z(n24938) );
  XOR U25157 ( .A(n24929), .B(n24930), .Z(n24915) );
  XOR U25158 ( .A(n24940), .B(n24941), .Z(n24930) );
  ANDN U25159 ( .B(n24942), .A(n24943), .Z(n24940) );
  XOR U25160 ( .A(n24941), .B(n24944), .Z(n24942) );
  XOR U25161 ( .A(n24945), .B(n24946), .Z(n24929) );
  XOR U25162 ( .A(n24947), .B(n24948), .Z(n24946) );
  ANDN U25163 ( .B(n24949), .A(n24950), .Z(n24947) );
  XOR U25164 ( .A(n24951), .B(n24948), .Z(n24949) );
  IV U25165 ( .A(n24927), .Z(n24945) );
  XOR U25166 ( .A(n24952), .B(n24953), .Z(n24927) );
  ANDN U25167 ( .B(n24954), .A(n24955), .Z(n24952) );
  XOR U25168 ( .A(n24953), .B(n24956), .Z(n24954) );
  IV U25169 ( .A(n24935), .Z(n24939) );
  XOR U25170 ( .A(n24935), .B(n24917), .Z(n24937) );
  XOR U25171 ( .A(n24957), .B(n24958), .Z(n24917) );
  AND U25172 ( .A(n1278), .B(n24959), .Z(n24957) );
  XOR U25173 ( .A(n24960), .B(n24958), .Z(n24959) );
  NANDN U25174 ( .A(n24919), .B(n24921), .Z(n24935) );
  XOR U25175 ( .A(n24961), .B(n24962), .Z(n24921) );
  AND U25176 ( .A(n1278), .B(n24963), .Z(n24961) );
  XOR U25177 ( .A(n24962), .B(n24964), .Z(n24963) );
  XOR U25178 ( .A(n24965), .B(n24966), .Z(n1278) );
  AND U25179 ( .A(n24967), .B(n24968), .Z(n24965) );
  XNOR U25180 ( .A(n24966), .B(n24932), .Z(n24968) );
  XNOR U25181 ( .A(n24969), .B(n24970), .Z(n24932) );
  ANDN U25182 ( .B(n24971), .A(n24972), .Z(n24969) );
  XOR U25183 ( .A(n24970), .B(n24973), .Z(n24971) );
  XOR U25184 ( .A(n24966), .B(n24934), .Z(n24967) );
  XOR U25185 ( .A(n24974), .B(n24975), .Z(n24934) );
  AND U25186 ( .A(n1282), .B(n24976), .Z(n24974) );
  XOR U25187 ( .A(n24977), .B(n24975), .Z(n24976) );
  XNOR U25188 ( .A(n24978), .B(n24979), .Z(n24966) );
  NAND U25189 ( .A(n24980), .B(n24981), .Z(n24979) );
  XOR U25190 ( .A(n24982), .B(n24958), .Z(n24981) );
  XOR U25191 ( .A(n24972), .B(n24973), .Z(n24958) );
  XOR U25192 ( .A(n24983), .B(n24984), .Z(n24973) );
  ANDN U25193 ( .B(n24985), .A(n24986), .Z(n24983) );
  XOR U25194 ( .A(n24984), .B(n24987), .Z(n24985) );
  XOR U25195 ( .A(n24988), .B(n24989), .Z(n24972) );
  XOR U25196 ( .A(n24990), .B(n24991), .Z(n24989) );
  ANDN U25197 ( .B(n24992), .A(n24993), .Z(n24990) );
  XOR U25198 ( .A(n24994), .B(n24991), .Z(n24992) );
  IV U25199 ( .A(n24970), .Z(n24988) );
  XOR U25200 ( .A(n24995), .B(n24996), .Z(n24970) );
  ANDN U25201 ( .B(n24997), .A(n24998), .Z(n24995) );
  XOR U25202 ( .A(n24996), .B(n24999), .Z(n24997) );
  IV U25203 ( .A(n24978), .Z(n24982) );
  XOR U25204 ( .A(n24978), .B(n24960), .Z(n24980) );
  XOR U25205 ( .A(n25000), .B(n25001), .Z(n24960) );
  AND U25206 ( .A(n1282), .B(n25002), .Z(n25000) );
  XOR U25207 ( .A(n25003), .B(n25001), .Z(n25002) );
  NANDN U25208 ( .A(n24962), .B(n24964), .Z(n24978) );
  XOR U25209 ( .A(n25004), .B(n25005), .Z(n24964) );
  AND U25210 ( .A(n1282), .B(n25006), .Z(n25004) );
  XOR U25211 ( .A(n25005), .B(n25007), .Z(n25006) );
  XOR U25212 ( .A(n25008), .B(n25009), .Z(n1282) );
  AND U25213 ( .A(n25010), .B(n25011), .Z(n25008) );
  XNOR U25214 ( .A(n25009), .B(n24975), .Z(n25011) );
  XNOR U25215 ( .A(n25012), .B(n25013), .Z(n24975) );
  ANDN U25216 ( .B(n25014), .A(n25015), .Z(n25012) );
  XOR U25217 ( .A(n25013), .B(n25016), .Z(n25014) );
  XOR U25218 ( .A(n25009), .B(n24977), .Z(n25010) );
  XOR U25219 ( .A(n25017), .B(n25018), .Z(n24977) );
  AND U25220 ( .A(n1286), .B(n25019), .Z(n25017) );
  XOR U25221 ( .A(n25020), .B(n25018), .Z(n25019) );
  XNOR U25222 ( .A(n25021), .B(n25022), .Z(n25009) );
  NAND U25223 ( .A(n25023), .B(n25024), .Z(n25022) );
  XOR U25224 ( .A(n25025), .B(n25001), .Z(n25024) );
  XOR U25225 ( .A(n25015), .B(n25016), .Z(n25001) );
  XOR U25226 ( .A(n25026), .B(n25027), .Z(n25016) );
  ANDN U25227 ( .B(n25028), .A(n25029), .Z(n25026) );
  XOR U25228 ( .A(n25027), .B(n25030), .Z(n25028) );
  XOR U25229 ( .A(n25031), .B(n25032), .Z(n25015) );
  XOR U25230 ( .A(n25033), .B(n25034), .Z(n25032) );
  ANDN U25231 ( .B(n25035), .A(n25036), .Z(n25033) );
  XOR U25232 ( .A(n25037), .B(n25034), .Z(n25035) );
  IV U25233 ( .A(n25013), .Z(n25031) );
  XOR U25234 ( .A(n25038), .B(n25039), .Z(n25013) );
  ANDN U25235 ( .B(n25040), .A(n25041), .Z(n25038) );
  XOR U25236 ( .A(n25039), .B(n25042), .Z(n25040) );
  IV U25237 ( .A(n25021), .Z(n25025) );
  XOR U25238 ( .A(n25021), .B(n25003), .Z(n25023) );
  XOR U25239 ( .A(n25043), .B(n25044), .Z(n25003) );
  AND U25240 ( .A(n1286), .B(n25045), .Z(n25043) );
  XOR U25241 ( .A(n25046), .B(n25044), .Z(n25045) );
  NANDN U25242 ( .A(n25005), .B(n25007), .Z(n25021) );
  XOR U25243 ( .A(n25047), .B(n25048), .Z(n25007) );
  AND U25244 ( .A(n1286), .B(n25049), .Z(n25047) );
  XOR U25245 ( .A(n25048), .B(n25050), .Z(n25049) );
  XOR U25246 ( .A(n25051), .B(n25052), .Z(n1286) );
  AND U25247 ( .A(n25053), .B(n25054), .Z(n25051) );
  XNOR U25248 ( .A(n25052), .B(n25018), .Z(n25054) );
  XNOR U25249 ( .A(n25055), .B(n25056), .Z(n25018) );
  ANDN U25250 ( .B(n25057), .A(n25058), .Z(n25055) );
  XOR U25251 ( .A(n25056), .B(n25059), .Z(n25057) );
  XOR U25252 ( .A(n25052), .B(n25020), .Z(n25053) );
  XOR U25253 ( .A(n25060), .B(n25061), .Z(n25020) );
  AND U25254 ( .A(n1290), .B(n25062), .Z(n25060) );
  XOR U25255 ( .A(n25063), .B(n25061), .Z(n25062) );
  XNOR U25256 ( .A(n25064), .B(n25065), .Z(n25052) );
  NAND U25257 ( .A(n25066), .B(n25067), .Z(n25065) );
  XOR U25258 ( .A(n25068), .B(n25044), .Z(n25067) );
  XOR U25259 ( .A(n25058), .B(n25059), .Z(n25044) );
  XOR U25260 ( .A(n25069), .B(n25070), .Z(n25059) );
  ANDN U25261 ( .B(n25071), .A(n25072), .Z(n25069) );
  XOR U25262 ( .A(n25070), .B(n25073), .Z(n25071) );
  XOR U25263 ( .A(n25074), .B(n25075), .Z(n25058) );
  XOR U25264 ( .A(n25076), .B(n25077), .Z(n25075) );
  ANDN U25265 ( .B(n25078), .A(n25079), .Z(n25076) );
  XOR U25266 ( .A(n25080), .B(n25077), .Z(n25078) );
  IV U25267 ( .A(n25056), .Z(n25074) );
  XOR U25268 ( .A(n25081), .B(n25082), .Z(n25056) );
  ANDN U25269 ( .B(n25083), .A(n25084), .Z(n25081) );
  XOR U25270 ( .A(n25082), .B(n25085), .Z(n25083) );
  IV U25271 ( .A(n25064), .Z(n25068) );
  XOR U25272 ( .A(n25064), .B(n25046), .Z(n25066) );
  XOR U25273 ( .A(n25086), .B(n25087), .Z(n25046) );
  AND U25274 ( .A(n1290), .B(n25088), .Z(n25086) );
  XOR U25275 ( .A(n25089), .B(n25087), .Z(n25088) );
  NANDN U25276 ( .A(n25048), .B(n25050), .Z(n25064) );
  XOR U25277 ( .A(n25090), .B(n25091), .Z(n25050) );
  AND U25278 ( .A(n1290), .B(n25092), .Z(n25090) );
  XOR U25279 ( .A(n25091), .B(n25093), .Z(n25092) );
  XOR U25280 ( .A(n25094), .B(n25095), .Z(n1290) );
  AND U25281 ( .A(n25096), .B(n25097), .Z(n25094) );
  XNOR U25282 ( .A(n25095), .B(n25061), .Z(n25097) );
  XNOR U25283 ( .A(n25098), .B(n25099), .Z(n25061) );
  ANDN U25284 ( .B(n25100), .A(n25101), .Z(n25098) );
  XOR U25285 ( .A(n25099), .B(n25102), .Z(n25100) );
  XOR U25286 ( .A(n25095), .B(n25063), .Z(n25096) );
  XOR U25287 ( .A(n25103), .B(n25104), .Z(n25063) );
  AND U25288 ( .A(n1294), .B(n25105), .Z(n25103) );
  XOR U25289 ( .A(n25106), .B(n25104), .Z(n25105) );
  XNOR U25290 ( .A(n25107), .B(n25108), .Z(n25095) );
  NAND U25291 ( .A(n25109), .B(n25110), .Z(n25108) );
  XOR U25292 ( .A(n25111), .B(n25087), .Z(n25110) );
  XOR U25293 ( .A(n25101), .B(n25102), .Z(n25087) );
  XOR U25294 ( .A(n25112), .B(n25113), .Z(n25102) );
  ANDN U25295 ( .B(n25114), .A(n25115), .Z(n25112) );
  XOR U25296 ( .A(n25113), .B(n25116), .Z(n25114) );
  XOR U25297 ( .A(n25117), .B(n25118), .Z(n25101) );
  XOR U25298 ( .A(n25119), .B(n25120), .Z(n25118) );
  ANDN U25299 ( .B(n25121), .A(n25122), .Z(n25119) );
  XOR U25300 ( .A(n25123), .B(n25120), .Z(n25121) );
  IV U25301 ( .A(n25099), .Z(n25117) );
  XOR U25302 ( .A(n25124), .B(n25125), .Z(n25099) );
  ANDN U25303 ( .B(n25126), .A(n25127), .Z(n25124) );
  XOR U25304 ( .A(n25125), .B(n25128), .Z(n25126) );
  IV U25305 ( .A(n25107), .Z(n25111) );
  XOR U25306 ( .A(n25107), .B(n25089), .Z(n25109) );
  XOR U25307 ( .A(n25129), .B(n25130), .Z(n25089) );
  AND U25308 ( .A(n1294), .B(n25131), .Z(n25129) );
  XOR U25309 ( .A(n25132), .B(n25130), .Z(n25131) );
  NANDN U25310 ( .A(n25091), .B(n25093), .Z(n25107) );
  XOR U25311 ( .A(n25133), .B(n25134), .Z(n25093) );
  AND U25312 ( .A(n1294), .B(n25135), .Z(n25133) );
  XOR U25313 ( .A(n25134), .B(n25136), .Z(n25135) );
  XOR U25314 ( .A(n25137), .B(n25138), .Z(n1294) );
  AND U25315 ( .A(n25139), .B(n25140), .Z(n25137) );
  XNOR U25316 ( .A(n25138), .B(n25104), .Z(n25140) );
  XNOR U25317 ( .A(n25141), .B(n25142), .Z(n25104) );
  ANDN U25318 ( .B(n25143), .A(n25144), .Z(n25141) );
  XOR U25319 ( .A(n25142), .B(n25145), .Z(n25143) );
  XOR U25320 ( .A(n25138), .B(n25106), .Z(n25139) );
  XOR U25321 ( .A(n25146), .B(n25147), .Z(n25106) );
  AND U25322 ( .A(n1298), .B(n25148), .Z(n25146) );
  XOR U25323 ( .A(n25149), .B(n25147), .Z(n25148) );
  XNOR U25324 ( .A(n25150), .B(n25151), .Z(n25138) );
  NAND U25325 ( .A(n25152), .B(n25153), .Z(n25151) );
  XOR U25326 ( .A(n25154), .B(n25130), .Z(n25153) );
  XOR U25327 ( .A(n25144), .B(n25145), .Z(n25130) );
  XOR U25328 ( .A(n25155), .B(n25156), .Z(n25145) );
  ANDN U25329 ( .B(n25157), .A(n25158), .Z(n25155) );
  XOR U25330 ( .A(n25156), .B(n25159), .Z(n25157) );
  XOR U25331 ( .A(n25160), .B(n25161), .Z(n25144) );
  XOR U25332 ( .A(n25162), .B(n25163), .Z(n25161) );
  ANDN U25333 ( .B(n25164), .A(n25165), .Z(n25162) );
  XOR U25334 ( .A(n25166), .B(n25163), .Z(n25164) );
  IV U25335 ( .A(n25142), .Z(n25160) );
  XOR U25336 ( .A(n25167), .B(n25168), .Z(n25142) );
  ANDN U25337 ( .B(n25169), .A(n25170), .Z(n25167) );
  XOR U25338 ( .A(n25168), .B(n25171), .Z(n25169) );
  IV U25339 ( .A(n25150), .Z(n25154) );
  XOR U25340 ( .A(n25150), .B(n25132), .Z(n25152) );
  XOR U25341 ( .A(n25172), .B(n25173), .Z(n25132) );
  AND U25342 ( .A(n1298), .B(n25174), .Z(n25172) );
  XOR U25343 ( .A(n25175), .B(n25173), .Z(n25174) );
  NANDN U25344 ( .A(n25134), .B(n25136), .Z(n25150) );
  XOR U25345 ( .A(n25176), .B(n25177), .Z(n25136) );
  AND U25346 ( .A(n1298), .B(n25178), .Z(n25176) );
  XOR U25347 ( .A(n25177), .B(n25179), .Z(n25178) );
  XOR U25348 ( .A(n25180), .B(n25181), .Z(n1298) );
  AND U25349 ( .A(n25182), .B(n25183), .Z(n25180) );
  XNOR U25350 ( .A(n25181), .B(n25147), .Z(n25183) );
  XNOR U25351 ( .A(n25184), .B(n25185), .Z(n25147) );
  ANDN U25352 ( .B(n25186), .A(n25187), .Z(n25184) );
  XOR U25353 ( .A(n25185), .B(n25188), .Z(n25186) );
  XOR U25354 ( .A(n25181), .B(n25149), .Z(n25182) );
  XOR U25355 ( .A(n25189), .B(n25190), .Z(n25149) );
  AND U25356 ( .A(n1302), .B(n25191), .Z(n25189) );
  XOR U25357 ( .A(n25192), .B(n25190), .Z(n25191) );
  XNOR U25358 ( .A(n25193), .B(n25194), .Z(n25181) );
  NAND U25359 ( .A(n25195), .B(n25196), .Z(n25194) );
  XOR U25360 ( .A(n25197), .B(n25173), .Z(n25196) );
  XOR U25361 ( .A(n25187), .B(n25188), .Z(n25173) );
  XOR U25362 ( .A(n25198), .B(n25199), .Z(n25188) );
  ANDN U25363 ( .B(n25200), .A(n25201), .Z(n25198) );
  XOR U25364 ( .A(n25199), .B(n25202), .Z(n25200) );
  XOR U25365 ( .A(n25203), .B(n25204), .Z(n25187) );
  XOR U25366 ( .A(n25205), .B(n25206), .Z(n25204) );
  ANDN U25367 ( .B(n25207), .A(n25208), .Z(n25205) );
  XOR U25368 ( .A(n25209), .B(n25206), .Z(n25207) );
  IV U25369 ( .A(n25185), .Z(n25203) );
  XOR U25370 ( .A(n25210), .B(n25211), .Z(n25185) );
  ANDN U25371 ( .B(n25212), .A(n25213), .Z(n25210) );
  XOR U25372 ( .A(n25211), .B(n25214), .Z(n25212) );
  IV U25373 ( .A(n25193), .Z(n25197) );
  XOR U25374 ( .A(n25193), .B(n25175), .Z(n25195) );
  XOR U25375 ( .A(n25215), .B(n25216), .Z(n25175) );
  AND U25376 ( .A(n1302), .B(n25217), .Z(n25215) );
  XOR U25377 ( .A(n25218), .B(n25216), .Z(n25217) );
  NANDN U25378 ( .A(n25177), .B(n25179), .Z(n25193) );
  XOR U25379 ( .A(n25219), .B(n25220), .Z(n25179) );
  AND U25380 ( .A(n1302), .B(n25221), .Z(n25219) );
  XOR U25381 ( .A(n25220), .B(n25222), .Z(n25221) );
  XOR U25382 ( .A(n25223), .B(n25224), .Z(n1302) );
  AND U25383 ( .A(n25225), .B(n25226), .Z(n25223) );
  XNOR U25384 ( .A(n25224), .B(n25190), .Z(n25226) );
  XNOR U25385 ( .A(n25227), .B(n25228), .Z(n25190) );
  ANDN U25386 ( .B(n25229), .A(n25230), .Z(n25227) );
  XOR U25387 ( .A(n25228), .B(n25231), .Z(n25229) );
  XOR U25388 ( .A(n25224), .B(n25192), .Z(n25225) );
  XOR U25389 ( .A(n25232), .B(n25233), .Z(n25192) );
  AND U25390 ( .A(n1306), .B(n25234), .Z(n25232) );
  XOR U25391 ( .A(n25235), .B(n25233), .Z(n25234) );
  XNOR U25392 ( .A(n25236), .B(n25237), .Z(n25224) );
  NAND U25393 ( .A(n25238), .B(n25239), .Z(n25237) );
  XOR U25394 ( .A(n25240), .B(n25216), .Z(n25239) );
  XOR U25395 ( .A(n25230), .B(n25231), .Z(n25216) );
  XOR U25396 ( .A(n25241), .B(n25242), .Z(n25231) );
  ANDN U25397 ( .B(n25243), .A(n25244), .Z(n25241) );
  XOR U25398 ( .A(n25242), .B(n25245), .Z(n25243) );
  XOR U25399 ( .A(n25246), .B(n25247), .Z(n25230) );
  XOR U25400 ( .A(n25248), .B(n25249), .Z(n25247) );
  ANDN U25401 ( .B(n25250), .A(n25251), .Z(n25248) );
  XOR U25402 ( .A(n25252), .B(n25249), .Z(n25250) );
  IV U25403 ( .A(n25228), .Z(n25246) );
  XOR U25404 ( .A(n25253), .B(n25254), .Z(n25228) );
  ANDN U25405 ( .B(n25255), .A(n25256), .Z(n25253) );
  XOR U25406 ( .A(n25254), .B(n25257), .Z(n25255) );
  IV U25407 ( .A(n25236), .Z(n25240) );
  XOR U25408 ( .A(n25236), .B(n25218), .Z(n25238) );
  XOR U25409 ( .A(n25258), .B(n25259), .Z(n25218) );
  AND U25410 ( .A(n1306), .B(n25260), .Z(n25258) );
  XOR U25411 ( .A(n25261), .B(n25259), .Z(n25260) );
  NANDN U25412 ( .A(n25220), .B(n25222), .Z(n25236) );
  XOR U25413 ( .A(n25262), .B(n25263), .Z(n25222) );
  AND U25414 ( .A(n1306), .B(n25264), .Z(n25262) );
  XOR U25415 ( .A(n25263), .B(n25265), .Z(n25264) );
  XOR U25416 ( .A(n25266), .B(n25267), .Z(n1306) );
  AND U25417 ( .A(n25268), .B(n25269), .Z(n25266) );
  XNOR U25418 ( .A(n25267), .B(n25233), .Z(n25269) );
  XNOR U25419 ( .A(n25270), .B(n25271), .Z(n25233) );
  ANDN U25420 ( .B(n25272), .A(n25273), .Z(n25270) );
  XOR U25421 ( .A(n25271), .B(n25274), .Z(n25272) );
  XOR U25422 ( .A(n25267), .B(n25235), .Z(n25268) );
  XOR U25423 ( .A(n25275), .B(n25276), .Z(n25235) );
  AND U25424 ( .A(n1310), .B(n25277), .Z(n25275) );
  XOR U25425 ( .A(n25278), .B(n25276), .Z(n25277) );
  XNOR U25426 ( .A(n25279), .B(n25280), .Z(n25267) );
  NAND U25427 ( .A(n25281), .B(n25282), .Z(n25280) );
  XOR U25428 ( .A(n25283), .B(n25259), .Z(n25282) );
  XOR U25429 ( .A(n25273), .B(n25274), .Z(n25259) );
  XOR U25430 ( .A(n25284), .B(n25285), .Z(n25274) );
  ANDN U25431 ( .B(n25286), .A(n25287), .Z(n25284) );
  XOR U25432 ( .A(n25285), .B(n25288), .Z(n25286) );
  XOR U25433 ( .A(n25289), .B(n25290), .Z(n25273) );
  XOR U25434 ( .A(n25291), .B(n25292), .Z(n25290) );
  ANDN U25435 ( .B(n25293), .A(n25294), .Z(n25291) );
  XOR U25436 ( .A(n25295), .B(n25292), .Z(n25293) );
  IV U25437 ( .A(n25271), .Z(n25289) );
  XOR U25438 ( .A(n25296), .B(n25297), .Z(n25271) );
  ANDN U25439 ( .B(n25298), .A(n25299), .Z(n25296) );
  XOR U25440 ( .A(n25297), .B(n25300), .Z(n25298) );
  IV U25441 ( .A(n25279), .Z(n25283) );
  XOR U25442 ( .A(n25279), .B(n25261), .Z(n25281) );
  XOR U25443 ( .A(n25301), .B(n25302), .Z(n25261) );
  AND U25444 ( .A(n1310), .B(n25303), .Z(n25301) );
  XOR U25445 ( .A(n25304), .B(n25302), .Z(n25303) );
  NANDN U25446 ( .A(n25263), .B(n25265), .Z(n25279) );
  XOR U25447 ( .A(n25305), .B(n25306), .Z(n25265) );
  AND U25448 ( .A(n1310), .B(n25307), .Z(n25305) );
  XOR U25449 ( .A(n25306), .B(n25308), .Z(n25307) );
  XOR U25450 ( .A(n25309), .B(n25310), .Z(n1310) );
  AND U25451 ( .A(n25311), .B(n25312), .Z(n25309) );
  XNOR U25452 ( .A(n25310), .B(n25276), .Z(n25312) );
  XNOR U25453 ( .A(n25313), .B(n25314), .Z(n25276) );
  ANDN U25454 ( .B(n25315), .A(n25316), .Z(n25313) );
  XOR U25455 ( .A(n25314), .B(n25317), .Z(n25315) );
  XOR U25456 ( .A(n25310), .B(n25278), .Z(n25311) );
  XOR U25457 ( .A(n25318), .B(n25319), .Z(n25278) );
  AND U25458 ( .A(n1314), .B(n25320), .Z(n25318) );
  XOR U25459 ( .A(n25321), .B(n25319), .Z(n25320) );
  XNOR U25460 ( .A(n25322), .B(n25323), .Z(n25310) );
  NAND U25461 ( .A(n25324), .B(n25325), .Z(n25323) );
  XOR U25462 ( .A(n25326), .B(n25302), .Z(n25325) );
  XOR U25463 ( .A(n25316), .B(n25317), .Z(n25302) );
  XOR U25464 ( .A(n25327), .B(n25328), .Z(n25317) );
  ANDN U25465 ( .B(n25329), .A(n25330), .Z(n25327) );
  XOR U25466 ( .A(n25328), .B(n25331), .Z(n25329) );
  XOR U25467 ( .A(n25332), .B(n25333), .Z(n25316) );
  XOR U25468 ( .A(n25334), .B(n25335), .Z(n25333) );
  ANDN U25469 ( .B(n25336), .A(n25337), .Z(n25334) );
  XOR U25470 ( .A(n25338), .B(n25335), .Z(n25336) );
  IV U25471 ( .A(n25314), .Z(n25332) );
  XOR U25472 ( .A(n25339), .B(n25340), .Z(n25314) );
  ANDN U25473 ( .B(n25341), .A(n25342), .Z(n25339) );
  XOR U25474 ( .A(n25340), .B(n25343), .Z(n25341) );
  IV U25475 ( .A(n25322), .Z(n25326) );
  XOR U25476 ( .A(n25322), .B(n25304), .Z(n25324) );
  XOR U25477 ( .A(n25344), .B(n25345), .Z(n25304) );
  AND U25478 ( .A(n1314), .B(n25346), .Z(n25344) );
  XOR U25479 ( .A(n25347), .B(n25345), .Z(n25346) );
  NANDN U25480 ( .A(n25306), .B(n25308), .Z(n25322) );
  XOR U25481 ( .A(n25348), .B(n25349), .Z(n25308) );
  AND U25482 ( .A(n1314), .B(n25350), .Z(n25348) );
  XOR U25483 ( .A(n25349), .B(n25351), .Z(n25350) );
  XOR U25484 ( .A(n25352), .B(n25353), .Z(n1314) );
  AND U25485 ( .A(n25354), .B(n25355), .Z(n25352) );
  XNOR U25486 ( .A(n25353), .B(n25319), .Z(n25355) );
  XNOR U25487 ( .A(n25356), .B(n25357), .Z(n25319) );
  ANDN U25488 ( .B(n25358), .A(n25359), .Z(n25356) );
  XOR U25489 ( .A(n25357), .B(n25360), .Z(n25358) );
  XOR U25490 ( .A(n25353), .B(n25321), .Z(n25354) );
  XOR U25491 ( .A(n25361), .B(n25362), .Z(n25321) );
  AND U25492 ( .A(n1318), .B(n25363), .Z(n25361) );
  XOR U25493 ( .A(n25364), .B(n25362), .Z(n25363) );
  XNOR U25494 ( .A(n25365), .B(n25366), .Z(n25353) );
  NAND U25495 ( .A(n25367), .B(n25368), .Z(n25366) );
  XOR U25496 ( .A(n25369), .B(n25345), .Z(n25368) );
  XOR U25497 ( .A(n25359), .B(n25360), .Z(n25345) );
  XOR U25498 ( .A(n25370), .B(n25371), .Z(n25360) );
  ANDN U25499 ( .B(n25372), .A(n25373), .Z(n25370) );
  XOR U25500 ( .A(n25371), .B(n25374), .Z(n25372) );
  XOR U25501 ( .A(n25375), .B(n25376), .Z(n25359) );
  XOR U25502 ( .A(n25377), .B(n25378), .Z(n25376) );
  ANDN U25503 ( .B(n25379), .A(n25380), .Z(n25377) );
  XOR U25504 ( .A(n25381), .B(n25378), .Z(n25379) );
  IV U25505 ( .A(n25357), .Z(n25375) );
  XOR U25506 ( .A(n25382), .B(n25383), .Z(n25357) );
  ANDN U25507 ( .B(n25384), .A(n25385), .Z(n25382) );
  XOR U25508 ( .A(n25383), .B(n25386), .Z(n25384) );
  IV U25509 ( .A(n25365), .Z(n25369) );
  XOR U25510 ( .A(n25365), .B(n25347), .Z(n25367) );
  XOR U25511 ( .A(n25387), .B(n25388), .Z(n25347) );
  AND U25512 ( .A(n1318), .B(n25389), .Z(n25387) );
  XOR U25513 ( .A(n25390), .B(n25388), .Z(n25389) );
  NANDN U25514 ( .A(n25349), .B(n25351), .Z(n25365) );
  XOR U25515 ( .A(n25391), .B(n25392), .Z(n25351) );
  AND U25516 ( .A(n1318), .B(n25393), .Z(n25391) );
  XOR U25517 ( .A(n25392), .B(n25394), .Z(n25393) );
  XOR U25518 ( .A(n25395), .B(n25396), .Z(n1318) );
  AND U25519 ( .A(n25397), .B(n25398), .Z(n25395) );
  XNOR U25520 ( .A(n25396), .B(n25362), .Z(n25398) );
  XNOR U25521 ( .A(n25399), .B(n25400), .Z(n25362) );
  ANDN U25522 ( .B(n25401), .A(n25402), .Z(n25399) );
  XOR U25523 ( .A(n25400), .B(n25403), .Z(n25401) );
  XOR U25524 ( .A(n25396), .B(n25364), .Z(n25397) );
  XOR U25525 ( .A(n25404), .B(n25405), .Z(n25364) );
  AND U25526 ( .A(n1322), .B(n25406), .Z(n25404) );
  XOR U25527 ( .A(n25407), .B(n25405), .Z(n25406) );
  XNOR U25528 ( .A(n25408), .B(n25409), .Z(n25396) );
  NAND U25529 ( .A(n25410), .B(n25411), .Z(n25409) );
  XOR U25530 ( .A(n25412), .B(n25388), .Z(n25411) );
  XOR U25531 ( .A(n25402), .B(n25403), .Z(n25388) );
  XOR U25532 ( .A(n25413), .B(n25414), .Z(n25403) );
  ANDN U25533 ( .B(n25415), .A(n25416), .Z(n25413) );
  XOR U25534 ( .A(n25414), .B(n25417), .Z(n25415) );
  XOR U25535 ( .A(n25418), .B(n25419), .Z(n25402) );
  XOR U25536 ( .A(n25420), .B(n25421), .Z(n25419) );
  ANDN U25537 ( .B(n25422), .A(n25423), .Z(n25420) );
  XOR U25538 ( .A(n25424), .B(n25421), .Z(n25422) );
  IV U25539 ( .A(n25400), .Z(n25418) );
  XOR U25540 ( .A(n25425), .B(n25426), .Z(n25400) );
  ANDN U25541 ( .B(n25427), .A(n25428), .Z(n25425) );
  XOR U25542 ( .A(n25426), .B(n25429), .Z(n25427) );
  IV U25543 ( .A(n25408), .Z(n25412) );
  XOR U25544 ( .A(n25408), .B(n25390), .Z(n25410) );
  XOR U25545 ( .A(n25430), .B(n25431), .Z(n25390) );
  AND U25546 ( .A(n1322), .B(n25432), .Z(n25430) );
  XOR U25547 ( .A(n25433), .B(n25431), .Z(n25432) );
  NANDN U25548 ( .A(n25392), .B(n25394), .Z(n25408) );
  XOR U25549 ( .A(n25434), .B(n25435), .Z(n25394) );
  AND U25550 ( .A(n1322), .B(n25436), .Z(n25434) );
  XOR U25551 ( .A(n25435), .B(n25437), .Z(n25436) );
  XOR U25552 ( .A(n25438), .B(n25439), .Z(n1322) );
  AND U25553 ( .A(n25440), .B(n25441), .Z(n25438) );
  XNOR U25554 ( .A(n25439), .B(n25405), .Z(n25441) );
  XNOR U25555 ( .A(n25442), .B(n25443), .Z(n25405) );
  ANDN U25556 ( .B(n25444), .A(n25445), .Z(n25442) );
  XOR U25557 ( .A(n25443), .B(n25446), .Z(n25444) );
  XOR U25558 ( .A(n25439), .B(n25407), .Z(n25440) );
  XOR U25559 ( .A(n25447), .B(n25448), .Z(n25407) );
  AND U25560 ( .A(n1326), .B(n25449), .Z(n25447) );
  XOR U25561 ( .A(n25450), .B(n25448), .Z(n25449) );
  XNOR U25562 ( .A(n25451), .B(n25452), .Z(n25439) );
  NAND U25563 ( .A(n25453), .B(n25454), .Z(n25452) );
  XOR U25564 ( .A(n25455), .B(n25431), .Z(n25454) );
  XOR U25565 ( .A(n25445), .B(n25446), .Z(n25431) );
  XOR U25566 ( .A(n25456), .B(n25457), .Z(n25446) );
  ANDN U25567 ( .B(n25458), .A(n25459), .Z(n25456) );
  XOR U25568 ( .A(n25457), .B(n25460), .Z(n25458) );
  XOR U25569 ( .A(n25461), .B(n25462), .Z(n25445) );
  XOR U25570 ( .A(n25463), .B(n25464), .Z(n25462) );
  ANDN U25571 ( .B(n25465), .A(n25466), .Z(n25463) );
  XOR U25572 ( .A(n25467), .B(n25464), .Z(n25465) );
  IV U25573 ( .A(n25443), .Z(n25461) );
  XOR U25574 ( .A(n25468), .B(n25469), .Z(n25443) );
  ANDN U25575 ( .B(n25470), .A(n25471), .Z(n25468) );
  XOR U25576 ( .A(n25469), .B(n25472), .Z(n25470) );
  IV U25577 ( .A(n25451), .Z(n25455) );
  XOR U25578 ( .A(n25451), .B(n25433), .Z(n25453) );
  XOR U25579 ( .A(n25473), .B(n25474), .Z(n25433) );
  AND U25580 ( .A(n1326), .B(n25475), .Z(n25473) );
  XOR U25581 ( .A(n25476), .B(n25474), .Z(n25475) );
  NANDN U25582 ( .A(n25435), .B(n25437), .Z(n25451) );
  XOR U25583 ( .A(n25477), .B(n25478), .Z(n25437) );
  AND U25584 ( .A(n1326), .B(n25479), .Z(n25477) );
  XOR U25585 ( .A(n25478), .B(n25480), .Z(n25479) );
  XOR U25586 ( .A(n25481), .B(n25482), .Z(n1326) );
  AND U25587 ( .A(n25483), .B(n25484), .Z(n25481) );
  XNOR U25588 ( .A(n25482), .B(n25448), .Z(n25484) );
  XNOR U25589 ( .A(n25485), .B(n25486), .Z(n25448) );
  ANDN U25590 ( .B(n25487), .A(n25488), .Z(n25485) );
  XOR U25591 ( .A(n25486), .B(n25489), .Z(n25487) );
  XOR U25592 ( .A(n25482), .B(n25450), .Z(n25483) );
  XOR U25593 ( .A(n25490), .B(n25491), .Z(n25450) );
  AND U25594 ( .A(n1330), .B(n25492), .Z(n25490) );
  XOR U25595 ( .A(n25493), .B(n25491), .Z(n25492) );
  XNOR U25596 ( .A(n25494), .B(n25495), .Z(n25482) );
  NAND U25597 ( .A(n25496), .B(n25497), .Z(n25495) );
  XOR U25598 ( .A(n25498), .B(n25474), .Z(n25497) );
  XOR U25599 ( .A(n25488), .B(n25489), .Z(n25474) );
  XOR U25600 ( .A(n25499), .B(n25500), .Z(n25489) );
  ANDN U25601 ( .B(n25501), .A(n25502), .Z(n25499) );
  XOR U25602 ( .A(n25500), .B(n25503), .Z(n25501) );
  XOR U25603 ( .A(n25504), .B(n25505), .Z(n25488) );
  XOR U25604 ( .A(n25506), .B(n25507), .Z(n25505) );
  ANDN U25605 ( .B(n25508), .A(n25509), .Z(n25506) );
  XOR U25606 ( .A(n25510), .B(n25507), .Z(n25508) );
  IV U25607 ( .A(n25486), .Z(n25504) );
  XOR U25608 ( .A(n25511), .B(n25512), .Z(n25486) );
  ANDN U25609 ( .B(n25513), .A(n25514), .Z(n25511) );
  XOR U25610 ( .A(n25512), .B(n25515), .Z(n25513) );
  IV U25611 ( .A(n25494), .Z(n25498) );
  XOR U25612 ( .A(n25494), .B(n25476), .Z(n25496) );
  XOR U25613 ( .A(n25516), .B(n25517), .Z(n25476) );
  AND U25614 ( .A(n1330), .B(n25518), .Z(n25516) );
  XOR U25615 ( .A(n25519), .B(n25517), .Z(n25518) );
  NANDN U25616 ( .A(n25478), .B(n25480), .Z(n25494) );
  XOR U25617 ( .A(n25520), .B(n25521), .Z(n25480) );
  AND U25618 ( .A(n1330), .B(n25522), .Z(n25520) );
  XOR U25619 ( .A(n25521), .B(n25523), .Z(n25522) );
  XOR U25620 ( .A(n25524), .B(n25525), .Z(n1330) );
  AND U25621 ( .A(n25526), .B(n25527), .Z(n25524) );
  XNOR U25622 ( .A(n25525), .B(n25491), .Z(n25527) );
  XNOR U25623 ( .A(n25528), .B(n25529), .Z(n25491) );
  ANDN U25624 ( .B(n25530), .A(n25531), .Z(n25528) );
  XOR U25625 ( .A(n25529), .B(n25532), .Z(n25530) );
  XOR U25626 ( .A(n25525), .B(n25493), .Z(n25526) );
  XOR U25627 ( .A(n25533), .B(n25534), .Z(n25493) );
  AND U25628 ( .A(n1334), .B(n25535), .Z(n25533) );
  XOR U25629 ( .A(n25536), .B(n25534), .Z(n25535) );
  XNOR U25630 ( .A(n25537), .B(n25538), .Z(n25525) );
  NAND U25631 ( .A(n25539), .B(n25540), .Z(n25538) );
  XOR U25632 ( .A(n25541), .B(n25517), .Z(n25540) );
  XOR U25633 ( .A(n25531), .B(n25532), .Z(n25517) );
  XOR U25634 ( .A(n25542), .B(n25543), .Z(n25532) );
  ANDN U25635 ( .B(n25544), .A(n25545), .Z(n25542) );
  XOR U25636 ( .A(n25543), .B(n25546), .Z(n25544) );
  XOR U25637 ( .A(n25547), .B(n25548), .Z(n25531) );
  XOR U25638 ( .A(n25549), .B(n25550), .Z(n25548) );
  ANDN U25639 ( .B(n25551), .A(n25552), .Z(n25549) );
  XOR U25640 ( .A(n25553), .B(n25550), .Z(n25551) );
  IV U25641 ( .A(n25529), .Z(n25547) );
  XOR U25642 ( .A(n25554), .B(n25555), .Z(n25529) );
  ANDN U25643 ( .B(n25556), .A(n25557), .Z(n25554) );
  XOR U25644 ( .A(n25555), .B(n25558), .Z(n25556) );
  IV U25645 ( .A(n25537), .Z(n25541) );
  XOR U25646 ( .A(n25537), .B(n25519), .Z(n25539) );
  XOR U25647 ( .A(n25559), .B(n25560), .Z(n25519) );
  AND U25648 ( .A(n1334), .B(n25561), .Z(n25559) );
  XOR U25649 ( .A(n25562), .B(n25560), .Z(n25561) );
  NANDN U25650 ( .A(n25521), .B(n25523), .Z(n25537) );
  XOR U25651 ( .A(n25563), .B(n25564), .Z(n25523) );
  AND U25652 ( .A(n1334), .B(n25565), .Z(n25563) );
  XOR U25653 ( .A(n25564), .B(n25566), .Z(n25565) );
  XOR U25654 ( .A(n25567), .B(n25568), .Z(n1334) );
  AND U25655 ( .A(n25569), .B(n25570), .Z(n25567) );
  XNOR U25656 ( .A(n25568), .B(n25534), .Z(n25570) );
  XNOR U25657 ( .A(n25571), .B(n25572), .Z(n25534) );
  ANDN U25658 ( .B(n25573), .A(n25574), .Z(n25571) );
  XOR U25659 ( .A(n25572), .B(n25575), .Z(n25573) );
  XOR U25660 ( .A(n25568), .B(n25536), .Z(n25569) );
  XOR U25661 ( .A(n25576), .B(n25577), .Z(n25536) );
  AND U25662 ( .A(n1338), .B(n25578), .Z(n25576) );
  XOR U25663 ( .A(n25579), .B(n25577), .Z(n25578) );
  XNOR U25664 ( .A(n25580), .B(n25581), .Z(n25568) );
  NAND U25665 ( .A(n25582), .B(n25583), .Z(n25581) );
  XOR U25666 ( .A(n25584), .B(n25560), .Z(n25583) );
  XOR U25667 ( .A(n25574), .B(n25575), .Z(n25560) );
  XOR U25668 ( .A(n25585), .B(n25586), .Z(n25575) );
  ANDN U25669 ( .B(n25587), .A(n25588), .Z(n25585) );
  XOR U25670 ( .A(n25586), .B(n25589), .Z(n25587) );
  XOR U25671 ( .A(n25590), .B(n25591), .Z(n25574) );
  XOR U25672 ( .A(n25592), .B(n25593), .Z(n25591) );
  ANDN U25673 ( .B(n25594), .A(n25595), .Z(n25592) );
  XOR U25674 ( .A(n25596), .B(n25593), .Z(n25594) );
  IV U25675 ( .A(n25572), .Z(n25590) );
  XOR U25676 ( .A(n25597), .B(n25598), .Z(n25572) );
  ANDN U25677 ( .B(n25599), .A(n25600), .Z(n25597) );
  XOR U25678 ( .A(n25598), .B(n25601), .Z(n25599) );
  IV U25679 ( .A(n25580), .Z(n25584) );
  XOR U25680 ( .A(n25580), .B(n25562), .Z(n25582) );
  XOR U25681 ( .A(n25602), .B(n25603), .Z(n25562) );
  AND U25682 ( .A(n1338), .B(n25604), .Z(n25602) );
  XOR U25683 ( .A(n25605), .B(n25603), .Z(n25604) );
  NANDN U25684 ( .A(n25564), .B(n25566), .Z(n25580) );
  XOR U25685 ( .A(n25606), .B(n25607), .Z(n25566) );
  AND U25686 ( .A(n1338), .B(n25608), .Z(n25606) );
  XOR U25687 ( .A(n25607), .B(n25609), .Z(n25608) );
  XOR U25688 ( .A(n25610), .B(n25611), .Z(n1338) );
  AND U25689 ( .A(n25612), .B(n25613), .Z(n25610) );
  XNOR U25690 ( .A(n25611), .B(n25577), .Z(n25613) );
  XNOR U25691 ( .A(n25614), .B(n25615), .Z(n25577) );
  ANDN U25692 ( .B(n25616), .A(n25617), .Z(n25614) );
  XOR U25693 ( .A(n25615), .B(n25618), .Z(n25616) );
  XOR U25694 ( .A(n25611), .B(n25579), .Z(n25612) );
  XOR U25695 ( .A(n25619), .B(n25620), .Z(n25579) );
  AND U25696 ( .A(n1342), .B(n25621), .Z(n25619) );
  XOR U25697 ( .A(n25622), .B(n25620), .Z(n25621) );
  XNOR U25698 ( .A(n25623), .B(n25624), .Z(n25611) );
  NAND U25699 ( .A(n25625), .B(n25626), .Z(n25624) );
  XOR U25700 ( .A(n25627), .B(n25603), .Z(n25626) );
  XOR U25701 ( .A(n25617), .B(n25618), .Z(n25603) );
  XOR U25702 ( .A(n25628), .B(n25629), .Z(n25618) );
  ANDN U25703 ( .B(n25630), .A(n25631), .Z(n25628) );
  XOR U25704 ( .A(n25629), .B(n25632), .Z(n25630) );
  XOR U25705 ( .A(n25633), .B(n25634), .Z(n25617) );
  XOR U25706 ( .A(n25635), .B(n25636), .Z(n25634) );
  ANDN U25707 ( .B(n25637), .A(n25638), .Z(n25635) );
  XOR U25708 ( .A(n25639), .B(n25636), .Z(n25637) );
  IV U25709 ( .A(n25615), .Z(n25633) );
  XOR U25710 ( .A(n25640), .B(n25641), .Z(n25615) );
  ANDN U25711 ( .B(n25642), .A(n25643), .Z(n25640) );
  XOR U25712 ( .A(n25641), .B(n25644), .Z(n25642) );
  IV U25713 ( .A(n25623), .Z(n25627) );
  XOR U25714 ( .A(n25623), .B(n25605), .Z(n25625) );
  XOR U25715 ( .A(n25645), .B(n25646), .Z(n25605) );
  AND U25716 ( .A(n1342), .B(n25647), .Z(n25645) );
  XOR U25717 ( .A(n25648), .B(n25646), .Z(n25647) );
  NANDN U25718 ( .A(n25607), .B(n25609), .Z(n25623) );
  XOR U25719 ( .A(n25649), .B(n25650), .Z(n25609) );
  AND U25720 ( .A(n1342), .B(n25651), .Z(n25649) );
  XOR U25721 ( .A(n25650), .B(n25652), .Z(n25651) );
  XOR U25722 ( .A(n25653), .B(n25654), .Z(n1342) );
  AND U25723 ( .A(n25655), .B(n25656), .Z(n25653) );
  XNOR U25724 ( .A(n25654), .B(n25620), .Z(n25656) );
  XNOR U25725 ( .A(n25657), .B(n25658), .Z(n25620) );
  ANDN U25726 ( .B(n25659), .A(n25660), .Z(n25657) );
  XOR U25727 ( .A(n25658), .B(n25661), .Z(n25659) );
  XOR U25728 ( .A(n25654), .B(n25622), .Z(n25655) );
  XOR U25729 ( .A(n25662), .B(n25663), .Z(n25622) );
  AND U25730 ( .A(n1346), .B(n25664), .Z(n25662) );
  XOR U25731 ( .A(n25665), .B(n25663), .Z(n25664) );
  XNOR U25732 ( .A(n25666), .B(n25667), .Z(n25654) );
  NAND U25733 ( .A(n25668), .B(n25669), .Z(n25667) );
  XOR U25734 ( .A(n25670), .B(n25646), .Z(n25669) );
  XOR U25735 ( .A(n25660), .B(n25661), .Z(n25646) );
  XOR U25736 ( .A(n25671), .B(n25672), .Z(n25661) );
  ANDN U25737 ( .B(n25673), .A(n25674), .Z(n25671) );
  XOR U25738 ( .A(n25672), .B(n25675), .Z(n25673) );
  XOR U25739 ( .A(n25676), .B(n25677), .Z(n25660) );
  XOR U25740 ( .A(n25678), .B(n25679), .Z(n25677) );
  ANDN U25741 ( .B(n25680), .A(n25681), .Z(n25678) );
  XOR U25742 ( .A(n25682), .B(n25679), .Z(n25680) );
  IV U25743 ( .A(n25658), .Z(n25676) );
  XOR U25744 ( .A(n25683), .B(n25684), .Z(n25658) );
  ANDN U25745 ( .B(n25685), .A(n25686), .Z(n25683) );
  XOR U25746 ( .A(n25684), .B(n25687), .Z(n25685) );
  IV U25747 ( .A(n25666), .Z(n25670) );
  XOR U25748 ( .A(n25666), .B(n25648), .Z(n25668) );
  XOR U25749 ( .A(n25688), .B(n25689), .Z(n25648) );
  AND U25750 ( .A(n1346), .B(n25690), .Z(n25688) );
  XOR U25751 ( .A(n25691), .B(n25689), .Z(n25690) );
  NANDN U25752 ( .A(n25650), .B(n25652), .Z(n25666) );
  XOR U25753 ( .A(n25692), .B(n25693), .Z(n25652) );
  AND U25754 ( .A(n1346), .B(n25694), .Z(n25692) );
  XOR U25755 ( .A(n25693), .B(n25695), .Z(n25694) );
  XOR U25756 ( .A(n25696), .B(n25697), .Z(n1346) );
  AND U25757 ( .A(n25698), .B(n25699), .Z(n25696) );
  XNOR U25758 ( .A(n25697), .B(n25663), .Z(n25699) );
  XNOR U25759 ( .A(n25700), .B(n25701), .Z(n25663) );
  ANDN U25760 ( .B(n25702), .A(n25703), .Z(n25700) );
  XOR U25761 ( .A(n25701), .B(n25704), .Z(n25702) );
  XOR U25762 ( .A(n25697), .B(n25665), .Z(n25698) );
  XOR U25763 ( .A(n25705), .B(n25706), .Z(n25665) );
  AND U25764 ( .A(n1350), .B(n25707), .Z(n25705) );
  XOR U25765 ( .A(n25708), .B(n25706), .Z(n25707) );
  XNOR U25766 ( .A(n25709), .B(n25710), .Z(n25697) );
  NAND U25767 ( .A(n25711), .B(n25712), .Z(n25710) );
  XOR U25768 ( .A(n25713), .B(n25689), .Z(n25712) );
  XOR U25769 ( .A(n25703), .B(n25704), .Z(n25689) );
  XOR U25770 ( .A(n25714), .B(n25715), .Z(n25704) );
  ANDN U25771 ( .B(n25716), .A(n25717), .Z(n25714) );
  XOR U25772 ( .A(n25715), .B(n25718), .Z(n25716) );
  XOR U25773 ( .A(n25719), .B(n25720), .Z(n25703) );
  XOR U25774 ( .A(n25721), .B(n25722), .Z(n25720) );
  ANDN U25775 ( .B(n25723), .A(n25724), .Z(n25721) );
  XOR U25776 ( .A(n25725), .B(n25722), .Z(n25723) );
  IV U25777 ( .A(n25701), .Z(n25719) );
  XOR U25778 ( .A(n25726), .B(n25727), .Z(n25701) );
  ANDN U25779 ( .B(n25728), .A(n25729), .Z(n25726) );
  XOR U25780 ( .A(n25727), .B(n25730), .Z(n25728) );
  IV U25781 ( .A(n25709), .Z(n25713) );
  XOR U25782 ( .A(n25709), .B(n25691), .Z(n25711) );
  XOR U25783 ( .A(n25731), .B(n25732), .Z(n25691) );
  AND U25784 ( .A(n1350), .B(n25733), .Z(n25731) );
  XOR U25785 ( .A(n25734), .B(n25732), .Z(n25733) );
  NANDN U25786 ( .A(n25693), .B(n25695), .Z(n25709) );
  XOR U25787 ( .A(n25735), .B(n25736), .Z(n25695) );
  AND U25788 ( .A(n1350), .B(n25737), .Z(n25735) );
  XOR U25789 ( .A(n25736), .B(n25738), .Z(n25737) );
  XOR U25790 ( .A(n25739), .B(n25740), .Z(n1350) );
  AND U25791 ( .A(n25741), .B(n25742), .Z(n25739) );
  XNOR U25792 ( .A(n25740), .B(n25706), .Z(n25742) );
  XNOR U25793 ( .A(n25743), .B(n25744), .Z(n25706) );
  ANDN U25794 ( .B(n25745), .A(n25746), .Z(n25743) );
  XOR U25795 ( .A(n25744), .B(n25747), .Z(n25745) );
  XOR U25796 ( .A(n25740), .B(n25708), .Z(n25741) );
  XOR U25797 ( .A(n25748), .B(n25749), .Z(n25708) );
  AND U25798 ( .A(n1354), .B(n25750), .Z(n25748) );
  XOR U25799 ( .A(n25751), .B(n25749), .Z(n25750) );
  XNOR U25800 ( .A(n25752), .B(n25753), .Z(n25740) );
  NAND U25801 ( .A(n25754), .B(n25755), .Z(n25753) );
  XOR U25802 ( .A(n25756), .B(n25732), .Z(n25755) );
  XOR U25803 ( .A(n25746), .B(n25747), .Z(n25732) );
  XOR U25804 ( .A(n25757), .B(n25758), .Z(n25747) );
  ANDN U25805 ( .B(n25759), .A(n25760), .Z(n25757) );
  XOR U25806 ( .A(n25758), .B(n25761), .Z(n25759) );
  XOR U25807 ( .A(n25762), .B(n25763), .Z(n25746) );
  XOR U25808 ( .A(n25764), .B(n25765), .Z(n25763) );
  ANDN U25809 ( .B(n25766), .A(n25767), .Z(n25764) );
  XOR U25810 ( .A(n25768), .B(n25765), .Z(n25766) );
  IV U25811 ( .A(n25744), .Z(n25762) );
  XOR U25812 ( .A(n25769), .B(n25770), .Z(n25744) );
  ANDN U25813 ( .B(n25771), .A(n25772), .Z(n25769) );
  XOR U25814 ( .A(n25770), .B(n25773), .Z(n25771) );
  IV U25815 ( .A(n25752), .Z(n25756) );
  XOR U25816 ( .A(n25752), .B(n25734), .Z(n25754) );
  XOR U25817 ( .A(n25774), .B(n25775), .Z(n25734) );
  AND U25818 ( .A(n1354), .B(n25776), .Z(n25774) );
  XOR U25819 ( .A(n25777), .B(n25775), .Z(n25776) );
  NANDN U25820 ( .A(n25736), .B(n25738), .Z(n25752) );
  XOR U25821 ( .A(n25778), .B(n25779), .Z(n25738) );
  AND U25822 ( .A(n1354), .B(n25780), .Z(n25778) );
  XOR U25823 ( .A(n25779), .B(n25781), .Z(n25780) );
  XOR U25824 ( .A(n25782), .B(n25783), .Z(n1354) );
  AND U25825 ( .A(n25784), .B(n25785), .Z(n25782) );
  XNOR U25826 ( .A(n25783), .B(n25749), .Z(n25785) );
  XNOR U25827 ( .A(n25786), .B(n25787), .Z(n25749) );
  ANDN U25828 ( .B(n25788), .A(n25789), .Z(n25786) );
  XOR U25829 ( .A(n25787), .B(n25790), .Z(n25788) );
  XOR U25830 ( .A(n25783), .B(n25751), .Z(n25784) );
  XOR U25831 ( .A(n25791), .B(n25792), .Z(n25751) );
  AND U25832 ( .A(n1358), .B(n25793), .Z(n25791) );
  XOR U25833 ( .A(n25794), .B(n25792), .Z(n25793) );
  XNOR U25834 ( .A(n25795), .B(n25796), .Z(n25783) );
  NAND U25835 ( .A(n25797), .B(n25798), .Z(n25796) );
  XOR U25836 ( .A(n25799), .B(n25775), .Z(n25798) );
  XOR U25837 ( .A(n25789), .B(n25790), .Z(n25775) );
  XOR U25838 ( .A(n25800), .B(n25801), .Z(n25790) );
  ANDN U25839 ( .B(n25802), .A(n25803), .Z(n25800) );
  XOR U25840 ( .A(n25801), .B(n25804), .Z(n25802) );
  XOR U25841 ( .A(n25805), .B(n25806), .Z(n25789) );
  XOR U25842 ( .A(n25807), .B(n25808), .Z(n25806) );
  ANDN U25843 ( .B(n25809), .A(n25810), .Z(n25807) );
  XOR U25844 ( .A(n25811), .B(n25808), .Z(n25809) );
  IV U25845 ( .A(n25787), .Z(n25805) );
  XOR U25846 ( .A(n25812), .B(n25813), .Z(n25787) );
  ANDN U25847 ( .B(n25814), .A(n25815), .Z(n25812) );
  XOR U25848 ( .A(n25813), .B(n25816), .Z(n25814) );
  IV U25849 ( .A(n25795), .Z(n25799) );
  XOR U25850 ( .A(n25795), .B(n25777), .Z(n25797) );
  XOR U25851 ( .A(n25817), .B(n25818), .Z(n25777) );
  AND U25852 ( .A(n1358), .B(n25819), .Z(n25817) );
  XOR U25853 ( .A(n25820), .B(n25818), .Z(n25819) );
  NANDN U25854 ( .A(n25779), .B(n25781), .Z(n25795) );
  XOR U25855 ( .A(n25821), .B(n25822), .Z(n25781) );
  AND U25856 ( .A(n1358), .B(n25823), .Z(n25821) );
  XOR U25857 ( .A(n25822), .B(n25824), .Z(n25823) );
  XOR U25858 ( .A(n25825), .B(n25826), .Z(n1358) );
  AND U25859 ( .A(n25827), .B(n25828), .Z(n25825) );
  XNOR U25860 ( .A(n25826), .B(n25792), .Z(n25828) );
  XNOR U25861 ( .A(n25829), .B(n25830), .Z(n25792) );
  ANDN U25862 ( .B(n25831), .A(n25832), .Z(n25829) );
  XOR U25863 ( .A(n25830), .B(n25833), .Z(n25831) );
  XOR U25864 ( .A(n25826), .B(n25794), .Z(n25827) );
  XOR U25865 ( .A(n25834), .B(n25835), .Z(n25794) );
  AND U25866 ( .A(n1362), .B(n25836), .Z(n25834) );
  XOR U25867 ( .A(n25837), .B(n25835), .Z(n25836) );
  XNOR U25868 ( .A(n25838), .B(n25839), .Z(n25826) );
  NAND U25869 ( .A(n25840), .B(n25841), .Z(n25839) );
  XOR U25870 ( .A(n25842), .B(n25818), .Z(n25841) );
  XOR U25871 ( .A(n25832), .B(n25833), .Z(n25818) );
  XOR U25872 ( .A(n25843), .B(n25844), .Z(n25833) );
  ANDN U25873 ( .B(n25845), .A(n25846), .Z(n25843) );
  XOR U25874 ( .A(n25844), .B(n25847), .Z(n25845) );
  XOR U25875 ( .A(n25848), .B(n25849), .Z(n25832) );
  XOR U25876 ( .A(n25850), .B(n25851), .Z(n25849) );
  ANDN U25877 ( .B(n25852), .A(n25853), .Z(n25850) );
  XOR U25878 ( .A(n25854), .B(n25851), .Z(n25852) );
  IV U25879 ( .A(n25830), .Z(n25848) );
  XOR U25880 ( .A(n25855), .B(n25856), .Z(n25830) );
  ANDN U25881 ( .B(n25857), .A(n25858), .Z(n25855) );
  XOR U25882 ( .A(n25856), .B(n25859), .Z(n25857) );
  IV U25883 ( .A(n25838), .Z(n25842) );
  XOR U25884 ( .A(n25838), .B(n25820), .Z(n25840) );
  XOR U25885 ( .A(n25860), .B(n25861), .Z(n25820) );
  AND U25886 ( .A(n1362), .B(n25862), .Z(n25860) );
  XOR U25887 ( .A(n25863), .B(n25861), .Z(n25862) );
  NANDN U25888 ( .A(n25822), .B(n25824), .Z(n25838) );
  XOR U25889 ( .A(n25864), .B(n25865), .Z(n25824) );
  AND U25890 ( .A(n1362), .B(n25866), .Z(n25864) );
  XOR U25891 ( .A(n25865), .B(n25867), .Z(n25866) );
  XOR U25892 ( .A(n25868), .B(n25869), .Z(n1362) );
  AND U25893 ( .A(n25870), .B(n25871), .Z(n25868) );
  XNOR U25894 ( .A(n25869), .B(n25835), .Z(n25871) );
  XNOR U25895 ( .A(n25872), .B(n25873), .Z(n25835) );
  ANDN U25896 ( .B(n25874), .A(n25875), .Z(n25872) );
  XOR U25897 ( .A(n25873), .B(n25876), .Z(n25874) );
  XOR U25898 ( .A(n25869), .B(n25837), .Z(n25870) );
  XOR U25899 ( .A(n25877), .B(n25878), .Z(n25837) );
  AND U25900 ( .A(n1366), .B(n25879), .Z(n25877) );
  XOR U25901 ( .A(n25880), .B(n25878), .Z(n25879) );
  XNOR U25902 ( .A(n25881), .B(n25882), .Z(n25869) );
  NAND U25903 ( .A(n25883), .B(n25884), .Z(n25882) );
  XOR U25904 ( .A(n25885), .B(n25861), .Z(n25884) );
  XOR U25905 ( .A(n25875), .B(n25876), .Z(n25861) );
  XOR U25906 ( .A(n25886), .B(n25887), .Z(n25876) );
  ANDN U25907 ( .B(n25888), .A(n25889), .Z(n25886) );
  XOR U25908 ( .A(n25887), .B(n25890), .Z(n25888) );
  XOR U25909 ( .A(n25891), .B(n25892), .Z(n25875) );
  XOR U25910 ( .A(n25893), .B(n25894), .Z(n25892) );
  ANDN U25911 ( .B(n25895), .A(n25896), .Z(n25893) );
  XOR U25912 ( .A(n25897), .B(n25894), .Z(n25895) );
  IV U25913 ( .A(n25873), .Z(n25891) );
  XOR U25914 ( .A(n25898), .B(n25899), .Z(n25873) );
  ANDN U25915 ( .B(n25900), .A(n25901), .Z(n25898) );
  XOR U25916 ( .A(n25899), .B(n25902), .Z(n25900) );
  IV U25917 ( .A(n25881), .Z(n25885) );
  XOR U25918 ( .A(n25881), .B(n25863), .Z(n25883) );
  XOR U25919 ( .A(n25903), .B(n25904), .Z(n25863) );
  AND U25920 ( .A(n1366), .B(n25905), .Z(n25903) );
  XOR U25921 ( .A(n25906), .B(n25904), .Z(n25905) );
  NANDN U25922 ( .A(n25865), .B(n25867), .Z(n25881) );
  XOR U25923 ( .A(n25907), .B(n25908), .Z(n25867) );
  AND U25924 ( .A(n1366), .B(n25909), .Z(n25907) );
  XOR U25925 ( .A(n25908), .B(n25910), .Z(n25909) );
  XOR U25926 ( .A(n25911), .B(n25912), .Z(n1366) );
  AND U25927 ( .A(n25913), .B(n25914), .Z(n25911) );
  XNOR U25928 ( .A(n25912), .B(n25878), .Z(n25914) );
  XNOR U25929 ( .A(n25915), .B(n25916), .Z(n25878) );
  ANDN U25930 ( .B(n25917), .A(n25918), .Z(n25915) );
  XOR U25931 ( .A(n25916), .B(n25919), .Z(n25917) );
  XOR U25932 ( .A(n25912), .B(n25880), .Z(n25913) );
  XOR U25933 ( .A(n25920), .B(n25921), .Z(n25880) );
  AND U25934 ( .A(n1370), .B(n25922), .Z(n25920) );
  XOR U25935 ( .A(n25923), .B(n25921), .Z(n25922) );
  XNOR U25936 ( .A(n25924), .B(n25925), .Z(n25912) );
  NAND U25937 ( .A(n25926), .B(n25927), .Z(n25925) );
  XOR U25938 ( .A(n25928), .B(n25904), .Z(n25927) );
  XOR U25939 ( .A(n25918), .B(n25919), .Z(n25904) );
  XOR U25940 ( .A(n25929), .B(n25930), .Z(n25919) );
  ANDN U25941 ( .B(n25931), .A(n25932), .Z(n25929) );
  XOR U25942 ( .A(n25930), .B(n25933), .Z(n25931) );
  XOR U25943 ( .A(n25934), .B(n25935), .Z(n25918) );
  XOR U25944 ( .A(n25936), .B(n25937), .Z(n25935) );
  ANDN U25945 ( .B(n25938), .A(n25939), .Z(n25936) );
  XOR U25946 ( .A(n25940), .B(n25937), .Z(n25938) );
  IV U25947 ( .A(n25916), .Z(n25934) );
  XOR U25948 ( .A(n25941), .B(n25942), .Z(n25916) );
  ANDN U25949 ( .B(n25943), .A(n25944), .Z(n25941) );
  XOR U25950 ( .A(n25942), .B(n25945), .Z(n25943) );
  IV U25951 ( .A(n25924), .Z(n25928) );
  XOR U25952 ( .A(n25924), .B(n25906), .Z(n25926) );
  XOR U25953 ( .A(n25946), .B(n25947), .Z(n25906) );
  AND U25954 ( .A(n1370), .B(n25948), .Z(n25946) );
  XOR U25955 ( .A(n25949), .B(n25947), .Z(n25948) );
  NANDN U25956 ( .A(n25908), .B(n25910), .Z(n25924) );
  XOR U25957 ( .A(n25950), .B(n25951), .Z(n25910) );
  AND U25958 ( .A(n1370), .B(n25952), .Z(n25950) );
  XOR U25959 ( .A(n25951), .B(n25953), .Z(n25952) );
  XOR U25960 ( .A(n25954), .B(n25955), .Z(n1370) );
  AND U25961 ( .A(n25956), .B(n25957), .Z(n25954) );
  XNOR U25962 ( .A(n25955), .B(n25921), .Z(n25957) );
  XNOR U25963 ( .A(n25958), .B(n25959), .Z(n25921) );
  ANDN U25964 ( .B(n25960), .A(n25961), .Z(n25958) );
  XOR U25965 ( .A(n25959), .B(n25962), .Z(n25960) );
  XOR U25966 ( .A(n25955), .B(n25923), .Z(n25956) );
  XOR U25967 ( .A(n25963), .B(n25964), .Z(n25923) );
  AND U25968 ( .A(n1374), .B(n25965), .Z(n25963) );
  XOR U25969 ( .A(n25966), .B(n25964), .Z(n25965) );
  XNOR U25970 ( .A(n25967), .B(n25968), .Z(n25955) );
  NAND U25971 ( .A(n25969), .B(n25970), .Z(n25968) );
  XOR U25972 ( .A(n25971), .B(n25947), .Z(n25970) );
  XOR U25973 ( .A(n25961), .B(n25962), .Z(n25947) );
  XOR U25974 ( .A(n25972), .B(n25973), .Z(n25962) );
  ANDN U25975 ( .B(n25974), .A(n25975), .Z(n25972) );
  XOR U25976 ( .A(n25973), .B(n25976), .Z(n25974) );
  XOR U25977 ( .A(n25977), .B(n25978), .Z(n25961) );
  XOR U25978 ( .A(n25979), .B(n25980), .Z(n25978) );
  ANDN U25979 ( .B(n25981), .A(n25982), .Z(n25979) );
  XOR U25980 ( .A(n25983), .B(n25980), .Z(n25981) );
  IV U25981 ( .A(n25959), .Z(n25977) );
  XOR U25982 ( .A(n25984), .B(n25985), .Z(n25959) );
  ANDN U25983 ( .B(n25986), .A(n25987), .Z(n25984) );
  XOR U25984 ( .A(n25985), .B(n25988), .Z(n25986) );
  IV U25985 ( .A(n25967), .Z(n25971) );
  XOR U25986 ( .A(n25967), .B(n25949), .Z(n25969) );
  XOR U25987 ( .A(n25989), .B(n25990), .Z(n25949) );
  AND U25988 ( .A(n1374), .B(n25991), .Z(n25989) );
  XOR U25989 ( .A(n25992), .B(n25990), .Z(n25991) );
  NANDN U25990 ( .A(n25951), .B(n25953), .Z(n25967) );
  XOR U25991 ( .A(n25993), .B(n25994), .Z(n25953) );
  AND U25992 ( .A(n1374), .B(n25995), .Z(n25993) );
  XOR U25993 ( .A(n25994), .B(n25996), .Z(n25995) );
  XOR U25994 ( .A(n25997), .B(n25998), .Z(n1374) );
  AND U25995 ( .A(n25999), .B(n26000), .Z(n25997) );
  XNOR U25996 ( .A(n25998), .B(n25964), .Z(n26000) );
  XNOR U25997 ( .A(n26001), .B(n26002), .Z(n25964) );
  ANDN U25998 ( .B(n26003), .A(n26004), .Z(n26001) );
  XOR U25999 ( .A(n26002), .B(n26005), .Z(n26003) );
  XOR U26000 ( .A(n25998), .B(n25966), .Z(n25999) );
  XOR U26001 ( .A(n26006), .B(n26007), .Z(n25966) );
  AND U26002 ( .A(n1378), .B(n26008), .Z(n26006) );
  XOR U26003 ( .A(n26009), .B(n26007), .Z(n26008) );
  XNOR U26004 ( .A(n26010), .B(n26011), .Z(n25998) );
  NAND U26005 ( .A(n26012), .B(n26013), .Z(n26011) );
  XOR U26006 ( .A(n26014), .B(n25990), .Z(n26013) );
  XOR U26007 ( .A(n26004), .B(n26005), .Z(n25990) );
  XOR U26008 ( .A(n26015), .B(n26016), .Z(n26005) );
  ANDN U26009 ( .B(n26017), .A(n26018), .Z(n26015) );
  XOR U26010 ( .A(n26016), .B(n26019), .Z(n26017) );
  XOR U26011 ( .A(n26020), .B(n26021), .Z(n26004) );
  XOR U26012 ( .A(n26022), .B(n26023), .Z(n26021) );
  ANDN U26013 ( .B(n26024), .A(n26025), .Z(n26022) );
  XOR U26014 ( .A(n26026), .B(n26023), .Z(n26024) );
  IV U26015 ( .A(n26002), .Z(n26020) );
  XOR U26016 ( .A(n26027), .B(n26028), .Z(n26002) );
  ANDN U26017 ( .B(n26029), .A(n26030), .Z(n26027) );
  XOR U26018 ( .A(n26028), .B(n26031), .Z(n26029) );
  IV U26019 ( .A(n26010), .Z(n26014) );
  XOR U26020 ( .A(n26010), .B(n25992), .Z(n26012) );
  XOR U26021 ( .A(n26032), .B(n26033), .Z(n25992) );
  AND U26022 ( .A(n1378), .B(n26034), .Z(n26032) );
  XOR U26023 ( .A(n26035), .B(n26033), .Z(n26034) );
  NANDN U26024 ( .A(n25994), .B(n25996), .Z(n26010) );
  XOR U26025 ( .A(n26036), .B(n26037), .Z(n25996) );
  AND U26026 ( .A(n1378), .B(n26038), .Z(n26036) );
  XOR U26027 ( .A(n26037), .B(n26039), .Z(n26038) );
  XOR U26028 ( .A(n26040), .B(n26041), .Z(n1378) );
  AND U26029 ( .A(n26042), .B(n26043), .Z(n26040) );
  XNOR U26030 ( .A(n26041), .B(n26007), .Z(n26043) );
  XNOR U26031 ( .A(n26044), .B(n26045), .Z(n26007) );
  ANDN U26032 ( .B(n26046), .A(n26047), .Z(n26044) );
  XOR U26033 ( .A(n26045), .B(n26048), .Z(n26046) );
  XOR U26034 ( .A(n26041), .B(n26009), .Z(n26042) );
  XOR U26035 ( .A(n26049), .B(n26050), .Z(n26009) );
  AND U26036 ( .A(n1382), .B(n26051), .Z(n26049) );
  XOR U26037 ( .A(n26052), .B(n26050), .Z(n26051) );
  XNOR U26038 ( .A(n26053), .B(n26054), .Z(n26041) );
  NAND U26039 ( .A(n26055), .B(n26056), .Z(n26054) );
  XOR U26040 ( .A(n26057), .B(n26033), .Z(n26056) );
  XOR U26041 ( .A(n26047), .B(n26048), .Z(n26033) );
  XOR U26042 ( .A(n26058), .B(n26059), .Z(n26048) );
  ANDN U26043 ( .B(n26060), .A(n26061), .Z(n26058) );
  XOR U26044 ( .A(n26059), .B(n26062), .Z(n26060) );
  XOR U26045 ( .A(n26063), .B(n26064), .Z(n26047) );
  XOR U26046 ( .A(n26065), .B(n26066), .Z(n26064) );
  ANDN U26047 ( .B(n26067), .A(n26068), .Z(n26065) );
  XOR U26048 ( .A(n26069), .B(n26066), .Z(n26067) );
  IV U26049 ( .A(n26045), .Z(n26063) );
  XOR U26050 ( .A(n26070), .B(n26071), .Z(n26045) );
  ANDN U26051 ( .B(n26072), .A(n26073), .Z(n26070) );
  XOR U26052 ( .A(n26071), .B(n26074), .Z(n26072) );
  IV U26053 ( .A(n26053), .Z(n26057) );
  XOR U26054 ( .A(n26053), .B(n26035), .Z(n26055) );
  XOR U26055 ( .A(n26075), .B(n26076), .Z(n26035) );
  AND U26056 ( .A(n1382), .B(n26077), .Z(n26075) );
  XOR U26057 ( .A(n26078), .B(n26076), .Z(n26077) );
  NANDN U26058 ( .A(n26037), .B(n26039), .Z(n26053) );
  XOR U26059 ( .A(n26079), .B(n26080), .Z(n26039) );
  AND U26060 ( .A(n1382), .B(n26081), .Z(n26079) );
  XOR U26061 ( .A(n26080), .B(n26082), .Z(n26081) );
  XOR U26062 ( .A(n26083), .B(n26084), .Z(n1382) );
  AND U26063 ( .A(n26085), .B(n26086), .Z(n26083) );
  XNOR U26064 ( .A(n26084), .B(n26050), .Z(n26086) );
  XNOR U26065 ( .A(n26087), .B(n26088), .Z(n26050) );
  ANDN U26066 ( .B(n26089), .A(n26090), .Z(n26087) );
  XOR U26067 ( .A(n26088), .B(n26091), .Z(n26089) );
  XOR U26068 ( .A(n26084), .B(n26052), .Z(n26085) );
  XOR U26069 ( .A(n26092), .B(n26093), .Z(n26052) );
  AND U26070 ( .A(n1386), .B(n26094), .Z(n26092) );
  XOR U26071 ( .A(n26095), .B(n26093), .Z(n26094) );
  XNOR U26072 ( .A(n26096), .B(n26097), .Z(n26084) );
  NAND U26073 ( .A(n26098), .B(n26099), .Z(n26097) );
  XOR U26074 ( .A(n26100), .B(n26076), .Z(n26099) );
  XOR U26075 ( .A(n26090), .B(n26091), .Z(n26076) );
  XOR U26076 ( .A(n26101), .B(n26102), .Z(n26091) );
  ANDN U26077 ( .B(n26103), .A(n26104), .Z(n26101) );
  XOR U26078 ( .A(n26102), .B(n26105), .Z(n26103) );
  XOR U26079 ( .A(n26106), .B(n26107), .Z(n26090) );
  XOR U26080 ( .A(n26108), .B(n26109), .Z(n26107) );
  ANDN U26081 ( .B(n26110), .A(n26111), .Z(n26108) );
  XOR U26082 ( .A(n26112), .B(n26109), .Z(n26110) );
  IV U26083 ( .A(n26088), .Z(n26106) );
  XOR U26084 ( .A(n26113), .B(n26114), .Z(n26088) );
  ANDN U26085 ( .B(n26115), .A(n26116), .Z(n26113) );
  XOR U26086 ( .A(n26114), .B(n26117), .Z(n26115) );
  IV U26087 ( .A(n26096), .Z(n26100) );
  XOR U26088 ( .A(n26096), .B(n26078), .Z(n26098) );
  XOR U26089 ( .A(n26118), .B(n26119), .Z(n26078) );
  AND U26090 ( .A(n1386), .B(n26120), .Z(n26118) );
  XOR U26091 ( .A(n26121), .B(n26119), .Z(n26120) );
  NANDN U26092 ( .A(n26080), .B(n26082), .Z(n26096) );
  XOR U26093 ( .A(n26122), .B(n26123), .Z(n26082) );
  AND U26094 ( .A(n1386), .B(n26124), .Z(n26122) );
  XOR U26095 ( .A(n26123), .B(n26125), .Z(n26124) );
  XOR U26096 ( .A(n26126), .B(n26127), .Z(n1386) );
  AND U26097 ( .A(n26128), .B(n26129), .Z(n26126) );
  XNOR U26098 ( .A(n26127), .B(n26093), .Z(n26129) );
  XNOR U26099 ( .A(n26130), .B(n26131), .Z(n26093) );
  ANDN U26100 ( .B(n26132), .A(n26133), .Z(n26130) );
  XOR U26101 ( .A(n26131), .B(n26134), .Z(n26132) );
  XOR U26102 ( .A(n26127), .B(n26095), .Z(n26128) );
  XOR U26103 ( .A(n26135), .B(n26136), .Z(n26095) );
  AND U26104 ( .A(n1390), .B(n26137), .Z(n26135) );
  XOR U26105 ( .A(n26138), .B(n26136), .Z(n26137) );
  XNOR U26106 ( .A(n26139), .B(n26140), .Z(n26127) );
  NAND U26107 ( .A(n26141), .B(n26142), .Z(n26140) );
  XOR U26108 ( .A(n26143), .B(n26119), .Z(n26142) );
  XOR U26109 ( .A(n26133), .B(n26134), .Z(n26119) );
  XOR U26110 ( .A(n26144), .B(n26145), .Z(n26134) );
  ANDN U26111 ( .B(n26146), .A(n26147), .Z(n26144) );
  XOR U26112 ( .A(n26145), .B(n26148), .Z(n26146) );
  XOR U26113 ( .A(n26149), .B(n26150), .Z(n26133) );
  XOR U26114 ( .A(n26151), .B(n26152), .Z(n26150) );
  ANDN U26115 ( .B(n26153), .A(n26154), .Z(n26151) );
  XOR U26116 ( .A(n26155), .B(n26152), .Z(n26153) );
  IV U26117 ( .A(n26131), .Z(n26149) );
  XOR U26118 ( .A(n26156), .B(n26157), .Z(n26131) );
  ANDN U26119 ( .B(n26158), .A(n26159), .Z(n26156) );
  XOR U26120 ( .A(n26157), .B(n26160), .Z(n26158) );
  IV U26121 ( .A(n26139), .Z(n26143) );
  XOR U26122 ( .A(n26139), .B(n26121), .Z(n26141) );
  XOR U26123 ( .A(n26161), .B(n26162), .Z(n26121) );
  AND U26124 ( .A(n1390), .B(n26163), .Z(n26161) );
  XOR U26125 ( .A(n26164), .B(n26162), .Z(n26163) );
  NANDN U26126 ( .A(n26123), .B(n26125), .Z(n26139) );
  XOR U26127 ( .A(n26165), .B(n26166), .Z(n26125) );
  AND U26128 ( .A(n1390), .B(n26167), .Z(n26165) );
  XOR U26129 ( .A(n26166), .B(n26168), .Z(n26167) );
  XOR U26130 ( .A(n26169), .B(n26170), .Z(n1390) );
  AND U26131 ( .A(n26171), .B(n26172), .Z(n26169) );
  XNOR U26132 ( .A(n26170), .B(n26136), .Z(n26172) );
  XNOR U26133 ( .A(n26173), .B(n26174), .Z(n26136) );
  ANDN U26134 ( .B(n26175), .A(n26176), .Z(n26173) );
  XOR U26135 ( .A(n26174), .B(n26177), .Z(n26175) );
  XOR U26136 ( .A(n26170), .B(n26138), .Z(n26171) );
  XOR U26137 ( .A(n26178), .B(n26179), .Z(n26138) );
  AND U26138 ( .A(n1394), .B(n26180), .Z(n26178) );
  XOR U26139 ( .A(n26181), .B(n26179), .Z(n26180) );
  XNOR U26140 ( .A(n26182), .B(n26183), .Z(n26170) );
  NAND U26141 ( .A(n26184), .B(n26185), .Z(n26183) );
  XOR U26142 ( .A(n26186), .B(n26162), .Z(n26185) );
  XOR U26143 ( .A(n26176), .B(n26177), .Z(n26162) );
  XOR U26144 ( .A(n26187), .B(n26188), .Z(n26177) );
  ANDN U26145 ( .B(n26189), .A(n26190), .Z(n26187) );
  XOR U26146 ( .A(n26188), .B(n26191), .Z(n26189) );
  XOR U26147 ( .A(n26192), .B(n26193), .Z(n26176) );
  XOR U26148 ( .A(n26194), .B(n26195), .Z(n26193) );
  ANDN U26149 ( .B(n26196), .A(n26197), .Z(n26194) );
  XOR U26150 ( .A(n26198), .B(n26195), .Z(n26196) );
  IV U26151 ( .A(n26174), .Z(n26192) );
  XOR U26152 ( .A(n26199), .B(n26200), .Z(n26174) );
  ANDN U26153 ( .B(n26201), .A(n26202), .Z(n26199) );
  XOR U26154 ( .A(n26200), .B(n26203), .Z(n26201) );
  IV U26155 ( .A(n26182), .Z(n26186) );
  XOR U26156 ( .A(n26182), .B(n26164), .Z(n26184) );
  XOR U26157 ( .A(n26204), .B(n26205), .Z(n26164) );
  AND U26158 ( .A(n1394), .B(n26206), .Z(n26204) );
  XOR U26159 ( .A(n26207), .B(n26205), .Z(n26206) );
  NANDN U26160 ( .A(n26166), .B(n26168), .Z(n26182) );
  XOR U26161 ( .A(n26208), .B(n26209), .Z(n26168) );
  AND U26162 ( .A(n1394), .B(n26210), .Z(n26208) );
  XOR U26163 ( .A(n26209), .B(n26211), .Z(n26210) );
  XOR U26164 ( .A(n26212), .B(n26213), .Z(n1394) );
  AND U26165 ( .A(n26214), .B(n26215), .Z(n26212) );
  XNOR U26166 ( .A(n26213), .B(n26179), .Z(n26215) );
  XNOR U26167 ( .A(n26216), .B(n26217), .Z(n26179) );
  ANDN U26168 ( .B(n26218), .A(n26219), .Z(n26216) );
  XOR U26169 ( .A(n26217), .B(n26220), .Z(n26218) );
  XOR U26170 ( .A(n26213), .B(n26181), .Z(n26214) );
  XOR U26171 ( .A(n26221), .B(n26222), .Z(n26181) );
  AND U26172 ( .A(n1398), .B(n26223), .Z(n26221) );
  XOR U26173 ( .A(n26224), .B(n26222), .Z(n26223) );
  XNOR U26174 ( .A(n26225), .B(n26226), .Z(n26213) );
  NAND U26175 ( .A(n26227), .B(n26228), .Z(n26226) );
  XOR U26176 ( .A(n26229), .B(n26205), .Z(n26228) );
  XOR U26177 ( .A(n26219), .B(n26220), .Z(n26205) );
  XOR U26178 ( .A(n26230), .B(n26231), .Z(n26220) );
  ANDN U26179 ( .B(n26232), .A(n26233), .Z(n26230) );
  XOR U26180 ( .A(n26231), .B(n26234), .Z(n26232) );
  XOR U26181 ( .A(n26235), .B(n26236), .Z(n26219) );
  XOR U26182 ( .A(n26237), .B(n26238), .Z(n26236) );
  ANDN U26183 ( .B(n26239), .A(n26240), .Z(n26237) );
  XOR U26184 ( .A(n26241), .B(n26238), .Z(n26239) );
  IV U26185 ( .A(n26217), .Z(n26235) );
  XOR U26186 ( .A(n26242), .B(n26243), .Z(n26217) );
  ANDN U26187 ( .B(n26244), .A(n26245), .Z(n26242) );
  XOR U26188 ( .A(n26243), .B(n26246), .Z(n26244) );
  IV U26189 ( .A(n26225), .Z(n26229) );
  XOR U26190 ( .A(n26225), .B(n26207), .Z(n26227) );
  XOR U26191 ( .A(n26247), .B(n26248), .Z(n26207) );
  AND U26192 ( .A(n1398), .B(n26249), .Z(n26247) );
  XOR U26193 ( .A(n26250), .B(n26248), .Z(n26249) );
  NANDN U26194 ( .A(n26209), .B(n26211), .Z(n26225) );
  XOR U26195 ( .A(n26251), .B(n26252), .Z(n26211) );
  AND U26196 ( .A(n1398), .B(n26253), .Z(n26251) );
  XOR U26197 ( .A(n26252), .B(n26254), .Z(n26253) );
  XOR U26198 ( .A(n26255), .B(n26256), .Z(n1398) );
  AND U26199 ( .A(n26257), .B(n26258), .Z(n26255) );
  XNOR U26200 ( .A(n26256), .B(n26222), .Z(n26258) );
  XNOR U26201 ( .A(n26259), .B(n26260), .Z(n26222) );
  ANDN U26202 ( .B(n26261), .A(n26262), .Z(n26259) );
  XOR U26203 ( .A(n26260), .B(n26263), .Z(n26261) );
  XOR U26204 ( .A(n26256), .B(n26224), .Z(n26257) );
  XOR U26205 ( .A(n26264), .B(n26265), .Z(n26224) );
  AND U26206 ( .A(n1402), .B(n26266), .Z(n26264) );
  XOR U26207 ( .A(n26267), .B(n26265), .Z(n26266) );
  XNOR U26208 ( .A(n26268), .B(n26269), .Z(n26256) );
  NAND U26209 ( .A(n26270), .B(n26271), .Z(n26269) );
  XOR U26210 ( .A(n26272), .B(n26248), .Z(n26271) );
  XOR U26211 ( .A(n26262), .B(n26263), .Z(n26248) );
  XOR U26212 ( .A(n26273), .B(n26274), .Z(n26263) );
  ANDN U26213 ( .B(n26275), .A(n26276), .Z(n26273) );
  XOR U26214 ( .A(n26274), .B(n26277), .Z(n26275) );
  XOR U26215 ( .A(n26278), .B(n26279), .Z(n26262) );
  XOR U26216 ( .A(n26280), .B(n26281), .Z(n26279) );
  ANDN U26217 ( .B(n26282), .A(n26283), .Z(n26280) );
  XOR U26218 ( .A(n26284), .B(n26281), .Z(n26282) );
  IV U26219 ( .A(n26260), .Z(n26278) );
  XOR U26220 ( .A(n26285), .B(n26286), .Z(n26260) );
  ANDN U26221 ( .B(n26287), .A(n26288), .Z(n26285) );
  XOR U26222 ( .A(n26286), .B(n26289), .Z(n26287) );
  IV U26223 ( .A(n26268), .Z(n26272) );
  XOR U26224 ( .A(n26268), .B(n26250), .Z(n26270) );
  XOR U26225 ( .A(n26290), .B(n26291), .Z(n26250) );
  AND U26226 ( .A(n1402), .B(n26292), .Z(n26290) );
  XOR U26227 ( .A(n26293), .B(n26291), .Z(n26292) );
  NANDN U26228 ( .A(n26252), .B(n26254), .Z(n26268) );
  XOR U26229 ( .A(n26294), .B(n26295), .Z(n26254) );
  AND U26230 ( .A(n1402), .B(n26296), .Z(n26294) );
  XOR U26231 ( .A(n26295), .B(n26297), .Z(n26296) );
  XOR U26232 ( .A(n26298), .B(n26299), .Z(n1402) );
  AND U26233 ( .A(n26300), .B(n26301), .Z(n26298) );
  XNOR U26234 ( .A(n26299), .B(n26265), .Z(n26301) );
  XNOR U26235 ( .A(n26302), .B(n26303), .Z(n26265) );
  ANDN U26236 ( .B(n26304), .A(n26305), .Z(n26302) );
  XOR U26237 ( .A(n26303), .B(n26306), .Z(n26304) );
  XOR U26238 ( .A(n26299), .B(n26267), .Z(n26300) );
  XOR U26239 ( .A(n26307), .B(n26308), .Z(n26267) );
  AND U26240 ( .A(n1406), .B(n26309), .Z(n26307) );
  XOR U26241 ( .A(n26310), .B(n26308), .Z(n26309) );
  XNOR U26242 ( .A(n26311), .B(n26312), .Z(n26299) );
  NAND U26243 ( .A(n26313), .B(n26314), .Z(n26312) );
  XOR U26244 ( .A(n26315), .B(n26291), .Z(n26314) );
  XOR U26245 ( .A(n26305), .B(n26306), .Z(n26291) );
  XOR U26246 ( .A(n26316), .B(n26317), .Z(n26306) );
  ANDN U26247 ( .B(n26318), .A(n26319), .Z(n26316) );
  XOR U26248 ( .A(n26317), .B(n26320), .Z(n26318) );
  XOR U26249 ( .A(n26321), .B(n26322), .Z(n26305) );
  XOR U26250 ( .A(n26323), .B(n26324), .Z(n26322) );
  ANDN U26251 ( .B(n26325), .A(n26326), .Z(n26323) );
  XOR U26252 ( .A(n26327), .B(n26324), .Z(n26325) );
  IV U26253 ( .A(n26303), .Z(n26321) );
  XOR U26254 ( .A(n26328), .B(n26329), .Z(n26303) );
  ANDN U26255 ( .B(n26330), .A(n26331), .Z(n26328) );
  XOR U26256 ( .A(n26329), .B(n26332), .Z(n26330) );
  IV U26257 ( .A(n26311), .Z(n26315) );
  XOR U26258 ( .A(n26311), .B(n26293), .Z(n26313) );
  XOR U26259 ( .A(n26333), .B(n26334), .Z(n26293) );
  AND U26260 ( .A(n1406), .B(n26335), .Z(n26333) );
  XOR U26261 ( .A(n26336), .B(n26334), .Z(n26335) );
  NANDN U26262 ( .A(n26295), .B(n26297), .Z(n26311) );
  XOR U26263 ( .A(n26337), .B(n26338), .Z(n26297) );
  AND U26264 ( .A(n1406), .B(n26339), .Z(n26337) );
  XOR U26265 ( .A(n26338), .B(n26340), .Z(n26339) );
  XOR U26266 ( .A(n26341), .B(n26342), .Z(n1406) );
  AND U26267 ( .A(n26343), .B(n26344), .Z(n26341) );
  XNOR U26268 ( .A(n26342), .B(n26308), .Z(n26344) );
  XNOR U26269 ( .A(n26345), .B(n26346), .Z(n26308) );
  ANDN U26270 ( .B(n26347), .A(n26348), .Z(n26345) );
  XOR U26271 ( .A(n26346), .B(n26349), .Z(n26347) );
  XOR U26272 ( .A(n26342), .B(n26310), .Z(n26343) );
  XOR U26273 ( .A(n26350), .B(n26351), .Z(n26310) );
  AND U26274 ( .A(n1410), .B(n26352), .Z(n26350) );
  XOR U26275 ( .A(n26353), .B(n26351), .Z(n26352) );
  XNOR U26276 ( .A(n26354), .B(n26355), .Z(n26342) );
  NAND U26277 ( .A(n26356), .B(n26357), .Z(n26355) );
  XOR U26278 ( .A(n26358), .B(n26334), .Z(n26357) );
  XOR U26279 ( .A(n26348), .B(n26349), .Z(n26334) );
  XOR U26280 ( .A(n26359), .B(n26360), .Z(n26349) );
  ANDN U26281 ( .B(n26361), .A(n26362), .Z(n26359) );
  XOR U26282 ( .A(n26360), .B(n26363), .Z(n26361) );
  XOR U26283 ( .A(n26364), .B(n26365), .Z(n26348) );
  XOR U26284 ( .A(n26366), .B(n26367), .Z(n26365) );
  ANDN U26285 ( .B(n26368), .A(n26369), .Z(n26366) );
  XOR U26286 ( .A(n26370), .B(n26367), .Z(n26368) );
  IV U26287 ( .A(n26346), .Z(n26364) );
  XOR U26288 ( .A(n26371), .B(n26372), .Z(n26346) );
  ANDN U26289 ( .B(n26373), .A(n26374), .Z(n26371) );
  XOR U26290 ( .A(n26372), .B(n26375), .Z(n26373) );
  IV U26291 ( .A(n26354), .Z(n26358) );
  XOR U26292 ( .A(n26354), .B(n26336), .Z(n26356) );
  XOR U26293 ( .A(n26376), .B(n26377), .Z(n26336) );
  AND U26294 ( .A(n1410), .B(n26378), .Z(n26376) );
  XOR U26295 ( .A(n26379), .B(n26377), .Z(n26378) );
  NANDN U26296 ( .A(n26338), .B(n26340), .Z(n26354) );
  XOR U26297 ( .A(n26380), .B(n26381), .Z(n26340) );
  AND U26298 ( .A(n1410), .B(n26382), .Z(n26380) );
  XOR U26299 ( .A(n26381), .B(n26383), .Z(n26382) );
  XOR U26300 ( .A(n26384), .B(n26385), .Z(n1410) );
  AND U26301 ( .A(n26386), .B(n26387), .Z(n26384) );
  XNOR U26302 ( .A(n26385), .B(n26351), .Z(n26387) );
  XNOR U26303 ( .A(n26388), .B(n26389), .Z(n26351) );
  ANDN U26304 ( .B(n26390), .A(n26391), .Z(n26388) );
  XOR U26305 ( .A(n26389), .B(n26392), .Z(n26390) );
  XOR U26306 ( .A(n26385), .B(n26353), .Z(n26386) );
  XOR U26307 ( .A(n26393), .B(n26394), .Z(n26353) );
  AND U26308 ( .A(n1414), .B(n26395), .Z(n26393) );
  XOR U26309 ( .A(n26396), .B(n26394), .Z(n26395) );
  XNOR U26310 ( .A(n26397), .B(n26398), .Z(n26385) );
  NAND U26311 ( .A(n26399), .B(n26400), .Z(n26398) );
  XOR U26312 ( .A(n26401), .B(n26377), .Z(n26400) );
  XOR U26313 ( .A(n26391), .B(n26392), .Z(n26377) );
  XOR U26314 ( .A(n26402), .B(n26403), .Z(n26392) );
  ANDN U26315 ( .B(n26404), .A(n26405), .Z(n26402) );
  XOR U26316 ( .A(n26403), .B(n26406), .Z(n26404) );
  XOR U26317 ( .A(n26407), .B(n26408), .Z(n26391) );
  XOR U26318 ( .A(n26409), .B(n26410), .Z(n26408) );
  ANDN U26319 ( .B(n26411), .A(n26412), .Z(n26409) );
  XOR U26320 ( .A(n26413), .B(n26410), .Z(n26411) );
  IV U26321 ( .A(n26389), .Z(n26407) );
  XOR U26322 ( .A(n26414), .B(n26415), .Z(n26389) );
  ANDN U26323 ( .B(n26416), .A(n26417), .Z(n26414) );
  XOR U26324 ( .A(n26415), .B(n26418), .Z(n26416) );
  IV U26325 ( .A(n26397), .Z(n26401) );
  XOR U26326 ( .A(n26397), .B(n26379), .Z(n26399) );
  XOR U26327 ( .A(n26419), .B(n26420), .Z(n26379) );
  AND U26328 ( .A(n1414), .B(n26421), .Z(n26419) );
  XOR U26329 ( .A(n26422), .B(n26420), .Z(n26421) );
  NANDN U26330 ( .A(n26381), .B(n26383), .Z(n26397) );
  XOR U26331 ( .A(n26423), .B(n26424), .Z(n26383) );
  AND U26332 ( .A(n1414), .B(n26425), .Z(n26423) );
  XOR U26333 ( .A(n26424), .B(n26426), .Z(n26425) );
  XOR U26334 ( .A(n26427), .B(n26428), .Z(n1414) );
  AND U26335 ( .A(n26429), .B(n26430), .Z(n26427) );
  XNOR U26336 ( .A(n26428), .B(n26394), .Z(n26430) );
  XNOR U26337 ( .A(n26431), .B(n26432), .Z(n26394) );
  ANDN U26338 ( .B(n26433), .A(n26434), .Z(n26431) );
  XOR U26339 ( .A(n26432), .B(n26435), .Z(n26433) );
  XOR U26340 ( .A(n26428), .B(n26396), .Z(n26429) );
  XOR U26341 ( .A(n26436), .B(n26437), .Z(n26396) );
  AND U26342 ( .A(n1418), .B(n26438), .Z(n26436) );
  XOR U26343 ( .A(n26439), .B(n26437), .Z(n26438) );
  XNOR U26344 ( .A(n26440), .B(n26441), .Z(n26428) );
  NAND U26345 ( .A(n26442), .B(n26443), .Z(n26441) );
  XOR U26346 ( .A(n26444), .B(n26420), .Z(n26443) );
  XOR U26347 ( .A(n26434), .B(n26435), .Z(n26420) );
  XOR U26348 ( .A(n26445), .B(n26446), .Z(n26435) );
  ANDN U26349 ( .B(n26447), .A(n26448), .Z(n26445) );
  XOR U26350 ( .A(n26446), .B(n26449), .Z(n26447) );
  XOR U26351 ( .A(n26450), .B(n26451), .Z(n26434) );
  XOR U26352 ( .A(n26452), .B(n26453), .Z(n26451) );
  ANDN U26353 ( .B(n26454), .A(n26455), .Z(n26452) );
  XOR U26354 ( .A(n26456), .B(n26453), .Z(n26454) );
  IV U26355 ( .A(n26432), .Z(n26450) );
  XOR U26356 ( .A(n26457), .B(n26458), .Z(n26432) );
  ANDN U26357 ( .B(n26459), .A(n26460), .Z(n26457) );
  XOR U26358 ( .A(n26458), .B(n26461), .Z(n26459) );
  IV U26359 ( .A(n26440), .Z(n26444) );
  XOR U26360 ( .A(n26440), .B(n26422), .Z(n26442) );
  XOR U26361 ( .A(n26462), .B(n26463), .Z(n26422) );
  AND U26362 ( .A(n1418), .B(n26464), .Z(n26462) );
  XOR U26363 ( .A(n26465), .B(n26463), .Z(n26464) );
  NANDN U26364 ( .A(n26424), .B(n26426), .Z(n26440) );
  XOR U26365 ( .A(n26466), .B(n26467), .Z(n26426) );
  AND U26366 ( .A(n1418), .B(n26468), .Z(n26466) );
  XOR U26367 ( .A(n26467), .B(n26469), .Z(n26468) );
  XOR U26368 ( .A(n26470), .B(n26471), .Z(n1418) );
  AND U26369 ( .A(n26472), .B(n26473), .Z(n26470) );
  XNOR U26370 ( .A(n26471), .B(n26437), .Z(n26473) );
  XNOR U26371 ( .A(n26474), .B(n26475), .Z(n26437) );
  ANDN U26372 ( .B(n26476), .A(n26477), .Z(n26474) );
  XOR U26373 ( .A(n26475), .B(n26478), .Z(n26476) );
  XOR U26374 ( .A(n26471), .B(n26439), .Z(n26472) );
  XOR U26375 ( .A(n26479), .B(n26480), .Z(n26439) );
  AND U26376 ( .A(n1422), .B(n26481), .Z(n26479) );
  XOR U26377 ( .A(n26482), .B(n26480), .Z(n26481) );
  XNOR U26378 ( .A(n26483), .B(n26484), .Z(n26471) );
  NAND U26379 ( .A(n26485), .B(n26486), .Z(n26484) );
  XOR U26380 ( .A(n26487), .B(n26463), .Z(n26486) );
  XOR U26381 ( .A(n26477), .B(n26478), .Z(n26463) );
  XOR U26382 ( .A(n26488), .B(n26489), .Z(n26478) );
  ANDN U26383 ( .B(n26490), .A(n26491), .Z(n26488) );
  XOR U26384 ( .A(n26489), .B(n26492), .Z(n26490) );
  XOR U26385 ( .A(n26493), .B(n26494), .Z(n26477) );
  XOR U26386 ( .A(n26495), .B(n26496), .Z(n26494) );
  ANDN U26387 ( .B(n26497), .A(n26498), .Z(n26495) );
  XOR U26388 ( .A(n26499), .B(n26496), .Z(n26497) );
  IV U26389 ( .A(n26475), .Z(n26493) );
  XOR U26390 ( .A(n26500), .B(n26501), .Z(n26475) );
  ANDN U26391 ( .B(n26502), .A(n26503), .Z(n26500) );
  XOR U26392 ( .A(n26501), .B(n26504), .Z(n26502) );
  IV U26393 ( .A(n26483), .Z(n26487) );
  XOR U26394 ( .A(n26483), .B(n26465), .Z(n26485) );
  XOR U26395 ( .A(n26505), .B(n26506), .Z(n26465) );
  AND U26396 ( .A(n1422), .B(n26507), .Z(n26505) );
  XOR U26397 ( .A(n26508), .B(n26506), .Z(n26507) );
  NANDN U26398 ( .A(n26467), .B(n26469), .Z(n26483) );
  XOR U26399 ( .A(n26509), .B(n26510), .Z(n26469) );
  AND U26400 ( .A(n1422), .B(n26511), .Z(n26509) );
  XOR U26401 ( .A(n26510), .B(n26512), .Z(n26511) );
  XOR U26402 ( .A(n26513), .B(n26514), .Z(n1422) );
  AND U26403 ( .A(n26515), .B(n26516), .Z(n26513) );
  XNOR U26404 ( .A(n26514), .B(n26480), .Z(n26516) );
  XNOR U26405 ( .A(n26517), .B(n26518), .Z(n26480) );
  ANDN U26406 ( .B(n26519), .A(n26520), .Z(n26517) );
  XOR U26407 ( .A(n26518), .B(n26521), .Z(n26519) );
  XOR U26408 ( .A(n26514), .B(n26482), .Z(n26515) );
  XOR U26409 ( .A(n26522), .B(n26523), .Z(n26482) );
  AND U26410 ( .A(n1426), .B(n26524), .Z(n26522) );
  XOR U26411 ( .A(n26525), .B(n26523), .Z(n26524) );
  XNOR U26412 ( .A(n26526), .B(n26527), .Z(n26514) );
  NAND U26413 ( .A(n26528), .B(n26529), .Z(n26527) );
  XOR U26414 ( .A(n26530), .B(n26506), .Z(n26529) );
  XOR U26415 ( .A(n26520), .B(n26521), .Z(n26506) );
  XOR U26416 ( .A(n26531), .B(n26532), .Z(n26521) );
  ANDN U26417 ( .B(n26533), .A(n26534), .Z(n26531) );
  XOR U26418 ( .A(n26532), .B(n26535), .Z(n26533) );
  XOR U26419 ( .A(n26536), .B(n26537), .Z(n26520) );
  XOR U26420 ( .A(n26538), .B(n26539), .Z(n26537) );
  ANDN U26421 ( .B(n26540), .A(n26541), .Z(n26538) );
  XOR U26422 ( .A(n26542), .B(n26539), .Z(n26540) );
  IV U26423 ( .A(n26518), .Z(n26536) );
  XOR U26424 ( .A(n26543), .B(n26544), .Z(n26518) );
  ANDN U26425 ( .B(n26545), .A(n26546), .Z(n26543) );
  XOR U26426 ( .A(n26544), .B(n26547), .Z(n26545) );
  IV U26427 ( .A(n26526), .Z(n26530) );
  XOR U26428 ( .A(n26526), .B(n26508), .Z(n26528) );
  XOR U26429 ( .A(n26548), .B(n26549), .Z(n26508) );
  AND U26430 ( .A(n1426), .B(n26550), .Z(n26548) );
  XOR U26431 ( .A(n26551), .B(n26549), .Z(n26550) );
  NANDN U26432 ( .A(n26510), .B(n26512), .Z(n26526) );
  XOR U26433 ( .A(n26552), .B(n26553), .Z(n26512) );
  AND U26434 ( .A(n1426), .B(n26554), .Z(n26552) );
  XOR U26435 ( .A(n26553), .B(n26555), .Z(n26554) );
  XOR U26436 ( .A(n26556), .B(n26557), .Z(n1426) );
  AND U26437 ( .A(n26558), .B(n26559), .Z(n26556) );
  XNOR U26438 ( .A(n26557), .B(n26523), .Z(n26559) );
  XNOR U26439 ( .A(n26560), .B(n26561), .Z(n26523) );
  ANDN U26440 ( .B(n26562), .A(n26563), .Z(n26560) );
  XOR U26441 ( .A(n26561), .B(n26564), .Z(n26562) );
  XOR U26442 ( .A(n26557), .B(n26525), .Z(n26558) );
  XOR U26443 ( .A(n26565), .B(n26566), .Z(n26525) );
  AND U26444 ( .A(n1430), .B(n26567), .Z(n26565) );
  XOR U26445 ( .A(n26568), .B(n26566), .Z(n26567) );
  XNOR U26446 ( .A(n26569), .B(n26570), .Z(n26557) );
  NAND U26447 ( .A(n26571), .B(n26572), .Z(n26570) );
  XOR U26448 ( .A(n26573), .B(n26549), .Z(n26572) );
  XOR U26449 ( .A(n26563), .B(n26564), .Z(n26549) );
  XOR U26450 ( .A(n26574), .B(n26575), .Z(n26564) );
  ANDN U26451 ( .B(n26576), .A(n26577), .Z(n26574) );
  XOR U26452 ( .A(n26575), .B(n26578), .Z(n26576) );
  XOR U26453 ( .A(n26579), .B(n26580), .Z(n26563) );
  XOR U26454 ( .A(n26581), .B(n26582), .Z(n26580) );
  ANDN U26455 ( .B(n26583), .A(n26584), .Z(n26581) );
  XOR U26456 ( .A(n26585), .B(n26582), .Z(n26583) );
  IV U26457 ( .A(n26561), .Z(n26579) );
  XOR U26458 ( .A(n26586), .B(n26587), .Z(n26561) );
  ANDN U26459 ( .B(n26588), .A(n26589), .Z(n26586) );
  XOR U26460 ( .A(n26587), .B(n26590), .Z(n26588) );
  IV U26461 ( .A(n26569), .Z(n26573) );
  XOR U26462 ( .A(n26569), .B(n26551), .Z(n26571) );
  XOR U26463 ( .A(n26591), .B(n26592), .Z(n26551) );
  AND U26464 ( .A(n1430), .B(n26593), .Z(n26591) );
  XOR U26465 ( .A(n26594), .B(n26592), .Z(n26593) );
  NANDN U26466 ( .A(n26553), .B(n26555), .Z(n26569) );
  XOR U26467 ( .A(n26595), .B(n26596), .Z(n26555) );
  AND U26468 ( .A(n1430), .B(n26597), .Z(n26595) );
  XOR U26469 ( .A(n26596), .B(n26598), .Z(n26597) );
  XOR U26470 ( .A(n26599), .B(n26600), .Z(n1430) );
  AND U26471 ( .A(n26601), .B(n26602), .Z(n26599) );
  XNOR U26472 ( .A(n26600), .B(n26566), .Z(n26602) );
  XNOR U26473 ( .A(n26603), .B(n26604), .Z(n26566) );
  ANDN U26474 ( .B(n26605), .A(n26606), .Z(n26603) );
  XOR U26475 ( .A(n26604), .B(n26607), .Z(n26605) );
  XOR U26476 ( .A(n26600), .B(n26568), .Z(n26601) );
  XOR U26477 ( .A(n26608), .B(n26609), .Z(n26568) );
  AND U26478 ( .A(n1434), .B(n26610), .Z(n26608) );
  XOR U26479 ( .A(n26611), .B(n26609), .Z(n26610) );
  XNOR U26480 ( .A(n26612), .B(n26613), .Z(n26600) );
  NAND U26481 ( .A(n26614), .B(n26615), .Z(n26613) );
  XOR U26482 ( .A(n26616), .B(n26592), .Z(n26615) );
  XOR U26483 ( .A(n26606), .B(n26607), .Z(n26592) );
  XOR U26484 ( .A(n26617), .B(n26618), .Z(n26607) );
  ANDN U26485 ( .B(n26619), .A(n26620), .Z(n26617) );
  XOR U26486 ( .A(n26618), .B(n26621), .Z(n26619) );
  XOR U26487 ( .A(n26622), .B(n26623), .Z(n26606) );
  XOR U26488 ( .A(n26624), .B(n26625), .Z(n26623) );
  ANDN U26489 ( .B(n26626), .A(n26627), .Z(n26624) );
  XOR U26490 ( .A(n26628), .B(n26625), .Z(n26626) );
  IV U26491 ( .A(n26604), .Z(n26622) );
  XOR U26492 ( .A(n26629), .B(n26630), .Z(n26604) );
  ANDN U26493 ( .B(n26631), .A(n26632), .Z(n26629) );
  XOR U26494 ( .A(n26630), .B(n26633), .Z(n26631) );
  IV U26495 ( .A(n26612), .Z(n26616) );
  XOR U26496 ( .A(n26612), .B(n26594), .Z(n26614) );
  XOR U26497 ( .A(n26634), .B(n26635), .Z(n26594) );
  AND U26498 ( .A(n1434), .B(n26636), .Z(n26634) );
  XOR U26499 ( .A(n26637), .B(n26635), .Z(n26636) );
  NANDN U26500 ( .A(n26596), .B(n26598), .Z(n26612) );
  XOR U26501 ( .A(n26638), .B(n26639), .Z(n26598) );
  AND U26502 ( .A(n1434), .B(n26640), .Z(n26638) );
  XOR U26503 ( .A(n26639), .B(n26641), .Z(n26640) );
  XOR U26504 ( .A(n26642), .B(n26643), .Z(n1434) );
  AND U26505 ( .A(n26644), .B(n26645), .Z(n26642) );
  XNOR U26506 ( .A(n26643), .B(n26609), .Z(n26645) );
  XNOR U26507 ( .A(n26646), .B(n26647), .Z(n26609) );
  ANDN U26508 ( .B(n26648), .A(n26649), .Z(n26646) );
  XOR U26509 ( .A(n26647), .B(n26650), .Z(n26648) );
  XOR U26510 ( .A(n26643), .B(n26611), .Z(n26644) );
  XOR U26511 ( .A(n26651), .B(n26652), .Z(n26611) );
  AND U26512 ( .A(n1438), .B(n26653), .Z(n26651) );
  XOR U26513 ( .A(n26654), .B(n26652), .Z(n26653) );
  XNOR U26514 ( .A(n26655), .B(n26656), .Z(n26643) );
  NAND U26515 ( .A(n26657), .B(n26658), .Z(n26656) );
  XOR U26516 ( .A(n26659), .B(n26635), .Z(n26658) );
  XOR U26517 ( .A(n26649), .B(n26650), .Z(n26635) );
  XOR U26518 ( .A(n26660), .B(n26661), .Z(n26650) );
  ANDN U26519 ( .B(n26662), .A(n26663), .Z(n26660) );
  XOR U26520 ( .A(n26661), .B(n26664), .Z(n26662) );
  XOR U26521 ( .A(n26665), .B(n26666), .Z(n26649) );
  XOR U26522 ( .A(n26667), .B(n26668), .Z(n26666) );
  ANDN U26523 ( .B(n26669), .A(n26670), .Z(n26667) );
  XOR U26524 ( .A(n26671), .B(n26668), .Z(n26669) );
  IV U26525 ( .A(n26647), .Z(n26665) );
  XOR U26526 ( .A(n26672), .B(n26673), .Z(n26647) );
  ANDN U26527 ( .B(n26674), .A(n26675), .Z(n26672) );
  XOR U26528 ( .A(n26673), .B(n26676), .Z(n26674) );
  IV U26529 ( .A(n26655), .Z(n26659) );
  XOR U26530 ( .A(n26655), .B(n26637), .Z(n26657) );
  XOR U26531 ( .A(n26677), .B(n26678), .Z(n26637) );
  AND U26532 ( .A(n1438), .B(n26679), .Z(n26677) );
  XOR U26533 ( .A(n26680), .B(n26678), .Z(n26679) );
  NANDN U26534 ( .A(n26639), .B(n26641), .Z(n26655) );
  XOR U26535 ( .A(n26681), .B(n26682), .Z(n26641) );
  AND U26536 ( .A(n1438), .B(n26683), .Z(n26681) );
  XOR U26537 ( .A(n26682), .B(n26684), .Z(n26683) );
  XOR U26538 ( .A(n26685), .B(n26686), .Z(n1438) );
  AND U26539 ( .A(n26687), .B(n26688), .Z(n26685) );
  XNOR U26540 ( .A(n26686), .B(n26652), .Z(n26688) );
  XNOR U26541 ( .A(n26689), .B(n26690), .Z(n26652) );
  ANDN U26542 ( .B(n26691), .A(n26692), .Z(n26689) );
  XOR U26543 ( .A(n26690), .B(n26693), .Z(n26691) );
  XOR U26544 ( .A(n26686), .B(n26654), .Z(n26687) );
  XOR U26545 ( .A(n26694), .B(n26695), .Z(n26654) );
  AND U26546 ( .A(n1442), .B(n26696), .Z(n26694) );
  XOR U26547 ( .A(n26697), .B(n26695), .Z(n26696) );
  XNOR U26548 ( .A(n26698), .B(n26699), .Z(n26686) );
  NAND U26549 ( .A(n26700), .B(n26701), .Z(n26699) );
  XOR U26550 ( .A(n26702), .B(n26678), .Z(n26701) );
  XOR U26551 ( .A(n26692), .B(n26693), .Z(n26678) );
  XOR U26552 ( .A(n26703), .B(n26704), .Z(n26693) );
  ANDN U26553 ( .B(n26705), .A(n26706), .Z(n26703) );
  XOR U26554 ( .A(n26704), .B(n26707), .Z(n26705) );
  XOR U26555 ( .A(n26708), .B(n26709), .Z(n26692) );
  XOR U26556 ( .A(n26710), .B(n26711), .Z(n26709) );
  ANDN U26557 ( .B(n26712), .A(n26713), .Z(n26710) );
  XOR U26558 ( .A(n26714), .B(n26711), .Z(n26712) );
  IV U26559 ( .A(n26690), .Z(n26708) );
  XOR U26560 ( .A(n26715), .B(n26716), .Z(n26690) );
  ANDN U26561 ( .B(n26717), .A(n26718), .Z(n26715) );
  XOR U26562 ( .A(n26716), .B(n26719), .Z(n26717) );
  IV U26563 ( .A(n26698), .Z(n26702) );
  XOR U26564 ( .A(n26698), .B(n26680), .Z(n26700) );
  XOR U26565 ( .A(n26720), .B(n26721), .Z(n26680) );
  AND U26566 ( .A(n1442), .B(n26722), .Z(n26720) );
  XOR U26567 ( .A(n26723), .B(n26721), .Z(n26722) );
  NANDN U26568 ( .A(n26682), .B(n26684), .Z(n26698) );
  XOR U26569 ( .A(n26724), .B(n26725), .Z(n26684) );
  AND U26570 ( .A(n1442), .B(n26726), .Z(n26724) );
  XOR U26571 ( .A(n26725), .B(n26727), .Z(n26726) );
  XOR U26572 ( .A(n26728), .B(n26729), .Z(n1442) );
  AND U26573 ( .A(n26730), .B(n26731), .Z(n26728) );
  XNOR U26574 ( .A(n26729), .B(n26695), .Z(n26731) );
  XNOR U26575 ( .A(n26732), .B(n26733), .Z(n26695) );
  ANDN U26576 ( .B(n26734), .A(n26735), .Z(n26732) );
  XOR U26577 ( .A(n26733), .B(n26736), .Z(n26734) );
  XOR U26578 ( .A(n26729), .B(n26697), .Z(n26730) );
  XOR U26579 ( .A(n26737), .B(n26738), .Z(n26697) );
  AND U26580 ( .A(n1446), .B(n26739), .Z(n26737) );
  XOR U26581 ( .A(n26740), .B(n26738), .Z(n26739) );
  XNOR U26582 ( .A(n26741), .B(n26742), .Z(n26729) );
  NAND U26583 ( .A(n26743), .B(n26744), .Z(n26742) );
  XOR U26584 ( .A(n26745), .B(n26721), .Z(n26744) );
  XOR U26585 ( .A(n26735), .B(n26736), .Z(n26721) );
  XOR U26586 ( .A(n26746), .B(n26747), .Z(n26736) );
  ANDN U26587 ( .B(n26748), .A(n26749), .Z(n26746) );
  XOR U26588 ( .A(n26747), .B(n26750), .Z(n26748) );
  XOR U26589 ( .A(n26751), .B(n26752), .Z(n26735) );
  XOR U26590 ( .A(n26753), .B(n26754), .Z(n26752) );
  ANDN U26591 ( .B(n26755), .A(n26756), .Z(n26753) );
  XOR U26592 ( .A(n26757), .B(n26754), .Z(n26755) );
  IV U26593 ( .A(n26733), .Z(n26751) );
  XOR U26594 ( .A(n26758), .B(n26759), .Z(n26733) );
  ANDN U26595 ( .B(n26760), .A(n26761), .Z(n26758) );
  XOR U26596 ( .A(n26759), .B(n26762), .Z(n26760) );
  IV U26597 ( .A(n26741), .Z(n26745) );
  XOR U26598 ( .A(n26741), .B(n26723), .Z(n26743) );
  XOR U26599 ( .A(n26763), .B(n26764), .Z(n26723) );
  AND U26600 ( .A(n1446), .B(n26765), .Z(n26763) );
  XOR U26601 ( .A(n26766), .B(n26764), .Z(n26765) );
  NANDN U26602 ( .A(n26725), .B(n26727), .Z(n26741) );
  XOR U26603 ( .A(n26767), .B(n26768), .Z(n26727) );
  AND U26604 ( .A(n1446), .B(n26769), .Z(n26767) );
  XOR U26605 ( .A(n26768), .B(n26770), .Z(n26769) );
  XOR U26606 ( .A(n26771), .B(n26772), .Z(n1446) );
  AND U26607 ( .A(n26773), .B(n26774), .Z(n26771) );
  XNOR U26608 ( .A(n26772), .B(n26738), .Z(n26774) );
  XNOR U26609 ( .A(n26775), .B(n26776), .Z(n26738) );
  ANDN U26610 ( .B(n26777), .A(n26778), .Z(n26775) );
  XOR U26611 ( .A(n26776), .B(n26779), .Z(n26777) );
  XOR U26612 ( .A(n26772), .B(n26740), .Z(n26773) );
  XOR U26613 ( .A(n26780), .B(n26781), .Z(n26740) );
  AND U26614 ( .A(n1450), .B(n26782), .Z(n26780) );
  XOR U26615 ( .A(n26783), .B(n26781), .Z(n26782) );
  XNOR U26616 ( .A(n26784), .B(n26785), .Z(n26772) );
  NAND U26617 ( .A(n26786), .B(n26787), .Z(n26785) );
  XOR U26618 ( .A(n26788), .B(n26764), .Z(n26787) );
  XOR U26619 ( .A(n26778), .B(n26779), .Z(n26764) );
  XOR U26620 ( .A(n26789), .B(n26790), .Z(n26779) );
  ANDN U26621 ( .B(n26791), .A(n26792), .Z(n26789) );
  XOR U26622 ( .A(n26790), .B(n26793), .Z(n26791) );
  XOR U26623 ( .A(n26794), .B(n26795), .Z(n26778) );
  XOR U26624 ( .A(n26796), .B(n26797), .Z(n26795) );
  ANDN U26625 ( .B(n26798), .A(n26799), .Z(n26796) );
  XOR U26626 ( .A(n26800), .B(n26797), .Z(n26798) );
  IV U26627 ( .A(n26776), .Z(n26794) );
  XOR U26628 ( .A(n26801), .B(n26802), .Z(n26776) );
  ANDN U26629 ( .B(n26803), .A(n26804), .Z(n26801) );
  XOR U26630 ( .A(n26802), .B(n26805), .Z(n26803) );
  IV U26631 ( .A(n26784), .Z(n26788) );
  XOR U26632 ( .A(n26784), .B(n26766), .Z(n26786) );
  XOR U26633 ( .A(n26806), .B(n26807), .Z(n26766) );
  AND U26634 ( .A(n1450), .B(n26808), .Z(n26806) );
  XOR U26635 ( .A(n26809), .B(n26807), .Z(n26808) );
  NANDN U26636 ( .A(n26768), .B(n26770), .Z(n26784) );
  XOR U26637 ( .A(n26810), .B(n26811), .Z(n26770) );
  AND U26638 ( .A(n1450), .B(n26812), .Z(n26810) );
  XOR U26639 ( .A(n26811), .B(n26813), .Z(n26812) );
  XOR U26640 ( .A(n26814), .B(n26815), .Z(n1450) );
  AND U26641 ( .A(n26816), .B(n26817), .Z(n26814) );
  XNOR U26642 ( .A(n26815), .B(n26781), .Z(n26817) );
  XNOR U26643 ( .A(n26818), .B(n26819), .Z(n26781) );
  ANDN U26644 ( .B(n26820), .A(n26821), .Z(n26818) );
  XOR U26645 ( .A(n26819), .B(n26822), .Z(n26820) );
  XOR U26646 ( .A(n26815), .B(n26783), .Z(n26816) );
  XOR U26647 ( .A(n26823), .B(n26824), .Z(n26783) );
  AND U26648 ( .A(n1454), .B(n26825), .Z(n26823) );
  XOR U26649 ( .A(n26826), .B(n26824), .Z(n26825) );
  XNOR U26650 ( .A(n26827), .B(n26828), .Z(n26815) );
  NAND U26651 ( .A(n26829), .B(n26830), .Z(n26828) );
  XOR U26652 ( .A(n26831), .B(n26807), .Z(n26830) );
  XOR U26653 ( .A(n26821), .B(n26822), .Z(n26807) );
  XOR U26654 ( .A(n26832), .B(n26833), .Z(n26822) );
  ANDN U26655 ( .B(n26834), .A(n26835), .Z(n26832) );
  XOR U26656 ( .A(n26833), .B(n26836), .Z(n26834) );
  XOR U26657 ( .A(n26837), .B(n26838), .Z(n26821) );
  XOR U26658 ( .A(n26839), .B(n26840), .Z(n26838) );
  ANDN U26659 ( .B(n26841), .A(n26842), .Z(n26839) );
  XOR U26660 ( .A(n26843), .B(n26840), .Z(n26841) );
  IV U26661 ( .A(n26819), .Z(n26837) );
  XOR U26662 ( .A(n26844), .B(n26845), .Z(n26819) );
  ANDN U26663 ( .B(n26846), .A(n26847), .Z(n26844) );
  XOR U26664 ( .A(n26845), .B(n26848), .Z(n26846) );
  IV U26665 ( .A(n26827), .Z(n26831) );
  XOR U26666 ( .A(n26827), .B(n26809), .Z(n26829) );
  XOR U26667 ( .A(n26849), .B(n26850), .Z(n26809) );
  AND U26668 ( .A(n1454), .B(n26851), .Z(n26849) );
  XOR U26669 ( .A(n26852), .B(n26850), .Z(n26851) );
  NANDN U26670 ( .A(n26811), .B(n26813), .Z(n26827) );
  XOR U26671 ( .A(n26853), .B(n26854), .Z(n26813) );
  AND U26672 ( .A(n1454), .B(n26855), .Z(n26853) );
  XOR U26673 ( .A(n26854), .B(n26856), .Z(n26855) );
  XOR U26674 ( .A(n26857), .B(n26858), .Z(n1454) );
  AND U26675 ( .A(n26859), .B(n26860), .Z(n26857) );
  XNOR U26676 ( .A(n26858), .B(n26824), .Z(n26860) );
  XNOR U26677 ( .A(n26861), .B(n26862), .Z(n26824) );
  ANDN U26678 ( .B(n26863), .A(n26864), .Z(n26861) );
  XOR U26679 ( .A(n26862), .B(n26865), .Z(n26863) );
  XOR U26680 ( .A(n26858), .B(n26826), .Z(n26859) );
  XOR U26681 ( .A(n26866), .B(n26867), .Z(n26826) );
  AND U26682 ( .A(n1458), .B(n26868), .Z(n26866) );
  XOR U26683 ( .A(n26869), .B(n26867), .Z(n26868) );
  XNOR U26684 ( .A(n26870), .B(n26871), .Z(n26858) );
  NAND U26685 ( .A(n26872), .B(n26873), .Z(n26871) );
  XOR U26686 ( .A(n26874), .B(n26850), .Z(n26873) );
  XOR U26687 ( .A(n26864), .B(n26865), .Z(n26850) );
  XOR U26688 ( .A(n26875), .B(n26876), .Z(n26865) );
  ANDN U26689 ( .B(n26877), .A(n26878), .Z(n26875) );
  XOR U26690 ( .A(n26876), .B(n26879), .Z(n26877) );
  XOR U26691 ( .A(n26880), .B(n26881), .Z(n26864) );
  XOR U26692 ( .A(n26882), .B(n26883), .Z(n26881) );
  ANDN U26693 ( .B(n26884), .A(n26885), .Z(n26882) );
  XOR U26694 ( .A(n26886), .B(n26883), .Z(n26884) );
  IV U26695 ( .A(n26862), .Z(n26880) );
  XOR U26696 ( .A(n26887), .B(n26888), .Z(n26862) );
  ANDN U26697 ( .B(n26889), .A(n26890), .Z(n26887) );
  XOR U26698 ( .A(n26888), .B(n26891), .Z(n26889) );
  IV U26699 ( .A(n26870), .Z(n26874) );
  XOR U26700 ( .A(n26870), .B(n26852), .Z(n26872) );
  XOR U26701 ( .A(n26892), .B(n26893), .Z(n26852) );
  AND U26702 ( .A(n1458), .B(n26894), .Z(n26892) );
  XOR U26703 ( .A(n26895), .B(n26893), .Z(n26894) );
  NANDN U26704 ( .A(n26854), .B(n26856), .Z(n26870) );
  XOR U26705 ( .A(n26896), .B(n26897), .Z(n26856) );
  AND U26706 ( .A(n1458), .B(n26898), .Z(n26896) );
  XOR U26707 ( .A(n26897), .B(n26899), .Z(n26898) );
  XOR U26708 ( .A(n26900), .B(n26901), .Z(n1458) );
  AND U26709 ( .A(n26902), .B(n26903), .Z(n26900) );
  XNOR U26710 ( .A(n26901), .B(n26867), .Z(n26903) );
  XNOR U26711 ( .A(n26904), .B(n26905), .Z(n26867) );
  ANDN U26712 ( .B(n26906), .A(n26907), .Z(n26904) );
  XOR U26713 ( .A(n26905), .B(n26908), .Z(n26906) );
  XOR U26714 ( .A(n26901), .B(n26869), .Z(n26902) );
  XOR U26715 ( .A(n26909), .B(n26910), .Z(n26869) );
  AND U26716 ( .A(n1462), .B(n26911), .Z(n26909) );
  XOR U26717 ( .A(n26912), .B(n26910), .Z(n26911) );
  XNOR U26718 ( .A(n26913), .B(n26914), .Z(n26901) );
  NAND U26719 ( .A(n26915), .B(n26916), .Z(n26914) );
  XOR U26720 ( .A(n26917), .B(n26893), .Z(n26916) );
  XOR U26721 ( .A(n26907), .B(n26908), .Z(n26893) );
  XOR U26722 ( .A(n26918), .B(n26919), .Z(n26908) );
  ANDN U26723 ( .B(n26920), .A(n26921), .Z(n26918) );
  XOR U26724 ( .A(n26919), .B(n26922), .Z(n26920) );
  XOR U26725 ( .A(n26923), .B(n26924), .Z(n26907) );
  XOR U26726 ( .A(n26925), .B(n26926), .Z(n26924) );
  ANDN U26727 ( .B(n26927), .A(n26928), .Z(n26925) );
  XOR U26728 ( .A(n26929), .B(n26926), .Z(n26927) );
  IV U26729 ( .A(n26905), .Z(n26923) );
  XOR U26730 ( .A(n26930), .B(n26931), .Z(n26905) );
  ANDN U26731 ( .B(n26932), .A(n26933), .Z(n26930) );
  XOR U26732 ( .A(n26931), .B(n26934), .Z(n26932) );
  IV U26733 ( .A(n26913), .Z(n26917) );
  XOR U26734 ( .A(n26913), .B(n26895), .Z(n26915) );
  XOR U26735 ( .A(n26935), .B(n26936), .Z(n26895) );
  AND U26736 ( .A(n1462), .B(n26937), .Z(n26935) );
  XOR U26737 ( .A(n26938), .B(n26936), .Z(n26937) );
  NANDN U26738 ( .A(n26897), .B(n26899), .Z(n26913) );
  XOR U26739 ( .A(n26939), .B(n26940), .Z(n26899) );
  AND U26740 ( .A(n1462), .B(n26941), .Z(n26939) );
  XOR U26741 ( .A(n26940), .B(n26942), .Z(n26941) );
  XOR U26742 ( .A(n26943), .B(n26944), .Z(n1462) );
  AND U26743 ( .A(n26945), .B(n26946), .Z(n26943) );
  XNOR U26744 ( .A(n26944), .B(n26910), .Z(n26946) );
  XNOR U26745 ( .A(n26947), .B(n26948), .Z(n26910) );
  ANDN U26746 ( .B(n26949), .A(n26950), .Z(n26947) );
  XOR U26747 ( .A(n26948), .B(n26951), .Z(n26949) );
  XOR U26748 ( .A(n26944), .B(n26912), .Z(n26945) );
  XOR U26749 ( .A(n26952), .B(n26953), .Z(n26912) );
  AND U26750 ( .A(n1466), .B(n26954), .Z(n26952) );
  XOR U26751 ( .A(n26955), .B(n26953), .Z(n26954) );
  XNOR U26752 ( .A(n26956), .B(n26957), .Z(n26944) );
  NAND U26753 ( .A(n26958), .B(n26959), .Z(n26957) );
  XOR U26754 ( .A(n26960), .B(n26936), .Z(n26959) );
  XOR U26755 ( .A(n26950), .B(n26951), .Z(n26936) );
  XOR U26756 ( .A(n26961), .B(n26962), .Z(n26951) );
  ANDN U26757 ( .B(n26963), .A(n26964), .Z(n26961) );
  XOR U26758 ( .A(n26962), .B(n26965), .Z(n26963) );
  XOR U26759 ( .A(n26966), .B(n26967), .Z(n26950) );
  XOR U26760 ( .A(n26968), .B(n26969), .Z(n26967) );
  ANDN U26761 ( .B(n26970), .A(n26971), .Z(n26968) );
  XOR U26762 ( .A(n26972), .B(n26969), .Z(n26970) );
  IV U26763 ( .A(n26948), .Z(n26966) );
  XOR U26764 ( .A(n26973), .B(n26974), .Z(n26948) );
  ANDN U26765 ( .B(n26975), .A(n26976), .Z(n26973) );
  XOR U26766 ( .A(n26974), .B(n26977), .Z(n26975) );
  IV U26767 ( .A(n26956), .Z(n26960) );
  XOR U26768 ( .A(n26956), .B(n26938), .Z(n26958) );
  XOR U26769 ( .A(n26978), .B(n26979), .Z(n26938) );
  AND U26770 ( .A(n1466), .B(n26980), .Z(n26978) );
  XOR U26771 ( .A(n26981), .B(n26979), .Z(n26980) );
  NANDN U26772 ( .A(n26940), .B(n26942), .Z(n26956) );
  XOR U26773 ( .A(n26982), .B(n26983), .Z(n26942) );
  AND U26774 ( .A(n1466), .B(n26984), .Z(n26982) );
  XOR U26775 ( .A(n26983), .B(n26985), .Z(n26984) );
  XOR U26776 ( .A(n26986), .B(n26987), .Z(n1466) );
  AND U26777 ( .A(n26988), .B(n26989), .Z(n26986) );
  XNOR U26778 ( .A(n26987), .B(n26953), .Z(n26989) );
  XNOR U26779 ( .A(n26990), .B(n26991), .Z(n26953) );
  ANDN U26780 ( .B(n26992), .A(n26993), .Z(n26990) );
  XOR U26781 ( .A(n26991), .B(n26994), .Z(n26992) );
  XOR U26782 ( .A(n26987), .B(n26955), .Z(n26988) );
  XOR U26783 ( .A(n26995), .B(n26996), .Z(n26955) );
  AND U26784 ( .A(n1470), .B(n26997), .Z(n26995) );
  XOR U26785 ( .A(n26998), .B(n26996), .Z(n26997) );
  XNOR U26786 ( .A(n26999), .B(n27000), .Z(n26987) );
  NAND U26787 ( .A(n27001), .B(n27002), .Z(n27000) );
  XOR U26788 ( .A(n27003), .B(n26979), .Z(n27002) );
  XOR U26789 ( .A(n26993), .B(n26994), .Z(n26979) );
  XOR U26790 ( .A(n27004), .B(n27005), .Z(n26994) );
  ANDN U26791 ( .B(n27006), .A(n27007), .Z(n27004) );
  XOR U26792 ( .A(n27005), .B(n27008), .Z(n27006) );
  XOR U26793 ( .A(n27009), .B(n27010), .Z(n26993) );
  XOR U26794 ( .A(n27011), .B(n27012), .Z(n27010) );
  ANDN U26795 ( .B(n27013), .A(n27014), .Z(n27011) );
  XOR U26796 ( .A(n27015), .B(n27012), .Z(n27013) );
  IV U26797 ( .A(n26991), .Z(n27009) );
  XOR U26798 ( .A(n27016), .B(n27017), .Z(n26991) );
  ANDN U26799 ( .B(n27018), .A(n27019), .Z(n27016) );
  XOR U26800 ( .A(n27017), .B(n27020), .Z(n27018) );
  IV U26801 ( .A(n26999), .Z(n27003) );
  XOR U26802 ( .A(n26999), .B(n26981), .Z(n27001) );
  XOR U26803 ( .A(n27021), .B(n27022), .Z(n26981) );
  AND U26804 ( .A(n1470), .B(n27023), .Z(n27021) );
  XOR U26805 ( .A(n27024), .B(n27022), .Z(n27023) );
  NANDN U26806 ( .A(n26983), .B(n26985), .Z(n26999) );
  XOR U26807 ( .A(n27025), .B(n27026), .Z(n26985) );
  AND U26808 ( .A(n1470), .B(n27027), .Z(n27025) );
  XOR U26809 ( .A(n27026), .B(n27028), .Z(n27027) );
  XOR U26810 ( .A(n27029), .B(n27030), .Z(n1470) );
  AND U26811 ( .A(n27031), .B(n27032), .Z(n27029) );
  XNOR U26812 ( .A(n27030), .B(n26996), .Z(n27032) );
  XNOR U26813 ( .A(n27033), .B(n27034), .Z(n26996) );
  ANDN U26814 ( .B(n27035), .A(n27036), .Z(n27033) );
  XOR U26815 ( .A(n27034), .B(n27037), .Z(n27035) );
  XOR U26816 ( .A(n27030), .B(n26998), .Z(n27031) );
  XOR U26817 ( .A(n27038), .B(n27039), .Z(n26998) );
  AND U26818 ( .A(n1474), .B(n27040), .Z(n27038) );
  XOR U26819 ( .A(n27041), .B(n27039), .Z(n27040) );
  XNOR U26820 ( .A(n27042), .B(n27043), .Z(n27030) );
  NAND U26821 ( .A(n27044), .B(n27045), .Z(n27043) );
  XOR U26822 ( .A(n27046), .B(n27022), .Z(n27045) );
  XOR U26823 ( .A(n27036), .B(n27037), .Z(n27022) );
  XOR U26824 ( .A(n27047), .B(n27048), .Z(n27037) );
  ANDN U26825 ( .B(n27049), .A(n27050), .Z(n27047) );
  XOR U26826 ( .A(n27048), .B(n27051), .Z(n27049) );
  XOR U26827 ( .A(n27052), .B(n27053), .Z(n27036) );
  XOR U26828 ( .A(n27054), .B(n27055), .Z(n27053) );
  ANDN U26829 ( .B(n27056), .A(n27057), .Z(n27054) );
  XOR U26830 ( .A(n27058), .B(n27055), .Z(n27056) );
  IV U26831 ( .A(n27034), .Z(n27052) );
  XOR U26832 ( .A(n27059), .B(n27060), .Z(n27034) );
  ANDN U26833 ( .B(n27061), .A(n27062), .Z(n27059) );
  XOR U26834 ( .A(n27060), .B(n27063), .Z(n27061) );
  IV U26835 ( .A(n27042), .Z(n27046) );
  XOR U26836 ( .A(n27042), .B(n27024), .Z(n27044) );
  XOR U26837 ( .A(n27064), .B(n27065), .Z(n27024) );
  AND U26838 ( .A(n1474), .B(n27066), .Z(n27064) );
  XOR U26839 ( .A(n27067), .B(n27065), .Z(n27066) );
  NANDN U26840 ( .A(n27026), .B(n27028), .Z(n27042) );
  XOR U26841 ( .A(n27068), .B(n27069), .Z(n27028) );
  AND U26842 ( .A(n1474), .B(n27070), .Z(n27068) );
  XOR U26843 ( .A(n27069), .B(n27071), .Z(n27070) );
  XOR U26844 ( .A(n27072), .B(n27073), .Z(n1474) );
  AND U26845 ( .A(n27074), .B(n27075), .Z(n27072) );
  XNOR U26846 ( .A(n27073), .B(n27039), .Z(n27075) );
  XNOR U26847 ( .A(n27076), .B(n27077), .Z(n27039) );
  ANDN U26848 ( .B(n27078), .A(n27079), .Z(n27076) );
  XOR U26849 ( .A(n27077), .B(n27080), .Z(n27078) );
  XOR U26850 ( .A(n27073), .B(n27041), .Z(n27074) );
  XOR U26851 ( .A(n27081), .B(n27082), .Z(n27041) );
  AND U26852 ( .A(n1478), .B(n27083), .Z(n27081) );
  XOR U26853 ( .A(n27084), .B(n27082), .Z(n27083) );
  XNOR U26854 ( .A(n27085), .B(n27086), .Z(n27073) );
  NAND U26855 ( .A(n27087), .B(n27088), .Z(n27086) );
  XOR U26856 ( .A(n27089), .B(n27065), .Z(n27088) );
  XOR U26857 ( .A(n27079), .B(n27080), .Z(n27065) );
  XOR U26858 ( .A(n27090), .B(n27091), .Z(n27080) );
  ANDN U26859 ( .B(n27092), .A(n27093), .Z(n27090) );
  XOR U26860 ( .A(n27091), .B(n27094), .Z(n27092) );
  XOR U26861 ( .A(n27095), .B(n27096), .Z(n27079) );
  XOR U26862 ( .A(n27097), .B(n27098), .Z(n27096) );
  ANDN U26863 ( .B(n27099), .A(n27100), .Z(n27097) );
  XOR U26864 ( .A(n27101), .B(n27098), .Z(n27099) );
  IV U26865 ( .A(n27077), .Z(n27095) );
  XOR U26866 ( .A(n27102), .B(n27103), .Z(n27077) );
  ANDN U26867 ( .B(n27104), .A(n27105), .Z(n27102) );
  XOR U26868 ( .A(n27103), .B(n27106), .Z(n27104) );
  IV U26869 ( .A(n27085), .Z(n27089) );
  XOR U26870 ( .A(n27085), .B(n27067), .Z(n27087) );
  XOR U26871 ( .A(n27107), .B(n27108), .Z(n27067) );
  AND U26872 ( .A(n1478), .B(n27109), .Z(n27107) );
  XOR U26873 ( .A(n27110), .B(n27108), .Z(n27109) );
  NANDN U26874 ( .A(n27069), .B(n27071), .Z(n27085) );
  XOR U26875 ( .A(n27111), .B(n27112), .Z(n27071) );
  AND U26876 ( .A(n1478), .B(n27113), .Z(n27111) );
  XOR U26877 ( .A(n27112), .B(n27114), .Z(n27113) );
  XOR U26878 ( .A(n27115), .B(n27116), .Z(n1478) );
  AND U26879 ( .A(n27117), .B(n27118), .Z(n27115) );
  XNOR U26880 ( .A(n27116), .B(n27082), .Z(n27118) );
  XNOR U26881 ( .A(n27119), .B(n27120), .Z(n27082) );
  ANDN U26882 ( .B(n27121), .A(n27122), .Z(n27119) );
  XOR U26883 ( .A(n27120), .B(n27123), .Z(n27121) );
  XOR U26884 ( .A(n27116), .B(n27084), .Z(n27117) );
  XOR U26885 ( .A(n27124), .B(n27125), .Z(n27084) );
  AND U26886 ( .A(n1482), .B(n27126), .Z(n27124) );
  XOR U26887 ( .A(n27127), .B(n27125), .Z(n27126) );
  XNOR U26888 ( .A(n27128), .B(n27129), .Z(n27116) );
  NAND U26889 ( .A(n27130), .B(n27131), .Z(n27129) );
  XOR U26890 ( .A(n27132), .B(n27108), .Z(n27131) );
  XOR U26891 ( .A(n27122), .B(n27123), .Z(n27108) );
  XOR U26892 ( .A(n27133), .B(n27134), .Z(n27123) );
  ANDN U26893 ( .B(n27135), .A(n27136), .Z(n27133) );
  XOR U26894 ( .A(n27134), .B(n27137), .Z(n27135) );
  XOR U26895 ( .A(n27138), .B(n27139), .Z(n27122) );
  XOR U26896 ( .A(n27140), .B(n27141), .Z(n27139) );
  ANDN U26897 ( .B(n27142), .A(n27143), .Z(n27140) );
  XOR U26898 ( .A(n27144), .B(n27141), .Z(n27142) );
  IV U26899 ( .A(n27120), .Z(n27138) );
  XOR U26900 ( .A(n27145), .B(n27146), .Z(n27120) );
  ANDN U26901 ( .B(n27147), .A(n27148), .Z(n27145) );
  XOR U26902 ( .A(n27146), .B(n27149), .Z(n27147) );
  IV U26903 ( .A(n27128), .Z(n27132) );
  XOR U26904 ( .A(n27128), .B(n27110), .Z(n27130) );
  XOR U26905 ( .A(n27150), .B(n27151), .Z(n27110) );
  AND U26906 ( .A(n1482), .B(n27152), .Z(n27150) );
  XOR U26907 ( .A(n27153), .B(n27151), .Z(n27152) );
  NANDN U26908 ( .A(n27112), .B(n27114), .Z(n27128) );
  XOR U26909 ( .A(n27154), .B(n27155), .Z(n27114) );
  AND U26910 ( .A(n1482), .B(n27156), .Z(n27154) );
  XOR U26911 ( .A(n27155), .B(n27157), .Z(n27156) );
  XOR U26912 ( .A(n27158), .B(n27159), .Z(n1482) );
  AND U26913 ( .A(n27160), .B(n27161), .Z(n27158) );
  XNOR U26914 ( .A(n27159), .B(n27125), .Z(n27161) );
  XNOR U26915 ( .A(n27162), .B(n27163), .Z(n27125) );
  ANDN U26916 ( .B(n27164), .A(n27165), .Z(n27162) );
  XOR U26917 ( .A(n27163), .B(n27166), .Z(n27164) );
  XOR U26918 ( .A(n27159), .B(n27127), .Z(n27160) );
  XOR U26919 ( .A(n27167), .B(n27168), .Z(n27127) );
  AND U26920 ( .A(n1486), .B(n27169), .Z(n27167) );
  XOR U26921 ( .A(n27170), .B(n27168), .Z(n27169) );
  XNOR U26922 ( .A(n27171), .B(n27172), .Z(n27159) );
  NAND U26923 ( .A(n27173), .B(n27174), .Z(n27172) );
  XOR U26924 ( .A(n27175), .B(n27151), .Z(n27174) );
  XOR U26925 ( .A(n27165), .B(n27166), .Z(n27151) );
  XOR U26926 ( .A(n27176), .B(n27177), .Z(n27166) );
  ANDN U26927 ( .B(n27178), .A(n27179), .Z(n27176) );
  XOR U26928 ( .A(n27177), .B(n27180), .Z(n27178) );
  XOR U26929 ( .A(n27181), .B(n27182), .Z(n27165) );
  XOR U26930 ( .A(n27183), .B(n27184), .Z(n27182) );
  ANDN U26931 ( .B(n27185), .A(n27186), .Z(n27183) );
  XOR U26932 ( .A(n27187), .B(n27184), .Z(n27185) );
  IV U26933 ( .A(n27163), .Z(n27181) );
  XOR U26934 ( .A(n27188), .B(n27189), .Z(n27163) );
  ANDN U26935 ( .B(n27190), .A(n27191), .Z(n27188) );
  XOR U26936 ( .A(n27189), .B(n27192), .Z(n27190) );
  IV U26937 ( .A(n27171), .Z(n27175) );
  XOR U26938 ( .A(n27171), .B(n27153), .Z(n27173) );
  XOR U26939 ( .A(n27193), .B(n27194), .Z(n27153) );
  AND U26940 ( .A(n1486), .B(n27195), .Z(n27193) );
  XOR U26941 ( .A(n27196), .B(n27194), .Z(n27195) );
  NANDN U26942 ( .A(n27155), .B(n27157), .Z(n27171) );
  XOR U26943 ( .A(n27197), .B(n27198), .Z(n27157) );
  AND U26944 ( .A(n1486), .B(n27199), .Z(n27197) );
  XOR U26945 ( .A(n27198), .B(n27200), .Z(n27199) );
  XOR U26946 ( .A(n27201), .B(n27202), .Z(n1486) );
  AND U26947 ( .A(n27203), .B(n27204), .Z(n27201) );
  XNOR U26948 ( .A(n27202), .B(n27168), .Z(n27204) );
  XNOR U26949 ( .A(n27205), .B(n27206), .Z(n27168) );
  ANDN U26950 ( .B(n27207), .A(n27208), .Z(n27205) );
  XOR U26951 ( .A(n27206), .B(n27209), .Z(n27207) );
  XOR U26952 ( .A(n27202), .B(n27170), .Z(n27203) );
  XOR U26953 ( .A(n27210), .B(n27211), .Z(n27170) );
  AND U26954 ( .A(n1490), .B(n27212), .Z(n27210) );
  XOR U26955 ( .A(n27213), .B(n27211), .Z(n27212) );
  XNOR U26956 ( .A(n27214), .B(n27215), .Z(n27202) );
  NAND U26957 ( .A(n27216), .B(n27217), .Z(n27215) );
  XOR U26958 ( .A(n27218), .B(n27194), .Z(n27217) );
  XOR U26959 ( .A(n27208), .B(n27209), .Z(n27194) );
  XOR U26960 ( .A(n27219), .B(n27220), .Z(n27209) );
  ANDN U26961 ( .B(n27221), .A(n27222), .Z(n27219) );
  XOR U26962 ( .A(n27220), .B(n27223), .Z(n27221) );
  XOR U26963 ( .A(n27224), .B(n27225), .Z(n27208) );
  XOR U26964 ( .A(n27226), .B(n27227), .Z(n27225) );
  ANDN U26965 ( .B(n27228), .A(n27229), .Z(n27226) );
  XOR U26966 ( .A(n27230), .B(n27227), .Z(n27228) );
  IV U26967 ( .A(n27206), .Z(n27224) );
  XOR U26968 ( .A(n27231), .B(n27232), .Z(n27206) );
  ANDN U26969 ( .B(n27233), .A(n27234), .Z(n27231) );
  XOR U26970 ( .A(n27232), .B(n27235), .Z(n27233) );
  IV U26971 ( .A(n27214), .Z(n27218) );
  XOR U26972 ( .A(n27214), .B(n27196), .Z(n27216) );
  XOR U26973 ( .A(n27236), .B(n27237), .Z(n27196) );
  AND U26974 ( .A(n1490), .B(n27238), .Z(n27236) );
  XOR U26975 ( .A(n27239), .B(n27237), .Z(n27238) );
  NANDN U26976 ( .A(n27198), .B(n27200), .Z(n27214) );
  XOR U26977 ( .A(n27240), .B(n27241), .Z(n27200) );
  AND U26978 ( .A(n1490), .B(n27242), .Z(n27240) );
  XOR U26979 ( .A(n27241), .B(n27243), .Z(n27242) );
  XOR U26980 ( .A(n27244), .B(n27245), .Z(n1490) );
  AND U26981 ( .A(n27246), .B(n27247), .Z(n27244) );
  XNOR U26982 ( .A(n27245), .B(n27211), .Z(n27247) );
  XNOR U26983 ( .A(n27248), .B(n27249), .Z(n27211) );
  ANDN U26984 ( .B(n27250), .A(n27251), .Z(n27248) );
  XOR U26985 ( .A(n27249), .B(n27252), .Z(n27250) );
  XOR U26986 ( .A(n27245), .B(n27213), .Z(n27246) );
  XOR U26987 ( .A(n27253), .B(n27254), .Z(n27213) );
  AND U26988 ( .A(n1494), .B(n27255), .Z(n27253) );
  XOR U26989 ( .A(n27256), .B(n27254), .Z(n27255) );
  XNOR U26990 ( .A(n27257), .B(n27258), .Z(n27245) );
  NAND U26991 ( .A(n27259), .B(n27260), .Z(n27258) );
  XOR U26992 ( .A(n27261), .B(n27237), .Z(n27260) );
  XOR U26993 ( .A(n27251), .B(n27252), .Z(n27237) );
  XOR U26994 ( .A(n27262), .B(n27263), .Z(n27252) );
  ANDN U26995 ( .B(n27264), .A(n27265), .Z(n27262) );
  XOR U26996 ( .A(n27263), .B(n27266), .Z(n27264) );
  XOR U26997 ( .A(n27267), .B(n27268), .Z(n27251) );
  XOR U26998 ( .A(n27269), .B(n27270), .Z(n27268) );
  ANDN U26999 ( .B(n27271), .A(n27272), .Z(n27269) );
  XOR U27000 ( .A(n27273), .B(n27270), .Z(n27271) );
  IV U27001 ( .A(n27249), .Z(n27267) );
  XOR U27002 ( .A(n27274), .B(n27275), .Z(n27249) );
  ANDN U27003 ( .B(n27276), .A(n27277), .Z(n27274) );
  XOR U27004 ( .A(n27275), .B(n27278), .Z(n27276) );
  IV U27005 ( .A(n27257), .Z(n27261) );
  XOR U27006 ( .A(n27257), .B(n27239), .Z(n27259) );
  XOR U27007 ( .A(n27279), .B(n27280), .Z(n27239) );
  AND U27008 ( .A(n1494), .B(n27281), .Z(n27279) );
  XOR U27009 ( .A(n27282), .B(n27280), .Z(n27281) );
  NANDN U27010 ( .A(n27241), .B(n27243), .Z(n27257) );
  XOR U27011 ( .A(n27283), .B(n27284), .Z(n27243) );
  AND U27012 ( .A(n1494), .B(n27285), .Z(n27283) );
  XOR U27013 ( .A(n27284), .B(n27286), .Z(n27285) );
  XOR U27014 ( .A(n27287), .B(n27288), .Z(n1494) );
  AND U27015 ( .A(n27289), .B(n27290), .Z(n27287) );
  XNOR U27016 ( .A(n27288), .B(n27254), .Z(n27290) );
  XNOR U27017 ( .A(n27291), .B(n27292), .Z(n27254) );
  ANDN U27018 ( .B(n27293), .A(n27294), .Z(n27291) );
  XOR U27019 ( .A(n27292), .B(n27295), .Z(n27293) );
  XOR U27020 ( .A(n27288), .B(n27256), .Z(n27289) );
  XOR U27021 ( .A(n27296), .B(n27297), .Z(n27256) );
  AND U27022 ( .A(n1498), .B(n27298), .Z(n27296) );
  XOR U27023 ( .A(n27299), .B(n27297), .Z(n27298) );
  XNOR U27024 ( .A(n27300), .B(n27301), .Z(n27288) );
  NAND U27025 ( .A(n27302), .B(n27303), .Z(n27301) );
  XOR U27026 ( .A(n27304), .B(n27280), .Z(n27303) );
  XOR U27027 ( .A(n27294), .B(n27295), .Z(n27280) );
  XOR U27028 ( .A(n27305), .B(n27306), .Z(n27295) );
  ANDN U27029 ( .B(n27307), .A(n27308), .Z(n27305) );
  XOR U27030 ( .A(n27306), .B(n27309), .Z(n27307) );
  XOR U27031 ( .A(n27310), .B(n27311), .Z(n27294) );
  XOR U27032 ( .A(n27312), .B(n27313), .Z(n27311) );
  ANDN U27033 ( .B(n27314), .A(n27315), .Z(n27312) );
  XOR U27034 ( .A(n27316), .B(n27313), .Z(n27314) );
  IV U27035 ( .A(n27292), .Z(n27310) );
  XOR U27036 ( .A(n27317), .B(n27318), .Z(n27292) );
  ANDN U27037 ( .B(n27319), .A(n27320), .Z(n27317) );
  XOR U27038 ( .A(n27318), .B(n27321), .Z(n27319) );
  IV U27039 ( .A(n27300), .Z(n27304) );
  XOR U27040 ( .A(n27300), .B(n27282), .Z(n27302) );
  XOR U27041 ( .A(n27322), .B(n27323), .Z(n27282) );
  AND U27042 ( .A(n1498), .B(n27324), .Z(n27322) );
  XOR U27043 ( .A(n27325), .B(n27323), .Z(n27324) );
  NANDN U27044 ( .A(n27284), .B(n27286), .Z(n27300) );
  XOR U27045 ( .A(n27326), .B(n27327), .Z(n27286) );
  AND U27046 ( .A(n1498), .B(n27328), .Z(n27326) );
  XOR U27047 ( .A(n27327), .B(n27329), .Z(n27328) );
  XOR U27048 ( .A(n27330), .B(n27331), .Z(n1498) );
  AND U27049 ( .A(n27332), .B(n27333), .Z(n27330) );
  XNOR U27050 ( .A(n27331), .B(n27297), .Z(n27333) );
  XNOR U27051 ( .A(n27334), .B(n27335), .Z(n27297) );
  ANDN U27052 ( .B(n27336), .A(n27337), .Z(n27334) );
  XOR U27053 ( .A(n27335), .B(n27338), .Z(n27336) );
  XOR U27054 ( .A(n27331), .B(n27299), .Z(n27332) );
  XOR U27055 ( .A(n27339), .B(n27340), .Z(n27299) );
  AND U27056 ( .A(n1502), .B(n27341), .Z(n27339) );
  XOR U27057 ( .A(n27342), .B(n27340), .Z(n27341) );
  XNOR U27058 ( .A(n27343), .B(n27344), .Z(n27331) );
  NAND U27059 ( .A(n27345), .B(n27346), .Z(n27344) );
  XOR U27060 ( .A(n27347), .B(n27323), .Z(n27346) );
  XOR U27061 ( .A(n27337), .B(n27338), .Z(n27323) );
  XOR U27062 ( .A(n27348), .B(n27349), .Z(n27338) );
  ANDN U27063 ( .B(n27350), .A(n27351), .Z(n27348) );
  XOR U27064 ( .A(n27349), .B(n27352), .Z(n27350) );
  XOR U27065 ( .A(n27353), .B(n27354), .Z(n27337) );
  XOR U27066 ( .A(n27355), .B(n27356), .Z(n27354) );
  ANDN U27067 ( .B(n27357), .A(n27358), .Z(n27355) );
  XOR U27068 ( .A(n27359), .B(n27356), .Z(n27357) );
  IV U27069 ( .A(n27335), .Z(n27353) );
  XOR U27070 ( .A(n27360), .B(n27361), .Z(n27335) );
  ANDN U27071 ( .B(n27362), .A(n27363), .Z(n27360) );
  XOR U27072 ( .A(n27361), .B(n27364), .Z(n27362) );
  IV U27073 ( .A(n27343), .Z(n27347) );
  XOR U27074 ( .A(n27343), .B(n27325), .Z(n27345) );
  XOR U27075 ( .A(n27365), .B(n27366), .Z(n27325) );
  AND U27076 ( .A(n1502), .B(n27367), .Z(n27365) );
  XOR U27077 ( .A(n27368), .B(n27366), .Z(n27367) );
  NANDN U27078 ( .A(n27327), .B(n27329), .Z(n27343) );
  XOR U27079 ( .A(n27369), .B(n27370), .Z(n27329) );
  AND U27080 ( .A(n1502), .B(n27371), .Z(n27369) );
  XOR U27081 ( .A(n27370), .B(n27372), .Z(n27371) );
  XOR U27082 ( .A(n27373), .B(n27374), .Z(n1502) );
  AND U27083 ( .A(n27375), .B(n27376), .Z(n27373) );
  XNOR U27084 ( .A(n27374), .B(n27340), .Z(n27376) );
  XNOR U27085 ( .A(n27377), .B(n27378), .Z(n27340) );
  ANDN U27086 ( .B(n27379), .A(n27380), .Z(n27377) );
  XOR U27087 ( .A(n27378), .B(n27381), .Z(n27379) );
  XOR U27088 ( .A(n27374), .B(n27342), .Z(n27375) );
  XOR U27089 ( .A(n27382), .B(n27383), .Z(n27342) );
  AND U27090 ( .A(n1506), .B(n27384), .Z(n27382) );
  XOR U27091 ( .A(n27385), .B(n27383), .Z(n27384) );
  XNOR U27092 ( .A(n27386), .B(n27387), .Z(n27374) );
  NAND U27093 ( .A(n27388), .B(n27389), .Z(n27387) );
  XOR U27094 ( .A(n27390), .B(n27366), .Z(n27389) );
  XOR U27095 ( .A(n27380), .B(n27381), .Z(n27366) );
  XOR U27096 ( .A(n27391), .B(n27392), .Z(n27381) );
  ANDN U27097 ( .B(n27393), .A(n27394), .Z(n27391) );
  XOR U27098 ( .A(n27392), .B(n27395), .Z(n27393) );
  XOR U27099 ( .A(n27396), .B(n27397), .Z(n27380) );
  XOR U27100 ( .A(n27398), .B(n27399), .Z(n27397) );
  ANDN U27101 ( .B(n27400), .A(n27401), .Z(n27398) );
  XOR U27102 ( .A(n27402), .B(n27399), .Z(n27400) );
  IV U27103 ( .A(n27378), .Z(n27396) );
  XOR U27104 ( .A(n27403), .B(n27404), .Z(n27378) );
  ANDN U27105 ( .B(n27405), .A(n27406), .Z(n27403) );
  XOR U27106 ( .A(n27404), .B(n27407), .Z(n27405) );
  IV U27107 ( .A(n27386), .Z(n27390) );
  XOR U27108 ( .A(n27386), .B(n27368), .Z(n27388) );
  XOR U27109 ( .A(n27408), .B(n27409), .Z(n27368) );
  AND U27110 ( .A(n1506), .B(n27410), .Z(n27408) );
  XOR U27111 ( .A(n27411), .B(n27409), .Z(n27410) );
  NANDN U27112 ( .A(n27370), .B(n27372), .Z(n27386) );
  XOR U27113 ( .A(n27412), .B(n27413), .Z(n27372) );
  AND U27114 ( .A(n1506), .B(n27414), .Z(n27412) );
  XOR U27115 ( .A(n27413), .B(n27415), .Z(n27414) );
  XOR U27116 ( .A(n27416), .B(n27417), .Z(n1506) );
  AND U27117 ( .A(n27418), .B(n27419), .Z(n27416) );
  XNOR U27118 ( .A(n27417), .B(n27383), .Z(n27419) );
  XNOR U27119 ( .A(n27420), .B(n27421), .Z(n27383) );
  ANDN U27120 ( .B(n27422), .A(n27423), .Z(n27420) );
  XOR U27121 ( .A(n27421), .B(n27424), .Z(n27422) );
  XOR U27122 ( .A(n27417), .B(n27385), .Z(n27418) );
  XOR U27123 ( .A(n27425), .B(n27426), .Z(n27385) );
  AND U27124 ( .A(n1510), .B(n27427), .Z(n27425) );
  XOR U27125 ( .A(n27428), .B(n27426), .Z(n27427) );
  XNOR U27126 ( .A(n27429), .B(n27430), .Z(n27417) );
  NAND U27127 ( .A(n27431), .B(n27432), .Z(n27430) );
  XOR U27128 ( .A(n27433), .B(n27409), .Z(n27432) );
  XOR U27129 ( .A(n27423), .B(n27424), .Z(n27409) );
  XOR U27130 ( .A(n27434), .B(n27435), .Z(n27424) );
  ANDN U27131 ( .B(n27436), .A(n27437), .Z(n27434) );
  XOR U27132 ( .A(n27435), .B(n27438), .Z(n27436) );
  XOR U27133 ( .A(n27439), .B(n27440), .Z(n27423) );
  XOR U27134 ( .A(n27441), .B(n27442), .Z(n27440) );
  ANDN U27135 ( .B(n27443), .A(n27444), .Z(n27441) );
  XOR U27136 ( .A(n27445), .B(n27442), .Z(n27443) );
  IV U27137 ( .A(n27421), .Z(n27439) );
  XOR U27138 ( .A(n27446), .B(n27447), .Z(n27421) );
  ANDN U27139 ( .B(n27448), .A(n27449), .Z(n27446) );
  XOR U27140 ( .A(n27447), .B(n27450), .Z(n27448) );
  IV U27141 ( .A(n27429), .Z(n27433) );
  XOR U27142 ( .A(n27429), .B(n27411), .Z(n27431) );
  XOR U27143 ( .A(n27451), .B(n27452), .Z(n27411) );
  AND U27144 ( .A(n1510), .B(n27453), .Z(n27451) );
  XOR U27145 ( .A(n27454), .B(n27452), .Z(n27453) );
  NANDN U27146 ( .A(n27413), .B(n27415), .Z(n27429) );
  XOR U27147 ( .A(n27455), .B(n27456), .Z(n27415) );
  AND U27148 ( .A(n1510), .B(n27457), .Z(n27455) );
  XOR U27149 ( .A(n27456), .B(n27458), .Z(n27457) );
  XOR U27150 ( .A(n27459), .B(n27460), .Z(n1510) );
  AND U27151 ( .A(n27461), .B(n27462), .Z(n27459) );
  XNOR U27152 ( .A(n27460), .B(n27426), .Z(n27462) );
  XNOR U27153 ( .A(n27463), .B(n27464), .Z(n27426) );
  ANDN U27154 ( .B(n27465), .A(n27466), .Z(n27463) );
  XOR U27155 ( .A(n27464), .B(n27467), .Z(n27465) );
  XOR U27156 ( .A(n27460), .B(n27428), .Z(n27461) );
  XOR U27157 ( .A(n27468), .B(n27469), .Z(n27428) );
  AND U27158 ( .A(n1514), .B(n27470), .Z(n27468) );
  XOR U27159 ( .A(n27471), .B(n27469), .Z(n27470) );
  XNOR U27160 ( .A(n27472), .B(n27473), .Z(n27460) );
  NAND U27161 ( .A(n27474), .B(n27475), .Z(n27473) );
  XOR U27162 ( .A(n27476), .B(n27452), .Z(n27475) );
  XOR U27163 ( .A(n27466), .B(n27467), .Z(n27452) );
  XOR U27164 ( .A(n27477), .B(n27478), .Z(n27467) );
  ANDN U27165 ( .B(n27479), .A(n27480), .Z(n27477) );
  XOR U27166 ( .A(n27478), .B(n27481), .Z(n27479) );
  XOR U27167 ( .A(n27482), .B(n27483), .Z(n27466) );
  XOR U27168 ( .A(n27484), .B(n27485), .Z(n27483) );
  ANDN U27169 ( .B(n27486), .A(n27487), .Z(n27484) );
  XOR U27170 ( .A(n27488), .B(n27485), .Z(n27486) );
  IV U27171 ( .A(n27464), .Z(n27482) );
  XOR U27172 ( .A(n27489), .B(n27490), .Z(n27464) );
  ANDN U27173 ( .B(n27491), .A(n27492), .Z(n27489) );
  XOR U27174 ( .A(n27490), .B(n27493), .Z(n27491) );
  IV U27175 ( .A(n27472), .Z(n27476) );
  XOR U27176 ( .A(n27472), .B(n27454), .Z(n27474) );
  XOR U27177 ( .A(n27494), .B(n27495), .Z(n27454) );
  AND U27178 ( .A(n1514), .B(n27496), .Z(n27494) );
  XOR U27179 ( .A(n27497), .B(n27495), .Z(n27496) );
  NANDN U27180 ( .A(n27456), .B(n27458), .Z(n27472) );
  XOR U27181 ( .A(n27498), .B(n27499), .Z(n27458) );
  AND U27182 ( .A(n1514), .B(n27500), .Z(n27498) );
  XOR U27183 ( .A(n27499), .B(n27501), .Z(n27500) );
  XOR U27184 ( .A(n27502), .B(n27503), .Z(n1514) );
  AND U27185 ( .A(n27504), .B(n27505), .Z(n27502) );
  XNOR U27186 ( .A(n27503), .B(n27469), .Z(n27505) );
  XNOR U27187 ( .A(n27506), .B(n27507), .Z(n27469) );
  ANDN U27188 ( .B(n27508), .A(n27509), .Z(n27506) );
  XOR U27189 ( .A(n27507), .B(n27510), .Z(n27508) );
  XOR U27190 ( .A(n27503), .B(n27471), .Z(n27504) );
  XOR U27191 ( .A(n27511), .B(n27512), .Z(n27471) );
  AND U27192 ( .A(n1518), .B(n27513), .Z(n27511) );
  XOR U27193 ( .A(n27514), .B(n27512), .Z(n27513) );
  XNOR U27194 ( .A(n27515), .B(n27516), .Z(n27503) );
  NAND U27195 ( .A(n27517), .B(n27518), .Z(n27516) );
  XOR U27196 ( .A(n27519), .B(n27495), .Z(n27518) );
  XOR U27197 ( .A(n27509), .B(n27510), .Z(n27495) );
  XOR U27198 ( .A(n27520), .B(n27521), .Z(n27510) );
  ANDN U27199 ( .B(n27522), .A(n27523), .Z(n27520) );
  XOR U27200 ( .A(n27521), .B(n27524), .Z(n27522) );
  XOR U27201 ( .A(n27525), .B(n27526), .Z(n27509) );
  XOR U27202 ( .A(n27527), .B(n27528), .Z(n27526) );
  ANDN U27203 ( .B(n27529), .A(n27530), .Z(n27527) );
  XOR U27204 ( .A(n27531), .B(n27528), .Z(n27529) );
  IV U27205 ( .A(n27507), .Z(n27525) );
  XOR U27206 ( .A(n27532), .B(n27533), .Z(n27507) );
  ANDN U27207 ( .B(n27534), .A(n27535), .Z(n27532) );
  XOR U27208 ( .A(n27533), .B(n27536), .Z(n27534) );
  IV U27209 ( .A(n27515), .Z(n27519) );
  XOR U27210 ( .A(n27515), .B(n27497), .Z(n27517) );
  XOR U27211 ( .A(n27537), .B(n27538), .Z(n27497) );
  AND U27212 ( .A(n1518), .B(n27539), .Z(n27537) );
  XOR U27213 ( .A(n27540), .B(n27538), .Z(n27539) );
  NANDN U27214 ( .A(n27499), .B(n27501), .Z(n27515) );
  XOR U27215 ( .A(n27541), .B(n27542), .Z(n27501) );
  AND U27216 ( .A(n1518), .B(n27543), .Z(n27541) );
  XOR U27217 ( .A(n27542), .B(n27544), .Z(n27543) );
  XOR U27218 ( .A(n27545), .B(n27546), .Z(n1518) );
  AND U27219 ( .A(n27547), .B(n27548), .Z(n27545) );
  XNOR U27220 ( .A(n27546), .B(n27512), .Z(n27548) );
  XNOR U27221 ( .A(n27549), .B(n27550), .Z(n27512) );
  ANDN U27222 ( .B(n27551), .A(n27552), .Z(n27549) );
  XOR U27223 ( .A(n27550), .B(n27553), .Z(n27551) );
  XOR U27224 ( .A(n27546), .B(n27514), .Z(n27547) );
  XOR U27225 ( .A(n27554), .B(n27555), .Z(n27514) );
  AND U27226 ( .A(n1522), .B(n27556), .Z(n27554) );
  XOR U27227 ( .A(n27557), .B(n27555), .Z(n27556) );
  XNOR U27228 ( .A(n27558), .B(n27559), .Z(n27546) );
  NAND U27229 ( .A(n27560), .B(n27561), .Z(n27559) );
  XOR U27230 ( .A(n27562), .B(n27538), .Z(n27561) );
  XOR U27231 ( .A(n27552), .B(n27553), .Z(n27538) );
  XOR U27232 ( .A(n27563), .B(n27564), .Z(n27553) );
  ANDN U27233 ( .B(n27565), .A(n27566), .Z(n27563) );
  XOR U27234 ( .A(n27564), .B(n27567), .Z(n27565) );
  XOR U27235 ( .A(n27568), .B(n27569), .Z(n27552) );
  XOR U27236 ( .A(n27570), .B(n27571), .Z(n27569) );
  ANDN U27237 ( .B(n27572), .A(n27573), .Z(n27570) );
  XOR U27238 ( .A(n27574), .B(n27571), .Z(n27572) );
  IV U27239 ( .A(n27550), .Z(n27568) );
  XOR U27240 ( .A(n27575), .B(n27576), .Z(n27550) );
  ANDN U27241 ( .B(n27577), .A(n27578), .Z(n27575) );
  XOR U27242 ( .A(n27576), .B(n27579), .Z(n27577) );
  IV U27243 ( .A(n27558), .Z(n27562) );
  XOR U27244 ( .A(n27558), .B(n27540), .Z(n27560) );
  XOR U27245 ( .A(n27580), .B(n27581), .Z(n27540) );
  AND U27246 ( .A(n1522), .B(n27582), .Z(n27580) );
  XOR U27247 ( .A(n27583), .B(n27581), .Z(n27582) );
  NANDN U27248 ( .A(n27542), .B(n27544), .Z(n27558) );
  XOR U27249 ( .A(n27584), .B(n27585), .Z(n27544) );
  AND U27250 ( .A(n1522), .B(n27586), .Z(n27584) );
  XOR U27251 ( .A(n27585), .B(n27587), .Z(n27586) );
  XOR U27252 ( .A(n27588), .B(n27589), .Z(n1522) );
  AND U27253 ( .A(n27590), .B(n27591), .Z(n27588) );
  XNOR U27254 ( .A(n27589), .B(n27555), .Z(n27591) );
  XNOR U27255 ( .A(n27592), .B(n27593), .Z(n27555) );
  ANDN U27256 ( .B(n27594), .A(n27595), .Z(n27592) );
  XOR U27257 ( .A(n27593), .B(n27596), .Z(n27594) );
  XOR U27258 ( .A(n27589), .B(n27557), .Z(n27590) );
  XOR U27259 ( .A(n27597), .B(n27598), .Z(n27557) );
  AND U27260 ( .A(n1526), .B(n27599), .Z(n27597) );
  XOR U27261 ( .A(n27600), .B(n27598), .Z(n27599) );
  XNOR U27262 ( .A(n27601), .B(n27602), .Z(n27589) );
  NAND U27263 ( .A(n27603), .B(n27604), .Z(n27602) );
  XOR U27264 ( .A(n27605), .B(n27581), .Z(n27604) );
  XOR U27265 ( .A(n27595), .B(n27596), .Z(n27581) );
  XOR U27266 ( .A(n27606), .B(n27607), .Z(n27596) );
  ANDN U27267 ( .B(n27608), .A(n27609), .Z(n27606) );
  XOR U27268 ( .A(n27607), .B(n27610), .Z(n27608) );
  XOR U27269 ( .A(n27611), .B(n27612), .Z(n27595) );
  XOR U27270 ( .A(n27613), .B(n27614), .Z(n27612) );
  ANDN U27271 ( .B(n27615), .A(n27616), .Z(n27613) );
  XOR U27272 ( .A(n27617), .B(n27614), .Z(n27615) );
  IV U27273 ( .A(n27593), .Z(n27611) );
  XOR U27274 ( .A(n27618), .B(n27619), .Z(n27593) );
  ANDN U27275 ( .B(n27620), .A(n27621), .Z(n27618) );
  XOR U27276 ( .A(n27619), .B(n27622), .Z(n27620) );
  IV U27277 ( .A(n27601), .Z(n27605) );
  XOR U27278 ( .A(n27601), .B(n27583), .Z(n27603) );
  XOR U27279 ( .A(n27623), .B(n27624), .Z(n27583) );
  AND U27280 ( .A(n1526), .B(n27625), .Z(n27623) );
  XOR U27281 ( .A(n27626), .B(n27624), .Z(n27625) );
  NANDN U27282 ( .A(n27585), .B(n27587), .Z(n27601) );
  XOR U27283 ( .A(n27627), .B(n27628), .Z(n27587) );
  AND U27284 ( .A(n1526), .B(n27629), .Z(n27627) );
  XOR U27285 ( .A(n27628), .B(n27630), .Z(n27629) );
  XOR U27286 ( .A(n27631), .B(n27632), .Z(n1526) );
  AND U27287 ( .A(n27633), .B(n27634), .Z(n27631) );
  XNOR U27288 ( .A(n27632), .B(n27598), .Z(n27634) );
  XNOR U27289 ( .A(n27635), .B(n27636), .Z(n27598) );
  ANDN U27290 ( .B(n27637), .A(n27638), .Z(n27635) );
  XOR U27291 ( .A(n27636), .B(n27639), .Z(n27637) );
  XOR U27292 ( .A(n27632), .B(n27600), .Z(n27633) );
  XOR U27293 ( .A(n27640), .B(n27641), .Z(n27600) );
  AND U27294 ( .A(n1530), .B(n27642), .Z(n27640) );
  XOR U27295 ( .A(n27643), .B(n27641), .Z(n27642) );
  XNOR U27296 ( .A(n27644), .B(n27645), .Z(n27632) );
  NAND U27297 ( .A(n27646), .B(n27647), .Z(n27645) );
  XOR U27298 ( .A(n27648), .B(n27624), .Z(n27647) );
  XOR U27299 ( .A(n27638), .B(n27639), .Z(n27624) );
  XOR U27300 ( .A(n27649), .B(n27650), .Z(n27639) );
  ANDN U27301 ( .B(n27651), .A(n27652), .Z(n27649) );
  XOR U27302 ( .A(n27650), .B(n27653), .Z(n27651) );
  XOR U27303 ( .A(n27654), .B(n27655), .Z(n27638) );
  XOR U27304 ( .A(n27656), .B(n27657), .Z(n27655) );
  ANDN U27305 ( .B(n27658), .A(n27659), .Z(n27656) );
  XOR U27306 ( .A(n27660), .B(n27657), .Z(n27658) );
  IV U27307 ( .A(n27636), .Z(n27654) );
  XOR U27308 ( .A(n27661), .B(n27662), .Z(n27636) );
  ANDN U27309 ( .B(n27663), .A(n27664), .Z(n27661) );
  XOR U27310 ( .A(n27662), .B(n27665), .Z(n27663) );
  IV U27311 ( .A(n27644), .Z(n27648) );
  XOR U27312 ( .A(n27644), .B(n27626), .Z(n27646) );
  XOR U27313 ( .A(n27666), .B(n27667), .Z(n27626) );
  AND U27314 ( .A(n1530), .B(n27668), .Z(n27666) );
  XOR U27315 ( .A(n27669), .B(n27667), .Z(n27668) );
  NANDN U27316 ( .A(n27628), .B(n27630), .Z(n27644) );
  XOR U27317 ( .A(n27670), .B(n27671), .Z(n27630) );
  AND U27318 ( .A(n1530), .B(n27672), .Z(n27670) );
  XOR U27319 ( .A(n27671), .B(n27673), .Z(n27672) );
  XOR U27320 ( .A(n27674), .B(n27675), .Z(n1530) );
  AND U27321 ( .A(n27676), .B(n27677), .Z(n27674) );
  XNOR U27322 ( .A(n27675), .B(n27641), .Z(n27677) );
  XNOR U27323 ( .A(n27678), .B(n27679), .Z(n27641) );
  ANDN U27324 ( .B(n27680), .A(n27681), .Z(n27678) );
  XOR U27325 ( .A(n27679), .B(n27682), .Z(n27680) );
  XOR U27326 ( .A(n27675), .B(n27643), .Z(n27676) );
  XOR U27327 ( .A(n27683), .B(n27684), .Z(n27643) );
  AND U27328 ( .A(n1534), .B(n27685), .Z(n27683) );
  XOR U27329 ( .A(n27686), .B(n27684), .Z(n27685) );
  XNOR U27330 ( .A(n27687), .B(n27688), .Z(n27675) );
  NAND U27331 ( .A(n27689), .B(n27690), .Z(n27688) );
  XOR U27332 ( .A(n27691), .B(n27667), .Z(n27690) );
  XOR U27333 ( .A(n27681), .B(n27682), .Z(n27667) );
  XOR U27334 ( .A(n27692), .B(n27693), .Z(n27682) );
  ANDN U27335 ( .B(n27694), .A(n27695), .Z(n27692) );
  XOR U27336 ( .A(n27693), .B(n27696), .Z(n27694) );
  XOR U27337 ( .A(n27697), .B(n27698), .Z(n27681) );
  XOR U27338 ( .A(n27699), .B(n27700), .Z(n27698) );
  ANDN U27339 ( .B(n27701), .A(n27702), .Z(n27699) );
  XOR U27340 ( .A(n27703), .B(n27700), .Z(n27701) );
  IV U27341 ( .A(n27679), .Z(n27697) );
  XOR U27342 ( .A(n27704), .B(n27705), .Z(n27679) );
  ANDN U27343 ( .B(n27706), .A(n27707), .Z(n27704) );
  XOR U27344 ( .A(n27705), .B(n27708), .Z(n27706) );
  IV U27345 ( .A(n27687), .Z(n27691) );
  XOR U27346 ( .A(n27687), .B(n27669), .Z(n27689) );
  XOR U27347 ( .A(n27709), .B(n27710), .Z(n27669) );
  AND U27348 ( .A(n1534), .B(n27711), .Z(n27709) );
  XOR U27349 ( .A(n27712), .B(n27710), .Z(n27711) );
  NANDN U27350 ( .A(n27671), .B(n27673), .Z(n27687) );
  XOR U27351 ( .A(n27713), .B(n27714), .Z(n27673) );
  AND U27352 ( .A(n1534), .B(n27715), .Z(n27713) );
  XOR U27353 ( .A(n27714), .B(n27716), .Z(n27715) );
  XOR U27354 ( .A(n27717), .B(n27718), .Z(n1534) );
  AND U27355 ( .A(n27719), .B(n27720), .Z(n27717) );
  XNOR U27356 ( .A(n27718), .B(n27684), .Z(n27720) );
  XNOR U27357 ( .A(n27721), .B(n27722), .Z(n27684) );
  ANDN U27358 ( .B(n27723), .A(n27724), .Z(n27721) );
  XOR U27359 ( .A(n27722), .B(n27725), .Z(n27723) );
  XOR U27360 ( .A(n27718), .B(n27686), .Z(n27719) );
  XOR U27361 ( .A(n27726), .B(n27727), .Z(n27686) );
  AND U27362 ( .A(n1538), .B(n27728), .Z(n27726) );
  XOR U27363 ( .A(n27729), .B(n27727), .Z(n27728) );
  XNOR U27364 ( .A(n27730), .B(n27731), .Z(n27718) );
  NAND U27365 ( .A(n27732), .B(n27733), .Z(n27731) );
  XOR U27366 ( .A(n27734), .B(n27710), .Z(n27733) );
  XOR U27367 ( .A(n27724), .B(n27725), .Z(n27710) );
  XOR U27368 ( .A(n27735), .B(n27736), .Z(n27725) );
  ANDN U27369 ( .B(n27737), .A(n27738), .Z(n27735) );
  XOR U27370 ( .A(n27736), .B(n27739), .Z(n27737) );
  XOR U27371 ( .A(n27740), .B(n27741), .Z(n27724) );
  XOR U27372 ( .A(n27742), .B(n27743), .Z(n27741) );
  ANDN U27373 ( .B(n27744), .A(n27745), .Z(n27742) );
  XOR U27374 ( .A(n27746), .B(n27743), .Z(n27744) );
  IV U27375 ( .A(n27722), .Z(n27740) );
  XOR U27376 ( .A(n27747), .B(n27748), .Z(n27722) );
  ANDN U27377 ( .B(n27749), .A(n27750), .Z(n27747) );
  XOR U27378 ( .A(n27748), .B(n27751), .Z(n27749) );
  IV U27379 ( .A(n27730), .Z(n27734) );
  XOR U27380 ( .A(n27730), .B(n27712), .Z(n27732) );
  XOR U27381 ( .A(n27752), .B(n27753), .Z(n27712) );
  AND U27382 ( .A(n1538), .B(n27754), .Z(n27752) );
  XOR U27383 ( .A(n27755), .B(n27753), .Z(n27754) );
  NANDN U27384 ( .A(n27714), .B(n27716), .Z(n27730) );
  XOR U27385 ( .A(n27756), .B(n27757), .Z(n27716) );
  AND U27386 ( .A(n1538), .B(n27758), .Z(n27756) );
  XOR U27387 ( .A(n27757), .B(n27759), .Z(n27758) );
  XOR U27388 ( .A(n27760), .B(n27761), .Z(n1538) );
  AND U27389 ( .A(n27762), .B(n27763), .Z(n27760) );
  XNOR U27390 ( .A(n27761), .B(n27727), .Z(n27763) );
  XNOR U27391 ( .A(n27764), .B(n27765), .Z(n27727) );
  ANDN U27392 ( .B(n27766), .A(n27767), .Z(n27764) );
  XOR U27393 ( .A(n27765), .B(n27768), .Z(n27766) );
  XOR U27394 ( .A(n27761), .B(n27729), .Z(n27762) );
  XOR U27395 ( .A(n27769), .B(n27770), .Z(n27729) );
  AND U27396 ( .A(n1542), .B(n27771), .Z(n27769) );
  XOR U27397 ( .A(n27772), .B(n27770), .Z(n27771) );
  XNOR U27398 ( .A(n27773), .B(n27774), .Z(n27761) );
  NAND U27399 ( .A(n27775), .B(n27776), .Z(n27774) );
  XOR U27400 ( .A(n27777), .B(n27753), .Z(n27776) );
  XOR U27401 ( .A(n27767), .B(n27768), .Z(n27753) );
  XOR U27402 ( .A(n27778), .B(n27779), .Z(n27768) );
  ANDN U27403 ( .B(n27780), .A(n27781), .Z(n27778) );
  XOR U27404 ( .A(n27779), .B(n27782), .Z(n27780) );
  XOR U27405 ( .A(n27783), .B(n27784), .Z(n27767) );
  XOR U27406 ( .A(n27785), .B(n27786), .Z(n27784) );
  ANDN U27407 ( .B(n27787), .A(n27788), .Z(n27785) );
  XOR U27408 ( .A(n27789), .B(n27786), .Z(n27787) );
  IV U27409 ( .A(n27765), .Z(n27783) );
  XOR U27410 ( .A(n27790), .B(n27791), .Z(n27765) );
  ANDN U27411 ( .B(n27792), .A(n27793), .Z(n27790) );
  XOR U27412 ( .A(n27791), .B(n27794), .Z(n27792) );
  IV U27413 ( .A(n27773), .Z(n27777) );
  XOR U27414 ( .A(n27773), .B(n27755), .Z(n27775) );
  XOR U27415 ( .A(n27795), .B(n27796), .Z(n27755) );
  AND U27416 ( .A(n1542), .B(n27797), .Z(n27795) );
  XOR U27417 ( .A(n27798), .B(n27796), .Z(n27797) );
  NANDN U27418 ( .A(n27757), .B(n27759), .Z(n27773) );
  XOR U27419 ( .A(n27799), .B(n27800), .Z(n27759) );
  AND U27420 ( .A(n1542), .B(n27801), .Z(n27799) );
  XOR U27421 ( .A(n27800), .B(n27802), .Z(n27801) );
  XOR U27422 ( .A(n27803), .B(n27804), .Z(n1542) );
  AND U27423 ( .A(n27805), .B(n27806), .Z(n27803) );
  XNOR U27424 ( .A(n27804), .B(n27770), .Z(n27806) );
  XNOR U27425 ( .A(n27807), .B(n27808), .Z(n27770) );
  ANDN U27426 ( .B(n27809), .A(n27810), .Z(n27807) );
  XOR U27427 ( .A(n27808), .B(n27811), .Z(n27809) );
  XOR U27428 ( .A(n27804), .B(n27772), .Z(n27805) );
  XOR U27429 ( .A(n27812), .B(n27813), .Z(n27772) );
  AND U27430 ( .A(n1546), .B(n27814), .Z(n27812) );
  XOR U27431 ( .A(n27815), .B(n27813), .Z(n27814) );
  XNOR U27432 ( .A(n27816), .B(n27817), .Z(n27804) );
  NAND U27433 ( .A(n27818), .B(n27819), .Z(n27817) );
  XOR U27434 ( .A(n27820), .B(n27796), .Z(n27819) );
  XOR U27435 ( .A(n27810), .B(n27811), .Z(n27796) );
  XOR U27436 ( .A(n27821), .B(n27822), .Z(n27811) );
  ANDN U27437 ( .B(n27823), .A(n27824), .Z(n27821) );
  XOR U27438 ( .A(n27822), .B(n27825), .Z(n27823) );
  XOR U27439 ( .A(n27826), .B(n27827), .Z(n27810) );
  XOR U27440 ( .A(n27828), .B(n27829), .Z(n27827) );
  ANDN U27441 ( .B(n27830), .A(n27831), .Z(n27828) );
  XOR U27442 ( .A(n27832), .B(n27829), .Z(n27830) );
  IV U27443 ( .A(n27808), .Z(n27826) );
  XOR U27444 ( .A(n27833), .B(n27834), .Z(n27808) );
  ANDN U27445 ( .B(n27835), .A(n27836), .Z(n27833) );
  XOR U27446 ( .A(n27834), .B(n27837), .Z(n27835) );
  IV U27447 ( .A(n27816), .Z(n27820) );
  XOR U27448 ( .A(n27816), .B(n27798), .Z(n27818) );
  XOR U27449 ( .A(n27838), .B(n27839), .Z(n27798) );
  AND U27450 ( .A(n1546), .B(n27840), .Z(n27838) );
  XOR U27451 ( .A(n27841), .B(n27839), .Z(n27840) );
  NANDN U27452 ( .A(n27800), .B(n27802), .Z(n27816) );
  XOR U27453 ( .A(n27842), .B(n27843), .Z(n27802) );
  AND U27454 ( .A(n1546), .B(n27844), .Z(n27842) );
  XOR U27455 ( .A(n27843), .B(n27845), .Z(n27844) );
  XOR U27456 ( .A(n27846), .B(n27847), .Z(n1546) );
  AND U27457 ( .A(n27848), .B(n27849), .Z(n27846) );
  XNOR U27458 ( .A(n27847), .B(n27813), .Z(n27849) );
  XNOR U27459 ( .A(n27850), .B(n27851), .Z(n27813) );
  ANDN U27460 ( .B(n27852), .A(n27853), .Z(n27850) );
  XOR U27461 ( .A(n27851), .B(n27854), .Z(n27852) );
  XOR U27462 ( .A(n27847), .B(n27815), .Z(n27848) );
  XOR U27463 ( .A(n27855), .B(n27856), .Z(n27815) );
  AND U27464 ( .A(n1550), .B(n27857), .Z(n27855) );
  XOR U27465 ( .A(n27858), .B(n27856), .Z(n27857) );
  XNOR U27466 ( .A(n27859), .B(n27860), .Z(n27847) );
  NAND U27467 ( .A(n27861), .B(n27862), .Z(n27860) );
  XOR U27468 ( .A(n27863), .B(n27839), .Z(n27862) );
  XOR U27469 ( .A(n27853), .B(n27854), .Z(n27839) );
  XOR U27470 ( .A(n27864), .B(n27865), .Z(n27854) );
  ANDN U27471 ( .B(n27866), .A(n27867), .Z(n27864) );
  XOR U27472 ( .A(n27865), .B(n27868), .Z(n27866) );
  XOR U27473 ( .A(n27869), .B(n27870), .Z(n27853) );
  XOR U27474 ( .A(n27871), .B(n27872), .Z(n27870) );
  ANDN U27475 ( .B(n27873), .A(n27874), .Z(n27871) );
  XOR U27476 ( .A(n27875), .B(n27872), .Z(n27873) );
  IV U27477 ( .A(n27851), .Z(n27869) );
  XOR U27478 ( .A(n27876), .B(n27877), .Z(n27851) );
  ANDN U27479 ( .B(n27878), .A(n27879), .Z(n27876) );
  XOR U27480 ( .A(n27877), .B(n27880), .Z(n27878) );
  IV U27481 ( .A(n27859), .Z(n27863) );
  XOR U27482 ( .A(n27859), .B(n27841), .Z(n27861) );
  XOR U27483 ( .A(n27881), .B(n27882), .Z(n27841) );
  AND U27484 ( .A(n1550), .B(n27883), .Z(n27881) );
  XOR U27485 ( .A(n27884), .B(n27882), .Z(n27883) );
  NANDN U27486 ( .A(n27843), .B(n27845), .Z(n27859) );
  XOR U27487 ( .A(n27885), .B(n27886), .Z(n27845) );
  AND U27488 ( .A(n1550), .B(n27887), .Z(n27885) );
  XOR U27489 ( .A(n27886), .B(n27888), .Z(n27887) );
  XOR U27490 ( .A(n27889), .B(n27890), .Z(n1550) );
  AND U27491 ( .A(n27891), .B(n27892), .Z(n27889) );
  XNOR U27492 ( .A(n27890), .B(n27856), .Z(n27892) );
  XNOR U27493 ( .A(n27893), .B(n27894), .Z(n27856) );
  ANDN U27494 ( .B(n27895), .A(n27896), .Z(n27893) );
  XOR U27495 ( .A(n27894), .B(n27897), .Z(n27895) );
  XOR U27496 ( .A(n27890), .B(n27858), .Z(n27891) );
  XOR U27497 ( .A(n27898), .B(n27899), .Z(n27858) );
  AND U27498 ( .A(n1554), .B(n27900), .Z(n27898) );
  XOR U27499 ( .A(n27901), .B(n27899), .Z(n27900) );
  XNOR U27500 ( .A(n27902), .B(n27903), .Z(n27890) );
  NAND U27501 ( .A(n27904), .B(n27905), .Z(n27903) );
  XOR U27502 ( .A(n27906), .B(n27882), .Z(n27905) );
  XOR U27503 ( .A(n27896), .B(n27897), .Z(n27882) );
  XOR U27504 ( .A(n27907), .B(n27908), .Z(n27897) );
  ANDN U27505 ( .B(n27909), .A(n27910), .Z(n27907) );
  XOR U27506 ( .A(n27908), .B(n27911), .Z(n27909) );
  XOR U27507 ( .A(n27912), .B(n27913), .Z(n27896) );
  XOR U27508 ( .A(n27914), .B(n27915), .Z(n27913) );
  ANDN U27509 ( .B(n27916), .A(n27917), .Z(n27914) );
  XOR U27510 ( .A(n27918), .B(n27915), .Z(n27916) );
  IV U27511 ( .A(n27894), .Z(n27912) );
  XOR U27512 ( .A(n27919), .B(n27920), .Z(n27894) );
  ANDN U27513 ( .B(n27921), .A(n27922), .Z(n27919) );
  XOR U27514 ( .A(n27920), .B(n27923), .Z(n27921) );
  IV U27515 ( .A(n27902), .Z(n27906) );
  XOR U27516 ( .A(n27902), .B(n27884), .Z(n27904) );
  XOR U27517 ( .A(n27924), .B(n27925), .Z(n27884) );
  AND U27518 ( .A(n1554), .B(n27926), .Z(n27924) );
  XOR U27519 ( .A(n27927), .B(n27925), .Z(n27926) );
  NANDN U27520 ( .A(n27886), .B(n27888), .Z(n27902) );
  XOR U27521 ( .A(n27928), .B(n27929), .Z(n27888) );
  AND U27522 ( .A(n1554), .B(n27930), .Z(n27928) );
  XOR U27523 ( .A(n27929), .B(n27931), .Z(n27930) );
  XOR U27524 ( .A(n27932), .B(n27933), .Z(n1554) );
  AND U27525 ( .A(n27934), .B(n27935), .Z(n27932) );
  XNOR U27526 ( .A(n27933), .B(n27899), .Z(n27935) );
  XNOR U27527 ( .A(n27936), .B(n27937), .Z(n27899) );
  ANDN U27528 ( .B(n27938), .A(n27939), .Z(n27936) );
  XOR U27529 ( .A(n27937), .B(n27940), .Z(n27938) );
  XOR U27530 ( .A(n27933), .B(n27901), .Z(n27934) );
  XOR U27531 ( .A(n27941), .B(n27942), .Z(n27901) );
  AND U27532 ( .A(n1558), .B(n27943), .Z(n27941) );
  XOR U27533 ( .A(n27944), .B(n27942), .Z(n27943) );
  XNOR U27534 ( .A(n27945), .B(n27946), .Z(n27933) );
  NAND U27535 ( .A(n27947), .B(n27948), .Z(n27946) );
  XOR U27536 ( .A(n27949), .B(n27925), .Z(n27948) );
  XOR U27537 ( .A(n27939), .B(n27940), .Z(n27925) );
  XOR U27538 ( .A(n27950), .B(n27951), .Z(n27940) );
  ANDN U27539 ( .B(n27952), .A(n27953), .Z(n27950) );
  XOR U27540 ( .A(n27951), .B(n27954), .Z(n27952) );
  XOR U27541 ( .A(n27955), .B(n27956), .Z(n27939) );
  XOR U27542 ( .A(n27957), .B(n27958), .Z(n27956) );
  ANDN U27543 ( .B(n27959), .A(n27960), .Z(n27957) );
  XOR U27544 ( .A(n27961), .B(n27958), .Z(n27959) );
  IV U27545 ( .A(n27937), .Z(n27955) );
  XOR U27546 ( .A(n27962), .B(n27963), .Z(n27937) );
  ANDN U27547 ( .B(n27964), .A(n27965), .Z(n27962) );
  XOR U27548 ( .A(n27963), .B(n27966), .Z(n27964) );
  IV U27549 ( .A(n27945), .Z(n27949) );
  XOR U27550 ( .A(n27945), .B(n27927), .Z(n27947) );
  XOR U27551 ( .A(n27967), .B(n27968), .Z(n27927) );
  AND U27552 ( .A(n1558), .B(n27969), .Z(n27967) );
  XOR U27553 ( .A(n27970), .B(n27968), .Z(n27969) );
  NANDN U27554 ( .A(n27929), .B(n27931), .Z(n27945) );
  XOR U27555 ( .A(n27971), .B(n27972), .Z(n27931) );
  AND U27556 ( .A(n1558), .B(n27973), .Z(n27971) );
  XOR U27557 ( .A(n27972), .B(n27974), .Z(n27973) );
  XOR U27558 ( .A(n27975), .B(n27976), .Z(n1558) );
  AND U27559 ( .A(n27977), .B(n27978), .Z(n27975) );
  XNOR U27560 ( .A(n27976), .B(n27942), .Z(n27978) );
  XNOR U27561 ( .A(n27979), .B(n27980), .Z(n27942) );
  ANDN U27562 ( .B(n27981), .A(n27982), .Z(n27979) );
  XOR U27563 ( .A(n27980), .B(n27983), .Z(n27981) );
  XOR U27564 ( .A(n27976), .B(n27944), .Z(n27977) );
  XOR U27565 ( .A(n27984), .B(n27985), .Z(n27944) );
  AND U27566 ( .A(n1562), .B(n27986), .Z(n27984) );
  XOR U27567 ( .A(n27987), .B(n27985), .Z(n27986) );
  XNOR U27568 ( .A(n27988), .B(n27989), .Z(n27976) );
  NAND U27569 ( .A(n27990), .B(n27991), .Z(n27989) );
  XOR U27570 ( .A(n27992), .B(n27968), .Z(n27991) );
  XOR U27571 ( .A(n27982), .B(n27983), .Z(n27968) );
  XOR U27572 ( .A(n27993), .B(n27994), .Z(n27983) );
  ANDN U27573 ( .B(n27995), .A(n27996), .Z(n27993) );
  XOR U27574 ( .A(n27994), .B(n27997), .Z(n27995) );
  XOR U27575 ( .A(n27998), .B(n27999), .Z(n27982) );
  XOR U27576 ( .A(n28000), .B(n28001), .Z(n27999) );
  ANDN U27577 ( .B(n28002), .A(n28003), .Z(n28000) );
  XOR U27578 ( .A(n28004), .B(n28001), .Z(n28002) );
  IV U27579 ( .A(n27980), .Z(n27998) );
  XOR U27580 ( .A(n28005), .B(n28006), .Z(n27980) );
  ANDN U27581 ( .B(n28007), .A(n28008), .Z(n28005) );
  XOR U27582 ( .A(n28006), .B(n28009), .Z(n28007) );
  IV U27583 ( .A(n27988), .Z(n27992) );
  XOR U27584 ( .A(n27988), .B(n27970), .Z(n27990) );
  XOR U27585 ( .A(n28010), .B(n28011), .Z(n27970) );
  AND U27586 ( .A(n1562), .B(n28012), .Z(n28010) );
  XOR U27587 ( .A(n28013), .B(n28011), .Z(n28012) );
  NANDN U27588 ( .A(n27972), .B(n27974), .Z(n27988) );
  XOR U27589 ( .A(n28014), .B(n28015), .Z(n27974) );
  AND U27590 ( .A(n1562), .B(n28016), .Z(n28014) );
  XOR U27591 ( .A(n28015), .B(n28017), .Z(n28016) );
  XOR U27592 ( .A(n28018), .B(n28019), .Z(n1562) );
  AND U27593 ( .A(n28020), .B(n28021), .Z(n28018) );
  XNOR U27594 ( .A(n28019), .B(n27985), .Z(n28021) );
  XNOR U27595 ( .A(n28022), .B(n28023), .Z(n27985) );
  ANDN U27596 ( .B(n28024), .A(n28025), .Z(n28022) );
  XOR U27597 ( .A(n28023), .B(n28026), .Z(n28024) );
  XOR U27598 ( .A(n28019), .B(n27987), .Z(n28020) );
  XOR U27599 ( .A(n28027), .B(n28028), .Z(n27987) );
  AND U27600 ( .A(n1566), .B(n28029), .Z(n28027) );
  XOR U27601 ( .A(n28030), .B(n28028), .Z(n28029) );
  XNOR U27602 ( .A(n28031), .B(n28032), .Z(n28019) );
  NAND U27603 ( .A(n28033), .B(n28034), .Z(n28032) );
  XOR U27604 ( .A(n28035), .B(n28011), .Z(n28034) );
  XOR U27605 ( .A(n28025), .B(n28026), .Z(n28011) );
  XOR U27606 ( .A(n28036), .B(n28037), .Z(n28026) );
  ANDN U27607 ( .B(n28038), .A(n28039), .Z(n28036) );
  XOR U27608 ( .A(n28037), .B(n28040), .Z(n28038) );
  XOR U27609 ( .A(n28041), .B(n28042), .Z(n28025) );
  XOR U27610 ( .A(n28043), .B(n28044), .Z(n28042) );
  ANDN U27611 ( .B(n28045), .A(n28046), .Z(n28043) );
  XOR U27612 ( .A(n28047), .B(n28044), .Z(n28045) );
  IV U27613 ( .A(n28023), .Z(n28041) );
  XOR U27614 ( .A(n28048), .B(n28049), .Z(n28023) );
  ANDN U27615 ( .B(n28050), .A(n28051), .Z(n28048) );
  XOR U27616 ( .A(n28049), .B(n28052), .Z(n28050) );
  IV U27617 ( .A(n28031), .Z(n28035) );
  XOR U27618 ( .A(n28031), .B(n28013), .Z(n28033) );
  XOR U27619 ( .A(n28053), .B(n28054), .Z(n28013) );
  AND U27620 ( .A(n1566), .B(n28055), .Z(n28053) );
  XOR U27621 ( .A(n28056), .B(n28054), .Z(n28055) );
  NANDN U27622 ( .A(n28015), .B(n28017), .Z(n28031) );
  XOR U27623 ( .A(n28057), .B(n28058), .Z(n28017) );
  AND U27624 ( .A(n1566), .B(n28059), .Z(n28057) );
  XOR U27625 ( .A(n28058), .B(n28060), .Z(n28059) );
  XOR U27626 ( .A(n28061), .B(n28062), .Z(n1566) );
  AND U27627 ( .A(n28063), .B(n28064), .Z(n28061) );
  XNOR U27628 ( .A(n28062), .B(n28028), .Z(n28064) );
  XNOR U27629 ( .A(n28065), .B(n28066), .Z(n28028) );
  ANDN U27630 ( .B(n28067), .A(n28068), .Z(n28065) );
  XOR U27631 ( .A(n28066), .B(n28069), .Z(n28067) );
  XOR U27632 ( .A(n28062), .B(n28030), .Z(n28063) );
  XOR U27633 ( .A(n28070), .B(n28071), .Z(n28030) );
  AND U27634 ( .A(n1570), .B(n28072), .Z(n28070) );
  XOR U27635 ( .A(n28073), .B(n28071), .Z(n28072) );
  XNOR U27636 ( .A(n28074), .B(n28075), .Z(n28062) );
  NAND U27637 ( .A(n28076), .B(n28077), .Z(n28075) );
  XOR U27638 ( .A(n28078), .B(n28054), .Z(n28077) );
  XOR U27639 ( .A(n28068), .B(n28069), .Z(n28054) );
  XOR U27640 ( .A(n28079), .B(n28080), .Z(n28069) );
  ANDN U27641 ( .B(n28081), .A(n28082), .Z(n28079) );
  XOR U27642 ( .A(n28080), .B(n28083), .Z(n28081) );
  XOR U27643 ( .A(n28084), .B(n28085), .Z(n28068) );
  XOR U27644 ( .A(n28086), .B(n28087), .Z(n28085) );
  ANDN U27645 ( .B(n28088), .A(n28089), .Z(n28086) );
  XOR U27646 ( .A(n28090), .B(n28087), .Z(n28088) );
  IV U27647 ( .A(n28066), .Z(n28084) );
  XOR U27648 ( .A(n28091), .B(n28092), .Z(n28066) );
  ANDN U27649 ( .B(n28093), .A(n28094), .Z(n28091) );
  XOR U27650 ( .A(n28092), .B(n28095), .Z(n28093) );
  IV U27651 ( .A(n28074), .Z(n28078) );
  XOR U27652 ( .A(n28074), .B(n28056), .Z(n28076) );
  XOR U27653 ( .A(n28096), .B(n28097), .Z(n28056) );
  AND U27654 ( .A(n1570), .B(n28098), .Z(n28096) );
  XOR U27655 ( .A(n28099), .B(n28097), .Z(n28098) );
  NANDN U27656 ( .A(n28058), .B(n28060), .Z(n28074) );
  XOR U27657 ( .A(n28100), .B(n28101), .Z(n28060) );
  AND U27658 ( .A(n1570), .B(n28102), .Z(n28100) );
  XOR U27659 ( .A(n28101), .B(n28103), .Z(n28102) );
  XOR U27660 ( .A(n28104), .B(n28105), .Z(n1570) );
  AND U27661 ( .A(n28106), .B(n28107), .Z(n28104) );
  XNOR U27662 ( .A(n28105), .B(n28071), .Z(n28107) );
  XNOR U27663 ( .A(n28108), .B(n28109), .Z(n28071) );
  ANDN U27664 ( .B(n28110), .A(n28111), .Z(n28108) );
  XOR U27665 ( .A(n28109), .B(n28112), .Z(n28110) );
  XOR U27666 ( .A(n28105), .B(n28073), .Z(n28106) );
  XOR U27667 ( .A(n28113), .B(n28114), .Z(n28073) );
  AND U27668 ( .A(n1574), .B(n28115), .Z(n28113) );
  XOR U27669 ( .A(n28116), .B(n28114), .Z(n28115) );
  XNOR U27670 ( .A(n28117), .B(n28118), .Z(n28105) );
  NAND U27671 ( .A(n28119), .B(n28120), .Z(n28118) );
  XOR U27672 ( .A(n28121), .B(n28097), .Z(n28120) );
  XOR U27673 ( .A(n28111), .B(n28112), .Z(n28097) );
  XOR U27674 ( .A(n28122), .B(n28123), .Z(n28112) );
  ANDN U27675 ( .B(n28124), .A(n28125), .Z(n28122) );
  XOR U27676 ( .A(n28123), .B(n28126), .Z(n28124) );
  XOR U27677 ( .A(n28127), .B(n28128), .Z(n28111) );
  XOR U27678 ( .A(n28129), .B(n28130), .Z(n28128) );
  ANDN U27679 ( .B(n28131), .A(n28132), .Z(n28129) );
  XOR U27680 ( .A(n28133), .B(n28130), .Z(n28131) );
  IV U27681 ( .A(n28109), .Z(n28127) );
  XOR U27682 ( .A(n28134), .B(n28135), .Z(n28109) );
  ANDN U27683 ( .B(n28136), .A(n28137), .Z(n28134) );
  XOR U27684 ( .A(n28135), .B(n28138), .Z(n28136) );
  IV U27685 ( .A(n28117), .Z(n28121) );
  XOR U27686 ( .A(n28117), .B(n28099), .Z(n28119) );
  XOR U27687 ( .A(n28139), .B(n28140), .Z(n28099) );
  AND U27688 ( .A(n1574), .B(n28141), .Z(n28139) );
  XOR U27689 ( .A(n28142), .B(n28140), .Z(n28141) );
  NANDN U27690 ( .A(n28101), .B(n28103), .Z(n28117) );
  XOR U27691 ( .A(n28143), .B(n28144), .Z(n28103) );
  AND U27692 ( .A(n1574), .B(n28145), .Z(n28143) );
  XOR U27693 ( .A(n28144), .B(n28146), .Z(n28145) );
  XOR U27694 ( .A(n28147), .B(n28148), .Z(n1574) );
  AND U27695 ( .A(n28149), .B(n28150), .Z(n28147) );
  XNOR U27696 ( .A(n28148), .B(n28114), .Z(n28150) );
  XNOR U27697 ( .A(n28151), .B(n28152), .Z(n28114) );
  ANDN U27698 ( .B(n28153), .A(n28154), .Z(n28151) );
  XOR U27699 ( .A(n28152), .B(n28155), .Z(n28153) );
  XOR U27700 ( .A(n28148), .B(n28116), .Z(n28149) );
  XOR U27701 ( .A(n28156), .B(n28157), .Z(n28116) );
  AND U27702 ( .A(n1578), .B(n28158), .Z(n28156) );
  XOR U27703 ( .A(n28159), .B(n28157), .Z(n28158) );
  XNOR U27704 ( .A(n28160), .B(n28161), .Z(n28148) );
  NAND U27705 ( .A(n28162), .B(n28163), .Z(n28161) );
  XOR U27706 ( .A(n28164), .B(n28140), .Z(n28163) );
  XOR U27707 ( .A(n28154), .B(n28155), .Z(n28140) );
  XOR U27708 ( .A(n28165), .B(n28166), .Z(n28155) );
  ANDN U27709 ( .B(n28167), .A(n28168), .Z(n28165) );
  XOR U27710 ( .A(n28166), .B(n28169), .Z(n28167) );
  XOR U27711 ( .A(n28170), .B(n28171), .Z(n28154) );
  XOR U27712 ( .A(n28172), .B(n28173), .Z(n28171) );
  ANDN U27713 ( .B(n28174), .A(n28175), .Z(n28172) );
  XOR U27714 ( .A(n28176), .B(n28173), .Z(n28174) );
  IV U27715 ( .A(n28152), .Z(n28170) );
  XOR U27716 ( .A(n28177), .B(n28178), .Z(n28152) );
  ANDN U27717 ( .B(n28179), .A(n28180), .Z(n28177) );
  XOR U27718 ( .A(n28178), .B(n28181), .Z(n28179) );
  IV U27719 ( .A(n28160), .Z(n28164) );
  XOR U27720 ( .A(n28160), .B(n28142), .Z(n28162) );
  XOR U27721 ( .A(n28182), .B(n28183), .Z(n28142) );
  AND U27722 ( .A(n1578), .B(n28184), .Z(n28182) );
  XOR U27723 ( .A(n28185), .B(n28183), .Z(n28184) );
  NANDN U27724 ( .A(n28144), .B(n28146), .Z(n28160) );
  XOR U27725 ( .A(n28186), .B(n28187), .Z(n28146) );
  AND U27726 ( .A(n1578), .B(n28188), .Z(n28186) );
  XOR U27727 ( .A(n28187), .B(n28189), .Z(n28188) );
  XOR U27728 ( .A(n28190), .B(n28191), .Z(n1578) );
  AND U27729 ( .A(n28192), .B(n28193), .Z(n28190) );
  XNOR U27730 ( .A(n28191), .B(n28157), .Z(n28193) );
  XNOR U27731 ( .A(n28194), .B(n28195), .Z(n28157) );
  ANDN U27732 ( .B(n28196), .A(n28197), .Z(n28194) );
  XOR U27733 ( .A(n28195), .B(n28198), .Z(n28196) );
  XOR U27734 ( .A(n28191), .B(n28159), .Z(n28192) );
  XOR U27735 ( .A(n28199), .B(n28200), .Z(n28159) );
  AND U27736 ( .A(n1582), .B(n28201), .Z(n28199) );
  XOR U27737 ( .A(n28202), .B(n28200), .Z(n28201) );
  XNOR U27738 ( .A(n28203), .B(n28204), .Z(n28191) );
  NAND U27739 ( .A(n28205), .B(n28206), .Z(n28204) );
  XOR U27740 ( .A(n28207), .B(n28183), .Z(n28206) );
  XOR U27741 ( .A(n28197), .B(n28198), .Z(n28183) );
  XOR U27742 ( .A(n28208), .B(n28209), .Z(n28198) );
  ANDN U27743 ( .B(n28210), .A(n28211), .Z(n28208) );
  XOR U27744 ( .A(n28209), .B(n28212), .Z(n28210) );
  XOR U27745 ( .A(n28213), .B(n28214), .Z(n28197) );
  XOR U27746 ( .A(n28215), .B(n28216), .Z(n28214) );
  ANDN U27747 ( .B(n28217), .A(n28218), .Z(n28215) );
  XOR U27748 ( .A(n28219), .B(n28216), .Z(n28217) );
  IV U27749 ( .A(n28195), .Z(n28213) );
  XOR U27750 ( .A(n28220), .B(n28221), .Z(n28195) );
  ANDN U27751 ( .B(n28222), .A(n28223), .Z(n28220) );
  XOR U27752 ( .A(n28221), .B(n28224), .Z(n28222) );
  IV U27753 ( .A(n28203), .Z(n28207) );
  XOR U27754 ( .A(n28203), .B(n28185), .Z(n28205) );
  XOR U27755 ( .A(n28225), .B(n28226), .Z(n28185) );
  AND U27756 ( .A(n1582), .B(n28227), .Z(n28225) );
  XOR U27757 ( .A(n28228), .B(n28226), .Z(n28227) );
  NANDN U27758 ( .A(n28187), .B(n28189), .Z(n28203) );
  XOR U27759 ( .A(n28229), .B(n28230), .Z(n28189) );
  AND U27760 ( .A(n1582), .B(n28231), .Z(n28229) );
  XOR U27761 ( .A(n28230), .B(n28232), .Z(n28231) );
  XOR U27762 ( .A(n28233), .B(n28234), .Z(n1582) );
  AND U27763 ( .A(n28235), .B(n28236), .Z(n28233) );
  XNOR U27764 ( .A(n28234), .B(n28200), .Z(n28236) );
  XNOR U27765 ( .A(n28237), .B(n28238), .Z(n28200) );
  ANDN U27766 ( .B(n28239), .A(n28240), .Z(n28237) );
  XOR U27767 ( .A(n28238), .B(n28241), .Z(n28239) );
  XOR U27768 ( .A(n28234), .B(n28202), .Z(n28235) );
  XOR U27769 ( .A(n28242), .B(n28243), .Z(n28202) );
  AND U27770 ( .A(n1586), .B(n28244), .Z(n28242) );
  XOR U27771 ( .A(n28245), .B(n28243), .Z(n28244) );
  XNOR U27772 ( .A(n28246), .B(n28247), .Z(n28234) );
  NAND U27773 ( .A(n28248), .B(n28249), .Z(n28247) );
  XOR U27774 ( .A(n28250), .B(n28226), .Z(n28249) );
  XOR U27775 ( .A(n28240), .B(n28241), .Z(n28226) );
  XOR U27776 ( .A(n28251), .B(n28252), .Z(n28241) );
  ANDN U27777 ( .B(n28253), .A(n28254), .Z(n28251) );
  XOR U27778 ( .A(n28252), .B(n28255), .Z(n28253) );
  XOR U27779 ( .A(n28256), .B(n28257), .Z(n28240) );
  XOR U27780 ( .A(n28258), .B(n28259), .Z(n28257) );
  ANDN U27781 ( .B(n28260), .A(n28261), .Z(n28258) );
  XOR U27782 ( .A(n28262), .B(n28259), .Z(n28260) );
  IV U27783 ( .A(n28238), .Z(n28256) );
  XOR U27784 ( .A(n28263), .B(n28264), .Z(n28238) );
  ANDN U27785 ( .B(n28265), .A(n28266), .Z(n28263) );
  XOR U27786 ( .A(n28264), .B(n28267), .Z(n28265) );
  IV U27787 ( .A(n28246), .Z(n28250) );
  XOR U27788 ( .A(n28246), .B(n28228), .Z(n28248) );
  XOR U27789 ( .A(n28268), .B(n28269), .Z(n28228) );
  AND U27790 ( .A(n1586), .B(n28270), .Z(n28268) );
  XOR U27791 ( .A(n28271), .B(n28269), .Z(n28270) );
  NANDN U27792 ( .A(n28230), .B(n28232), .Z(n28246) );
  XOR U27793 ( .A(n28272), .B(n28273), .Z(n28232) );
  AND U27794 ( .A(n1586), .B(n28274), .Z(n28272) );
  XOR U27795 ( .A(n28273), .B(n28275), .Z(n28274) );
  XOR U27796 ( .A(n28276), .B(n28277), .Z(n1586) );
  AND U27797 ( .A(n28278), .B(n28279), .Z(n28276) );
  XNOR U27798 ( .A(n28277), .B(n28243), .Z(n28279) );
  XNOR U27799 ( .A(n28280), .B(n28281), .Z(n28243) );
  ANDN U27800 ( .B(n28282), .A(n28283), .Z(n28280) );
  XOR U27801 ( .A(n28281), .B(n28284), .Z(n28282) );
  XOR U27802 ( .A(n28277), .B(n28245), .Z(n28278) );
  XOR U27803 ( .A(n28285), .B(n28286), .Z(n28245) );
  AND U27804 ( .A(n1590), .B(n28287), .Z(n28285) );
  XOR U27805 ( .A(n28288), .B(n28286), .Z(n28287) );
  XNOR U27806 ( .A(n28289), .B(n28290), .Z(n28277) );
  NAND U27807 ( .A(n28291), .B(n28292), .Z(n28290) );
  XOR U27808 ( .A(n28293), .B(n28269), .Z(n28292) );
  XOR U27809 ( .A(n28283), .B(n28284), .Z(n28269) );
  XOR U27810 ( .A(n28294), .B(n28295), .Z(n28284) );
  ANDN U27811 ( .B(n28296), .A(n28297), .Z(n28294) );
  XOR U27812 ( .A(n28295), .B(n28298), .Z(n28296) );
  XOR U27813 ( .A(n28299), .B(n28300), .Z(n28283) );
  XOR U27814 ( .A(n28301), .B(n28302), .Z(n28300) );
  ANDN U27815 ( .B(n28303), .A(n28304), .Z(n28301) );
  XOR U27816 ( .A(n28305), .B(n28302), .Z(n28303) );
  IV U27817 ( .A(n28281), .Z(n28299) );
  XOR U27818 ( .A(n28306), .B(n28307), .Z(n28281) );
  ANDN U27819 ( .B(n28308), .A(n28309), .Z(n28306) );
  XOR U27820 ( .A(n28307), .B(n28310), .Z(n28308) );
  IV U27821 ( .A(n28289), .Z(n28293) );
  XOR U27822 ( .A(n28289), .B(n28271), .Z(n28291) );
  XOR U27823 ( .A(n28311), .B(n28312), .Z(n28271) );
  AND U27824 ( .A(n1590), .B(n28313), .Z(n28311) );
  XOR U27825 ( .A(n28314), .B(n28312), .Z(n28313) );
  NANDN U27826 ( .A(n28273), .B(n28275), .Z(n28289) );
  XOR U27827 ( .A(n28315), .B(n28316), .Z(n28275) );
  AND U27828 ( .A(n1590), .B(n28317), .Z(n28315) );
  XOR U27829 ( .A(n28316), .B(n28318), .Z(n28317) );
  XOR U27830 ( .A(n28319), .B(n28320), .Z(n1590) );
  AND U27831 ( .A(n28321), .B(n28322), .Z(n28319) );
  XNOR U27832 ( .A(n28320), .B(n28286), .Z(n28322) );
  XNOR U27833 ( .A(n28323), .B(n28324), .Z(n28286) );
  ANDN U27834 ( .B(n28325), .A(n28326), .Z(n28323) );
  XOR U27835 ( .A(n28324), .B(n28327), .Z(n28325) );
  XOR U27836 ( .A(n28320), .B(n28288), .Z(n28321) );
  XOR U27837 ( .A(n28328), .B(n28329), .Z(n28288) );
  AND U27838 ( .A(n1594), .B(n28330), .Z(n28328) );
  XOR U27839 ( .A(n28331), .B(n28329), .Z(n28330) );
  XNOR U27840 ( .A(n28332), .B(n28333), .Z(n28320) );
  NAND U27841 ( .A(n28334), .B(n28335), .Z(n28333) );
  XOR U27842 ( .A(n28336), .B(n28312), .Z(n28335) );
  XOR U27843 ( .A(n28326), .B(n28327), .Z(n28312) );
  XOR U27844 ( .A(n28337), .B(n28338), .Z(n28327) );
  ANDN U27845 ( .B(n28339), .A(n28340), .Z(n28337) );
  XOR U27846 ( .A(n28338), .B(n28341), .Z(n28339) );
  XOR U27847 ( .A(n28342), .B(n28343), .Z(n28326) );
  XOR U27848 ( .A(n28344), .B(n28345), .Z(n28343) );
  ANDN U27849 ( .B(n28346), .A(n28347), .Z(n28344) );
  XOR U27850 ( .A(n28348), .B(n28345), .Z(n28346) );
  IV U27851 ( .A(n28324), .Z(n28342) );
  XOR U27852 ( .A(n28349), .B(n28350), .Z(n28324) );
  ANDN U27853 ( .B(n28351), .A(n28352), .Z(n28349) );
  XOR U27854 ( .A(n28350), .B(n28353), .Z(n28351) );
  IV U27855 ( .A(n28332), .Z(n28336) );
  XOR U27856 ( .A(n28332), .B(n28314), .Z(n28334) );
  XOR U27857 ( .A(n28354), .B(n28355), .Z(n28314) );
  AND U27858 ( .A(n1594), .B(n28356), .Z(n28354) );
  XOR U27859 ( .A(n28357), .B(n28355), .Z(n28356) );
  NANDN U27860 ( .A(n28316), .B(n28318), .Z(n28332) );
  XOR U27861 ( .A(n28358), .B(n28359), .Z(n28318) );
  AND U27862 ( .A(n1594), .B(n28360), .Z(n28358) );
  XOR U27863 ( .A(n28359), .B(n28361), .Z(n28360) );
  XOR U27864 ( .A(n28362), .B(n28363), .Z(n1594) );
  AND U27865 ( .A(n28364), .B(n28365), .Z(n28362) );
  XNOR U27866 ( .A(n28363), .B(n28329), .Z(n28365) );
  XNOR U27867 ( .A(n28366), .B(n28367), .Z(n28329) );
  ANDN U27868 ( .B(n28368), .A(n28369), .Z(n28366) );
  XOR U27869 ( .A(n28367), .B(n28370), .Z(n28368) );
  XOR U27870 ( .A(n28363), .B(n28331), .Z(n28364) );
  XOR U27871 ( .A(n28371), .B(n28372), .Z(n28331) );
  AND U27872 ( .A(n1598), .B(n28373), .Z(n28371) );
  XOR U27873 ( .A(n28374), .B(n28372), .Z(n28373) );
  XNOR U27874 ( .A(n28375), .B(n28376), .Z(n28363) );
  NAND U27875 ( .A(n28377), .B(n28378), .Z(n28376) );
  XOR U27876 ( .A(n28379), .B(n28355), .Z(n28378) );
  XOR U27877 ( .A(n28369), .B(n28370), .Z(n28355) );
  XOR U27878 ( .A(n28380), .B(n28381), .Z(n28370) );
  ANDN U27879 ( .B(n28382), .A(n28383), .Z(n28380) );
  XOR U27880 ( .A(n28381), .B(n28384), .Z(n28382) );
  XOR U27881 ( .A(n28385), .B(n28386), .Z(n28369) );
  XOR U27882 ( .A(n28387), .B(n28388), .Z(n28386) );
  ANDN U27883 ( .B(n28389), .A(n28390), .Z(n28387) );
  XOR U27884 ( .A(n28391), .B(n28388), .Z(n28389) );
  IV U27885 ( .A(n28367), .Z(n28385) );
  XOR U27886 ( .A(n28392), .B(n28393), .Z(n28367) );
  ANDN U27887 ( .B(n28394), .A(n28395), .Z(n28392) );
  XOR U27888 ( .A(n28393), .B(n28396), .Z(n28394) );
  IV U27889 ( .A(n28375), .Z(n28379) );
  XOR U27890 ( .A(n28375), .B(n28357), .Z(n28377) );
  XOR U27891 ( .A(n28397), .B(n28398), .Z(n28357) );
  AND U27892 ( .A(n1598), .B(n28399), .Z(n28397) );
  XOR U27893 ( .A(n28400), .B(n28398), .Z(n28399) );
  NANDN U27894 ( .A(n28359), .B(n28361), .Z(n28375) );
  XOR U27895 ( .A(n28401), .B(n28402), .Z(n28361) );
  AND U27896 ( .A(n1598), .B(n28403), .Z(n28401) );
  XOR U27897 ( .A(n28402), .B(n28404), .Z(n28403) );
  XOR U27898 ( .A(n28405), .B(n28406), .Z(n1598) );
  AND U27899 ( .A(n28407), .B(n28408), .Z(n28405) );
  XNOR U27900 ( .A(n28406), .B(n28372), .Z(n28408) );
  XNOR U27901 ( .A(n28409), .B(n28410), .Z(n28372) );
  ANDN U27902 ( .B(n28411), .A(n28412), .Z(n28409) );
  XOR U27903 ( .A(n28410), .B(n28413), .Z(n28411) );
  XOR U27904 ( .A(n28406), .B(n28374), .Z(n28407) );
  XOR U27905 ( .A(n28414), .B(n28415), .Z(n28374) );
  AND U27906 ( .A(n1602), .B(n28416), .Z(n28414) );
  XOR U27907 ( .A(n28417), .B(n28415), .Z(n28416) );
  XNOR U27908 ( .A(n28418), .B(n28419), .Z(n28406) );
  NAND U27909 ( .A(n28420), .B(n28421), .Z(n28419) );
  XOR U27910 ( .A(n28422), .B(n28398), .Z(n28421) );
  XOR U27911 ( .A(n28412), .B(n28413), .Z(n28398) );
  XOR U27912 ( .A(n28423), .B(n28424), .Z(n28413) );
  ANDN U27913 ( .B(n28425), .A(n28426), .Z(n28423) );
  XOR U27914 ( .A(n28424), .B(n28427), .Z(n28425) );
  XOR U27915 ( .A(n28428), .B(n28429), .Z(n28412) );
  XOR U27916 ( .A(n28430), .B(n28431), .Z(n28429) );
  ANDN U27917 ( .B(n28432), .A(n28433), .Z(n28430) );
  XOR U27918 ( .A(n28434), .B(n28431), .Z(n28432) );
  IV U27919 ( .A(n28410), .Z(n28428) );
  XOR U27920 ( .A(n28435), .B(n28436), .Z(n28410) );
  ANDN U27921 ( .B(n28437), .A(n28438), .Z(n28435) );
  XOR U27922 ( .A(n28436), .B(n28439), .Z(n28437) );
  IV U27923 ( .A(n28418), .Z(n28422) );
  XOR U27924 ( .A(n28418), .B(n28400), .Z(n28420) );
  XOR U27925 ( .A(n28440), .B(n28441), .Z(n28400) );
  AND U27926 ( .A(n1602), .B(n28442), .Z(n28440) );
  XOR U27927 ( .A(n28443), .B(n28441), .Z(n28442) );
  NANDN U27928 ( .A(n28402), .B(n28404), .Z(n28418) );
  XOR U27929 ( .A(n28444), .B(n28445), .Z(n28404) );
  AND U27930 ( .A(n1602), .B(n28446), .Z(n28444) );
  XOR U27931 ( .A(n28445), .B(n28447), .Z(n28446) );
  XOR U27932 ( .A(n28448), .B(n28449), .Z(n1602) );
  AND U27933 ( .A(n28450), .B(n28451), .Z(n28448) );
  XNOR U27934 ( .A(n28449), .B(n28415), .Z(n28451) );
  XNOR U27935 ( .A(n28452), .B(n28453), .Z(n28415) );
  ANDN U27936 ( .B(n28454), .A(n28455), .Z(n28452) );
  XOR U27937 ( .A(n28453), .B(n28456), .Z(n28454) );
  XOR U27938 ( .A(n28449), .B(n28417), .Z(n28450) );
  XOR U27939 ( .A(n28457), .B(n28458), .Z(n28417) );
  AND U27940 ( .A(n1606), .B(n28459), .Z(n28457) );
  XOR U27941 ( .A(n28460), .B(n28458), .Z(n28459) );
  XNOR U27942 ( .A(n28461), .B(n28462), .Z(n28449) );
  NAND U27943 ( .A(n28463), .B(n28464), .Z(n28462) );
  XOR U27944 ( .A(n28465), .B(n28441), .Z(n28464) );
  XOR U27945 ( .A(n28455), .B(n28456), .Z(n28441) );
  XOR U27946 ( .A(n28466), .B(n28467), .Z(n28456) );
  ANDN U27947 ( .B(n28468), .A(n28469), .Z(n28466) );
  XOR U27948 ( .A(n28467), .B(n28470), .Z(n28468) );
  XOR U27949 ( .A(n28471), .B(n28472), .Z(n28455) );
  XOR U27950 ( .A(n28473), .B(n28474), .Z(n28472) );
  ANDN U27951 ( .B(n28475), .A(n28476), .Z(n28473) );
  XOR U27952 ( .A(n28477), .B(n28474), .Z(n28475) );
  IV U27953 ( .A(n28453), .Z(n28471) );
  XOR U27954 ( .A(n28478), .B(n28479), .Z(n28453) );
  ANDN U27955 ( .B(n28480), .A(n28481), .Z(n28478) );
  XOR U27956 ( .A(n28479), .B(n28482), .Z(n28480) );
  IV U27957 ( .A(n28461), .Z(n28465) );
  XOR U27958 ( .A(n28461), .B(n28443), .Z(n28463) );
  XOR U27959 ( .A(n28483), .B(n28484), .Z(n28443) );
  AND U27960 ( .A(n1606), .B(n28485), .Z(n28483) );
  XOR U27961 ( .A(n28486), .B(n28484), .Z(n28485) );
  NANDN U27962 ( .A(n28445), .B(n28447), .Z(n28461) );
  XOR U27963 ( .A(n28487), .B(n28488), .Z(n28447) );
  AND U27964 ( .A(n1606), .B(n28489), .Z(n28487) );
  XOR U27965 ( .A(n28488), .B(n28490), .Z(n28489) );
  XOR U27966 ( .A(n28491), .B(n28492), .Z(n1606) );
  AND U27967 ( .A(n28493), .B(n28494), .Z(n28491) );
  XNOR U27968 ( .A(n28492), .B(n28458), .Z(n28494) );
  XNOR U27969 ( .A(n28495), .B(n28496), .Z(n28458) );
  ANDN U27970 ( .B(n28497), .A(n28498), .Z(n28495) );
  XOR U27971 ( .A(n28496), .B(n28499), .Z(n28497) );
  XOR U27972 ( .A(n28492), .B(n28460), .Z(n28493) );
  XOR U27973 ( .A(n28500), .B(n28501), .Z(n28460) );
  AND U27974 ( .A(n1610), .B(n28502), .Z(n28500) );
  XOR U27975 ( .A(n28503), .B(n28501), .Z(n28502) );
  XNOR U27976 ( .A(n28504), .B(n28505), .Z(n28492) );
  NAND U27977 ( .A(n28506), .B(n28507), .Z(n28505) );
  XOR U27978 ( .A(n28508), .B(n28484), .Z(n28507) );
  XOR U27979 ( .A(n28498), .B(n28499), .Z(n28484) );
  XOR U27980 ( .A(n28509), .B(n28510), .Z(n28499) );
  ANDN U27981 ( .B(n28511), .A(n28512), .Z(n28509) );
  XOR U27982 ( .A(n28510), .B(n28513), .Z(n28511) );
  XOR U27983 ( .A(n28514), .B(n28515), .Z(n28498) );
  XOR U27984 ( .A(n28516), .B(n28517), .Z(n28515) );
  ANDN U27985 ( .B(n28518), .A(n28519), .Z(n28516) );
  XOR U27986 ( .A(n28520), .B(n28517), .Z(n28518) );
  IV U27987 ( .A(n28496), .Z(n28514) );
  XOR U27988 ( .A(n28521), .B(n28522), .Z(n28496) );
  ANDN U27989 ( .B(n28523), .A(n28524), .Z(n28521) );
  XOR U27990 ( .A(n28522), .B(n28525), .Z(n28523) );
  IV U27991 ( .A(n28504), .Z(n28508) );
  XOR U27992 ( .A(n28504), .B(n28486), .Z(n28506) );
  XOR U27993 ( .A(n28526), .B(n28527), .Z(n28486) );
  AND U27994 ( .A(n1610), .B(n28528), .Z(n28526) );
  XOR U27995 ( .A(n28529), .B(n28527), .Z(n28528) );
  NANDN U27996 ( .A(n28488), .B(n28490), .Z(n28504) );
  XOR U27997 ( .A(n28530), .B(n28531), .Z(n28490) );
  AND U27998 ( .A(n1610), .B(n28532), .Z(n28530) );
  XOR U27999 ( .A(n28531), .B(n28533), .Z(n28532) );
  XOR U28000 ( .A(n28534), .B(n28535), .Z(n1610) );
  AND U28001 ( .A(n28536), .B(n28537), .Z(n28534) );
  XNOR U28002 ( .A(n28535), .B(n28501), .Z(n28537) );
  XNOR U28003 ( .A(n28538), .B(n28539), .Z(n28501) );
  ANDN U28004 ( .B(n28540), .A(n28541), .Z(n28538) );
  XOR U28005 ( .A(n28539), .B(n28542), .Z(n28540) );
  XOR U28006 ( .A(n28535), .B(n28503), .Z(n28536) );
  XOR U28007 ( .A(n28543), .B(n28544), .Z(n28503) );
  AND U28008 ( .A(n1614), .B(n28545), .Z(n28543) );
  XOR U28009 ( .A(n28546), .B(n28544), .Z(n28545) );
  XNOR U28010 ( .A(n28547), .B(n28548), .Z(n28535) );
  NAND U28011 ( .A(n28549), .B(n28550), .Z(n28548) );
  XOR U28012 ( .A(n28551), .B(n28527), .Z(n28550) );
  XOR U28013 ( .A(n28541), .B(n28542), .Z(n28527) );
  XOR U28014 ( .A(n28552), .B(n28553), .Z(n28542) );
  ANDN U28015 ( .B(n28554), .A(n28555), .Z(n28552) );
  XOR U28016 ( .A(n28553), .B(n28556), .Z(n28554) );
  XOR U28017 ( .A(n28557), .B(n28558), .Z(n28541) );
  XOR U28018 ( .A(n28559), .B(n28560), .Z(n28558) );
  ANDN U28019 ( .B(n28561), .A(n28562), .Z(n28559) );
  XOR U28020 ( .A(n28563), .B(n28560), .Z(n28561) );
  IV U28021 ( .A(n28539), .Z(n28557) );
  XOR U28022 ( .A(n28564), .B(n28565), .Z(n28539) );
  ANDN U28023 ( .B(n28566), .A(n28567), .Z(n28564) );
  XOR U28024 ( .A(n28565), .B(n28568), .Z(n28566) );
  IV U28025 ( .A(n28547), .Z(n28551) );
  XOR U28026 ( .A(n28547), .B(n28529), .Z(n28549) );
  XOR U28027 ( .A(n28569), .B(n28570), .Z(n28529) );
  AND U28028 ( .A(n1614), .B(n28571), .Z(n28569) );
  XOR U28029 ( .A(n28572), .B(n28570), .Z(n28571) );
  NANDN U28030 ( .A(n28531), .B(n28533), .Z(n28547) );
  XOR U28031 ( .A(n28573), .B(n28574), .Z(n28533) );
  AND U28032 ( .A(n1614), .B(n28575), .Z(n28573) );
  XOR U28033 ( .A(n28574), .B(n28576), .Z(n28575) );
  XOR U28034 ( .A(n28577), .B(n28578), .Z(n1614) );
  AND U28035 ( .A(n28579), .B(n28580), .Z(n28577) );
  XNOR U28036 ( .A(n28578), .B(n28544), .Z(n28580) );
  XNOR U28037 ( .A(n28581), .B(n28582), .Z(n28544) );
  ANDN U28038 ( .B(n28583), .A(n28584), .Z(n28581) );
  XOR U28039 ( .A(n28582), .B(n28585), .Z(n28583) );
  XOR U28040 ( .A(n28578), .B(n28546), .Z(n28579) );
  XOR U28041 ( .A(n28586), .B(n28587), .Z(n28546) );
  AND U28042 ( .A(n1618), .B(n28588), .Z(n28586) );
  XOR U28043 ( .A(n28589), .B(n28587), .Z(n28588) );
  XNOR U28044 ( .A(n28590), .B(n28591), .Z(n28578) );
  NAND U28045 ( .A(n28592), .B(n28593), .Z(n28591) );
  XOR U28046 ( .A(n28594), .B(n28570), .Z(n28593) );
  XOR U28047 ( .A(n28584), .B(n28585), .Z(n28570) );
  XOR U28048 ( .A(n28595), .B(n28596), .Z(n28585) );
  ANDN U28049 ( .B(n28597), .A(n28598), .Z(n28595) );
  XOR U28050 ( .A(n28596), .B(n28599), .Z(n28597) );
  XOR U28051 ( .A(n28600), .B(n28601), .Z(n28584) );
  XOR U28052 ( .A(n28602), .B(n28603), .Z(n28601) );
  ANDN U28053 ( .B(n28604), .A(n28605), .Z(n28602) );
  XOR U28054 ( .A(n28606), .B(n28603), .Z(n28604) );
  IV U28055 ( .A(n28582), .Z(n28600) );
  XOR U28056 ( .A(n28607), .B(n28608), .Z(n28582) );
  ANDN U28057 ( .B(n28609), .A(n28610), .Z(n28607) );
  XOR U28058 ( .A(n28608), .B(n28611), .Z(n28609) );
  IV U28059 ( .A(n28590), .Z(n28594) );
  XOR U28060 ( .A(n28590), .B(n28572), .Z(n28592) );
  XOR U28061 ( .A(n28612), .B(n28613), .Z(n28572) );
  AND U28062 ( .A(n1618), .B(n28614), .Z(n28612) );
  XOR U28063 ( .A(n28615), .B(n28613), .Z(n28614) );
  NANDN U28064 ( .A(n28574), .B(n28576), .Z(n28590) );
  XOR U28065 ( .A(n28616), .B(n28617), .Z(n28576) );
  AND U28066 ( .A(n1618), .B(n28618), .Z(n28616) );
  XOR U28067 ( .A(n28617), .B(n28619), .Z(n28618) );
  XOR U28068 ( .A(n28620), .B(n28621), .Z(n1618) );
  AND U28069 ( .A(n28622), .B(n28623), .Z(n28620) );
  XNOR U28070 ( .A(n28621), .B(n28587), .Z(n28623) );
  XNOR U28071 ( .A(n28624), .B(n28625), .Z(n28587) );
  ANDN U28072 ( .B(n28626), .A(n28627), .Z(n28624) );
  XOR U28073 ( .A(n28625), .B(n28628), .Z(n28626) );
  XOR U28074 ( .A(n28621), .B(n28589), .Z(n28622) );
  XOR U28075 ( .A(n28629), .B(n28630), .Z(n28589) );
  AND U28076 ( .A(n1622), .B(n28631), .Z(n28629) );
  XOR U28077 ( .A(n28632), .B(n28630), .Z(n28631) );
  XNOR U28078 ( .A(n28633), .B(n28634), .Z(n28621) );
  NAND U28079 ( .A(n28635), .B(n28636), .Z(n28634) );
  XOR U28080 ( .A(n28637), .B(n28613), .Z(n28636) );
  XOR U28081 ( .A(n28627), .B(n28628), .Z(n28613) );
  XOR U28082 ( .A(n28638), .B(n28639), .Z(n28628) );
  ANDN U28083 ( .B(n28640), .A(n28641), .Z(n28638) );
  XOR U28084 ( .A(n28639), .B(n28642), .Z(n28640) );
  XOR U28085 ( .A(n28643), .B(n28644), .Z(n28627) );
  XOR U28086 ( .A(n28645), .B(n28646), .Z(n28644) );
  ANDN U28087 ( .B(n28647), .A(n28648), .Z(n28645) );
  XOR U28088 ( .A(n28649), .B(n28646), .Z(n28647) );
  IV U28089 ( .A(n28625), .Z(n28643) );
  XOR U28090 ( .A(n28650), .B(n28651), .Z(n28625) );
  ANDN U28091 ( .B(n28652), .A(n28653), .Z(n28650) );
  XOR U28092 ( .A(n28651), .B(n28654), .Z(n28652) );
  IV U28093 ( .A(n28633), .Z(n28637) );
  XOR U28094 ( .A(n28633), .B(n28615), .Z(n28635) );
  XOR U28095 ( .A(n28655), .B(n28656), .Z(n28615) );
  AND U28096 ( .A(n1622), .B(n28657), .Z(n28655) );
  XOR U28097 ( .A(n28658), .B(n28656), .Z(n28657) );
  NANDN U28098 ( .A(n28617), .B(n28619), .Z(n28633) );
  XOR U28099 ( .A(n28659), .B(n28660), .Z(n28619) );
  AND U28100 ( .A(n1622), .B(n28661), .Z(n28659) );
  XOR U28101 ( .A(n28660), .B(n28662), .Z(n28661) );
  XOR U28102 ( .A(n28663), .B(n28664), .Z(n1622) );
  AND U28103 ( .A(n28665), .B(n28666), .Z(n28663) );
  XNOR U28104 ( .A(n28664), .B(n28630), .Z(n28666) );
  XNOR U28105 ( .A(n28667), .B(n28668), .Z(n28630) );
  ANDN U28106 ( .B(n28669), .A(n28670), .Z(n28667) );
  XOR U28107 ( .A(n28668), .B(n28671), .Z(n28669) );
  XOR U28108 ( .A(n28664), .B(n28632), .Z(n28665) );
  XOR U28109 ( .A(n28672), .B(n28673), .Z(n28632) );
  AND U28110 ( .A(n1626), .B(n28674), .Z(n28672) );
  XOR U28111 ( .A(n28675), .B(n28673), .Z(n28674) );
  XNOR U28112 ( .A(n28676), .B(n28677), .Z(n28664) );
  NAND U28113 ( .A(n28678), .B(n28679), .Z(n28677) );
  XOR U28114 ( .A(n28680), .B(n28656), .Z(n28679) );
  XOR U28115 ( .A(n28670), .B(n28671), .Z(n28656) );
  XOR U28116 ( .A(n28681), .B(n28682), .Z(n28671) );
  ANDN U28117 ( .B(n28683), .A(n28684), .Z(n28681) );
  XOR U28118 ( .A(n28682), .B(n28685), .Z(n28683) );
  XOR U28119 ( .A(n28686), .B(n28687), .Z(n28670) );
  XOR U28120 ( .A(n28688), .B(n28689), .Z(n28687) );
  ANDN U28121 ( .B(n28690), .A(n28691), .Z(n28688) );
  XOR U28122 ( .A(n28692), .B(n28689), .Z(n28690) );
  IV U28123 ( .A(n28668), .Z(n28686) );
  XOR U28124 ( .A(n28693), .B(n28694), .Z(n28668) );
  ANDN U28125 ( .B(n28695), .A(n28696), .Z(n28693) );
  XOR U28126 ( .A(n28694), .B(n28697), .Z(n28695) );
  IV U28127 ( .A(n28676), .Z(n28680) );
  XOR U28128 ( .A(n28676), .B(n28658), .Z(n28678) );
  XOR U28129 ( .A(n28698), .B(n28699), .Z(n28658) );
  AND U28130 ( .A(n1626), .B(n28700), .Z(n28698) );
  XOR U28131 ( .A(n28701), .B(n28699), .Z(n28700) );
  NANDN U28132 ( .A(n28660), .B(n28662), .Z(n28676) );
  XOR U28133 ( .A(n28702), .B(n28703), .Z(n28662) );
  AND U28134 ( .A(n1626), .B(n28704), .Z(n28702) );
  XOR U28135 ( .A(n28703), .B(n28705), .Z(n28704) );
  XOR U28136 ( .A(n28706), .B(n28707), .Z(n1626) );
  AND U28137 ( .A(n28708), .B(n28709), .Z(n28706) );
  XNOR U28138 ( .A(n28707), .B(n28673), .Z(n28709) );
  XNOR U28139 ( .A(n28710), .B(n28711), .Z(n28673) );
  ANDN U28140 ( .B(n28712), .A(n28713), .Z(n28710) );
  XOR U28141 ( .A(n28711), .B(n28714), .Z(n28712) );
  XOR U28142 ( .A(n28707), .B(n28675), .Z(n28708) );
  XOR U28143 ( .A(n28715), .B(n28716), .Z(n28675) );
  AND U28144 ( .A(n1630), .B(n28717), .Z(n28715) );
  XOR U28145 ( .A(n28718), .B(n28716), .Z(n28717) );
  XNOR U28146 ( .A(n28719), .B(n28720), .Z(n28707) );
  NAND U28147 ( .A(n28721), .B(n28722), .Z(n28720) );
  XOR U28148 ( .A(n28723), .B(n28699), .Z(n28722) );
  XOR U28149 ( .A(n28713), .B(n28714), .Z(n28699) );
  XOR U28150 ( .A(n28724), .B(n28725), .Z(n28714) );
  ANDN U28151 ( .B(n28726), .A(n28727), .Z(n28724) );
  XOR U28152 ( .A(n28725), .B(n28728), .Z(n28726) );
  XOR U28153 ( .A(n28729), .B(n28730), .Z(n28713) );
  XOR U28154 ( .A(n28731), .B(n28732), .Z(n28730) );
  ANDN U28155 ( .B(n28733), .A(n28734), .Z(n28731) );
  XOR U28156 ( .A(n28735), .B(n28732), .Z(n28733) );
  IV U28157 ( .A(n28711), .Z(n28729) );
  XOR U28158 ( .A(n28736), .B(n28737), .Z(n28711) );
  ANDN U28159 ( .B(n28738), .A(n28739), .Z(n28736) );
  XOR U28160 ( .A(n28737), .B(n28740), .Z(n28738) );
  IV U28161 ( .A(n28719), .Z(n28723) );
  XOR U28162 ( .A(n28719), .B(n28701), .Z(n28721) );
  XOR U28163 ( .A(n28741), .B(n28742), .Z(n28701) );
  AND U28164 ( .A(n1630), .B(n28743), .Z(n28741) );
  XOR U28165 ( .A(n28744), .B(n28742), .Z(n28743) );
  NANDN U28166 ( .A(n28703), .B(n28705), .Z(n28719) );
  XOR U28167 ( .A(n28745), .B(n28746), .Z(n28705) );
  AND U28168 ( .A(n1630), .B(n28747), .Z(n28745) );
  XOR U28169 ( .A(n28746), .B(n28748), .Z(n28747) );
  XOR U28170 ( .A(n28749), .B(n28750), .Z(n1630) );
  AND U28171 ( .A(n28751), .B(n28752), .Z(n28749) );
  XNOR U28172 ( .A(n28750), .B(n28716), .Z(n28752) );
  XNOR U28173 ( .A(n28753), .B(n28754), .Z(n28716) );
  ANDN U28174 ( .B(n28755), .A(n28756), .Z(n28753) );
  XOR U28175 ( .A(n28754), .B(n28757), .Z(n28755) );
  XOR U28176 ( .A(n28750), .B(n28718), .Z(n28751) );
  XOR U28177 ( .A(n28758), .B(n28759), .Z(n28718) );
  AND U28178 ( .A(n1634), .B(n28760), .Z(n28758) );
  XOR U28179 ( .A(n28761), .B(n28759), .Z(n28760) );
  XNOR U28180 ( .A(n28762), .B(n28763), .Z(n28750) );
  NAND U28181 ( .A(n28764), .B(n28765), .Z(n28763) );
  XOR U28182 ( .A(n28766), .B(n28742), .Z(n28765) );
  XOR U28183 ( .A(n28756), .B(n28757), .Z(n28742) );
  XOR U28184 ( .A(n28767), .B(n28768), .Z(n28757) );
  ANDN U28185 ( .B(n28769), .A(n28770), .Z(n28767) );
  XOR U28186 ( .A(n28768), .B(n28771), .Z(n28769) );
  XOR U28187 ( .A(n28772), .B(n28773), .Z(n28756) );
  XOR U28188 ( .A(n28774), .B(n28775), .Z(n28773) );
  ANDN U28189 ( .B(n28776), .A(n28777), .Z(n28774) );
  XOR U28190 ( .A(n28778), .B(n28775), .Z(n28776) );
  IV U28191 ( .A(n28754), .Z(n28772) );
  XOR U28192 ( .A(n28779), .B(n28780), .Z(n28754) );
  ANDN U28193 ( .B(n28781), .A(n28782), .Z(n28779) );
  XOR U28194 ( .A(n28780), .B(n28783), .Z(n28781) );
  IV U28195 ( .A(n28762), .Z(n28766) );
  XOR U28196 ( .A(n28762), .B(n28744), .Z(n28764) );
  XOR U28197 ( .A(n28784), .B(n28785), .Z(n28744) );
  AND U28198 ( .A(n1634), .B(n28786), .Z(n28784) );
  XOR U28199 ( .A(n28787), .B(n28785), .Z(n28786) );
  NANDN U28200 ( .A(n28746), .B(n28748), .Z(n28762) );
  XOR U28201 ( .A(n28788), .B(n28789), .Z(n28748) );
  AND U28202 ( .A(n1634), .B(n28790), .Z(n28788) );
  XOR U28203 ( .A(n28789), .B(n28791), .Z(n28790) );
  XOR U28204 ( .A(n28792), .B(n28793), .Z(n1634) );
  AND U28205 ( .A(n28794), .B(n28795), .Z(n28792) );
  XNOR U28206 ( .A(n28793), .B(n28759), .Z(n28795) );
  XNOR U28207 ( .A(n28796), .B(n28797), .Z(n28759) );
  ANDN U28208 ( .B(n28798), .A(n28799), .Z(n28796) );
  XOR U28209 ( .A(n28797), .B(n28800), .Z(n28798) );
  XOR U28210 ( .A(n28793), .B(n28761), .Z(n28794) );
  XOR U28211 ( .A(n28801), .B(n28802), .Z(n28761) );
  AND U28212 ( .A(n1638), .B(n28803), .Z(n28801) );
  XOR U28213 ( .A(n28804), .B(n28802), .Z(n28803) );
  XNOR U28214 ( .A(n28805), .B(n28806), .Z(n28793) );
  NAND U28215 ( .A(n28807), .B(n28808), .Z(n28806) );
  XOR U28216 ( .A(n28809), .B(n28785), .Z(n28808) );
  XOR U28217 ( .A(n28799), .B(n28800), .Z(n28785) );
  XOR U28218 ( .A(n28810), .B(n28811), .Z(n28800) );
  ANDN U28219 ( .B(n28812), .A(n28813), .Z(n28810) );
  XOR U28220 ( .A(n28811), .B(n28814), .Z(n28812) );
  XOR U28221 ( .A(n28815), .B(n28816), .Z(n28799) );
  XOR U28222 ( .A(n28817), .B(n28818), .Z(n28816) );
  ANDN U28223 ( .B(n28819), .A(n28820), .Z(n28817) );
  XOR U28224 ( .A(n28821), .B(n28818), .Z(n28819) );
  IV U28225 ( .A(n28797), .Z(n28815) );
  XOR U28226 ( .A(n28822), .B(n28823), .Z(n28797) );
  ANDN U28227 ( .B(n28824), .A(n28825), .Z(n28822) );
  XOR U28228 ( .A(n28823), .B(n28826), .Z(n28824) );
  IV U28229 ( .A(n28805), .Z(n28809) );
  XOR U28230 ( .A(n28805), .B(n28787), .Z(n28807) );
  XOR U28231 ( .A(n28827), .B(n28828), .Z(n28787) );
  AND U28232 ( .A(n1638), .B(n28829), .Z(n28827) );
  XOR U28233 ( .A(n28830), .B(n28828), .Z(n28829) );
  NANDN U28234 ( .A(n28789), .B(n28791), .Z(n28805) );
  XOR U28235 ( .A(n28831), .B(n28832), .Z(n28791) );
  AND U28236 ( .A(n1638), .B(n28833), .Z(n28831) );
  XOR U28237 ( .A(n28832), .B(n28834), .Z(n28833) );
  XOR U28238 ( .A(n28835), .B(n28836), .Z(n1638) );
  AND U28239 ( .A(n28837), .B(n28838), .Z(n28835) );
  XNOR U28240 ( .A(n28836), .B(n28802), .Z(n28838) );
  XNOR U28241 ( .A(n28839), .B(n28840), .Z(n28802) );
  ANDN U28242 ( .B(n28841), .A(n28842), .Z(n28839) );
  XOR U28243 ( .A(n28840), .B(n28843), .Z(n28841) );
  XOR U28244 ( .A(n28836), .B(n28804), .Z(n28837) );
  XOR U28245 ( .A(n28844), .B(n28845), .Z(n28804) );
  AND U28246 ( .A(n1642), .B(n28846), .Z(n28844) );
  XOR U28247 ( .A(n28847), .B(n28845), .Z(n28846) );
  XNOR U28248 ( .A(n28848), .B(n28849), .Z(n28836) );
  NAND U28249 ( .A(n28850), .B(n28851), .Z(n28849) );
  XOR U28250 ( .A(n28852), .B(n28828), .Z(n28851) );
  XOR U28251 ( .A(n28842), .B(n28843), .Z(n28828) );
  XOR U28252 ( .A(n28853), .B(n28854), .Z(n28843) );
  ANDN U28253 ( .B(n28855), .A(n28856), .Z(n28853) );
  XOR U28254 ( .A(n28854), .B(n28857), .Z(n28855) );
  XOR U28255 ( .A(n28858), .B(n28859), .Z(n28842) );
  XOR U28256 ( .A(n28860), .B(n28861), .Z(n28859) );
  ANDN U28257 ( .B(n28862), .A(n28863), .Z(n28860) );
  XOR U28258 ( .A(n28864), .B(n28861), .Z(n28862) );
  IV U28259 ( .A(n28840), .Z(n28858) );
  XOR U28260 ( .A(n28865), .B(n28866), .Z(n28840) );
  ANDN U28261 ( .B(n28867), .A(n28868), .Z(n28865) );
  XOR U28262 ( .A(n28866), .B(n28869), .Z(n28867) );
  IV U28263 ( .A(n28848), .Z(n28852) );
  XOR U28264 ( .A(n28848), .B(n28830), .Z(n28850) );
  XOR U28265 ( .A(n28870), .B(n28871), .Z(n28830) );
  AND U28266 ( .A(n1642), .B(n28872), .Z(n28870) );
  XOR U28267 ( .A(n28873), .B(n28871), .Z(n28872) );
  NANDN U28268 ( .A(n28832), .B(n28834), .Z(n28848) );
  XOR U28269 ( .A(n28874), .B(n28875), .Z(n28834) );
  AND U28270 ( .A(n1642), .B(n28876), .Z(n28874) );
  XOR U28271 ( .A(n28875), .B(n28877), .Z(n28876) );
  XOR U28272 ( .A(n28878), .B(n28879), .Z(n1642) );
  AND U28273 ( .A(n28880), .B(n28881), .Z(n28878) );
  XNOR U28274 ( .A(n28879), .B(n28845), .Z(n28881) );
  XNOR U28275 ( .A(n28882), .B(n28883), .Z(n28845) );
  ANDN U28276 ( .B(n28884), .A(n28885), .Z(n28882) );
  XOR U28277 ( .A(n28883), .B(n28886), .Z(n28884) );
  XOR U28278 ( .A(n28879), .B(n28847), .Z(n28880) );
  XOR U28279 ( .A(n28887), .B(n28888), .Z(n28847) );
  AND U28280 ( .A(n1646), .B(n28889), .Z(n28887) );
  XOR U28281 ( .A(n28890), .B(n28888), .Z(n28889) );
  XNOR U28282 ( .A(n28891), .B(n28892), .Z(n28879) );
  NAND U28283 ( .A(n28893), .B(n28894), .Z(n28892) );
  XOR U28284 ( .A(n28895), .B(n28871), .Z(n28894) );
  XOR U28285 ( .A(n28885), .B(n28886), .Z(n28871) );
  XOR U28286 ( .A(n28896), .B(n28897), .Z(n28886) );
  ANDN U28287 ( .B(n28898), .A(n28899), .Z(n28896) );
  XOR U28288 ( .A(n28897), .B(n28900), .Z(n28898) );
  XOR U28289 ( .A(n28901), .B(n28902), .Z(n28885) );
  XOR U28290 ( .A(n28903), .B(n28904), .Z(n28902) );
  ANDN U28291 ( .B(n28905), .A(n28906), .Z(n28903) );
  XOR U28292 ( .A(n28907), .B(n28904), .Z(n28905) );
  IV U28293 ( .A(n28883), .Z(n28901) );
  XOR U28294 ( .A(n28908), .B(n28909), .Z(n28883) );
  ANDN U28295 ( .B(n28910), .A(n28911), .Z(n28908) );
  XOR U28296 ( .A(n28909), .B(n28912), .Z(n28910) );
  IV U28297 ( .A(n28891), .Z(n28895) );
  XOR U28298 ( .A(n28891), .B(n28873), .Z(n28893) );
  XOR U28299 ( .A(n28913), .B(n28914), .Z(n28873) );
  AND U28300 ( .A(n1646), .B(n28915), .Z(n28913) );
  XOR U28301 ( .A(n28916), .B(n28914), .Z(n28915) );
  NANDN U28302 ( .A(n28875), .B(n28877), .Z(n28891) );
  XOR U28303 ( .A(n28917), .B(n28918), .Z(n28877) );
  AND U28304 ( .A(n1646), .B(n28919), .Z(n28917) );
  XOR U28305 ( .A(n28918), .B(n28920), .Z(n28919) );
  XOR U28306 ( .A(n28921), .B(n28922), .Z(n1646) );
  AND U28307 ( .A(n28923), .B(n28924), .Z(n28921) );
  XNOR U28308 ( .A(n28922), .B(n28888), .Z(n28924) );
  XNOR U28309 ( .A(n28925), .B(n28926), .Z(n28888) );
  ANDN U28310 ( .B(n28927), .A(n28928), .Z(n28925) );
  XOR U28311 ( .A(n28926), .B(n28929), .Z(n28927) );
  XOR U28312 ( .A(n28922), .B(n28890), .Z(n28923) );
  XOR U28313 ( .A(n28930), .B(n28931), .Z(n28890) );
  AND U28314 ( .A(n1650), .B(n28932), .Z(n28930) );
  XOR U28315 ( .A(n28933), .B(n28931), .Z(n28932) );
  XNOR U28316 ( .A(n28934), .B(n28935), .Z(n28922) );
  NAND U28317 ( .A(n28936), .B(n28937), .Z(n28935) );
  XOR U28318 ( .A(n28938), .B(n28914), .Z(n28937) );
  XOR U28319 ( .A(n28928), .B(n28929), .Z(n28914) );
  XOR U28320 ( .A(n28939), .B(n28940), .Z(n28929) );
  ANDN U28321 ( .B(n28941), .A(n28942), .Z(n28939) );
  XOR U28322 ( .A(n28940), .B(n28943), .Z(n28941) );
  XOR U28323 ( .A(n28944), .B(n28945), .Z(n28928) );
  XOR U28324 ( .A(n28946), .B(n28947), .Z(n28945) );
  ANDN U28325 ( .B(n28948), .A(n28949), .Z(n28946) );
  XOR U28326 ( .A(n28950), .B(n28947), .Z(n28948) );
  IV U28327 ( .A(n28926), .Z(n28944) );
  XOR U28328 ( .A(n28951), .B(n28952), .Z(n28926) );
  ANDN U28329 ( .B(n28953), .A(n28954), .Z(n28951) );
  XOR U28330 ( .A(n28952), .B(n28955), .Z(n28953) );
  IV U28331 ( .A(n28934), .Z(n28938) );
  XOR U28332 ( .A(n28934), .B(n28916), .Z(n28936) );
  XOR U28333 ( .A(n28956), .B(n28957), .Z(n28916) );
  AND U28334 ( .A(n1650), .B(n28958), .Z(n28956) );
  XOR U28335 ( .A(n28959), .B(n28957), .Z(n28958) );
  NANDN U28336 ( .A(n28918), .B(n28920), .Z(n28934) );
  XOR U28337 ( .A(n28960), .B(n28961), .Z(n28920) );
  AND U28338 ( .A(n1650), .B(n28962), .Z(n28960) );
  XOR U28339 ( .A(n28961), .B(n28963), .Z(n28962) );
  XOR U28340 ( .A(n28964), .B(n28965), .Z(n1650) );
  AND U28341 ( .A(n28966), .B(n28967), .Z(n28964) );
  XNOR U28342 ( .A(n28965), .B(n28931), .Z(n28967) );
  XNOR U28343 ( .A(n28968), .B(n28969), .Z(n28931) );
  ANDN U28344 ( .B(n28970), .A(n28971), .Z(n28968) );
  XOR U28345 ( .A(n28969), .B(n28972), .Z(n28970) );
  XOR U28346 ( .A(n28965), .B(n28933), .Z(n28966) );
  XOR U28347 ( .A(n28973), .B(n28974), .Z(n28933) );
  AND U28348 ( .A(n1654), .B(n28975), .Z(n28973) );
  XOR U28349 ( .A(n28976), .B(n28974), .Z(n28975) );
  XNOR U28350 ( .A(n28977), .B(n28978), .Z(n28965) );
  NAND U28351 ( .A(n28979), .B(n28980), .Z(n28978) );
  XOR U28352 ( .A(n28981), .B(n28957), .Z(n28980) );
  XOR U28353 ( .A(n28971), .B(n28972), .Z(n28957) );
  XOR U28354 ( .A(n28982), .B(n28983), .Z(n28972) );
  ANDN U28355 ( .B(n28984), .A(n28985), .Z(n28982) );
  XOR U28356 ( .A(n28983), .B(n28986), .Z(n28984) );
  XOR U28357 ( .A(n28987), .B(n28988), .Z(n28971) );
  XOR U28358 ( .A(n28989), .B(n28990), .Z(n28988) );
  ANDN U28359 ( .B(n28991), .A(n28992), .Z(n28989) );
  XOR U28360 ( .A(n28993), .B(n28990), .Z(n28991) );
  IV U28361 ( .A(n28969), .Z(n28987) );
  XOR U28362 ( .A(n28994), .B(n28995), .Z(n28969) );
  ANDN U28363 ( .B(n28996), .A(n28997), .Z(n28994) );
  XOR U28364 ( .A(n28995), .B(n28998), .Z(n28996) );
  IV U28365 ( .A(n28977), .Z(n28981) );
  XOR U28366 ( .A(n28977), .B(n28959), .Z(n28979) );
  XOR U28367 ( .A(n28999), .B(n29000), .Z(n28959) );
  AND U28368 ( .A(n1654), .B(n29001), .Z(n28999) );
  XOR U28369 ( .A(n29002), .B(n29000), .Z(n29001) );
  NANDN U28370 ( .A(n28961), .B(n28963), .Z(n28977) );
  XOR U28371 ( .A(n29003), .B(n29004), .Z(n28963) );
  AND U28372 ( .A(n1654), .B(n29005), .Z(n29003) );
  XOR U28373 ( .A(n29004), .B(n29006), .Z(n29005) );
  XOR U28374 ( .A(n29007), .B(n29008), .Z(n1654) );
  AND U28375 ( .A(n29009), .B(n29010), .Z(n29007) );
  XNOR U28376 ( .A(n29008), .B(n28974), .Z(n29010) );
  XNOR U28377 ( .A(n29011), .B(n29012), .Z(n28974) );
  ANDN U28378 ( .B(n29013), .A(n29014), .Z(n29011) );
  XOR U28379 ( .A(n29012), .B(n29015), .Z(n29013) );
  XOR U28380 ( .A(n29008), .B(n28976), .Z(n29009) );
  XOR U28381 ( .A(n29016), .B(n29017), .Z(n28976) );
  AND U28382 ( .A(n1658), .B(n29018), .Z(n29016) );
  XOR U28383 ( .A(n29019), .B(n29017), .Z(n29018) );
  XNOR U28384 ( .A(n29020), .B(n29021), .Z(n29008) );
  NAND U28385 ( .A(n29022), .B(n29023), .Z(n29021) );
  XOR U28386 ( .A(n29024), .B(n29000), .Z(n29023) );
  XOR U28387 ( .A(n29014), .B(n29015), .Z(n29000) );
  XOR U28388 ( .A(n29025), .B(n29026), .Z(n29015) );
  ANDN U28389 ( .B(n29027), .A(n29028), .Z(n29025) );
  XOR U28390 ( .A(n29026), .B(n29029), .Z(n29027) );
  XOR U28391 ( .A(n29030), .B(n29031), .Z(n29014) );
  XOR U28392 ( .A(n29032), .B(n29033), .Z(n29031) );
  ANDN U28393 ( .B(n29034), .A(n29035), .Z(n29032) );
  XOR U28394 ( .A(n29036), .B(n29033), .Z(n29034) );
  IV U28395 ( .A(n29012), .Z(n29030) );
  XOR U28396 ( .A(n29037), .B(n29038), .Z(n29012) );
  ANDN U28397 ( .B(n29039), .A(n29040), .Z(n29037) );
  XOR U28398 ( .A(n29038), .B(n29041), .Z(n29039) );
  IV U28399 ( .A(n29020), .Z(n29024) );
  XOR U28400 ( .A(n29020), .B(n29002), .Z(n29022) );
  XOR U28401 ( .A(n29042), .B(n29043), .Z(n29002) );
  AND U28402 ( .A(n1658), .B(n29044), .Z(n29042) );
  XOR U28403 ( .A(n29045), .B(n29043), .Z(n29044) );
  NANDN U28404 ( .A(n29004), .B(n29006), .Z(n29020) );
  XOR U28405 ( .A(n29046), .B(n29047), .Z(n29006) );
  AND U28406 ( .A(n1658), .B(n29048), .Z(n29046) );
  XOR U28407 ( .A(n29047), .B(n29049), .Z(n29048) );
  XOR U28408 ( .A(n29050), .B(n29051), .Z(n1658) );
  AND U28409 ( .A(n29052), .B(n29053), .Z(n29050) );
  XNOR U28410 ( .A(n29051), .B(n29017), .Z(n29053) );
  XNOR U28411 ( .A(n29054), .B(n29055), .Z(n29017) );
  ANDN U28412 ( .B(n29056), .A(n29057), .Z(n29054) );
  XOR U28413 ( .A(n29055), .B(n29058), .Z(n29056) );
  XOR U28414 ( .A(n29051), .B(n29019), .Z(n29052) );
  XOR U28415 ( .A(n29059), .B(n29060), .Z(n29019) );
  AND U28416 ( .A(n1662), .B(n29061), .Z(n29059) );
  XOR U28417 ( .A(n29062), .B(n29060), .Z(n29061) );
  XNOR U28418 ( .A(n29063), .B(n29064), .Z(n29051) );
  NAND U28419 ( .A(n29065), .B(n29066), .Z(n29064) );
  XOR U28420 ( .A(n29067), .B(n29043), .Z(n29066) );
  XOR U28421 ( .A(n29057), .B(n29058), .Z(n29043) );
  XOR U28422 ( .A(n29068), .B(n29069), .Z(n29058) );
  ANDN U28423 ( .B(n29070), .A(n29071), .Z(n29068) );
  XOR U28424 ( .A(n29069), .B(n29072), .Z(n29070) );
  XOR U28425 ( .A(n29073), .B(n29074), .Z(n29057) );
  XOR U28426 ( .A(n29075), .B(n29076), .Z(n29074) );
  ANDN U28427 ( .B(n29077), .A(n29078), .Z(n29075) );
  XOR U28428 ( .A(n29079), .B(n29076), .Z(n29077) );
  IV U28429 ( .A(n29055), .Z(n29073) );
  XOR U28430 ( .A(n29080), .B(n29081), .Z(n29055) );
  ANDN U28431 ( .B(n29082), .A(n29083), .Z(n29080) );
  XOR U28432 ( .A(n29081), .B(n29084), .Z(n29082) );
  IV U28433 ( .A(n29063), .Z(n29067) );
  XOR U28434 ( .A(n29063), .B(n29045), .Z(n29065) );
  XOR U28435 ( .A(n29085), .B(n29086), .Z(n29045) );
  AND U28436 ( .A(n1662), .B(n29087), .Z(n29085) );
  XOR U28437 ( .A(n29088), .B(n29086), .Z(n29087) );
  NANDN U28438 ( .A(n29047), .B(n29049), .Z(n29063) );
  XOR U28439 ( .A(n29089), .B(n29090), .Z(n29049) );
  AND U28440 ( .A(n1662), .B(n29091), .Z(n29089) );
  XOR U28441 ( .A(n29090), .B(n29092), .Z(n29091) );
  XOR U28442 ( .A(n29093), .B(n29094), .Z(n1662) );
  AND U28443 ( .A(n29095), .B(n29096), .Z(n29093) );
  XNOR U28444 ( .A(n29094), .B(n29060), .Z(n29096) );
  XNOR U28445 ( .A(n29097), .B(n29098), .Z(n29060) );
  ANDN U28446 ( .B(n29099), .A(n29100), .Z(n29097) );
  XOR U28447 ( .A(n29098), .B(n29101), .Z(n29099) );
  XOR U28448 ( .A(n29094), .B(n29062), .Z(n29095) );
  XOR U28449 ( .A(n29102), .B(n29103), .Z(n29062) );
  AND U28450 ( .A(n1666), .B(n29104), .Z(n29102) );
  XOR U28451 ( .A(n29105), .B(n29103), .Z(n29104) );
  XNOR U28452 ( .A(n29106), .B(n29107), .Z(n29094) );
  NAND U28453 ( .A(n29108), .B(n29109), .Z(n29107) );
  XOR U28454 ( .A(n29110), .B(n29086), .Z(n29109) );
  XOR U28455 ( .A(n29100), .B(n29101), .Z(n29086) );
  XOR U28456 ( .A(n29111), .B(n29112), .Z(n29101) );
  ANDN U28457 ( .B(n29113), .A(n29114), .Z(n29111) );
  XOR U28458 ( .A(n29112), .B(n29115), .Z(n29113) );
  XOR U28459 ( .A(n29116), .B(n29117), .Z(n29100) );
  XOR U28460 ( .A(n29118), .B(n29119), .Z(n29117) );
  ANDN U28461 ( .B(n29120), .A(n29121), .Z(n29118) );
  XOR U28462 ( .A(n29122), .B(n29119), .Z(n29120) );
  IV U28463 ( .A(n29098), .Z(n29116) );
  XOR U28464 ( .A(n29123), .B(n29124), .Z(n29098) );
  ANDN U28465 ( .B(n29125), .A(n29126), .Z(n29123) );
  XOR U28466 ( .A(n29124), .B(n29127), .Z(n29125) );
  IV U28467 ( .A(n29106), .Z(n29110) );
  XOR U28468 ( .A(n29106), .B(n29088), .Z(n29108) );
  XOR U28469 ( .A(n29128), .B(n29129), .Z(n29088) );
  AND U28470 ( .A(n1666), .B(n29130), .Z(n29128) );
  XOR U28471 ( .A(n29131), .B(n29129), .Z(n29130) );
  NANDN U28472 ( .A(n29090), .B(n29092), .Z(n29106) );
  XOR U28473 ( .A(n29132), .B(n29133), .Z(n29092) );
  AND U28474 ( .A(n1666), .B(n29134), .Z(n29132) );
  XOR U28475 ( .A(n29133), .B(n29135), .Z(n29134) );
  XOR U28476 ( .A(n29136), .B(n29137), .Z(n1666) );
  AND U28477 ( .A(n29138), .B(n29139), .Z(n29136) );
  XNOR U28478 ( .A(n29137), .B(n29103), .Z(n29139) );
  XNOR U28479 ( .A(n29140), .B(n29141), .Z(n29103) );
  ANDN U28480 ( .B(n29142), .A(n29143), .Z(n29140) );
  XOR U28481 ( .A(n29141), .B(n29144), .Z(n29142) );
  XOR U28482 ( .A(n29137), .B(n29105), .Z(n29138) );
  XOR U28483 ( .A(n29145), .B(n29146), .Z(n29105) );
  AND U28484 ( .A(n1670), .B(n29147), .Z(n29145) );
  XOR U28485 ( .A(n29148), .B(n29146), .Z(n29147) );
  XNOR U28486 ( .A(n29149), .B(n29150), .Z(n29137) );
  NAND U28487 ( .A(n29151), .B(n29152), .Z(n29150) );
  XOR U28488 ( .A(n29153), .B(n29129), .Z(n29152) );
  XOR U28489 ( .A(n29143), .B(n29144), .Z(n29129) );
  XOR U28490 ( .A(n29154), .B(n29155), .Z(n29144) );
  ANDN U28491 ( .B(n29156), .A(n29157), .Z(n29154) );
  XOR U28492 ( .A(n29155), .B(n29158), .Z(n29156) );
  XOR U28493 ( .A(n29159), .B(n29160), .Z(n29143) );
  XOR U28494 ( .A(n29161), .B(n29162), .Z(n29160) );
  ANDN U28495 ( .B(n29163), .A(n29164), .Z(n29161) );
  XOR U28496 ( .A(n29165), .B(n29162), .Z(n29163) );
  IV U28497 ( .A(n29141), .Z(n29159) );
  XOR U28498 ( .A(n29166), .B(n29167), .Z(n29141) );
  ANDN U28499 ( .B(n29168), .A(n29169), .Z(n29166) );
  XOR U28500 ( .A(n29167), .B(n29170), .Z(n29168) );
  IV U28501 ( .A(n29149), .Z(n29153) );
  XOR U28502 ( .A(n29149), .B(n29131), .Z(n29151) );
  XOR U28503 ( .A(n29171), .B(n29172), .Z(n29131) );
  AND U28504 ( .A(n1670), .B(n29173), .Z(n29171) );
  XOR U28505 ( .A(n29174), .B(n29172), .Z(n29173) );
  NANDN U28506 ( .A(n29133), .B(n29135), .Z(n29149) );
  XOR U28507 ( .A(n29175), .B(n29176), .Z(n29135) );
  AND U28508 ( .A(n1670), .B(n29177), .Z(n29175) );
  XOR U28509 ( .A(n29176), .B(n29178), .Z(n29177) );
  XOR U28510 ( .A(n29179), .B(n29180), .Z(n1670) );
  AND U28511 ( .A(n29181), .B(n29182), .Z(n29179) );
  XNOR U28512 ( .A(n29180), .B(n29146), .Z(n29182) );
  XNOR U28513 ( .A(n29183), .B(n29184), .Z(n29146) );
  ANDN U28514 ( .B(n29185), .A(n29186), .Z(n29183) );
  XOR U28515 ( .A(n29184), .B(n29187), .Z(n29185) );
  XOR U28516 ( .A(n29180), .B(n29148), .Z(n29181) );
  XOR U28517 ( .A(n29188), .B(n29189), .Z(n29148) );
  AND U28518 ( .A(n1674), .B(n29190), .Z(n29188) );
  XOR U28519 ( .A(n29191), .B(n29189), .Z(n29190) );
  XNOR U28520 ( .A(n29192), .B(n29193), .Z(n29180) );
  NAND U28521 ( .A(n29194), .B(n29195), .Z(n29193) );
  XOR U28522 ( .A(n29196), .B(n29172), .Z(n29195) );
  XOR U28523 ( .A(n29186), .B(n29187), .Z(n29172) );
  XOR U28524 ( .A(n29197), .B(n29198), .Z(n29187) );
  ANDN U28525 ( .B(n29199), .A(n29200), .Z(n29197) );
  XOR U28526 ( .A(n29198), .B(n29201), .Z(n29199) );
  XOR U28527 ( .A(n29202), .B(n29203), .Z(n29186) );
  XOR U28528 ( .A(n29204), .B(n29205), .Z(n29203) );
  ANDN U28529 ( .B(n29206), .A(n29207), .Z(n29204) );
  XOR U28530 ( .A(n29208), .B(n29205), .Z(n29206) );
  IV U28531 ( .A(n29184), .Z(n29202) );
  XOR U28532 ( .A(n29209), .B(n29210), .Z(n29184) );
  ANDN U28533 ( .B(n29211), .A(n29212), .Z(n29209) );
  XOR U28534 ( .A(n29210), .B(n29213), .Z(n29211) );
  IV U28535 ( .A(n29192), .Z(n29196) );
  XOR U28536 ( .A(n29192), .B(n29174), .Z(n29194) );
  XOR U28537 ( .A(n29214), .B(n29215), .Z(n29174) );
  AND U28538 ( .A(n1674), .B(n29216), .Z(n29214) );
  XOR U28539 ( .A(n29217), .B(n29215), .Z(n29216) );
  NANDN U28540 ( .A(n29176), .B(n29178), .Z(n29192) );
  XOR U28541 ( .A(n29218), .B(n29219), .Z(n29178) );
  AND U28542 ( .A(n1674), .B(n29220), .Z(n29218) );
  XOR U28543 ( .A(n29219), .B(n29221), .Z(n29220) );
  XOR U28544 ( .A(n29222), .B(n29223), .Z(n1674) );
  AND U28545 ( .A(n29224), .B(n29225), .Z(n29222) );
  XNOR U28546 ( .A(n29223), .B(n29189), .Z(n29225) );
  XNOR U28547 ( .A(n29226), .B(n29227), .Z(n29189) );
  ANDN U28548 ( .B(n29228), .A(n29229), .Z(n29226) );
  XOR U28549 ( .A(n29227), .B(n29230), .Z(n29228) );
  XOR U28550 ( .A(n29223), .B(n29191), .Z(n29224) );
  XOR U28551 ( .A(n29231), .B(n29232), .Z(n29191) );
  AND U28552 ( .A(n1678), .B(n29233), .Z(n29231) );
  XOR U28553 ( .A(n29234), .B(n29232), .Z(n29233) );
  XNOR U28554 ( .A(n29235), .B(n29236), .Z(n29223) );
  NAND U28555 ( .A(n29237), .B(n29238), .Z(n29236) );
  XOR U28556 ( .A(n29239), .B(n29215), .Z(n29238) );
  XOR U28557 ( .A(n29229), .B(n29230), .Z(n29215) );
  XOR U28558 ( .A(n29240), .B(n29241), .Z(n29230) );
  ANDN U28559 ( .B(n29242), .A(n29243), .Z(n29240) );
  XOR U28560 ( .A(n29241), .B(n29244), .Z(n29242) );
  XOR U28561 ( .A(n29245), .B(n29246), .Z(n29229) );
  XOR U28562 ( .A(n29247), .B(n29248), .Z(n29246) );
  ANDN U28563 ( .B(n29249), .A(n29250), .Z(n29247) );
  XOR U28564 ( .A(n29251), .B(n29248), .Z(n29249) );
  IV U28565 ( .A(n29227), .Z(n29245) );
  XOR U28566 ( .A(n29252), .B(n29253), .Z(n29227) );
  ANDN U28567 ( .B(n29254), .A(n29255), .Z(n29252) );
  XOR U28568 ( .A(n29253), .B(n29256), .Z(n29254) );
  IV U28569 ( .A(n29235), .Z(n29239) );
  XOR U28570 ( .A(n29235), .B(n29217), .Z(n29237) );
  XOR U28571 ( .A(n29257), .B(n29258), .Z(n29217) );
  AND U28572 ( .A(n1678), .B(n29259), .Z(n29257) );
  XOR U28573 ( .A(n29260), .B(n29258), .Z(n29259) );
  NANDN U28574 ( .A(n29219), .B(n29221), .Z(n29235) );
  XOR U28575 ( .A(n29261), .B(n29262), .Z(n29221) );
  AND U28576 ( .A(n1678), .B(n29263), .Z(n29261) );
  XOR U28577 ( .A(n29262), .B(n29264), .Z(n29263) );
  XOR U28578 ( .A(n29265), .B(n29266), .Z(n1678) );
  AND U28579 ( .A(n29267), .B(n29268), .Z(n29265) );
  XNOR U28580 ( .A(n29266), .B(n29232), .Z(n29268) );
  XNOR U28581 ( .A(n29269), .B(n29270), .Z(n29232) );
  ANDN U28582 ( .B(n29271), .A(n29272), .Z(n29269) );
  XOR U28583 ( .A(n29270), .B(n29273), .Z(n29271) );
  XOR U28584 ( .A(n29266), .B(n29234), .Z(n29267) );
  XOR U28585 ( .A(n29274), .B(n29275), .Z(n29234) );
  AND U28586 ( .A(n1682), .B(n29276), .Z(n29274) );
  XOR U28587 ( .A(n29277), .B(n29275), .Z(n29276) );
  XNOR U28588 ( .A(n29278), .B(n29279), .Z(n29266) );
  NAND U28589 ( .A(n29280), .B(n29281), .Z(n29279) );
  XOR U28590 ( .A(n29282), .B(n29258), .Z(n29281) );
  XOR U28591 ( .A(n29272), .B(n29273), .Z(n29258) );
  XOR U28592 ( .A(n29283), .B(n29284), .Z(n29273) );
  ANDN U28593 ( .B(n29285), .A(n29286), .Z(n29283) );
  XOR U28594 ( .A(n29284), .B(n29287), .Z(n29285) );
  XOR U28595 ( .A(n29288), .B(n29289), .Z(n29272) );
  XOR U28596 ( .A(n29290), .B(n29291), .Z(n29289) );
  ANDN U28597 ( .B(n29292), .A(n29293), .Z(n29290) );
  XOR U28598 ( .A(n29294), .B(n29291), .Z(n29292) );
  IV U28599 ( .A(n29270), .Z(n29288) );
  XOR U28600 ( .A(n29295), .B(n29296), .Z(n29270) );
  ANDN U28601 ( .B(n29297), .A(n29298), .Z(n29295) );
  XOR U28602 ( .A(n29296), .B(n29299), .Z(n29297) );
  IV U28603 ( .A(n29278), .Z(n29282) );
  XOR U28604 ( .A(n29278), .B(n29260), .Z(n29280) );
  XOR U28605 ( .A(n29300), .B(n29301), .Z(n29260) );
  AND U28606 ( .A(n1682), .B(n29302), .Z(n29300) );
  XOR U28607 ( .A(n29303), .B(n29301), .Z(n29302) );
  NANDN U28608 ( .A(n29262), .B(n29264), .Z(n29278) );
  XOR U28609 ( .A(n29304), .B(n29305), .Z(n29264) );
  AND U28610 ( .A(n1682), .B(n29306), .Z(n29304) );
  XOR U28611 ( .A(n29305), .B(n29307), .Z(n29306) );
  XOR U28612 ( .A(n29308), .B(n29309), .Z(n1682) );
  AND U28613 ( .A(n29310), .B(n29311), .Z(n29308) );
  XNOR U28614 ( .A(n29309), .B(n29275), .Z(n29311) );
  XNOR U28615 ( .A(n29312), .B(n29313), .Z(n29275) );
  ANDN U28616 ( .B(n29314), .A(n29315), .Z(n29312) );
  XOR U28617 ( .A(n29313), .B(n29316), .Z(n29314) );
  XOR U28618 ( .A(n29309), .B(n29277), .Z(n29310) );
  XOR U28619 ( .A(n29317), .B(n29318), .Z(n29277) );
  AND U28620 ( .A(n1686), .B(n29319), .Z(n29317) );
  XOR U28621 ( .A(n29320), .B(n29318), .Z(n29319) );
  XNOR U28622 ( .A(n29321), .B(n29322), .Z(n29309) );
  NAND U28623 ( .A(n29323), .B(n29324), .Z(n29322) );
  XOR U28624 ( .A(n29325), .B(n29301), .Z(n29324) );
  XOR U28625 ( .A(n29315), .B(n29316), .Z(n29301) );
  XOR U28626 ( .A(n29326), .B(n29327), .Z(n29316) );
  ANDN U28627 ( .B(n29328), .A(n29329), .Z(n29326) );
  XOR U28628 ( .A(n29327), .B(n29330), .Z(n29328) );
  XOR U28629 ( .A(n29331), .B(n29332), .Z(n29315) );
  XOR U28630 ( .A(n29333), .B(n29334), .Z(n29332) );
  ANDN U28631 ( .B(n29335), .A(n29336), .Z(n29333) );
  XOR U28632 ( .A(n29337), .B(n29334), .Z(n29335) );
  IV U28633 ( .A(n29313), .Z(n29331) );
  XOR U28634 ( .A(n29338), .B(n29339), .Z(n29313) );
  ANDN U28635 ( .B(n29340), .A(n29341), .Z(n29338) );
  XOR U28636 ( .A(n29339), .B(n29342), .Z(n29340) );
  IV U28637 ( .A(n29321), .Z(n29325) );
  XOR U28638 ( .A(n29321), .B(n29303), .Z(n29323) );
  XOR U28639 ( .A(n29343), .B(n29344), .Z(n29303) );
  AND U28640 ( .A(n1686), .B(n29345), .Z(n29343) );
  XOR U28641 ( .A(n29346), .B(n29344), .Z(n29345) );
  NANDN U28642 ( .A(n29305), .B(n29307), .Z(n29321) );
  XOR U28643 ( .A(n29347), .B(n29348), .Z(n29307) );
  AND U28644 ( .A(n1686), .B(n29349), .Z(n29347) );
  XOR U28645 ( .A(n29348), .B(n29350), .Z(n29349) );
  XOR U28646 ( .A(n29351), .B(n29352), .Z(n1686) );
  AND U28647 ( .A(n29353), .B(n29354), .Z(n29351) );
  XNOR U28648 ( .A(n29352), .B(n29318), .Z(n29354) );
  XNOR U28649 ( .A(n29355), .B(n29356), .Z(n29318) );
  ANDN U28650 ( .B(n29357), .A(n29358), .Z(n29355) );
  XOR U28651 ( .A(n29356), .B(n29359), .Z(n29357) );
  XOR U28652 ( .A(n29352), .B(n29320), .Z(n29353) );
  XOR U28653 ( .A(n29360), .B(n29361), .Z(n29320) );
  AND U28654 ( .A(n1690), .B(n29362), .Z(n29360) );
  XOR U28655 ( .A(n29363), .B(n29361), .Z(n29362) );
  XNOR U28656 ( .A(n29364), .B(n29365), .Z(n29352) );
  NAND U28657 ( .A(n29366), .B(n29367), .Z(n29365) );
  XOR U28658 ( .A(n29368), .B(n29344), .Z(n29367) );
  XOR U28659 ( .A(n29358), .B(n29359), .Z(n29344) );
  XOR U28660 ( .A(n29369), .B(n29370), .Z(n29359) );
  ANDN U28661 ( .B(n29371), .A(n29372), .Z(n29369) );
  XOR U28662 ( .A(n29370), .B(n29373), .Z(n29371) );
  XOR U28663 ( .A(n29374), .B(n29375), .Z(n29358) );
  XOR U28664 ( .A(n29376), .B(n29377), .Z(n29375) );
  ANDN U28665 ( .B(n29378), .A(n29379), .Z(n29376) );
  XOR U28666 ( .A(n29380), .B(n29377), .Z(n29378) );
  IV U28667 ( .A(n29356), .Z(n29374) );
  XOR U28668 ( .A(n29381), .B(n29382), .Z(n29356) );
  ANDN U28669 ( .B(n29383), .A(n29384), .Z(n29381) );
  XOR U28670 ( .A(n29382), .B(n29385), .Z(n29383) );
  IV U28671 ( .A(n29364), .Z(n29368) );
  XOR U28672 ( .A(n29364), .B(n29346), .Z(n29366) );
  XOR U28673 ( .A(n29386), .B(n29387), .Z(n29346) );
  AND U28674 ( .A(n1690), .B(n29388), .Z(n29386) );
  XOR U28675 ( .A(n29389), .B(n29387), .Z(n29388) );
  NANDN U28676 ( .A(n29348), .B(n29350), .Z(n29364) );
  XOR U28677 ( .A(n29390), .B(n29391), .Z(n29350) );
  AND U28678 ( .A(n1690), .B(n29392), .Z(n29390) );
  XOR U28679 ( .A(n29391), .B(n29393), .Z(n29392) );
  XOR U28680 ( .A(n29394), .B(n29395), .Z(n1690) );
  AND U28681 ( .A(n29396), .B(n29397), .Z(n29394) );
  XNOR U28682 ( .A(n29395), .B(n29361), .Z(n29397) );
  XNOR U28683 ( .A(n29398), .B(n29399), .Z(n29361) );
  ANDN U28684 ( .B(n29400), .A(n29401), .Z(n29398) );
  XOR U28685 ( .A(n29399), .B(n29402), .Z(n29400) );
  XOR U28686 ( .A(n29395), .B(n29363), .Z(n29396) );
  XOR U28687 ( .A(n29403), .B(n29404), .Z(n29363) );
  AND U28688 ( .A(n1694), .B(n29405), .Z(n29403) );
  XOR U28689 ( .A(n29406), .B(n29404), .Z(n29405) );
  XNOR U28690 ( .A(n29407), .B(n29408), .Z(n29395) );
  NAND U28691 ( .A(n29409), .B(n29410), .Z(n29408) );
  XOR U28692 ( .A(n29411), .B(n29387), .Z(n29410) );
  XOR U28693 ( .A(n29401), .B(n29402), .Z(n29387) );
  XOR U28694 ( .A(n29412), .B(n29413), .Z(n29402) );
  ANDN U28695 ( .B(n29414), .A(n29415), .Z(n29412) );
  XOR U28696 ( .A(n29413), .B(n29416), .Z(n29414) );
  XOR U28697 ( .A(n29417), .B(n29418), .Z(n29401) );
  XOR U28698 ( .A(n29419), .B(n29420), .Z(n29418) );
  ANDN U28699 ( .B(n29421), .A(n29422), .Z(n29419) );
  XOR U28700 ( .A(n29423), .B(n29420), .Z(n29421) );
  IV U28701 ( .A(n29399), .Z(n29417) );
  XOR U28702 ( .A(n29424), .B(n29425), .Z(n29399) );
  ANDN U28703 ( .B(n29426), .A(n29427), .Z(n29424) );
  XOR U28704 ( .A(n29425), .B(n29428), .Z(n29426) );
  IV U28705 ( .A(n29407), .Z(n29411) );
  XOR U28706 ( .A(n29407), .B(n29389), .Z(n29409) );
  XOR U28707 ( .A(n29429), .B(n29430), .Z(n29389) );
  AND U28708 ( .A(n1694), .B(n29431), .Z(n29429) );
  XOR U28709 ( .A(n29432), .B(n29430), .Z(n29431) );
  NANDN U28710 ( .A(n29391), .B(n29393), .Z(n29407) );
  XOR U28711 ( .A(n29433), .B(n29434), .Z(n29393) );
  AND U28712 ( .A(n1694), .B(n29435), .Z(n29433) );
  XOR U28713 ( .A(n29434), .B(n29436), .Z(n29435) );
  XOR U28714 ( .A(n29437), .B(n29438), .Z(n1694) );
  AND U28715 ( .A(n29439), .B(n29440), .Z(n29437) );
  XNOR U28716 ( .A(n29438), .B(n29404), .Z(n29440) );
  XNOR U28717 ( .A(n29441), .B(n29442), .Z(n29404) );
  ANDN U28718 ( .B(n29443), .A(n29444), .Z(n29441) );
  XOR U28719 ( .A(n29442), .B(n29445), .Z(n29443) );
  XOR U28720 ( .A(n29438), .B(n29406), .Z(n29439) );
  XOR U28721 ( .A(n29446), .B(n29447), .Z(n29406) );
  AND U28722 ( .A(n1698), .B(n29448), .Z(n29446) );
  XOR U28723 ( .A(n29449), .B(n29447), .Z(n29448) );
  XNOR U28724 ( .A(n29450), .B(n29451), .Z(n29438) );
  NAND U28725 ( .A(n29452), .B(n29453), .Z(n29451) );
  XOR U28726 ( .A(n29454), .B(n29430), .Z(n29453) );
  XOR U28727 ( .A(n29444), .B(n29445), .Z(n29430) );
  XOR U28728 ( .A(n29455), .B(n29456), .Z(n29445) );
  ANDN U28729 ( .B(n29457), .A(n29458), .Z(n29455) );
  XOR U28730 ( .A(n29456), .B(n29459), .Z(n29457) );
  XOR U28731 ( .A(n29460), .B(n29461), .Z(n29444) );
  XOR U28732 ( .A(n29462), .B(n29463), .Z(n29461) );
  ANDN U28733 ( .B(n29464), .A(n29465), .Z(n29462) );
  XOR U28734 ( .A(n29466), .B(n29463), .Z(n29464) );
  IV U28735 ( .A(n29442), .Z(n29460) );
  XOR U28736 ( .A(n29467), .B(n29468), .Z(n29442) );
  ANDN U28737 ( .B(n29469), .A(n29470), .Z(n29467) );
  XOR U28738 ( .A(n29468), .B(n29471), .Z(n29469) );
  IV U28739 ( .A(n29450), .Z(n29454) );
  XOR U28740 ( .A(n29450), .B(n29432), .Z(n29452) );
  XOR U28741 ( .A(n29472), .B(n29473), .Z(n29432) );
  AND U28742 ( .A(n1698), .B(n29474), .Z(n29472) );
  XOR U28743 ( .A(n29475), .B(n29473), .Z(n29474) );
  NANDN U28744 ( .A(n29434), .B(n29436), .Z(n29450) );
  XOR U28745 ( .A(n29476), .B(n29477), .Z(n29436) );
  AND U28746 ( .A(n1698), .B(n29478), .Z(n29476) );
  XOR U28747 ( .A(n29477), .B(n29479), .Z(n29478) );
  XOR U28748 ( .A(n29480), .B(n29481), .Z(n1698) );
  AND U28749 ( .A(n29482), .B(n29483), .Z(n29480) );
  XNOR U28750 ( .A(n29481), .B(n29447), .Z(n29483) );
  XNOR U28751 ( .A(n29484), .B(n29485), .Z(n29447) );
  ANDN U28752 ( .B(n29486), .A(n29487), .Z(n29484) );
  XOR U28753 ( .A(n29485), .B(n29488), .Z(n29486) );
  XOR U28754 ( .A(n29481), .B(n29449), .Z(n29482) );
  XOR U28755 ( .A(n29489), .B(n29490), .Z(n29449) );
  AND U28756 ( .A(n1702), .B(n29491), .Z(n29489) );
  XOR U28757 ( .A(n29492), .B(n29490), .Z(n29491) );
  XNOR U28758 ( .A(n29493), .B(n29494), .Z(n29481) );
  NAND U28759 ( .A(n29495), .B(n29496), .Z(n29494) );
  XOR U28760 ( .A(n29497), .B(n29473), .Z(n29496) );
  XOR U28761 ( .A(n29487), .B(n29488), .Z(n29473) );
  XOR U28762 ( .A(n29498), .B(n29499), .Z(n29488) );
  ANDN U28763 ( .B(n29500), .A(n29501), .Z(n29498) );
  XOR U28764 ( .A(n29499), .B(n29502), .Z(n29500) );
  XOR U28765 ( .A(n29503), .B(n29504), .Z(n29487) );
  XOR U28766 ( .A(n29505), .B(n29506), .Z(n29504) );
  ANDN U28767 ( .B(n29507), .A(n29508), .Z(n29505) );
  XOR U28768 ( .A(n29509), .B(n29506), .Z(n29507) );
  IV U28769 ( .A(n29485), .Z(n29503) );
  XOR U28770 ( .A(n29510), .B(n29511), .Z(n29485) );
  ANDN U28771 ( .B(n29512), .A(n29513), .Z(n29510) );
  XOR U28772 ( .A(n29511), .B(n29514), .Z(n29512) );
  IV U28773 ( .A(n29493), .Z(n29497) );
  XOR U28774 ( .A(n29493), .B(n29475), .Z(n29495) );
  XOR U28775 ( .A(n29515), .B(n29516), .Z(n29475) );
  AND U28776 ( .A(n1702), .B(n29517), .Z(n29515) );
  XOR U28777 ( .A(n29518), .B(n29516), .Z(n29517) );
  NANDN U28778 ( .A(n29477), .B(n29479), .Z(n29493) );
  XOR U28779 ( .A(n29519), .B(n29520), .Z(n29479) );
  AND U28780 ( .A(n1702), .B(n29521), .Z(n29519) );
  XOR U28781 ( .A(n29520), .B(n29522), .Z(n29521) );
  XOR U28782 ( .A(n29523), .B(n29524), .Z(n1702) );
  AND U28783 ( .A(n29525), .B(n29526), .Z(n29523) );
  XNOR U28784 ( .A(n29524), .B(n29490), .Z(n29526) );
  XNOR U28785 ( .A(n29527), .B(n29528), .Z(n29490) );
  ANDN U28786 ( .B(n29529), .A(n29530), .Z(n29527) );
  XOR U28787 ( .A(n29528), .B(n29531), .Z(n29529) );
  XOR U28788 ( .A(n29524), .B(n29492), .Z(n29525) );
  XOR U28789 ( .A(n29532), .B(n29533), .Z(n29492) );
  AND U28790 ( .A(n1706), .B(n29534), .Z(n29532) );
  XOR U28791 ( .A(n29535), .B(n29533), .Z(n29534) );
  XNOR U28792 ( .A(n29536), .B(n29537), .Z(n29524) );
  NAND U28793 ( .A(n29538), .B(n29539), .Z(n29537) );
  XOR U28794 ( .A(n29540), .B(n29516), .Z(n29539) );
  XOR U28795 ( .A(n29530), .B(n29531), .Z(n29516) );
  XOR U28796 ( .A(n29541), .B(n29542), .Z(n29531) );
  ANDN U28797 ( .B(n29543), .A(n29544), .Z(n29541) );
  XOR U28798 ( .A(n29542), .B(n29545), .Z(n29543) );
  XOR U28799 ( .A(n29546), .B(n29547), .Z(n29530) );
  XOR U28800 ( .A(n29548), .B(n29549), .Z(n29547) );
  ANDN U28801 ( .B(n29550), .A(n29551), .Z(n29548) );
  XOR U28802 ( .A(n29552), .B(n29549), .Z(n29550) );
  IV U28803 ( .A(n29528), .Z(n29546) );
  XOR U28804 ( .A(n29553), .B(n29554), .Z(n29528) );
  ANDN U28805 ( .B(n29555), .A(n29556), .Z(n29553) );
  XOR U28806 ( .A(n29554), .B(n29557), .Z(n29555) );
  IV U28807 ( .A(n29536), .Z(n29540) );
  XOR U28808 ( .A(n29536), .B(n29518), .Z(n29538) );
  XOR U28809 ( .A(n29558), .B(n29559), .Z(n29518) );
  AND U28810 ( .A(n1706), .B(n29560), .Z(n29558) );
  XOR U28811 ( .A(n29561), .B(n29559), .Z(n29560) );
  NANDN U28812 ( .A(n29520), .B(n29522), .Z(n29536) );
  XOR U28813 ( .A(n29562), .B(n29563), .Z(n29522) );
  AND U28814 ( .A(n1706), .B(n29564), .Z(n29562) );
  XOR U28815 ( .A(n29563), .B(n29565), .Z(n29564) );
  XOR U28816 ( .A(n29566), .B(n29567), .Z(n1706) );
  AND U28817 ( .A(n29568), .B(n29569), .Z(n29566) );
  XNOR U28818 ( .A(n29567), .B(n29533), .Z(n29569) );
  XNOR U28819 ( .A(n29570), .B(n29571), .Z(n29533) );
  ANDN U28820 ( .B(n29572), .A(n29573), .Z(n29570) );
  XOR U28821 ( .A(n29571), .B(n29574), .Z(n29572) );
  XOR U28822 ( .A(n29567), .B(n29535), .Z(n29568) );
  XOR U28823 ( .A(n29575), .B(n29576), .Z(n29535) );
  AND U28824 ( .A(n1710), .B(n29577), .Z(n29575) );
  XOR U28825 ( .A(n29578), .B(n29576), .Z(n29577) );
  XNOR U28826 ( .A(n29579), .B(n29580), .Z(n29567) );
  NAND U28827 ( .A(n29581), .B(n29582), .Z(n29580) );
  XOR U28828 ( .A(n29583), .B(n29559), .Z(n29582) );
  XOR U28829 ( .A(n29573), .B(n29574), .Z(n29559) );
  XOR U28830 ( .A(n29584), .B(n29585), .Z(n29574) );
  ANDN U28831 ( .B(n29586), .A(n29587), .Z(n29584) );
  XOR U28832 ( .A(n29585), .B(n29588), .Z(n29586) );
  XOR U28833 ( .A(n29589), .B(n29590), .Z(n29573) );
  XOR U28834 ( .A(n29591), .B(n29592), .Z(n29590) );
  ANDN U28835 ( .B(n29593), .A(n29594), .Z(n29591) );
  XOR U28836 ( .A(n29595), .B(n29592), .Z(n29593) );
  IV U28837 ( .A(n29571), .Z(n29589) );
  XOR U28838 ( .A(n29596), .B(n29597), .Z(n29571) );
  ANDN U28839 ( .B(n29598), .A(n29599), .Z(n29596) );
  XOR U28840 ( .A(n29597), .B(n29600), .Z(n29598) );
  IV U28841 ( .A(n29579), .Z(n29583) );
  XOR U28842 ( .A(n29579), .B(n29561), .Z(n29581) );
  XOR U28843 ( .A(n29601), .B(n29602), .Z(n29561) );
  AND U28844 ( .A(n1710), .B(n29603), .Z(n29601) );
  XOR U28845 ( .A(n29604), .B(n29602), .Z(n29603) );
  NANDN U28846 ( .A(n29563), .B(n29565), .Z(n29579) );
  XOR U28847 ( .A(n29605), .B(n29606), .Z(n29565) );
  AND U28848 ( .A(n1710), .B(n29607), .Z(n29605) );
  XOR U28849 ( .A(n29606), .B(n29608), .Z(n29607) );
  XOR U28850 ( .A(n29609), .B(n29610), .Z(n1710) );
  AND U28851 ( .A(n29611), .B(n29612), .Z(n29609) );
  XNOR U28852 ( .A(n29610), .B(n29576), .Z(n29612) );
  XNOR U28853 ( .A(n29613), .B(n29614), .Z(n29576) );
  ANDN U28854 ( .B(n29615), .A(n29616), .Z(n29613) );
  XOR U28855 ( .A(n29614), .B(n29617), .Z(n29615) );
  XOR U28856 ( .A(n29610), .B(n29578), .Z(n29611) );
  XOR U28857 ( .A(n29618), .B(n29619), .Z(n29578) );
  AND U28858 ( .A(n1714), .B(n29620), .Z(n29618) );
  XOR U28859 ( .A(n29621), .B(n29619), .Z(n29620) );
  XNOR U28860 ( .A(n29622), .B(n29623), .Z(n29610) );
  NAND U28861 ( .A(n29624), .B(n29625), .Z(n29623) );
  XOR U28862 ( .A(n29626), .B(n29602), .Z(n29625) );
  XOR U28863 ( .A(n29616), .B(n29617), .Z(n29602) );
  XOR U28864 ( .A(n29627), .B(n29628), .Z(n29617) );
  ANDN U28865 ( .B(n29629), .A(n29630), .Z(n29627) );
  XOR U28866 ( .A(n29628), .B(n29631), .Z(n29629) );
  XOR U28867 ( .A(n29632), .B(n29633), .Z(n29616) );
  XOR U28868 ( .A(n29634), .B(n29635), .Z(n29633) );
  ANDN U28869 ( .B(n29636), .A(n29637), .Z(n29634) );
  XOR U28870 ( .A(n29638), .B(n29635), .Z(n29636) );
  IV U28871 ( .A(n29614), .Z(n29632) );
  XOR U28872 ( .A(n29639), .B(n29640), .Z(n29614) );
  ANDN U28873 ( .B(n29641), .A(n29642), .Z(n29639) );
  XOR U28874 ( .A(n29640), .B(n29643), .Z(n29641) );
  IV U28875 ( .A(n29622), .Z(n29626) );
  XOR U28876 ( .A(n29622), .B(n29604), .Z(n29624) );
  XOR U28877 ( .A(n29644), .B(n29645), .Z(n29604) );
  AND U28878 ( .A(n1714), .B(n29646), .Z(n29644) );
  XOR U28879 ( .A(n29647), .B(n29645), .Z(n29646) );
  NANDN U28880 ( .A(n29606), .B(n29608), .Z(n29622) );
  XOR U28881 ( .A(n29648), .B(n29649), .Z(n29608) );
  AND U28882 ( .A(n1714), .B(n29650), .Z(n29648) );
  XOR U28883 ( .A(n29649), .B(n29651), .Z(n29650) );
  XOR U28884 ( .A(n29652), .B(n29653), .Z(n1714) );
  AND U28885 ( .A(n29654), .B(n29655), .Z(n29652) );
  XNOR U28886 ( .A(n29653), .B(n29619), .Z(n29655) );
  XNOR U28887 ( .A(n29656), .B(n29657), .Z(n29619) );
  ANDN U28888 ( .B(n29658), .A(n29659), .Z(n29656) );
  XOR U28889 ( .A(n29657), .B(n29660), .Z(n29658) );
  XOR U28890 ( .A(n29653), .B(n29621), .Z(n29654) );
  XOR U28891 ( .A(n29661), .B(n29662), .Z(n29621) );
  AND U28892 ( .A(n1718), .B(n29663), .Z(n29661) );
  XOR U28893 ( .A(n29664), .B(n29662), .Z(n29663) );
  XNOR U28894 ( .A(n29665), .B(n29666), .Z(n29653) );
  NAND U28895 ( .A(n29667), .B(n29668), .Z(n29666) );
  XOR U28896 ( .A(n29669), .B(n29645), .Z(n29668) );
  XOR U28897 ( .A(n29659), .B(n29660), .Z(n29645) );
  XOR U28898 ( .A(n29670), .B(n29671), .Z(n29660) );
  ANDN U28899 ( .B(n29672), .A(n29673), .Z(n29670) );
  XOR U28900 ( .A(n29671), .B(n29674), .Z(n29672) );
  XOR U28901 ( .A(n29675), .B(n29676), .Z(n29659) );
  XOR U28902 ( .A(n29677), .B(n29678), .Z(n29676) );
  ANDN U28903 ( .B(n29679), .A(n29680), .Z(n29677) );
  XOR U28904 ( .A(n29681), .B(n29678), .Z(n29679) );
  IV U28905 ( .A(n29657), .Z(n29675) );
  XOR U28906 ( .A(n29682), .B(n29683), .Z(n29657) );
  ANDN U28907 ( .B(n29684), .A(n29685), .Z(n29682) );
  XOR U28908 ( .A(n29683), .B(n29686), .Z(n29684) );
  IV U28909 ( .A(n29665), .Z(n29669) );
  XOR U28910 ( .A(n29665), .B(n29647), .Z(n29667) );
  XOR U28911 ( .A(n29687), .B(n29688), .Z(n29647) );
  AND U28912 ( .A(n1718), .B(n29689), .Z(n29687) );
  XOR U28913 ( .A(n29690), .B(n29688), .Z(n29689) );
  NANDN U28914 ( .A(n29649), .B(n29651), .Z(n29665) );
  XOR U28915 ( .A(n29691), .B(n29692), .Z(n29651) );
  AND U28916 ( .A(n1718), .B(n29693), .Z(n29691) );
  XOR U28917 ( .A(n29692), .B(n29694), .Z(n29693) );
  XOR U28918 ( .A(n29695), .B(n29696), .Z(n1718) );
  AND U28919 ( .A(n29697), .B(n29698), .Z(n29695) );
  XNOR U28920 ( .A(n29696), .B(n29662), .Z(n29698) );
  XNOR U28921 ( .A(n29699), .B(n29700), .Z(n29662) );
  ANDN U28922 ( .B(n29701), .A(n29702), .Z(n29699) );
  XOR U28923 ( .A(n29700), .B(n29703), .Z(n29701) );
  XOR U28924 ( .A(n29696), .B(n29664), .Z(n29697) );
  XOR U28925 ( .A(n29704), .B(n29705), .Z(n29664) );
  AND U28926 ( .A(n1722), .B(n29706), .Z(n29704) );
  XOR U28927 ( .A(n29707), .B(n29705), .Z(n29706) );
  XNOR U28928 ( .A(n29708), .B(n29709), .Z(n29696) );
  NAND U28929 ( .A(n29710), .B(n29711), .Z(n29709) );
  XOR U28930 ( .A(n29712), .B(n29688), .Z(n29711) );
  XOR U28931 ( .A(n29702), .B(n29703), .Z(n29688) );
  XOR U28932 ( .A(n29713), .B(n29714), .Z(n29703) );
  ANDN U28933 ( .B(n29715), .A(n29716), .Z(n29713) );
  XOR U28934 ( .A(n29714), .B(n29717), .Z(n29715) );
  XOR U28935 ( .A(n29718), .B(n29719), .Z(n29702) );
  XOR U28936 ( .A(n29720), .B(n29721), .Z(n29719) );
  ANDN U28937 ( .B(n29722), .A(n29723), .Z(n29720) );
  XOR U28938 ( .A(n29724), .B(n29721), .Z(n29722) );
  IV U28939 ( .A(n29700), .Z(n29718) );
  XOR U28940 ( .A(n29725), .B(n29726), .Z(n29700) );
  ANDN U28941 ( .B(n29727), .A(n29728), .Z(n29725) );
  XOR U28942 ( .A(n29726), .B(n29729), .Z(n29727) );
  IV U28943 ( .A(n29708), .Z(n29712) );
  XOR U28944 ( .A(n29708), .B(n29690), .Z(n29710) );
  XOR U28945 ( .A(n29730), .B(n29731), .Z(n29690) );
  AND U28946 ( .A(n1722), .B(n29732), .Z(n29730) );
  XOR U28947 ( .A(n29733), .B(n29731), .Z(n29732) );
  NANDN U28948 ( .A(n29692), .B(n29694), .Z(n29708) );
  XOR U28949 ( .A(n29734), .B(n29735), .Z(n29694) );
  AND U28950 ( .A(n1722), .B(n29736), .Z(n29734) );
  XOR U28951 ( .A(n29735), .B(n29737), .Z(n29736) );
  XOR U28952 ( .A(n29738), .B(n29739), .Z(n1722) );
  AND U28953 ( .A(n29740), .B(n29741), .Z(n29738) );
  XNOR U28954 ( .A(n29739), .B(n29705), .Z(n29741) );
  XNOR U28955 ( .A(n29742), .B(n29743), .Z(n29705) );
  ANDN U28956 ( .B(n29744), .A(n29745), .Z(n29742) );
  XOR U28957 ( .A(n29743), .B(n29746), .Z(n29744) );
  XOR U28958 ( .A(n29739), .B(n29707), .Z(n29740) );
  XOR U28959 ( .A(n29747), .B(n29748), .Z(n29707) );
  AND U28960 ( .A(n1726), .B(n29749), .Z(n29747) );
  XOR U28961 ( .A(n29750), .B(n29748), .Z(n29749) );
  XNOR U28962 ( .A(n29751), .B(n29752), .Z(n29739) );
  NAND U28963 ( .A(n29753), .B(n29754), .Z(n29752) );
  XOR U28964 ( .A(n29755), .B(n29731), .Z(n29754) );
  XOR U28965 ( .A(n29745), .B(n29746), .Z(n29731) );
  XOR U28966 ( .A(n29756), .B(n29757), .Z(n29746) );
  ANDN U28967 ( .B(n29758), .A(n29759), .Z(n29756) );
  XOR U28968 ( .A(n29757), .B(n29760), .Z(n29758) );
  XOR U28969 ( .A(n29761), .B(n29762), .Z(n29745) );
  XOR U28970 ( .A(n29763), .B(n29764), .Z(n29762) );
  ANDN U28971 ( .B(n29765), .A(n29766), .Z(n29763) );
  XOR U28972 ( .A(n29767), .B(n29764), .Z(n29765) );
  IV U28973 ( .A(n29743), .Z(n29761) );
  XOR U28974 ( .A(n29768), .B(n29769), .Z(n29743) );
  ANDN U28975 ( .B(n29770), .A(n29771), .Z(n29768) );
  XOR U28976 ( .A(n29769), .B(n29772), .Z(n29770) );
  IV U28977 ( .A(n29751), .Z(n29755) );
  XOR U28978 ( .A(n29751), .B(n29733), .Z(n29753) );
  XOR U28979 ( .A(n29773), .B(n29774), .Z(n29733) );
  AND U28980 ( .A(n1726), .B(n29775), .Z(n29773) );
  XOR U28981 ( .A(n29776), .B(n29774), .Z(n29775) );
  NANDN U28982 ( .A(n29735), .B(n29737), .Z(n29751) );
  XOR U28983 ( .A(n29777), .B(n29778), .Z(n29737) );
  AND U28984 ( .A(n1726), .B(n29779), .Z(n29777) );
  XOR U28985 ( .A(n29778), .B(n29780), .Z(n29779) );
  XOR U28986 ( .A(n29781), .B(n29782), .Z(n1726) );
  AND U28987 ( .A(n29783), .B(n29784), .Z(n29781) );
  XNOR U28988 ( .A(n29782), .B(n29748), .Z(n29784) );
  XNOR U28989 ( .A(n29785), .B(n29786), .Z(n29748) );
  ANDN U28990 ( .B(n29787), .A(n29788), .Z(n29785) );
  XOR U28991 ( .A(n29786), .B(n29789), .Z(n29787) );
  XOR U28992 ( .A(n29782), .B(n29750), .Z(n29783) );
  XOR U28993 ( .A(n29790), .B(n29791), .Z(n29750) );
  AND U28994 ( .A(n1730), .B(n29792), .Z(n29790) );
  XOR U28995 ( .A(n29793), .B(n29791), .Z(n29792) );
  XNOR U28996 ( .A(n29794), .B(n29795), .Z(n29782) );
  NAND U28997 ( .A(n29796), .B(n29797), .Z(n29795) );
  XOR U28998 ( .A(n29798), .B(n29774), .Z(n29797) );
  XOR U28999 ( .A(n29788), .B(n29789), .Z(n29774) );
  XOR U29000 ( .A(n29799), .B(n29800), .Z(n29789) );
  ANDN U29001 ( .B(n29801), .A(n29802), .Z(n29799) );
  XOR U29002 ( .A(n29800), .B(n29803), .Z(n29801) );
  XOR U29003 ( .A(n29804), .B(n29805), .Z(n29788) );
  XOR U29004 ( .A(n29806), .B(n29807), .Z(n29805) );
  ANDN U29005 ( .B(n29808), .A(n29809), .Z(n29806) );
  XOR U29006 ( .A(n29810), .B(n29807), .Z(n29808) );
  IV U29007 ( .A(n29786), .Z(n29804) );
  XOR U29008 ( .A(n29811), .B(n29812), .Z(n29786) );
  ANDN U29009 ( .B(n29813), .A(n29814), .Z(n29811) );
  XOR U29010 ( .A(n29812), .B(n29815), .Z(n29813) );
  IV U29011 ( .A(n29794), .Z(n29798) );
  XOR U29012 ( .A(n29794), .B(n29776), .Z(n29796) );
  XOR U29013 ( .A(n29816), .B(n29817), .Z(n29776) );
  AND U29014 ( .A(n1730), .B(n29818), .Z(n29816) );
  XOR U29015 ( .A(n29819), .B(n29817), .Z(n29818) );
  NANDN U29016 ( .A(n29778), .B(n29780), .Z(n29794) );
  XOR U29017 ( .A(n29820), .B(n29821), .Z(n29780) );
  AND U29018 ( .A(n1730), .B(n29822), .Z(n29820) );
  XOR U29019 ( .A(n29821), .B(n29823), .Z(n29822) );
  XOR U29020 ( .A(n29824), .B(n29825), .Z(n1730) );
  AND U29021 ( .A(n29826), .B(n29827), .Z(n29824) );
  XNOR U29022 ( .A(n29825), .B(n29791), .Z(n29827) );
  XNOR U29023 ( .A(n29828), .B(n29829), .Z(n29791) );
  ANDN U29024 ( .B(n29830), .A(n29831), .Z(n29828) );
  XOR U29025 ( .A(n29829), .B(n29832), .Z(n29830) );
  XOR U29026 ( .A(n29825), .B(n29793), .Z(n29826) );
  XOR U29027 ( .A(n29833), .B(n29834), .Z(n29793) );
  AND U29028 ( .A(n1734), .B(n29835), .Z(n29833) );
  XOR U29029 ( .A(n29836), .B(n29834), .Z(n29835) );
  XNOR U29030 ( .A(n29837), .B(n29838), .Z(n29825) );
  NAND U29031 ( .A(n29839), .B(n29840), .Z(n29838) );
  XOR U29032 ( .A(n29841), .B(n29817), .Z(n29840) );
  XOR U29033 ( .A(n29831), .B(n29832), .Z(n29817) );
  XOR U29034 ( .A(n29842), .B(n29843), .Z(n29832) );
  ANDN U29035 ( .B(n29844), .A(n29845), .Z(n29842) );
  XOR U29036 ( .A(n29843), .B(n29846), .Z(n29844) );
  XOR U29037 ( .A(n29847), .B(n29848), .Z(n29831) );
  XOR U29038 ( .A(n29849), .B(n29850), .Z(n29848) );
  ANDN U29039 ( .B(n29851), .A(n29852), .Z(n29849) );
  XOR U29040 ( .A(n29853), .B(n29850), .Z(n29851) );
  IV U29041 ( .A(n29829), .Z(n29847) );
  XOR U29042 ( .A(n29854), .B(n29855), .Z(n29829) );
  ANDN U29043 ( .B(n29856), .A(n29857), .Z(n29854) );
  XOR U29044 ( .A(n29855), .B(n29858), .Z(n29856) );
  IV U29045 ( .A(n29837), .Z(n29841) );
  XOR U29046 ( .A(n29837), .B(n29819), .Z(n29839) );
  XOR U29047 ( .A(n29859), .B(n29860), .Z(n29819) );
  AND U29048 ( .A(n1734), .B(n29861), .Z(n29859) );
  XOR U29049 ( .A(n29862), .B(n29860), .Z(n29861) );
  NANDN U29050 ( .A(n29821), .B(n29823), .Z(n29837) );
  XOR U29051 ( .A(n29863), .B(n29864), .Z(n29823) );
  AND U29052 ( .A(n1734), .B(n29865), .Z(n29863) );
  XOR U29053 ( .A(n29864), .B(n29866), .Z(n29865) );
  XOR U29054 ( .A(n29867), .B(n29868), .Z(n1734) );
  AND U29055 ( .A(n29869), .B(n29870), .Z(n29867) );
  XNOR U29056 ( .A(n29868), .B(n29834), .Z(n29870) );
  XNOR U29057 ( .A(n29871), .B(n29872), .Z(n29834) );
  ANDN U29058 ( .B(n29873), .A(n29874), .Z(n29871) );
  XOR U29059 ( .A(n29872), .B(n29875), .Z(n29873) );
  XOR U29060 ( .A(n29868), .B(n29836), .Z(n29869) );
  XOR U29061 ( .A(n29876), .B(n29877), .Z(n29836) );
  AND U29062 ( .A(n1738), .B(n29878), .Z(n29876) );
  XOR U29063 ( .A(n29879), .B(n29877), .Z(n29878) );
  XNOR U29064 ( .A(n29880), .B(n29881), .Z(n29868) );
  NAND U29065 ( .A(n29882), .B(n29883), .Z(n29881) );
  XOR U29066 ( .A(n29884), .B(n29860), .Z(n29883) );
  XOR U29067 ( .A(n29874), .B(n29875), .Z(n29860) );
  XOR U29068 ( .A(n29885), .B(n29886), .Z(n29875) );
  ANDN U29069 ( .B(n29887), .A(n29888), .Z(n29885) );
  XOR U29070 ( .A(n29886), .B(n29889), .Z(n29887) );
  XOR U29071 ( .A(n29890), .B(n29891), .Z(n29874) );
  XOR U29072 ( .A(n29892), .B(n29893), .Z(n29891) );
  ANDN U29073 ( .B(n29894), .A(n29895), .Z(n29892) );
  XOR U29074 ( .A(n29896), .B(n29893), .Z(n29894) );
  IV U29075 ( .A(n29872), .Z(n29890) );
  XOR U29076 ( .A(n29897), .B(n29898), .Z(n29872) );
  ANDN U29077 ( .B(n29899), .A(n29900), .Z(n29897) );
  XOR U29078 ( .A(n29898), .B(n29901), .Z(n29899) );
  IV U29079 ( .A(n29880), .Z(n29884) );
  XOR U29080 ( .A(n29880), .B(n29862), .Z(n29882) );
  XOR U29081 ( .A(n29902), .B(n29903), .Z(n29862) );
  AND U29082 ( .A(n1738), .B(n29904), .Z(n29902) );
  XOR U29083 ( .A(n29905), .B(n29903), .Z(n29904) );
  NANDN U29084 ( .A(n29864), .B(n29866), .Z(n29880) );
  XOR U29085 ( .A(n29906), .B(n29907), .Z(n29866) );
  AND U29086 ( .A(n1738), .B(n29908), .Z(n29906) );
  XOR U29087 ( .A(n29907), .B(n29909), .Z(n29908) );
  XOR U29088 ( .A(n29910), .B(n29911), .Z(n1738) );
  AND U29089 ( .A(n29912), .B(n29913), .Z(n29910) );
  XNOR U29090 ( .A(n29911), .B(n29877), .Z(n29913) );
  XNOR U29091 ( .A(n29914), .B(n29915), .Z(n29877) );
  ANDN U29092 ( .B(n29916), .A(n29917), .Z(n29914) );
  XOR U29093 ( .A(n29915), .B(n29918), .Z(n29916) );
  XOR U29094 ( .A(n29911), .B(n29879), .Z(n29912) );
  XOR U29095 ( .A(n29919), .B(n29920), .Z(n29879) );
  AND U29096 ( .A(n1742), .B(n29921), .Z(n29919) );
  XOR U29097 ( .A(n29922), .B(n29920), .Z(n29921) );
  XNOR U29098 ( .A(n29923), .B(n29924), .Z(n29911) );
  NAND U29099 ( .A(n29925), .B(n29926), .Z(n29924) );
  XOR U29100 ( .A(n29927), .B(n29903), .Z(n29926) );
  XOR U29101 ( .A(n29917), .B(n29918), .Z(n29903) );
  XOR U29102 ( .A(n29928), .B(n29929), .Z(n29918) );
  ANDN U29103 ( .B(n29930), .A(n29931), .Z(n29928) );
  XOR U29104 ( .A(n29929), .B(n29932), .Z(n29930) );
  XOR U29105 ( .A(n29933), .B(n29934), .Z(n29917) );
  XOR U29106 ( .A(n29935), .B(n29936), .Z(n29934) );
  ANDN U29107 ( .B(n29937), .A(n29938), .Z(n29935) );
  XOR U29108 ( .A(n29939), .B(n29936), .Z(n29937) );
  IV U29109 ( .A(n29915), .Z(n29933) );
  XOR U29110 ( .A(n29940), .B(n29941), .Z(n29915) );
  ANDN U29111 ( .B(n29942), .A(n29943), .Z(n29940) );
  XOR U29112 ( .A(n29941), .B(n29944), .Z(n29942) );
  IV U29113 ( .A(n29923), .Z(n29927) );
  XOR U29114 ( .A(n29923), .B(n29905), .Z(n29925) );
  XOR U29115 ( .A(n29945), .B(n29946), .Z(n29905) );
  AND U29116 ( .A(n1742), .B(n29947), .Z(n29945) );
  XOR U29117 ( .A(n29948), .B(n29946), .Z(n29947) );
  NANDN U29118 ( .A(n29907), .B(n29909), .Z(n29923) );
  XOR U29119 ( .A(n29949), .B(n29950), .Z(n29909) );
  AND U29120 ( .A(n1742), .B(n29951), .Z(n29949) );
  XOR U29121 ( .A(n29950), .B(n29952), .Z(n29951) );
  XOR U29122 ( .A(n29953), .B(n29954), .Z(n1742) );
  AND U29123 ( .A(n29955), .B(n29956), .Z(n29953) );
  XNOR U29124 ( .A(n29954), .B(n29920), .Z(n29956) );
  XNOR U29125 ( .A(n29957), .B(n29958), .Z(n29920) );
  ANDN U29126 ( .B(n29959), .A(n29960), .Z(n29957) );
  XOR U29127 ( .A(n29958), .B(n29961), .Z(n29959) );
  XOR U29128 ( .A(n29954), .B(n29922), .Z(n29955) );
  XOR U29129 ( .A(n29962), .B(n29963), .Z(n29922) );
  AND U29130 ( .A(n1746), .B(n29964), .Z(n29962) );
  XOR U29131 ( .A(n29965), .B(n29963), .Z(n29964) );
  XNOR U29132 ( .A(n29966), .B(n29967), .Z(n29954) );
  NAND U29133 ( .A(n29968), .B(n29969), .Z(n29967) );
  XOR U29134 ( .A(n29970), .B(n29946), .Z(n29969) );
  XOR U29135 ( .A(n29960), .B(n29961), .Z(n29946) );
  XOR U29136 ( .A(n29971), .B(n29972), .Z(n29961) );
  ANDN U29137 ( .B(n29973), .A(n29974), .Z(n29971) );
  XOR U29138 ( .A(n29972), .B(n29975), .Z(n29973) );
  XOR U29139 ( .A(n29976), .B(n29977), .Z(n29960) );
  XOR U29140 ( .A(n29978), .B(n29979), .Z(n29977) );
  ANDN U29141 ( .B(n29980), .A(n29981), .Z(n29978) );
  XOR U29142 ( .A(n29982), .B(n29979), .Z(n29980) );
  IV U29143 ( .A(n29958), .Z(n29976) );
  XOR U29144 ( .A(n29983), .B(n29984), .Z(n29958) );
  ANDN U29145 ( .B(n29985), .A(n29986), .Z(n29983) );
  XOR U29146 ( .A(n29984), .B(n29987), .Z(n29985) );
  IV U29147 ( .A(n29966), .Z(n29970) );
  XOR U29148 ( .A(n29966), .B(n29948), .Z(n29968) );
  XOR U29149 ( .A(n29988), .B(n29989), .Z(n29948) );
  AND U29150 ( .A(n1746), .B(n29990), .Z(n29988) );
  XOR U29151 ( .A(n29991), .B(n29989), .Z(n29990) );
  NANDN U29152 ( .A(n29950), .B(n29952), .Z(n29966) );
  XOR U29153 ( .A(n29992), .B(n29993), .Z(n29952) );
  AND U29154 ( .A(n1746), .B(n29994), .Z(n29992) );
  XOR U29155 ( .A(n29993), .B(n29995), .Z(n29994) );
  XOR U29156 ( .A(n29996), .B(n29997), .Z(n1746) );
  AND U29157 ( .A(n29998), .B(n29999), .Z(n29996) );
  XNOR U29158 ( .A(n29997), .B(n29963), .Z(n29999) );
  XNOR U29159 ( .A(n30000), .B(n30001), .Z(n29963) );
  ANDN U29160 ( .B(n30002), .A(n30003), .Z(n30000) );
  XOR U29161 ( .A(n30001), .B(n30004), .Z(n30002) );
  XOR U29162 ( .A(n29997), .B(n29965), .Z(n29998) );
  XOR U29163 ( .A(n30005), .B(n30006), .Z(n29965) );
  AND U29164 ( .A(n1750), .B(n30007), .Z(n30005) );
  XOR U29165 ( .A(n30008), .B(n30006), .Z(n30007) );
  XNOR U29166 ( .A(n30009), .B(n30010), .Z(n29997) );
  NAND U29167 ( .A(n30011), .B(n30012), .Z(n30010) );
  XOR U29168 ( .A(n30013), .B(n29989), .Z(n30012) );
  XOR U29169 ( .A(n30003), .B(n30004), .Z(n29989) );
  XOR U29170 ( .A(n30014), .B(n30015), .Z(n30004) );
  ANDN U29171 ( .B(n30016), .A(n30017), .Z(n30014) );
  XOR U29172 ( .A(n30015), .B(n30018), .Z(n30016) );
  XOR U29173 ( .A(n30019), .B(n30020), .Z(n30003) );
  XOR U29174 ( .A(n30021), .B(n30022), .Z(n30020) );
  ANDN U29175 ( .B(n30023), .A(n30024), .Z(n30021) );
  XOR U29176 ( .A(n30025), .B(n30022), .Z(n30023) );
  IV U29177 ( .A(n30001), .Z(n30019) );
  XOR U29178 ( .A(n30026), .B(n30027), .Z(n30001) );
  ANDN U29179 ( .B(n30028), .A(n30029), .Z(n30026) );
  XOR U29180 ( .A(n30027), .B(n30030), .Z(n30028) );
  IV U29181 ( .A(n30009), .Z(n30013) );
  XOR U29182 ( .A(n30009), .B(n29991), .Z(n30011) );
  XOR U29183 ( .A(n30031), .B(n30032), .Z(n29991) );
  AND U29184 ( .A(n1750), .B(n30033), .Z(n30031) );
  XOR U29185 ( .A(n30034), .B(n30032), .Z(n30033) );
  NANDN U29186 ( .A(n29993), .B(n29995), .Z(n30009) );
  XOR U29187 ( .A(n30035), .B(n30036), .Z(n29995) );
  AND U29188 ( .A(n1750), .B(n30037), .Z(n30035) );
  XOR U29189 ( .A(n30036), .B(n30038), .Z(n30037) );
  XOR U29190 ( .A(n30039), .B(n30040), .Z(n1750) );
  AND U29191 ( .A(n30041), .B(n30042), .Z(n30039) );
  XNOR U29192 ( .A(n30040), .B(n30006), .Z(n30042) );
  XNOR U29193 ( .A(n30043), .B(n30044), .Z(n30006) );
  ANDN U29194 ( .B(n30045), .A(n30046), .Z(n30043) );
  XOR U29195 ( .A(n30044), .B(n30047), .Z(n30045) );
  XOR U29196 ( .A(n30040), .B(n30008), .Z(n30041) );
  XOR U29197 ( .A(n30048), .B(n30049), .Z(n30008) );
  AND U29198 ( .A(n1754), .B(n30050), .Z(n30048) );
  XOR U29199 ( .A(n30051), .B(n30049), .Z(n30050) );
  XNOR U29200 ( .A(n30052), .B(n30053), .Z(n30040) );
  NAND U29201 ( .A(n30054), .B(n30055), .Z(n30053) );
  XOR U29202 ( .A(n30056), .B(n30032), .Z(n30055) );
  XOR U29203 ( .A(n30046), .B(n30047), .Z(n30032) );
  XOR U29204 ( .A(n30057), .B(n30058), .Z(n30047) );
  ANDN U29205 ( .B(n30059), .A(n30060), .Z(n30057) );
  XOR U29206 ( .A(n30058), .B(n30061), .Z(n30059) );
  XOR U29207 ( .A(n30062), .B(n30063), .Z(n30046) );
  XOR U29208 ( .A(n30064), .B(n30065), .Z(n30063) );
  ANDN U29209 ( .B(n30066), .A(n30067), .Z(n30064) );
  XOR U29210 ( .A(n30068), .B(n30065), .Z(n30066) );
  IV U29211 ( .A(n30044), .Z(n30062) );
  XOR U29212 ( .A(n30069), .B(n30070), .Z(n30044) );
  ANDN U29213 ( .B(n30071), .A(n30072), .Z(n30069) );
  XOR U29214 ( .A(n30070), .B(n30073), .Z(n30071) );
  IV U29215 ( .A(n30052), .Z(n30056) );
  XOR U29216 ( .A(n30052), .B(n30034), .Z(n30054) );
  XOR U29217 ( .A(n30074), .B(n30075), .Z(n30034) );
  AND U29218 ( .A(n1754), .B(n30076), .Z(n30074) );
  XOR U29219 ( .A(n30077), .B(n30075), .Z(n30076) );
  NANDN U29220 ( .A(n30036), .B(n30038), .Z(n30052) );
  XOR U29221 ( .A(n30078), .B(n30079), .Z(n30038) );
  AND U29222 ( .A(n1754), .B(n30080), .Z(n30078) );
  XOR U29223 ( .A(n30079), .B(n30081), .Z(n30080) );
  XOR U29224 ( .A(n30082), .B(n30083), .Z(n1754) );
  AND U29225 ( .A(n30084), .B(n30085), .Z(n30082) );
  XNOR U29226 ( .A(n30083), .B(n30049), .Z(n30085) );
  XNOR U29227 ( .A(n30086), .B(n30087), .Z(n30049) );
  ANDN U29228 ( .B(n30088), .A(n30089), .Z(n30086) );
  XOR U29229 ( .A(n30087), .B(n30090), .Z(n30088) );
  XOR U29230 ( .A(n30083), .B(n30051), .Z(n30084) );
  XOR U29231 ( .A(n30091), .B(n30092), .Z(n30051) );
  AND U29232 ( .A(n1758), .B(n30093), .Z(n30091) );
  XOR U29233 ( .A(n30094), .B(n30092), .Z(n30093) );
  XNOR U29234 ( .A(n30095), .B(n30096), .Z(n30083) );
  NAND U29235 ( .A(n30097), .B(n30098), .Z(n30096) );
  XOR U29236 ( .A(n30099), .B(n30075), .Z(n30098) );
  XOR U29237 ( .A(n30089), .B(n30090), .Z(n30075) );
  XOR U29238 ( .A(n30100), .B(n30101), .Z(n30090) );
  ANDN U29239 ( .B(n30102), .A(n30103), .Z(n30100) );
  XOR U29240 ( .A(n30101), .B(n30104), .Z(n30102) );
  XOR U29241 ( .A(n30105), .B(n30106), .Z(n30089) );
  XOR U29242 ( .A(n30107), .B(n30108), .Z(n30106) );
  ANDN U29243 ( .B(n30109), .A(n30110), .Z(n30107) );
  XOR U29244 ( .A(n30111), .B(n30108), .Z(n30109) );
  IV U29245 ( .A(n30087), .Z(n30105) );
  XOR U29246 ( .A(n30112), .B(n30113), .Z(n30087) );
  ANDN U29247 ( .B(n30114), .A(n30115), .Z(n30112) );
  XOR U29248 ( .A(n30113), .B(n30116), .Z(n30114) );
  IV U29249 ( .A(n30095), .Z(n30099) );
  XOR U29250 ( .A(n30095), .B(n30077), .Z(n30097) );
  XOR U29251 ( .A(n30117), .B(n30118), .Z(n30077) );
  AND U29252 ( .A(n1758), .B(n30119), .Z(n30117) );
  XOR U29253 ( .A(n30120), .B(n30118), .Z(n30119) );
  NANDN U29254 ( .A(n30079), .B(n30081), .Z(n30095) );
  XOR U29255 ( .A(n30121), .B(n30122), .Z(n30081) );
  AND U29256 ( .A(n1758), .B(n30123), .Z(n30121) );
  XOR U29257 ( .A(n30122), .B(n30124), .Z(n30123) );
  XOR U29258 ( .A(n30125), .B(n30126), .Z(n1758) );
  AND U29259 ( .A(n30127), .B(n30128), .Z(n30125) );
  XNOR U29260 ( .A(n30126), .B(n30092), .Z(n30128) );
  XNOR U29261 ( .A(n30129), .B(n30130), .Z(n30092) );
  ANDN U29262 ( .B(n30131), .A(n30132), .Z(n30129) );
  XOR U29263 ( .A(n30130), .B(n30133), .Z(n30131) );
  XOR U29264 ( .A(n30126), .B(n30094), .Z(n30127) );
  XOR U29265 ( .A(n30134), .B(n30135), .Z(n30094) );
  AND U29266 ( .A(n1762), .B(n30136), .Z(n30134) );
  XOR U29267 ( .A(n30137), .B(n30135), .Z(n30136) );
  XNOR U29268 ( .A(n30138), .B(n30139), .Z(n30126) );
  NAND U29269 ( .A(n30140), .B(n30141), .Z(n30139) );
  XOR U29270 ( .A(n30142), .B(n30118), .Z(n30141) );
  XOR U29271 ( .A(n30132), .B(n30133), .Z(n30118) );
  XOR U29272 ( .A(n30143), .B(n30144), .Z(n30133) );
  ANDN U29273 ( .B(n30145), .A(n30146), .Z(n30143) );
  XOR U29274 ( .A(n30144), .B(n30147), .Z(n30145) );
  XOR U29275 ( .A(n30148), .B(n30149), .Z(n30132) );
  XOR U29276 ( .A(n30150), .B(n30151), .Z(n30149) );
  ANDN U29277 ( .B(n30152), .A(n30153), .Z(n30150) );
  XOR U29278 ( .A(n30154), .B(n30151), .Z(n30152) );
  IV U29279 ( .A(n30130), .Z(n30148) );
  XOR U29280 ( .A(n30155), .B(n30156), .Z(n30130) );
  ANDN U29281 ( .B(n30157), .A(n30158), .Z(n30155) );
  XOR U29282 ( .A(n30156), .B(n30159), .Z(n30157) );
  IV U29283 ( .A(n30138), .Z(n30142) );
  XOR U29284 ( .A(n30138), .B(n30120), .Z(n30140) );
  XOR U29285 ( .A(n30160), .B(n30161), .Z(n30120) );
  AND U29286 ( .A(n1762), .B(n30162), .Z(n30160) );
  XOR U29287 ( .A(n30163), .B(n30161), .Z(n30162) );
  NANDN U29288 ( .A(n30122), .B(n30124), .Z(n30138) );
  XOR U29289 ( .A(n30164), .B(n30165), .Z(n30124) );
  AND U29290 ( .A(n1762), .B(n30166), .Z(n30164) );
  XOR U29291 ( .A(n30165), .B(n30167), .Z(n30166) );
  XOR U29292 ( .A(n30168), .B(n30169), .Z(n1762) );
  AND U29293 ( .A(n30170), .B(n30171), .Z(n30168) );
  XNOR U29294 ( .A(n30169), .B(n30135), .Z(n30171) );
  XNOR U29295 ( .A(n30172), .B(n30173), .Z(n30135) );
  ANDN U29296 ( .B(n30174), .A(n30175), .Z(n30172) );
  XOR U29297 ( .A(n30173), .B(n30176), .Z(n30174) );
  XOR U29298 ( .A(n30169), .B(n30137), .Z(n30170) );
  XOR U29299 ( .A(n30177), .B(n30178), .Z(n30137) );
  AND U29300 ( .A(n1766), .B(n30179), .Z(n30177) );
  XOR U29301 ( .A(n30180), .B(n30178), .Z(n30179) );
  XNOR U29302 ( .A(n30181), .B(n30182), .Z(n30169) );
  NAND U29303 ( .A(n30183), .B(n30184), .Z(n30182) );
  XOR U29304 ( .A(n30185), .B(n30161), .Z(n30184) );
  XOR U29305 ( .A(n30175), .B(n30176), .Z(n30161) );
  XOR U29306 ( .A(n30186), .B(n30187), .Z(n30176) );
  ANDN U29307 ( .B(n30188), .A(n30189), .Z(n30186) );
  XOR U29308 ( .A(n30187), .B(n30190), .Z(n30188) );
  XOR U29309 ( .A(n30191), .B(n30192), .Z(n30175) );
  XOR U29310 ( .A(n30193), .B(n30194), .Z(n30192) );
  ANDN U29311 ( .B(n30195), .A(n30196), .Z(n30193) );
  XOR U29312 ( .A(n30197), .B(n30194), .Z(n30195) );
  IV U29313 ( .A(n30173), .Z(n30191) );
  XOR U29314 ( .A(n30198), .B(n30199), .Z(n30173) );
  ANDN U29315 ( .B(n30200), .A(n30201), .Z(n30198) );
  XOR U29316 ( .A(n30199), .B(n30202), .Z(n30200) );
  IV U29317 ( .A(n30181), .Z(n30185) );
  XOR U29318 ( .A(n30181), .B(n30163), .Z(n30183) );
  XOR U29319 ( .A(n30203), .B(n30204), .Z(n30163) );
  AND U29320 ( .A(n1766), .B(n30205), .Z(n30203) );
  XOR U29321 ( .A(n30206), .B(n30204), .Z(n30205) );
  NANDN U29322 ( .A(n30165), .B(n30167), .Z(n30181) );
  XOR U29323 ( .A(n30207), .B(n30208), .Z(n30167) );
  AND U29324 ( .A(n1766), .B(n30209), .Z(n30207) );
  XOR U29325 ( .A(n30208), .B(n30210), .Z(n30209) );
  XOR U29326 ( .A(n30211), .B(n30212), .Z(n1766) );
  AND U29327 ( .A(n30213), .B(n30214), .Z(n30211) );
  XNOR U29328 ( .A(n30212), .B(n30178), .Z(n30214) );
  XNOR U29329 ( .A(n30215), .B(n30216), .Z(n30178) );
  ANDN U29330 ( .B(n30217), .A(n30218), .Z(n30215) );
  XOR U29331 ( .A(n30216), .B(n30219), .Z(n30217) );
  XOR U29332 ( .A(n30212), .B(n30180), .Z(n30213) );
  XOR U29333 ( .A(n30220), .B(n30221), .Z(n30180) );
  AND U29334 ( .A(n1770), .B(n30222), .Z(n30220) );
  XOR U29335 ( .A(n30223), .B(n30221), .Z(n30222) );
  XNOR U29336 ( .A(n30224), .B(n30225), .Z(n30212) );
  NAND U29337 ( .A(n30226), .B(n30227), .Z(n30225) );
  XOR U29338 ( .A(n30228), .B(n30204), .Z(n30227) );
  XOR U29339 ( .A(n30218), .B(n30219), .Z(n30204) );
  XOR U29340 ( .A(n30229), .B(n30230), .Z(n30219) );
  ANDN U29341 ( .B(n30231), .A(n30232), .Z(n30229) );
  XOR U29342 ( .A(n30230), .B(n30233), .Z(n30231) );
  XOR U29343 ( .A(n30234), .B(n30235), .Z(n30218) );
  XOR U29344 ( .A(n30236), .B(n30237), .Z(n30235) );
  ANDN U29345 ( .B(n30238), .A(n30239), .Z(n30236) );
  XOR U29346 ( .A(n30240), .B(n30237), .Z(n30238) );
  IV U29347 ( .A(n30216), .Z(n30234) );
  XOR U29348 ( .A(n30241), .B(n30242), .Z(n30216) );
  ANDN U29349 ( .B(n30243), .A(n30244), .Z(n30241) );
  XOR U29350 ( .A(n30242), .B(n30245), .Z(n30243) );
  IV U29351 ( .A(n30224), .Z(n30228) );
  XOR U29352 ( .A(n30224), .B(n30206), .Z(n30226) );
  XOR U29353 ( .A(n30246), .B(n30247), .Z(n30206) );
  AND U29354 ( .A(n1770), .B(n30248), .Z(n30246) );
  XOR U29355 ( .A(n30249), .B(n30247), .Z(n30248) );
  NANDN U29356 ( .A(n30208), .B(n30210), .Z(n30224) );
  XOR U29357 ( .A(n30250), .B(n30251), .Z(n30210) );
  AND U29358 ( .A(n1770), .B(n30252), .Z(n30250) );
  XOR U29359 ( .A(n30251), .B(n30253), .Z(n30252) );
  XOR U29360 ( .A(n30254), .B(n30255), .Z(n1770) );
  AND U29361 ( .A(n30256), .B(n30257), .Z(n30254) );
  XNOR U29362 ( .A(n30255), .B(n30221), .Z(n30257) );
  XNOR U29363 ( .A(n30258), .B(n30259), .Z(n30221) );
  ANDN U29364 ( .B(n30260), .A(n30261), .Z(n30258) );
  XOR U29365 ( .A(n30259), .B(n30262), .Z(n30260) );
  XOR U29366 ( .A(n30255), .B(n30223), .Z(n30256) );
  XOR U29367 ( .A(n30263), .B(n30264), .Z(n30223) );
  AND U29368 ( .A(n1774), .B(n30265), .Z(n30263) );
  XOR U29369 ( .A(n30266), .B(n30264), .Z(n30265) );
  XNOR U29370 ( .A(n30267), .B(n30268), .Z(n30255) );
  NAND U29371 ( .A(n30269), .B(n30270), .Z(n30268) );
  XOR U29372 ( .A(n30271), .B(n30247), .Z(n30270) );
  XOR U29373 ( .A(n30261), .B(n30262), .Z(n30247) );
  XOR U29374 ( .A(n30272), .B(n30273), .Z(n30262) );
  ANDN U29375 ( .B(n30274), .A(n30275), .Z(n30272) );
  XOR U29376 ( .A(n30273), .B(n30276), .Z(n30274) );
  XOR U29377 ( .A(n30277), .B(n30278), .Z(n30261) );
  XOR U29378 ( .A(n30279), .B(n30280), .Z(n30278) );
  ANDN U29379 ( .B(n30281), .A(n30282), .Z(n30279) );
  XOR U29380 ( .A(n30283), .B(n30280), .Z(n30281) );
  IV U29381 ( .A(n30259), .Z(n30277) );
  XOR U29382 ( .A(n30284), .B(n30285), .Z(n30259) );
  ANDN U29383 ( .B(n30286), .A(n30287), .Z(n30284) );
  XOR U29384 ( .A(n30285), .B(n30288), .Z(n30286) );
  IV U29385 ( .A(n30267), .Z(n30271) );
  XOR U29386 ( .A(n30267), .B(n30249), .Z(n30269) );
  XOR U29387 ( .A(n30289), .B(n30290), .Z(n30249) );
  AND U29388 ( .A(n1774), .B(n30291), .Z(n30289) );
  XOR U29389 ( .A(n30292), .B(n30290), .Z(n30291) );
  NANDN U29390 ( .A(n30251), .B(n30253), .Z(n30267) );
  XOR U29391 ( .A(n30293), .B(n30294), .Z(n30253) );
  AND U29392 ( .A(n1774), .B(n30295), .Z(n30293) );
  XOR U29393 ( .A(n30294), .B(n30296), .Z(n30295) );
  XOR U29394 ( .A(n30297), .B(n30298), .Z(n1774) );
  AND U29395 ( .A(n30299), .B(n30300), .Z(n30297) );
  XNOR U29396 ( .A(n30298), .B(n30264), .Z(n30300) );
  XNOR U29397 ( .A(n30301), .B(n30302), .Z(n30264) );
  ANDN U29398 ( .B(n30303), .A(n30304), .Z(n30301) );
  XOR U29399 ( .A(n30302), .B(n30305), .Z(n30303) );
  XOR U29400 ( .A(n30298), .B(n30266), .Z(n30299) );
  XOR U29401 ( .A(n30306), .B(n30307), .Z(n30266) );
  AND U29402 ( .A(n1778), .B(n30308), .Z(n30306) );
  XOR U29403 ( .A(n30309), .B(n30307), .Z(n30308) );
  XNOR U29404 ( .A(n30310), .B(n30311), .Z(n30298) );
  NAND U29405 ( .A(n30312), .B(n30313), .Z(n30311) );
  XOR U29406 ( .A(n30314), .B(n30290), .Z(n30313) );
  XOR U29407 ( .A(n30304), .B(n30305), .Z(n30290) );
  XOR U29408 ( .A(n30315), .B(n30316), .Z(n30305) );
  ANDN U29409 ( .B(n30317), .A(n30318), .Z(n30315) );
  XOR U29410 ( .A(n30316), .B(n30319), .Z(n30317) );
  XOR U29411 ( .A(n30320), .B(n30321), .Z(n30304) );
  XOR U29412 ( .A(n30322), .B(n30323), .Z(n30321) );
  ANDN U29413 ( .B(n30324), .A(n30325), .Z(n30322) );
  XOR U29414 ( .A(n30326), .B(n30323), .Z(n30324) );
  IV U29415 ( .A(n30302), .Z(n30320) );
  XOR U29416 ( .A(n30327), .B(n30328), .Z(n30302) );
  ANDN U29417 ( .B(n30329), .A(n30330), .Z(n30327) );
  XOR U29418 ( .A(n30328), .B(n30331), .Z(n30329) );
  IV U29419 ( .A(n30310), .Z(n30314) );
  XOR U29420 ( .A(n30310), .B(n30292), .Z(n30312) );
  XOR U29421 ( .A(n30332), .B(n30333), .Z(n30292) );
  AND U29422 ( .A(n1778), .B(n30334), .Z(n30332) );
  XOR U29423 ( .A(n30335), .B(n30333), .Z(n30334) );
  NANDN U29424 ( .A(n30294), .B(n30296), .Z(n30310) );
  XOR U29425 ( .A(n30336), .B(n30337), .Z(n30296) );
  AND U29426 ( .A(n1778), .B(n30338), .Z(n30336) );
  XOR U29427 ( .A(n30337), .B(n30339), .Z(n30338) );
  XOR U29428 ( .A(n30340), .B(n30341), .Z(n1778) );
  AND U29429 ( .A(n30342), .B(n30343), .Z(n30340) );
  XNOR U29430 ( .A(n30341), .B(n30307), .Z(n30343) );
  XNOR U29431 ( .A(n30344), .B(n30345), .Z(n30307) );
  ANDN U29432 ( .B(n30346), .A(n30347), .Z(n30344) );
  XOR U29433 ( .A(n30345), .B(n30348), .Z(n30346) );
  XOR U29434 ( .A(n30341), .B(n30309), .Z(n30342) );
  XOR U29435 ( .A(n30349), .B(n30350), .Z(n30309) );
  AND U29436 ( .A(n1782), .B(n30351), .Z(n30349) );
  XOR U29437 ( .A(n30352), .B(n30350), .Z(n30351) );
  XNOR U29438 ( .A(n30353), .B(n30354), .Z(n30341) );
  NAND U29439 ( .A(n30355), .B(n30356), .Z(n30354) );
  XOR U29440 ( .A(n30357), .B(n30333), .Z(n30356) );
  XOR U29441 ( .A(n30347), .B(n30348), .Z(n30333) );
  XOR U29442 ( .A(n30358), .B(n30359), .Z(n30348) );
  ANDN U29443 ( .B(n30360), .A(n30361), .Z(n30358) );
  XOR U29444 ( .A(n30359), .B(n30362), .Z(n30360) );
  XOR U29445 ( .A(n30363), .B(n30364), .Z(n30347) );
  XOR U29446 ( .A(n30365), .B(n30366), .Z(n30364) );
  ANDN U29447 ( .B(n30367), .A(n30368), .Z(n30365) );
  XOR U29448 ( .A(n30369), .B(n30366), .Z(n30367) );
  IV U29449 ( .A(n30345), .Z(n30363) );
  XOR U29450 ( .A(n30370), .B(n30371), .Z(n30345) );
  ANDN U29451 ( .B(n30372), .A(n30373), .Z(n30370) );
  XOR U29452 ( .A(n30371), .B(n30374), .Z(n30372) );
  IV U29453 ( .A(n30353), .Z(n30357) );
  XOR U29454 ( .A(n30353), .B(n30335), .Z(n30355) );
  XOR U29455 ( .A(n30375), .B(n30376), .Z(n30335) );
  AND U29456 ( .A(n1782), .B(n30377), .Z(n30375) );
  XOR U29457 ( .A(n30378), .B(n30376), .Z(n30377) );
  NANDN U29458 ( .A(n30337), .B(n30339), .Z(n30353) );
  XOR U29459 ( .A(n30379), .B(n30380), .Z(n30339) );
  AND U29460 ( .A(n1782), .B(n30381), .Z(n30379) );
  XOR U29461 ( .A(n30380), .B(n30382), .Z(n30381) );
  XOR U29462 ( .A(n30383), .B(n30384), .Z(n1782) );
  AND U29463 ( .A(n30385), .B(n30386), .Z(n30383) );
  XNOR U29464 ( .A(n30384), .B(n30350), .Z(n30386) );
  XNOR U29465 ( .A(n30387), .B(n30388), .Z(n30350) );
  ANDN U29466 ( .B(n30389), .A(n30390), .Z(n30387) );
  XOR U29467 ( .A(n30388), .B(n30391), .Z(n30389) );
  XOR U29468 ( .A(n30384), .B(n30352), .Z(n30385) );
  XOR U29469 ( .A(n30392), .B(n30393), .Z(n30352) );
  AND U29470 ( .A(n1786), .B(n30394), .Z(n30392) );
  XOR U29471 ( .A(n30395), .B(n30393), .Z(n30394) );
  XNOR U29472 ( .A(n30396), .B(n30397), .Z(n30384) );
  NAND U29473 ( .A(n30398), .B(n30399), .Z(n30397) );
  XOR U29474 ( .A(n30400), .B(n30376), .Z(n30399) );
  XOR U29475 ( .A(n30390), .B(n30391), .Z(n30376) );
  XOR U29476 ( .A(n30401), .B(n30402), .Z(n30391) );
  ANDN U29477 ( .B(n30403), .A(n30404), .Z(n30401) );
  XOR U29478 ( .A(n30402), .B(n30405), .Z(n30403) );
  XOR U29479 ( .A(n30406), .B(n30407), .Z(n30390) );
  XOR U29480 ( .A(n30408), .B(n30409), .Z(n30407) );
  ANDN U29481 ( .B(n30410), .A(n30411), .Z(n30408) );
  XOR U29482 ( .A(n30412), .B(n30409), .Z(n30410) );
  IV U29483 ( .A(n30388), .Z(n30406) );
  XOR U29484 ( .A(n30413), .B(n30414), .Z(n30388) );
  ANDN U29485 ( .B(n30415), .A(n30416), .Z(n30413) );
  XOR U29486 ( .A(n30414), .B(n30417), .Z(n30415) );
  IV U29487 ( .A(n30396), .Z(n30400) );
  XOR U29488 ( .A(n30396), .B(n30378), .Z(n30398) );
  XOR U29489 ( .A(n30418), .B(n30419), .Z(n30378) );
  AND U29490 ( .A(n1786), .B(n30420), .Z(n30418) );
  XOR U29491 ( .A(n30421), .B(n30419), .Z(n30420) );
  NANDN U29492 ( .A(n30380), .B(n30382), .Z(n30396) );
  XOR U29493 ( .A(n30422), .B(n30423), .Z(n30382) );
  AND U29494 ( .A(n1786), .B(n30424), .Z(n30422) );
  XOR U29495 ( .A(n30423), .B(n30425), .Z(n30424) );
  XOR U29496 ( .A(n30426), .B(n30427), .Z(n1786) );
  AND U29497 ( .A(n30428), .B(n30429), .Z(n30426) );
  XNOR U29498 ( .A(n30427), .B(n30393), .Z(n30429) );
  XNOR U29499 ( .A(n30430), .B(n30431), .Z(n30393) );
  ANDN U29500 ( .B(n30432), .A(n30433), .Z(n30430) );
  XOR U29501 ( .A(n30431), .B(n30434), .Z(n30432) );
  XOR U29502 ( .A(n30427), .B(n30395), .Z(n30428) );
  XOR U29503 ( .A(n30435), .B(n30436), .Z(n30395) );
  AND U29504 ( .A(n1790), .B(n30437), .Z(n30435) );
  XOR U29505 ( .A(n30438), .B(n30436), .Z(n30437) );
  XNOR U29506 ( .A(n30439), .B(n30440), .Z(n30427) );
  NAND U29507 ( .A(n30441), .B(n30442), .Z(n30440) );
  XOR U29508 ( .A(n30443), .B(n30419), .Z(n30442) );
  XOR U29509 ( .A(n30433), .B(n30434), .Z(n30419) );
  XOR U29510 ( .A(n30444), .B(n30445), .Z(n30434) );
  ANDN U29511 ( .B(n30446), .A(n30447), .Z(n30444) );
  XOR U29512 ( .A(n30445), .B(n30448), .Z(n30446) );
  XOR U29513 ( .A(n30449), .B(n30450), .Z(n30433) );
  XOR U29514 ( .A(n30451), .B(n30452), .Z(n30450) );
  ANDN U29515 ( .B(n30453), .A(n30454), .Z(n30451) );
  XOR U29516 ( .A(n30455), .B(n30452), .Z(n30453) );
  IV U29517 ( .A(n30431), .Z(n30449) );
  XOR U29518 ( .A(n30456), .B(n30457), .Z(n30431) );
  ANDN U29519 ( .B(n30458), .A(n30459), .Z(n30456) );
  XOR U29520 ( .A(n30457), .B(n30460), .Z(n30458) );
  IV U29521 ( .A(n30439), .Z(n30443) );
  XOR U29522 ( .A(n30439), .B(n30421), .Z(n30441) );
  XOR U29523 ( .A(n30461), .B(n30462), .Z(n30421) );
  AND U29524 ( .A(n1790), .B(n30463), .Z(n30461) );
  XOR U29525 ( .A(n30464), .B(n30462), .Z(n30463) );
  NANDN U29526 ( .A(n30423), .B(n30425), .Z(n30439) );
  XOR U29527 ( .A(n30465), .B(n30466), .Z(n30425) );
  AND U29528 ( .A(n1790), .B(n30467), .Z(n30465) );
  XOR U29529 ( .A(n30466), .B(n30468), .Z(n30467) );
  XOR U29530 ( .A(n30469), .B(n30470), .Z(n1790) );
  AND U29531 ( .A(n30471), .B(n30472), .Z(n30469) );
  XNOR U29532 ( .A(n30470), .B(n30436), .Z(n30472) );
  XNOR U29533 ( .A(n30473), .B(n30474), .Z(n30436) );
  ANDN U29534 ( .B(n30475), .A(n30476), .Z(n30473) );
  XOR U29535 ( .A(n30474), .B(n30477), .Z(n30475) );
  XOR U29536 ( .A(n30470), .B(n30438), .Z(n30471) );
  XOR U29537 ( .A(n30478), .B(n30479), .Z(n30438) );
  AND U29538 ( .A(n1794), .B(n30480), .Z(n30478) );
  XOR U29539 ( .A(n30481), .B(n30479), .Z(n30480) );
  XNOR U29540 ( .A(n30482), .B(n30483), .Z(n30470) );
  NAND U29541 ( .A(n30484), .B(n30485), .Z(n30483) );
  XOR U29542 ( .A(n30486), .B(n30462), .Z(n30485) );
  XOR U29543 ( .A(n30476), .B(n30477), .Z(n30462) );
  XOR U29544 ( .A(n30487), .B(n30488), .Z(n30477) );
  ANDN U29545 ( .B(n30489), .A(n30490), .Z(n30487) );
  XOR U29546 ( .A(n30488), .B(n30491), .Z(n30489) );
  XOR U29547 ( .A(n30492), .B(n30493), .Z(n30476) );
  XOR U29548 ( .A(n30494), .B(n30495), .Z(n30493) );
  ANDN U29549 ( .B(n30496), .A(n30497), .Z(n30494) );
  XOR U29550 ( .A(n30498), .B(n30495), .Z(n30496) );
  IV U29551 ( .A(n30474), .Z(n30492) );
  XOR U29552 ( .A(n30499), .B(n30500), .Z(n30474) );
  ANDN U29553 ( .B(n30501), .A(n30502), .Z(n30499) );
  XOR U29554 ( .A(n30500), .B(n30503), .Z(n30501) );
  IV U29555 ( .A(n30482), .Z(n30486) );
  XOR U29556 ( .A(n30482), .B(n30464), .Z(n30484) );
  XOR U29557 ( .A(n30504), .B(n30505), .Z(n30464) );
  AND U29558 ( .A(n1794), .B(n30506), .Z(n30504) );
  XOR U29559 ( .A(n30507), .B(n30505), .Z(n30506) );
  NANDN U29560 ( .A(n30466), .B(n30468), .Z(n30482) );
  XOR U29561 ( .A(n30508), .B(n30509), .Z(n30468) );
  AND U29562 ( .A(n1794), .B(n30510), .Z(n30508) );
  XOR U29563 ( .A(n30509), .B(n30511), .Z(n30510) );
  XOR U29564 ( .A(n30512), .B(n30513), .Z(n1794) );
  AND U29565 ( .A(n30514), .B(n30515), .Z(n30512) );
  XNOR U29566 ( .A(n30513), .B(n30479), .Z(n30515) );
  XNOR U29567 ( .A(n30516), .B(n30517), .Z(n30479) );
  ANDN U29568 ( .B(n30518), .A(n30519), .Z(n30516) );
  XOR U29569 ( .A(n30517), .B(n30520), .Z(n30518) );
  XOR U29570 ( .A(n30513), .B(n30481), .Z(n30514) );
  XOR U29571 ( .A(n30521), .B(n30522), .Z(n30481) );
  AND U29572 ( .A(n1798), .B(n30523), .Z(n30521) );
  XOR U29573 ( .A(n30524), .B(n30522), .Z(n30523) );
  XNOR U29574 ( .A(n30525), .B(n30526), .Z(n30513) );
  NAND U29575 ( .A(n30527), .B(n30528), .Z(n30526) );
  XOR U29576 ( .A(n30529), .B(n30505), .Z(n30528) );
  XOR U29577 ( .A(n30519), .B(n30520), .Z(n30505) );
  XOR U29578 ( .A(n30530), .B(n30531), .Z(n30520) );
  ANDN U29579 ( .B(n30532), .A(n30533), .Z(n30530) );
  XOR U29580 ( .A(n30531), .B(n30534), .Z(n30532) );
  XOR U29581 ( .A(n30535), .B(n30536), .Z(n30519) );
  XOR U29582 ( .A(n30537), .B(n30538), .Z(n30536) );
  ANDN U29583 ( .B(n30539), .A(n30540), .Z(n30537) );
  XOR U29584 ( .A(n30541), .B(n30538), .Z(n30539) );
  IV U29585 ( .A(n30517), .Z(n30535) );
  XOR U29586 ( .A(n30542), .B(n30543), .Z(n30517) );
  ANDN U29587 ( .B(n30544), .A(n30545), .Z(n30542) );
  XOR U29588 ( .A(n30543), .B(n30546), .Z(n30544) );
  IV U29589 ( .A(n30525), .Z(n30529) );
  XOR U29590 ( .A(n30525), .B(n30507), .Z(n30527) );
  XOR U29591 ( .A(n30547), .B(n30548), .Z(n30507) );
  AND U29592 ( .A(n1798), .B(n30549), .Z(n30547) );
  XOR U29593 ( .A(n30550), .B(n30548), .Z(n30549) );
  NANDN U29594 ( .A(n30509), .B(n30511), .Z(n30525) );
  XOR U29595 ( .A(n30551), .B(n30552), .Z(n30511) );
  AND U29596 ( .A(n1798), .B(n30553), .Z(n30551) );
  XOR U29597 ( .A(n30552), .B(n30554), .Z(n30553) );
  XOR U29598 ( .A(n30555), .B(n30556), .Z(n1798) );
  AND U29599 ( .A(n30557), .B(n30558), .Z(n30555) );
  XNOR U29600 ( .A(n30556), .B(n30522), .Z(n30558) );
  XNOR U29601 ( .A(n30559), .B(n30560), .Z(n30522) );
  ANDN U29602 ( .B(n30561), .A(n30562), .Z(n30559) );
  XOR U29603 ( .A(n30560), .B(n30563), .Z(n30561) );
  XOR U29604 ( .A(n30556), .B(n30524), .Z(n30557) );
  XOR U29605 ( .A(n30564), .B(n30565), .Z(n30524) );
  AND U29606 ( .A(n1802), .B(n30566), .Z(n30564) );
  XOR U29607 ( .A(n30567), .B(n30565), .Z(n30566) );
  XNOR U29608 ( .A(n30568), .B(n30569), .Z(n30556) );
  NAND U29609 ( .A(n30570), .B(n30571), .Z(n30569) );
  XOR U29610 ( .A(n30572), .B(n30548), .Z(n30571) );
  XOR U29611 ( .A(n30562), .B(n30563), .Z(n30548) );
  XOR U29612 ( .A(n30573), .B(n30574), .Z(n30563) );
  ANDN U29613 ( .B(n30575), .A(n30576), .Z(n30573) );
  XOR U29614 ( .A(n30574), .B(n30577), .Z(n30575) );
  XOR U29615 ( .A(n30578), .B(n30579), .Z(n30562) );
  XOR U29616 ( .A(n30580), .B(n30581), .Z(n30579) );
  ANDN U29617 ( .B(n30582), .A(n30583), .Z(n30580) );
  XOR U29618 ( .A(n30584), .B(n30581), .Z(n30582) );
  IV U29619 ( .A(n30560), .Z(n30578) );
  XOR U29620 ( .A(n30585), .B(n30586), .Z(n30560) );
  ANDN U29621 ( .B(n30587), .A(n30588), .Z(n30585) );
  XOR U29622 ( .A(n30586), .B(n30589), .Z(n30587) );
  IV U29623 ( .A(n30568), .Z(n30572) );
  XOR U29624 ( .A(n30568), .B(n30550), .Z(n30570) );
  XOR U29625 ( .A(n30590), .B(n30591), .Z(n30550) );
  AND U29626 ( .A(n1802), .B(n30592), .Z(n30590) );
  XOR U29627 ( .A(n30593), .B(n30591), .Z(n30592) );
  NANDN U29628 ( .A(n30552), .B(n30554), .Z(n30568) );
  XOR U29629 ( .A(n30594), .B(n30595), .Z(n30554) );
  AND U29630 ( .A(n1802), .B(n30596), .Z(n30594) );
  XOR U29631 ( .A(n30595), .B(n30597), .Z(n30596) );
  XOR U29632 ( .A(n30598), .B(n30599), .Z(n1802) );
  AND U29633 ( .A(n30600), .B(n30601), .Z(n30598) );
  XNOR U29634 ( .A(n30599), .B(n30565), .Z(n30601) );
  XNOR U29635 ( .A(n30602), .B(n30603), .Z(n30565) );
  ANDN U29636 ( .B(n30604), .A(n30605), .Z(n30602) );
  XOR U29637 ( .A(n30603), .B(n30606), .Z(n30604) );
  XOR U29638 ( .A(n30599), .B(n30567), .Z(n30600) );
  XOR U29639 ( .A(n30607), .B(n30608), .Z(n30567) );
  AND U29640 ( .A(n1806), .B(n30609), .Z(n30607) );
  XOR U29641 ( .A(n30610), .B(n30608), .Z(n30609) );
  XNOR U29642 ( .A(n30611), .B(n30612), .Z(n30599) );
  NAND U29643 ( .A(n30613), .B(n30614), .Z(n30612) );
  XOR U29644 ( .A(n30615), .B(n30591), .Z(n30614) );
  XOR U29645 ( .A(n30605), .B(n30606), .Z(n30591) );
  XOR U29646 ( .A(n30616), .B(n30617), .Z(n30606) );
  ANDN U29647 ( .B(n30618), .A(n30619), .Z(n30616) );
  XOR U29648 ( .A(n30617), .B(n30620), .Z(n30618) );
  XOR U29649 ( .A(n30621), .B(n30622), .Z(n30605) );
  XOR U29650 ( .A(n30623), .B(n30624), .Z(n30622) );
  ANDN U29651 ( .B(n30625), .A(n30626), .Z(n30623) );
  XOR U29652 ( .A(n30627), .B(n30624), .Z(n30625) );
  IV U29653 ( .A(n30603), .Z(n30621) );
  XOR U29654 ( .A(n30628), .B(n30629), .Z(n30603) );
  ANDN U29655 ( .B(n30630), .A(n30631), .Z(n30628) );
  XOR U29656 ( .A(n30629), .B(n30632), .Z(n30630) );
  IV U29657 ( .A(n30611), .Z(n30615) );
  XOR U29658 ( .A(n30611), .B(n30593), .Z(n30613) );
  XOR U29659 ( .A(n30633), .B(n30634), .Z(n30593) );
  AND U29660 ( .A(n1806), .B(n30635), .Z(n30633) );
  XOR U29661 ( .A(n30636), .B(n30634), .Z(n30635) );
  NANDN U29662 ( .A(n30595), .B(n30597), .Z(n30611) );
  XOR U29663 ( .A(n30637), .B(n30638), .Z(n30597) );
  AND U29664 ( .A(n1806), .B(n30639), .Z(n30637) );
  XOR U29665 ( .A(n30638), .B(n30640), .Z(n30639) );
  XOR U29666 ( .A(n30641), .B(n30642), .Z(n1806) );
  AND U29667 ( .A(n30643), .B(n30644), .Z(n30641) );
  XNOR U29668 ( .A(n30642), .B(n30608), .Z(n30644) );
  XNOR U29669 ( .A(n30645), .B(n30646), .Z(n30608) );
  ANDN U29670 ( .B(n30647), .A(n30648), .Z(n30645) );
  XOR U29671 ( .A(n30646), .B(n30649), .Z(n30647) );
  XOR U29672 ( .A(n30642), .B(n30610), .Z(n30643) );
  XOR U29673 ( .A(n30650), .B(n30651), .Z(n30610) );
  AND U29674 ( .A(n1810), .B(n30652), .Z(n30650) );
  XOR U29675 ( .A(n30653), .B(n30651), .Z(n30652) );
  XNOR U29676 ( .A(n30654), .B(n30655), .Z(n30642) );
  NAND U29677 ( .A(n30656), .B(n30657), .Z(n30655) );
  XOR U29678 ( .A(n30658), .B(n30634), .Z(n30657) );
  XOR U29679 ( .A(n30648), .B(n30649), .Z(n30634) );
  XOR U29680 ( .A(n30659), .B(n30660), .Z(n30649) );
  ANDN U29681 ( .B(n30661), .A(n30662), .Z(n30659) );
  XOR U29682 ( .A(n30660), .B(n30663), .Z(n30661) );
  XOR U29683 ( .A(n30664), .B(n30665), .Z(n30648) );
  XOR U29684 ( .A(n30666), .B(n30667), .Z(n30665) );
  ANDN U29685 ( .B(n30668), .A(n30669), .Z(n30666) );
  XOR U29686 ( .A(n30670), .B(n30667), .Z(n30668) );
  IV U29687 ( .A(n30646), .Z(n30664) );
  XOR U29688 ( .A(n30671), .B(n30672), .Z(n30646) );
  ANDN U29689 ( .B(n30673), .A(n30674), .Z(n30671) );
  XOR U29690 ( .A(n30672), .B(n30675), .Z(n30673) );
  IV U29691 ( .A(n30654), .Z(n30658) );
  XOR U29692 ( .A(n30654), .B(n30636), .Z(n30656) );
  XOR U29693 ( .A(n30676), .B(n30677), .Z(n30636) );
  AND U29694 ( .A(n1810), .B(n30678), .Z(n30676) );
  XOR U29695 ( .A(n30679), .B(n30677), .Z(n30678) );
  NANDN U29696 ( .A(n30638), .B(n30640), .Z(n30654) );
  XOR U29697 ( .A(n30680), .B(n30681), .Z(n30640) );
  AND U29698 ( .A(n1810), .B(n30682), .Z(n30680) );
  XOR U29699 ( .A(n30681), .B(n30683), .Z(n30682) );
  XOR U29700 ( .A(n30684), .B(n30685), .Z(n1810) );
  AND U29701 ( .A(n30686), .B(n30687), .Z(n30684) );
  XNOR U29702 ( .A(n30685), .B(n30651), .Z(n30687) );
  XNOR U29703 ( .A(n30688), .B(n30689), .Z(n30651) );
  ANDN U29704 ( .B(n30690), .A(n30691), .Z(n30688) );
  XOR U29705 ( .A(n30689), .B(n30692), .Z(n30690) );
  XOR U29706 ( .A(n30685), .B(n30653), .Z(n30686) );
  XOR U29707 ( .A(n30693), .B(n30694), .Z(n30653) );
  AND U29708 ( .A(n1814), .B(n30695), .Z(n30693) );
  XOR U29709 ( .A(n30696), .B(n30694), .Z(n30695) );
  XNOR U29710 ( .A(n30697), .B(n30698), .Z(n30685) );
  NAND U29711 ( .A(n30699), .B(n30700), .Z(n30698) );
  XOR U29712 ( .A(n30701), .B(n30677), .Z(n30700) );
  XOR U29713 ( .A(n30691), .B(n30692), .Z(n30677) );
  XOR U29714 ( .A(n30702), .B(n30703), .Z(n30692) );
  ANDN U29715 ( .B(n30704), .A(n30705), .Z(n30702) );
  XOR U29716 ( .A(n30703), .B(n30706), .Z(n30704) );
  XOR U29717 ( .A(n30707), .B(n30708), .Z(n30691) );
  XOR U29718 ( .A(n30709), .B(n30710), .Z(n30708) );
  ANDN U29719 ( .B(n30711), .A(n30712), .Z(n30709) );
  XOR U29720 ( .A(n30713), .B(n30710), .Z(n30711) );
  IV U29721 ( .A(n30689), .Z(n30707) );
  XOR U29722 ( .A(n30714), .B(n30715), .Z(n30689) );
  ANDN U29723 ( .B(n30716), .A(n30717), .Z(n30714) );
  XOR U29724 ( .A(n30715), .B(n30718), .Z(n30716) );
  IV U29725 ( .A(n30697), .Z(n30701) );
  XOR U29726 ( .A(n30697), .B(n30679), .Z(n30699) );
  XOR U29727 ( .A(n30719), .B(n30720), .Z(n30679) );
  AND U29728 ( .A(n1814), .B(n30721), .Z(n30719) );
  XOR U29729 ( .A(n30722), .B(n30720), .Z(n30721) );
  NANDN U29730 ( .A(n30681), .B(n30683), .Z(n30697) );
  XOR U29731 ( .A(n30723), .B(n30724), .Z(n30683) );
  AND U29732 ( .A(n1814), .B(n30725), .Z(n30723) );
  XOR U29733 ( .A(n30724), .B(n30726), .Z(n30725) );
  XOR U29734 ( .A(n30727), .B(n30728), .Z(n1814) );
  AND U29735 ( .A(n30729), .B(n30730), .Z(n30727) );
  XNOR U29736 ( .A(n30728), .B(n30694), .Z(n30730) );
  XNOR U29737 ( .A(n30731), .B(n30732), .Z(n30694) );
  ANDN U29738 ( .B(n30733), .A(n30734), .Z(n30731) );
  XOR U29739 ( .A(n30732), .B(n30735), .Z(n30733) );
  XOR U29740 ( .A(n30728), .B(n30696), .Z(n30729) );
  XOR U29741 ( .A(n30736), .B(n30737), .Z(n30696) );
  AND U29742 ( .A(n1818), .B(n30738), .Z(n30736) );
  XOR U29743 ( .A(n30739), .B(n30737), .Z(n30738) );
  XNOR U29744 ( .A(n30740), .B(n30741), .Z(n30728) );
  NAND U29745 ( .A(n30742), .B(n30743), .Z(n30741) );
  XOR U29746 ( .A(n30744), .B(n30720), .Z(n30743) );
  XOR U29747 ( .A(n30734), .B(n30735), .Z(n30720) );
  XOR U29748 ( .A(n30745), .B(n30746), .Z(n30735) );
  ANDN U29749 ( .B(n30747), .A(n30748), .Z(n30745) );
  XOR U29750 ( .A(n30746), .B(n30749), .Z(n30747) );
  XOR U29751 ( .A(n30750), .B(n30751), .Z(n30734) );
  XOR U29752 ( .A(n30752), .B(n30753), .Z(n30751) );
  ANDN U29753 ( .B(n30754), .A(n30755), .Z(n30752) );
  XOR U29754 ( .A(n30756), .B(n30753), .Z(n30754) );
  IV U29755 ( .A(n30732), .Z(n30750) );
  XOR U29756 ( .A(n30757), .B(n30758), .Z(n30732) );
  ANDN U29757 ( .B(n30759), .A(n30760), .Z(n30757) );
  XOR U29758 ( .A(n30758), .B(n30761), .Z(n30759) );
  IV U29759 ( .A(n30740), .Z(n30744) );
  XOR U29760 ( .A(n30740), .B(n30722), .Z(n30742) );
  XOR U29761 ( .A(n30762), .B(n30763), .Z(n30722) );
  AND U29762 ( .A(n1818), .B(n30764), .Z(n30762) );
  XOR U29763 ( .A(n30765), .B(n30763), .Z(n30764) );
  NANDN U29764 ( .A(n30724), .B(n30726), .Z(n30740) );
  XOR U29765 ( .A(n30766), .B(n30767), .Z(n30726) );
  AND U29766 ( .A(n1818), .B(n30768), .Z(n30766) );
  XOR U29767 ( .A(n30767), .B(n30769), .Z(n30768) );
  XOR U29768 ( .A(n30770), .B(n30771), .Z(n1818) );
  AND U29769 ( .A(n30772), .B(n30773), .Z(n30770) );
  XNOR U29770 ( .A(n30771), .B(n30737), .Z(n30773) );
  XNOR U29771 ( .A(n30774), .B(n30775), .Z(n30737) );
  ANDN U29772 ( .B(n30776), .A(n30777), .Z(n30774) );
  XOR U29773 ( .A(n30775), .B(n30778), .Z(n30776) );
  XOR U29774 ( .A(n30771), .B(n30739), .Z(n30772) );
  XOR U29775 ( .A(n30779), .B(n30780), .Z(n30739) );
  AND U29776 ( .A(n1822), .B(n30781), .Z(n30779) );
  XOR U29777 ( .A(n30782), .B(n30780), .Z(n30781) );
  XNOR U29778 ( .A(n30783), .B(n30784), .Z(n30771) );
  NAND U29779 ( .A(n30785), .B(n30786), .Z(n30784) );
  XOR U29780 ( .A(n30787), .B(n30763), .Z(n30786) );
  XOR U29781 ( .A(n30777), .B(n30778), .Z(n30763) );
  XOR U29782 ( .A(n30788), .B(n30789), .Z(n30778) );
  ANDN U29783 ( .B(n30790), .A(n30791), .Z(n30788) );
  XOR U29784 ( .A(n30789), .B(n30792), .Z(n30790) );
  XOR U29785 ( .A(n30793), .B(n30794), .Z(n30777) );
  XOR U29786 ( .A(n30795), .B(n30796), .Z(n30794) );
  ANDN U29787 ( .B(n30797), .A(n30798), .Z(n30795) );
  XOR U29788 ( .A(n30799), .B(n30796), .Z(n30797) );
  IV U29789 ( .A(n30775), .Z(n30793) );
  XOR U29790 ( .A(n30800), .B(n30801), .Z(n30775) );
  ANDN U29791 ( .B(n30802), .A(n30803), .Z(n30800) );
  XOR U29792 ( .A(n30801), .B(n30804), .Z(n30802) );
  IV U29793 ( .A(n30783), .Z(n30787) );
  XOR U29794 ( .A(n30783), .B(n30765), .Z(n30785) );
  XOR U29795 ( .A(n30805), .B(n30806), .Z(n30765) );
  AND U29796 ( .A(n1822), .B(n30807), .Z(n30805) );
  XOR U29797 ( .A(n30808), .B(n30806), .Z(n30807) );
  NANDN U29798 ( .A(n30767), .B(n30769), .Z(n30783) );
  XOR U29799 ( .A(n30809), .B(n30810), .Z(n30769) );
  AND U29800 ( .A(n1822), .B(n30811), .Z(n30809) );
  XOR U29801 ( .A(n30810), .B(n30812), .Z(n30811) );
  XOR U29802 ( .A(n30813), .B(n30814), .Z(n1822) );
  AND U29803 ( .A(n30815), .B(n30816), .Z(n30813) );
  XNOR U29804 ( .A(n30814), .B(n30780), .Z(n30816) );
  XNOR U29805 ( .A(n30817), .B(n30818), .Z(n30780) );
  ANDN U29806 ( .B(n30819), .A(n30820), .Z(n30817) );
  XOR U29807 ( .A(n30818), .B(n30821), .Z(n30819) );
  XOR U29808 ( .A(n30814), .B(n30782), .Z(n30815) );
  XOR U29809 ( .A(n30822), .B(n30823), .Z(n30782) );
  AND U29810 ( .A(n1826), .B(n30824), .Z(n30822) );
  XOR U29811 ( .A(n30825), .B(n30823), .Z(n30824) );
  XNOR U29812 ( .A(n30826), .B(n30827), .Z(n30814) );
  NAND U29813 ( .A(n30828), .B(n30829), .Z(n30827) );
  XOR U29814 ( .A(n30830), .B(n30806), .Z(n30829) );
  XOR U29815 ( .A(n30820), .B(n30821), .Z(n30806) );
  XOR U29816 ( .A(n30831), .B(n30832), .Z(n30821) );
  ANDN U29817 ( .B(n30833), .A(n30834), .Z(n30831) );
  XOR U29818 ( .A(n30832), .B(n30835), .Z(n30833) );
  XOR U29819 ( .A(n30836), .B(n30837), .Z(n30820) );
  XOR U29820 ( .A(n30838), .B(n30839), .Z(n30837) );
  ANDN U29821 ( .B(n30840), .A(n30841), .Z(n30838) );
  XOR U29822 ( .A(n30842), .B(n30839), .Z(n30840) );
  IV U29823 ( .A(n30818), .Z(n30836) );
  XOR U29824 ( .A(n30843), .B(n30844), .Z(n30818) );
  ANDN U29825 ( .B(n30845), .A(n30846), .Z(n30843) );
  XOR U29826 ( .A(n30844), .B(n30847), .Z(n30845) );
  IV U29827 ( .A(n30826), .Z(n30830) );
  XOR U29828 ( .A(n30826), .B(n30808), .Z(n30828) );
  XOR U29829 ( .A(n30848), .B(n30849), .Z(n30808) );
  AND U29830 ( .A(n1826), .B(n30850), .Z(n30848) );
  XOR U29831 ( .A(n30851), .B(n30849), .Z(n30850) );
  NANDN U29832 ( .A(n30810), .B(n30812), .Z(n30826) );
  XOR U29833 ( .A(n30852), .B(n30853), .Z(n30812) );
  AND U29834 ( .A(n1826), .B(n30854), .Z(n30852) );
  XOR U29835 ( .A(n30853), .B(n30855), .Z(n30854) );
  XOR U29836 ( .A(n30856), .B(n30857), .Z(n1826) );
  AND U29837 ( .A(n30858), .B(n30859), .Z(n30856) );
  XNOR U29838 ( .A(n30857), .B(n30823), .Z(n30859) );
  XNOR U29839 ( .A(n30860), .B(n30861), .Z(n30823) );
  ANDN U29840 ( .B(n30862), .A(n30863), .Z(n30860) );
  XOR U29841 ( .A(n30861), .B(n30864), .Z(n30862) );
  XOR U29842 ( .A(n30857), .B(n30825), .Z(n30858) );
  XOR U29843 ( .A(n30865), .B(n30866), .Z(n30825) );
  AND U29844 ( .A(n1830), .B(n30867), .Z(n30865) );
  XOR U29845 ( .A(n30868), .B(n30866), .Z(n30867) );
  XNOR U29846 ( .A(n30869), .B(n30870), .Z(n30857) );
  NAND U29847 ( .A(n30871), .B(n30872), .Z(n30870) );
  XOR U29848 ( .A(n30873), .B(n30849), .Z(n30872) );
  XOR U29849 ( .A(n30863), .B(n30864), .Z(n30849) );
  XOR U29850 ( .A(n30874), .B(n30875), .Z(n30864) );
  ANDN U29851 ( .B(n30876), .A(n30877), .Z(n30874) );
  XOR U29852 ( .A(n30875), .B(n30878), .Z(n30876) );
  XOR U29853 ( .A(n30879), .B(n30880), .Z(n30863) );
  XOR U29854 ( .A(n30881), .B(n30882), .Z(n30880) );
  ANDN U29855 ( .B(n30883), .A(n30884), .Z(n30881) );
  XOR U29856 ( .A(n30885), .B(n30882), .Z(n30883) );
  IV U29857 ( .A(n30861), .Z(n30879) );
  XOR U29858 ( .A(n30886), .B(n30887), .Z(n30861) );
  ANDN U29859 ( .B(n30888), .A(n30889), .Z(n30886) );
  XOR U29860 ( .A(n30887), .B(n30890), .Z(n30888) );
  IV U29861 ( .A(n30869), .Z(n30873) );
  XOR U29862 ( .A(n30869), .B(n30851), .Z(n30871) );
  XOR U29863 ( .A(n30891), .B(n30892), .Z(n30851) );
  AND U29864 ( .A(n1830), .B(n30893), .Z(n30891) );
  XOR U29865 ( .A(n30894), .B(n30892), .Z(n30893) );
  NANDN U29866 ( .A(n30853), .B(n30855), .Z(n30869) );
  XOR U29867 ( .A(n30895), .B(n30896), .Z(n30855) );
  AND U29868 ( .A(n1830), .B(n30897), .Z(n30895) );
  XOR U29869 ( .A(n30896), .B(n30898), .Z(n30897) );
  XOR U29870 ( .A(n30899), .B(n30900), .Z(n1830) );
  AND U29871 ( .A(n30901), .B(n30902), .Z(n30899) );
  XNOR U29872 ( .A(n30900), .B(n30866), .Z(n30902) );
  XNOR U29873 ( .A(n30903), .B(n30904), .Z(n30866) );
  ANDN U29874 ( .B(n30905), .A(n30906), .Z(n30903) );
  XOR U29875 ( .A(n30904), .B(n30907), .Z(n30905) );
  XOR U29876 ( .A(n30900), .B(n30868), .Z(n30901) );
  XOR U29877 ( .A(n30908), .B(n30909), .Z(n30868) );
  AND U29878 ( .A(n1834), .B(n30910), .Z(n30908) );
  XOR U29879 ( .A(n30911), .B(n30909), .Z(n30910) );
  XNOR U29880 ( .A(n30912), .B(n30913), .Z(n30900) );
  NAND U29881 ( .A(n30914), .B(n30915), .Z(n30913) );
  XOR U29882 ( .A(n30916), .B(n30892), .Z(n30915) );
  XOR U29883 ( .A(n30906), .B(n30907), .Z(n30892) );
  XOR U29884 ( .A(n30917), .B(n30918), .Z(n30907) );
  ANDN U29885 ( .B(n30919), .A(n30920), .Z(n30917) );
  XOR U29886 ( .A(n30918), .B(n30921), .Z(n30919) );
  XOR U29887 ( .A(n30922), .B(n30923), .Z(n30906) );
  XOR U29888 ( .A(n30924), .B(n30925), .Z(n30923) );
  ANDN U29889 ( .B(n30926), .A(n30927), .Z(n30924) );
  XOR U29890 ( .A(n30928), .B(n30925), .Z(n30926) );
  IV U29891 ( .A(n30904), .Z(n30922) );
  XOR U29892 ( .A(n30929), .B(n30930), .Z(n30904) );
  ANDN U29893 ( .B(n30931), .A(n30932), .Z(n30929) );
  XOR U29894 ( .A(n30930), .B(n30933), .Z(n30931) );
  IV U29895 ( .A(n30912), .Z(n30916) );
  XOR U29896 ( .A(n30912), .B(n30894), .Z(n30914) );
  XOR U29897 ( .A(n30934), .B(n30935), .Z(n30894) );
  AND U29898 ( .A(n1834), .B(n30936), .Z(n30934) );
  XOR U29899 ( .A(n30937), .B(n30935), .Z(n30936) );
  NANDN U29900 ( .A(n30896), .B(n30898), .Z(n30912) );
  XOR U29901 ( .A(n30938), .B(n30939), .Z(n30898) );
  AND U29902 ( .A(n1834), .B(n30940), .Z(n30938) );
  XOR U29903 ( .A(n30939), .B(n30941), .Z(n30940) );
  XOR U29904 ( .A(n30942), .B(n30943), .Z(n1834) );
  AND U29905 ( .A(n30944), .B(n30945), .Z(n30942) );
  XNOR U29906 ( .A(n30943), .B(n30909), .Z(n30945) );
  XNOR U29907 ( .A(n30946), .B(n30947), .Z(n30909) );
  ANDN U29908 ( .B(n30948), .A(n30949), .Z(n30946) );
  XOR U29909 ( .A(n30947), .B(n30950), .Z(n30948) );
  XOR U29910 ( .A(n30943), .B(n30911), .Z(n30944) );
  XOR U29911 ( .A(n30951), .B(n30952), .Z(n30911) );
  AND U29912 ( .A(n1838), .B(n30953), .Z(n30951) );
  XOR U29913 ( .A(n30954), .B(n30952), .Z(n30953) );
  XNOR U29914 ( .A(n30955), .B(n30956), .Z(n30943) );
  NAND U29915 ( .A(n30957), .B(n30958), .Z(n30956) );
  XOR U29916 ( .A(n30959), .B(n30935), .Z(n30958) );
  XOR U29917 ( .A(n30949), .B(n30950), .Z(n30935) );
  XOR U29918 ( .A(n30960), .B(n30961), .Z(n30950) );
  ANDN U29919 ( .B(n30962), .A(n30963), .Z(n30960) );
  XOR U29920 ( .A(n30961), .B(n30964), .Z(n30962) );
  XOR U29921 ( .A(n30965), .B(n30966), .Z(n30949) );
  XOR U29922 ( .A(n30967), .B(n30968), .Z(n30966) );
  ANDN U29923 ( .B(n30969), .A(n30970), .Z(n30967) );
  XOR U29924 ( .A(n30971), .B(n30968), .Z(n30969) );
  IV U29925 ( .A(n30947), .Z(n30965) );
  XOR U29926 ( .A(n30972), .B(n30973), .Z(n30947) );
  ANDN U29927 ( .B(n30974), .A(n30975), .Z(n30972) );
  XOR U29928 ( .A(n30973), .B(n30976), .Z(n30974) );
  IV U29929 ( .A(n30955), .Z(n30959) );
  XOR U29930 ( .A(n30955), .B(n30937), .Z(n30957) );
  XOR U29931 ( .A(n30977), .B(n30978), .Z(n30937) );
  AND U29932 ( .A(n1838), .B(n30979), .Z(n30977) );
  XOR U29933 ( .A(n30980), .B(n30978), .Z(n30979) );
  NANDN U29934 ( .A(n30939), .B(n30941), .Z(n30955) );
  XOR U29935 ( .A(n30981), .B(n30982), .Z(n30941) );
  AND U29936 ( .A(n1838), .B(n30983), .Z(n30981) );
  XOR U29937 ( .A(n30982), .B(n30984), .Z(n30983) );
  XOR U29938 ( .A(n30985), .B(n30986), .Z(n1838) );
  AND U29939 ( .A(n30987), .B(n30988), .Z(n30985) );
  XNOR U29940 ( .A(n30986), .B(n30952), .Z(n30988) );
  XNOR U29941 ( .A(n30989), .B(n30990), .Z(n30952) );
  ANDN U29942 ( .B(n30991), .A(n30992), .Z(n30989) );
  XOR U29943 ( .A(n30990), .B(n30993), .Z(n30991) );
  XOR U29944 ( .A(n30986), .B(n30954), .Z(n30987) );
  XOR U29945 ( .A(n30994), .B(n30995), .Z(n30954) );
  AND U29946 ( .A(n1842), .B(n30996), .Z(n30994) );
  XOR U29947 ( .A(n30997), .B(n30995), .Z(n30996) );
  XNOR U29948 ( .A(n30998), .B(n30999), .Z(n30986) );
  NAND U29949 ( .A(n31000), .B(n31001), .Z(n30999) );
  XOR U29950 ( .A(n31002), .B(n30978), .Z(n31001) );
  XOR U29951 ( .A(n30992), .B(n30993), .Z(n30978) );
  XOR U29952 ( .A(n31003), .B(n31004), .Z(n30993) );
  ANDN U29953 ( .B(n31005), .A(n31006), .Z(n31003) );
  XOR U29954 ( .A(n31004), .B(n31007), .Z(n31005) );
  XOR U29955 ( .A(n31008), .B(n31009), .Z(n30992) );
  XOR U29956 ( .A(n31010), .B(n31011), .Z(n31009) );
  ANDN U29957 ( .B(n31012), .A(n31013), .Z(n31010) );
  XOR U29958 ( .A(n31014), .B(n31011), .Z(n31012) );
  IV U29959 ( .A(n30990), .Z(n31008) );
  XOR U29960 ( .A(n31015), .B(n31016), .Z(n30990) );
  ANDN U29961 ( .B(n31017), .A(n31018), .Z(n31015) );
  XOR U29962 ( .A(n31016), .B(n31019), .Z(n31017) );
  IV U29963 ( .A(n30998), .Z(n31002) );
  XOR U29964 ( .A(n30998), .B(n30980), .Z(n31000) );
  XOR U29965 ( .A(n31020), .B(n31021), .Z(n30980) );
  AND U29966 ( .A(n1842), .B(n31022), .Z(n31020) );
  XOR U29967 ( .A(n31023), .B(n31021), .Z(n31022) );
  NANDN U29968 ( .A(n30982), .B(n30984), .Z(n30998) );
  XOR U29969 ( .A(n31024), .B(n31025), .Z(n30984) );
  AND U29970 ( .A(n1842), .B(n31026), .Z(n31024) );
  XOR U29971 ( .A(n31025), .B(n31027), .Z(n31026) );
  XOR U29972 ( .A(n31028), .B(n31029), .Z(n1842) );
  AND U29973 ( .A(n31030), .B(n31031), .Z(n31028) );
  XNOR U29974 ( .A(n31029), .B(n30995), .Z(n31031) );
  XNOR U29975 ( .A(n31032), .B(n31033), .Z(n30995) );
  ANDN U29976 ( .B(n31034), .A(n31035), .Z(n31032) );
  XOR U29977 ( .A(n31033), .B(n31036), .Z(n31034) );
  XOR U29978 ( .A(n31029), .B(n30997), .Z(n31030) );
  XOR U29979 ( .A(n31037), .B(n31038), .Z(n30997) );
  AND U29980 ( .A(n1846), .B(n31039), .Z(n31037) );
  XOR U29981 ( .A(n31040), .B(n31038), .Z(n31039) );
  XNOR U29982 ( .A(n31041), .B(n31042), .Z(n31029) );
  NAND U29983 ( .A(n31043), .B(n31044), .Z(n31042) );
  XOR U29984 ( .A(n31045), .B(n31021), .Z(n31044) );
  XOR U29985 ( .A(n31035), .B(n31036), .Z(n31021) );
  XOR U29986 ( .A(n31046), .B(n31047), .Z(n31036) );
  ANDN U29987 ( .B(n31048), .A(n31049), .Z(n31046) );
  XOR U29988 ( .A(n31047), .B(n31050), .Z(n31048) );
  XOR U29989 ( .A(n31051), .B(n31052), .Z(n31035) );
  XOR U29990 ( .A(n31053), .B(n31054), .Z(n31052) );
  ANDN U29991 ( .B(n31055), .A(n31056), .Z(n31053) );
  XOR U29992 ( .A(n31057), .B(n31054), .Z(n31055) );
  IV U29993 ( .A(n31033), .Z(n31051) );
  XOR U29994 ( .A(n31058), .B(n31059), .Z(n31033) );
  ANDN U29995 ( .B(n31060), .A(n31061), .Z(n31058) );
  XOR U29996 ( .A(n31059), .B(n31062), .Z(n31060) );
  IV U29997 ( .A(n31041), .Z(n31045) );
  XOR U29998 ( .A(n31041), .B(n31023), .Z(n31043) );
  XOR U29999 ( .A(n31063), .B(n31064), .Z(n31023) );
  AND U30000 ( .A(n1846), .B(n31065), .Z(n31063) );
  XOR U30001 ( .A(n31066), .B(n31064), .Z(n31065) );
  NANDN U30002 ( .A(n31025), .B(n31027), .Z(n31041) );
  XOR U30003 ( .A(n31067), .B(n31068), .Z(n31027) );
  AND U30004 ( .A(n1846), .B(n31069), .Z(n31067) );
  XOR U30005 ( .A(n31068), .B(n31070), .Z(n31069) );
  XOR U30006 ( .A(n31071), .B(n31072), .Z(n1846) );
  AND U30007 ( .A(n31073), .B(n31074), .Z(n31071) );
  XNOR U30008 ( .A(n31072), .B(n31038), .Z(n31074) );
  XNOR U30009 ( .A(n31075), .B(n31076), .Z(n31038) );
  ANDN U30010 ( .B(n31077), .A(n31078), .Z(n31075) );
  XOR U30011 ( .A(n31076), .B(n31079), .Z(n31077) );
  XOR U30012 ( .A(n31072), .B(n31040), .Z(n31073) );
  XOR U30013 ( .A(n31080), .B(n31081), .Z(n31040) );
  AND U30014 ( .A(n1850), .B(n31082), .Z(n31080) );
  XOR U30015 ( .A(n31083), .B(n31081), .Z(n31082) );
  XNOR U30016 ( .A(n31084), .B(n31085), .Z(n31072) );
  NAND U30017 ( .A(n31086), .B(n31087), .Z(n31085) );
  XOR U30018 ( .A(n31088), .B(n31064), .Z(n31087) );
  XOR U30019 ( .A(n31078), .B(n31079), .Z(n31064) );
  XOR U30020 ( .A(n31089), .B(n31090), .Z(n31079) );
  ANDN U30021 ( .B(n31091), .A(n31092), .Z(n31089) );
  XOR U30022 ( .A(n31090), .B(n31093), .Z(n31091) );
  XOR U30023 ( .A(n31094), .B(n31095), .Z(n31078) );
  XOR U30024 ( .A(n31096), .B(n31097), .Z(n31095) );
  ANDN U30025 ( .B(n31098), .A(n31099), .Z(n31096) );
  XOR U30026 ( .A(n31100), .B(n31097), .Z(n31098) );
  IV U30027 ( .A(n31076), .Z(n31094) );
  XOR U30028 ( .A(n31101), .B(n31102), .Z(n31076) );
  ANDN U30029 ( .B(n31103), .A(n31104), .Z(n31101) );
  XOR U30030 ( .A(n31102), .B(n31105), .Z(n31103) );
  IV U30031 ( .A(n31084), .Z(n31088) );
  XOR U30032 ( .A(n31084), .B(n31066), .Z(n31086) );
  XOR U30033 ( .A(n31106), .B(n31107), .Z(n31066) );
  AND U30034 ( .A(n1850), .B(n31108), .Z(n31106) );
  XOR U30035 ( .A(n31109), .B(n31107), .Z(n31108) );
  NANDN U30036 ( .A(n31068), .B(n31070), .Z(n31084) );
  XOR U30037 ( .A(n31110), .B(n31111), .Z(n31070) );
  AND U30038 ( .A(n1850), .B(n31112), .Z(n31110) );
  XOR U30039 ( .A(n31111), .B(n31113), .Z(n31112) );
  XOR U30040 ( .A(n31114), .B(n31115), .Z(n1850) );
  AND U30041 ( .A(n31116), .B(n31117), .Z(n31114) );
  XNOR U30042 ( .A(n31115), .B(n31081), .Z(n31117) );
  XNOR U30043 ( .A(n31118), .B(n31119), .Z(n31081) );
  ANDN U30044 ( .B(n31120), .A(n31121), .Z(n31118) );
  XOR U30045 ( .A(n31119), .B(n31122), .Z(n31120) );
  XOR U30046 ( .A(n31115), .B(n31083), .Z(n31116) );
  XOR U30047 ( .A(n31123), .B(n31124), .Z(n31083) );
  AND U30048 ( .A(n1854), .B(n31125), .Z(n31123) );
  XOR U30049 ( .A(n31126), .B(n31124), .Z(n31125) );
  XNOR U30050 ( .A(n31127), .B(n31128), .Z(n31115) );
  NAND U30051 ( .A(n31129), .B(n31130), .Z(n31128) );
  XOR U30052 ( .A(n31131), .B(n31107), .Z(n31130) );
  XOR U30053 ( .A(n31121), .B(n31122), .Z(n31107) );
  XOR U30054 ( .A(n31132), .B(n31133), .Z(n31122) );
  ANDN U30055 ( .B(n31134), .A(n31135), .Z(n31132) );
  XOR U30056 ( .A(n31133), .B(n31136), .Z(n31134) );
  XOR U30057 ( .A(n31137), .B(n31138), .Z(n31121) );
  XOR U30058 ( .A(n31139), .B(n31140), .Z(n31138) );
  ANDN U30059 ( .B(n31141), .A(n31142), .Z(n31139) );
  XOR U30060 ( .A(n31143), .B(n31140), .Z(n31141) );
  IV U30061 ( .A(n31119), .Z(n31137) );
  XOR U30062 ( .A(n31144), .B(n31145), .Z(n31119) );
  ANDN U30063 ( .B(n31146), .A(n31147), .Z(n31144) );
  XOR U30064 ( .A(n31145), .B(n31148), .Z(n31146) );
  IV U30065 ( .A(n31127), .Z(n31131) );
  XOR U30066 ( .A(n31127), .B(n31109), .Z(n31129) );
  XOR U30067 ( .A(n31149), .B(n31150), .Z(n31109) );
  AND U30068 ( .A(n1854), .B(n31151), .Z(n31149) );
  XOR U30069 ( .A(n31152), .B(n31150), .Z(n31151) );
  NANDN U30070 ( .A(n31111), .B(n31113), .Z(n31127) );
  XOR U30071 ( .A(n31153), .B(n31154), .Z(n31113) );
  AND U30072 ( .A(n1854), .B(n31155), .Z(n31153) );
  XOR U30073 ( .A(n31154), .B(n31156), .Z(n31155) );
  XOR U30074 ( .A(n31157), .B(n31158), .Z(n1854) );
  AND U30075 ( .A(n31159), .B(n31160), .Z(n31157) );
  XNOR U30076 ( .A(n31158), .B(n31124), .Z(n31160) );
  XNOR U30077 ( .A(n31161), .B(n31162), .Z(n31124) );
  ANDN U30078 ( .B(n31163), .A(n31164), .Z(n31161) );
  XOR U30079 ( .A(n31162), .B(n31165), .Z(n31163) );
  XOR U30080 ( .A(n31158), .B(n31126), .Z(n31159) );
  XOR U30081 ( .A(n31166), .B(n31167), .Z(n31126) );
  AND U30082 ( .A(n1858), .B(n31168), .Z(n31166) );
  XOR U30083 ( .A(n31169), .B(n31167), .Z(n31168) );
  XNOR U30084 ( .A(n31170), .B(n31171), .Z(n31158) );
  NAND U30085 ( .A(n31172), .B(n31173), .Z(n31171) );
  XOR U30086 ( .A(n31174), .B(n31150), .Z(n31173) );
  XOR U30087 ( .A(n31164), .B(n31165), .Z(n31150) );
  XOR U30088 ( .A(n31175), .B(n31176), .Z(n31165) );
  ANDN U30089 ( .B(n31177), .A(n31178), .Z(n31175) );
  XOR U30090 ( .A(n31176), .B(n31179), .Z(n31177) );
  XOR U30091 ( .A(n31180), .B(n31181), .Z(n31164) );
  XOR U30092 ( .A(n31182), .B(n31183), .Z(n31181) );
  ANDN U30093 ( .B(n31184), .A(n31185), .Z(n31182) );
  XOR U30094 ( .A(n31186), .B(n31183), .Z(n31184) );
  IV U30095 ( .A(n31162), .Z(n31180) );
  XOR U30096 ( .A(n31187), .B(n31188), .Z(n31162) );
  ANDN U30097 ( .B(n31189), .A(n31190), .Z(n31187) );
  XOR U30098 ( .A(n31188), .B(n31191), .Z(n31189) );
  IV U30099 ( .A(n31170), .Z(n31174) );
  XOR U30100 ( .A(n31170), .B(n31152), .Z(n31172) );
  XOR U30101 ( .A(n31192), .B(n31193), .Z(n31152) );
  AND U30102 ( .A(n1858), .B(n31194), .Z(n31192) );
  XOR U30103 ( .A(n31195), .B(n31193), .Z(n31194) );
  NANDN U30104 ( .A(n31154), .B(n31156), .Z(n31170) );
  XOR U30105 ( .A(n31196), .B(n31197), .Z(n31156) );
  AND U30106 ( .A(n1858), .B(n31198), .Z(n31196) );
  XOR U30107 ( .A(n31197), .B(n31199), .Z(n31198) );
  XOR U30108 ( .A(n31200), .B(n31201), .Z(n1858) );
  AND U30109 ( .A(n31202), .B(n31203), .Z(n31200) );
  XNOR U30110 ( .A(n31201), .B(n31167), .Z(n31203) );
  XNOR U30111 ( .A(n31204), .B(n31205), .Z(n31167) );
  ANDN U30112 ( .B(n31206), .A(n31207), .Z(n31204) );
  XOR U30113 ( .A(n31205), .B(n31208), .Z(n31206) );
  XOR U30114 ( .A(n31201), .B(n31169), .Z(n31202) );
  XOR U30115 ( .A(n31209), .B(n31210), .Z(n31169) );
  AND U30116 ( .A(n1862), .B(n31211), .Z(n31209) );
  XOR U30117 ( .A(n31212), .B(n31210), .Z(n31211) );
  XNOR U30118 ( .A(n31213), .B(n31214), .Z(n31201) );
  NAND U30119 ( .A(n31215), .B(n31216), .Z(n31214) );
  XOR U30120 ( .A(n31217), .B(n31193), .Z(n31216) );
  XOR U30121 ( .A(n31207), .B(n31208), .Z(n31193) );
  XOR U30122 ( .A(n31218), .B(n31219), .Z(n31208) );
  ANDN U30123 ( .B(n31220), .A(n31221), .Z(n31218) );
  XOR U30124 ( .A(n31219), .B(n31222), .Z(n31220) );
  XOR U30125 ( .A(n31223), .B(n31224), .Z(n31207) );
  XOR U30126 ( .A(n31225), .B(n31226), .Z(n31224) );
  ANDN U30127 ( .B(n31227), .A(n31228), .Z(n31225) );
  XOR U30128 ( .A(n31229), .B(n31226), .Z(n31227) );
  IV U30129 ( .A(n31205), .Z(n31223) );
  XOR U30130 ( .A(n31230), .B(n31231), .Z(n31205) );
  ANDN U30131 ( .B(n31232), .A(n31233), .Z(n31230) );
  XOR U30132 ( .A(n31231), .B(n31234), .Z(n31232) );
  IV U30133 ( .A(n31213), .Z(n31217) );
  XOR U30134 ( .A(n31213), .B(n31195), .Z(n31215) );
  XOR U30135 ( .A(n31235), .B(n31236), .Z(n31195) );
  AND U30136 ( .A(n1862), .B(n31237), .Z(n31235) );
  XOR U30137 ( .A(n31238), .B(n31236), .Z(n31237) );
  NANDN U30138 ( .A(n31197), .B(n31199), .Z(n31213) );
  XOR U30139 ( .A(n31239), .B(n31240), .Z(n31199) );
  AND U30140 ( .A(n1862), .B(n31241), .Z(n31239) );
  XOR U30141 ( .A(n31240), .B(n31242), .Z(n31241) );
  XOR U30142 ( .A(n31243), .B(n31244), .Z(n1862) );
  AND U30143 ( .A(n31245), .B(n31246), .Z(n31243) );
  XNOR U30144 ( .A(n31244), .B(n31210), .Z(n31246) );
  XNOR U30145 ( .A(n31247), .B(n31248), .Z(n31210) );
  ANDN U30146 ( .B(n31249), .A(n31250), .Z(n31247) );
  XOR U30147 ( .A(n31248), .B(n31251), .Z(n31249) );
  XOR U30148 ( .A(n31244), .B(n31212), .Z(n31245) );
  XOR U30149 ( .A(n31252), .B(n31253), .Z(n31212) );
  AND U30150 ( .A(n1866), .B(n31254), .Z(n31252) );
  XOR U30151 ( .A(n31255), .B(n31253), .Z(n31254) );
  XNOR U30152 ( .A(n31256), .B(n31257), .Z(n31244) );
  NAND U30153 ( .A(n31258), .B(n31259), .Z(n31257) );
  XOR U30154 ( .A(n31260), .B(n31236), .Z(n31259) );
  XOR U30155 ( .A(n31250), .B(n31251), .Z(n31236) );
  XOR U30156 ( .A(n31261), .B(n31262), .Z(n31251) );
  ANDN U30157 ( .B(n31263), .A(n31264), .Z(n31261) );
  XOR U30158 ( .A(n31262), .B(n31265), .Z(n31263) );
  XOR U30159 ( .A(n31266), .B(n31267), .Z(n31250) );
  XOR U30160 ( .A(n31268), .B(n31269), .Z(n31267) );
  ANDN U30161 ( .B(n31270), .A(n31271), .Z(n31268) );
  XOR U30162 ( .A(n31272), .B(n31269), .Z(n31270) );
  IV U30163 ( .A(n31248), .Z(n31266) );
  XOR U30164 ( .A(n31273), .B(n31274), .Z(n31248) );
  ANDN U30165 ( .B(n31275), .A(n31276), .Z(n31273) );
  XOR U30166 ( .A(n31274), .B(n31277), .Z(n31275) );
  IV U30167 ( .A(n31256), .Z(n31260) );
  XOR U30168 ( .A(n31256), .B(n31238), .Z(n31258) );
  XOR U30169 ( .A(n31278), .B(n31279), .Z(n31238) );
  AND U30170 ( .A(n1866), .B(n31280), .Z(n31278) );
  XOR U30171 ( .A(n31281), .B(n31279), .Z(n31280) );
  NANDN U30172 ( .A(n31240), .B(n31242), .Z(n31256) );
  XOR U30173 ( .A(n31282), .B(n31283), .Z(n31242) );
  AND U30174 ( .A(n1866), .B(n31284), .Z(n31282) );
  XOR U30175 ( .A(n31283), .B(n31285), .Z(n31284) );
  XOR U30176 ( .A(n31286), .B(n31287), .Z(n1866) );
  AND U30177 ( .A(n31288), .B(n31289), .Z(n31286) );
  XNOR U30178 ( .A(n31287), .B(n31253), .Z(n31289) );
  XNOR U30179 ( .A(n31290), .B(n31291), .Z(n31253) );
  ANDN U30180 ( .B(n31292), .A(n31293), .Z(n31290) );
  XOR U30181 ( .A(n31291), .B(n31294), .Z(n31292) );
  XOR U30182 ( .A(n31287), .B(n31255), .Z(n31288) );
  XOR U30183 ( .A(n31295), .B(n31296), .Z(n31255) );
  AND U30184 ( .A(n1870), .B(n31297), .Z(n31295) );
  XOR U30185 ( .A(n31298), .B(n31296), .Z(n31297) );
  XNOR U30186 ( .A(n31299), .B(n31300), .Z(n31287) );
  NAND U30187 ( .A(n31301), .B(n31302), .Z(n31300) );
  XOR U30188 ( .A(n31303), .B(n31279), .Z(n31302) );
  XOR U30189 ( .A(n31293), .B(n31294), .Z(n31279) );
  XOR U30190 ( .A(n31304), .B(n31305), .Z(n31294) );
  ANDN U30191 ( .B(n31306), .A(n31307), .Z(n31304) );
  XOR U30192 ( .A(n31305), .B(n31308), .Z(n31306) );
  XOR U30193 ( .A(n31309), .B(n31310), .Z(n31293) );
  XOR U30194 ( .A(n31311), .B(n31312), .Z(n31310) );
  ANDN U30195 ( .B(n31313), .A(n31314), .Z(n31311) );
  XOR U30196 ( .A(n31315), .B(n31312), .Z(n31313) );
  IV U30197 ( .A(n31291), .Z(n31309) );
  XOR U30198 ( .A(n31316), .B(n31317), .Z(n31291) );
  ANDN U30199 ( .B(n31318), .A(n31319), .Z(n31316) );
  XOR U30200 ( .A(n31317), .B(n31320), .Z(n31318) );
  IV U30201 ( .A(n31299), .Z(n31303) );
  XOR U30202 ( .A(n31299), .B(n31281), .Z(n31301) );
  XOR U30203 ( .A(n31321), .B(n31322), .Z(n31281) );
  AND U30204 ( .A(n1870), .B(n31323), .Z(n31321) );
  XOR U30205 ( .A(n31324), .B(n31322), .Z(n31323) );
  NANDN U30206 ( .A(n31283), .B(n31285), .Z(n31299) );
  XOR U30207 ( .A(n31325), .B(n31326), .Z(n31285) );
  AND U30208 ( .A(n1870), .B(n31327), .Z(n31325) );
  XOR U30209 ( .A(n31326), .B(n31328), .Z(n31327) );
  XOR U30210 ( .A(n31329), .B(n31330), .Z(n1870) );
  AND U30211 ( .A(n31331), .B(n31332), .Z(n31329) );
  XNOR U30212 ( .A(n31330), .B(n31296), .Z(n31332) );
  XNOR U30213 ( .A(n31333), .B(n31334), .Z(n31296) );
  ANDN U30214 ( .B(n31335), .A(n31336), .Z(n31333) );
  XOR U30215 ( .A(n31334), .B(n31337), .Z(n31335) );
  XOR U30216 ( .A(n31330), .B(n31298), .Z(n31331) );
  XOR U30217 ( .A(n31338), .B(n31339), .Z(n31298) );
  AND U30218 ( .A(n1874), .B(n31340), .Z(n31338) );
  XOR U30219 ( .A(n31341), .B(n31339), .Z(n31340) );
  XNOR U30220 ( .A(n31342), .B(n31343), .Z(n31330) );
  NAND U30221 ( .A(n31344), .B(n31345), .Z(n31343) );
  XOR U30222 ( .A(n31346), .B(n31322), .Z(n31345) );
  XOR U30223 ( .A(n31336), .B(n31337), .Z(n31322) );
  XOR U30224 ( .A(n31347), .B(n31348), .Z(n31337) );
  ANDN U30225 ( .B(n31349), .A(n31350), .Z(n31347) );
  XOR U30226 ( .A(n31348), .B(n31351), .Z(n31349) );
  XOR U30227 ( .A(n31352), .B(n31353), .Z(n31336) );
  XOR U30228 ( .A(n31354), .B(n31355), .Z(n31353) );
  ANDN U30229 ( .B(n31356), .A(n31357), .Z(n31354) );
  XOR U30230 ( .A(n31358), .B(n31355), .Z(n31356) );
  IV U30231 ( .A(n31334), .Z(n31352) );
  XOR U30232 ( .A(n31359), .B(n31360), .Z(n31334) );
  ANDN U30233 ( .B(n31361), .A(n31362), .Z(n31359) );
  XOR U30234 ( .A(n31360), .B(n31363), .Z(n31361) );
  IV U30235 ( .A(n31342), .Z(n31346) );
  XOR U30236 ( .A(n31342), .B(n31324), .Z(n31344) );
  XOR U30237 ( .A(n31364), .B(n31365), .Z(n31324) );
  AND U30238 ( .A(n1874), .B(n31366), .Z(n31364) );
  XOR U30239 ( .A(n31367), .B(n31365), .Z(n31366) );
  NANDN U30240 ( .A(n31326), .B(n31328), .Z(n31342) );
  XOR U30241 ( .A(n31368), .B(n31369), .Z(n31328) );
  AND U30242 ( .A(n1874), .B(n31370), .Z(n31368) );
  XOR U30243 ( .A(n31369), .B(n31371), .Z(n31370) );
  XOR U30244 ( .A(n31372), .B(n31373), .Z(n1874) );
  AND U30245 ( .A(n31374), .B(n31375), .Z(n31372) );
  XNOR U30246 ( .A(n31373), .B(n31339), .Z(n31375) );
  XNOR U30247 ( .A(n31376), .B(n31377), .Z(n31339) );
  ANDN U30248 ( .B(n31378), .A(n31379), .Z(n31376) );
  XOR U30249 ( .A(n31377), .B(n31380), .Z(n31378) );
  XOR U30250 ( .A(n31373), .B(n31341), .Z(n31374) );
  XOR U30251 ( .A(n31381), .B(n31382), .Z(n31341) );
  AND U30252 ( .A(n1878), .B(n31383), .Z(n31381) );
  XOR U30253 ( .A(n31384), .B(n31382), .Z(n31383) );
  XNOR U30254 ( .A(n31385), .B(n31386), .Z(n31373) );
  NAND U30255 ( .A(n31387), .B(n31388), .Z(n31386) );
  XOR U30256 ( .A(n31389), .B(n31365), .Z(n31388) );
  XOR U30257 ( .A(n31379), .B(n31380), .Z(n31365) );
  XOR U30258 ( .A(n31390), .B(n31391), .Z(n31380) );
  ANDN U30259 ( .B(n31392), .A(n31393), .Z(n31390) );
  XOR U30260 ( .A(n31391), .B(n31394), .Z(n31392) );
  XOR U30261 ( .A(n31395), .B(n31396), .Z(n31379) );
  XOR U30262 ( .A(n31397), .B(n31398), .Z(n31396) );
  ANDN U30263 ( .B(n31399), .A(n31400), .Z(n31397) );
  XOR U30264 ( .A(n31401), .B(n31398), .Z(n31399) );
  IV U30265 ( .A(n31377), .Z(n31395) );
  XOR U30266 ( .A(n31402), .B(n31403), .Z(n31377) );
  ANDN U30267 ( .B(n31404), .A(n31405), .Z(n31402) );
  XOR U30268 ( .A(n31403), .B(n31406), .Z(n31404) );
  IV U30269 ( .A(n31385), .Z(n31389) );
  XOR U30270 ( .A(n31385), .B(n31367), .Z(n31387) );
  XOR U30271 ( .A(n31407), .B(n31408), .Z(n31367) );
  AND U30272 ( .A(n1878), .B(n31409), .Z(n31407) );
  XOR U30273 ( .A(n31410), .B(n31408), .Z(n31409) );
  NANDN U30274 ( .A(n31369), .B(n31371), .Z(n31385) );
  XOR U30275 ( .A(n31411), .B(n31412), .Z(n31371) );
  AND U30276 ( .A(n1878), .B(n31413), .Z(n31411) );
  XOR U30277 ( .A(n31412), .B(n31414), .Z(n31413) );
  XOR U30278 ( .A(n31415), .B(n31416), .Z(n1878) );
  AND U30279 ( .A(n31417), .B(n31418), .Z(n31415) );
  XNOR U30280 ( .A(n31416), .B(n31382), .Z(n31418) );
  XNOR U30281 ( .A(n31419), .B(n31420), .Z(n31382) );
  ANDN U30282 ( .B(n31421), .A(n31422), .Z(n31419) );
  XOR U30283 ( .A(n31420), .B(n31423), .Z(n31421) );
  XOR U30284 ( .A(n31416), .B(n31384), .Z(n31417) );
  XOR U30285 ( .A(n31424), .B(n31425), .Z(n31384) );
  AND U30286 ( .A(n1882), .B(n31426), .Z(n31424) );
  XOR U30287 ( .A(n31427), .B(n31425), .Z(n31426) );
  XNOR U30288 ( .A(n31428), .B(n31429), .Z(n31416) );
  NAND U30289 ( .A(n31430), .B(n31431), .Z(n31429) );
  XOR U30290 ( .A(n31432), .B(n31408), .Z(n31431) );
  XOR U30291 ( .A(n31422), .B(n31423), .Z(n31408) );
  XOR U30292 ( .A(n31433), .B(n31434), .Z(n31423) );
  ANDN U30293 ( .B(n31435), .A(n31436), .Z(n31433) );
  XOR U30294 ( .A(n31434), .B(n31437), .Z(n31435) );
  XOR U30295 ( .A(n31438), .B(n31439), .Z(n31422) );
  XOR U30296 ( .A(n31440), .B(n31441), .Z(n31439) );
  ANDN U30297 ( .B(n31442), .A(n31443), .Z(n31440) );
  XOR U30298 ( .A(n31444), .B(n31441), .Z(n31442) );
  IV U30299 ( .A(n31420), .Z(n31438) );
  XOR U30300 ( .A(n31445), .B(n31446), .Z(n31420) );
  ANDN U30301 ( .B(n31447), .A(n31448), .Z(n31445) );
  XOR U30302 ( .A(n31446), .B(n31449), .Z(n31447) );
  IV U30303 ( .A(n31428), .Z(n31432) );
  XOR U30304 ( .A(n31428), .B(n31410), .Z(n31430) );
  XOR U30305 ( .A(n31450), .B(n31451), .Z(n31410) );
  AND U30306 ( .A(n1882), .B(n31452), .Z(n31450) );
  XOR U30307 ( .A(n31453), .B(n31451), .Z(n31452) );
  NANDN U30308 ( .A(n31412), .B(n31414), .Z(n31428) );
  XOR U30309 ( .A(n31454), .B(n31455), .Z(n31414) );
  AND U30310 ( .A(n1882), .B(n31456), .Z(n31454) );
  XOR U30311 ( .A(n31455), .B(n31457), .Z(n31456) );
  XOR U30312 ( .A(n31458), .B(n31459), .Z(n1882) );
  AND U30313 ( .A(n31460), .B(n31461), .Z(n31458) );
  XNOR U30314 ( .A(n31459), .B(n31425), .Z(n31461) );
  XNOR U30315 ( .A(n31462), .B(n31463), .Z(n31425) );
  ANDN U30316 ( .B(n31464), .A(n31465), .Z(n31462) );
  XOR U30317 ( .A(n31463), .B(n31466), .Z(n31464) );
  XOR U30318 ( .A(n31459), .B(n31427), .Z(n31460) );
  XOR U30319 ( .A(n31467), .B(n31468), .Z(n31427) );
  AND U30320 ( .A(n1886), .B(n31469), .Z(n31467) );
  XOR U30321 ( .A(n31470), .B(n31468), .Z(n31469) );
  XNOR U30322 ( .A(n31471), .B(n31472), .Z(n31459) );
  NAND U30323 ( .A(n31473), .B(n31474), .Z(n31472) );
  XOR U30324 ( .A(n31475), .B(n31451), .Z(n31474) );
  XOR U30325 ( .A(n31465), .B(n31466), .Z(n31451) );
  XOR U30326 ( .A(n31476), .B(n31477), .Z(n31466) );
  ANDN U30327 ( .B(n31478), .A(n31479), .Z(n31476) );
  XOR U30328 ( .A(n31477), .B(n31480), .Z(n31478) );
  XOR U30329 ( .A(n31481), .B(n31482), .Z(n31465) );
  XOR U30330 ( .A(n31483), .B(n31484), .Z(n31482) );
  ANDN U30331 ( .B(n31485), .A(n31486), .Z(n31483) );
  XOR U30332 ( .A(n31487), .B(n31484), .Z(n31485) );
  IV U30333 ( .A(n31463), .Z(n31481) );
  XOR U30334 ( .A(n31488), .B(n31489), .Z(n31463) );
  ANDN U30335 ( .B(n31490), .A(n31491), .Z(n31488) );
  XOR U30336 ( .A(n31489), .B(n31492), .Z(n31490) );
  IV U30337 ( .A(n31471), .Z(n31475) );
  XOR U30338 ( .A(n31471), .B(n31453), .Z(n31473) );
  XOR U30339 ( .A(n31493), .B(n31494), .Z(n31453) );
  AND U30340 ( .A(n1886), .B(n31495), .Z(n31493) );
  XOR U30341 ( .A(n31496), .B(n31494), .Z(n31495) );
  NANDN U30342 ( .A(n31455), .B(n31457), .Z(n31471) );
  XOR U30343 ( .A(n31497), .B(n31498), .Z(n31457) );
  AND U30344 ( .A(n1886), .B(n31499), .Z(n31497) );
  XOR U30345 ( .A(n31498), .B(n31500), .Z(n31499) );
  XOR U30346 ( .A(n31501), .B(n31502), .Z(n1886) );
  AND U30347 ( .A(n31503), .B(n31504), .Z(n31501) );
  XNOR U30348 ( .A(n31502), .B(n31468), .Z(n31504) );
  XNOR U30349 ( .A(n31505), .B(n31506), .Z(n31468) );
  ANDN U30350 ( .B(n31507), .A(n31508), .Z(n31505) );
  XOR U30351 ( .A(n31506), .B(n31509), .Z(n31507) );
  XOR U30352 ( .A(n31502), .B(n31470), .Z(n31503) );
  XOR U30353 ( .A(n31510), .B(n31511), .Z(n31470) );
  AND U30354 ( .A(n1890), .B(n31512), .Z(n31510) );
  XOR U30355 ( .A(n31513), .B(n31511), .Z(n31512) );
  XNOR U30356 ( .A(n31514), .B(n31515), .Z(n31502) );
  NAND U30357 ( .A(n31516), .B(n31517), .Z(n31515) );
  XOR U30358 ( .A(n31518), .B(n31494), .Z(n31517) );
  XOR U30359 ( .A(n31508), .B(n31509), .Z(n31494) );
  XOR U30360 ( .A(n31519), .B(n31520), .Z(n31509) );
  ANDN U30361 ( .B(n31521), .A(n31522), .Z(n31519) );
  XOR U30362 ( .A(n31520), .B(n31523), .Z(n31521) );
  XOR U30363 ( .A(n31524), .B(n31525), .Z(n31508) );
  XOR U30364 ( .A(n31526), .B(n31527), .Z(n31525) );
  ANDN U30365 ( .B(n31528), .A(n31529), .Z(n31526) );
  XOR U30366 ( .A(n31530), .B(n31527), .Z(n31528) );
  IV U30367 ( .A(n31506), .Z(n31524) );
  XOR U30368 ( .A(n31531), .B(n31532), .Z(n31506) );
  ANDN U30369 ( .B(n31533), .A(n31534), .Z(n31531) );
  XOR U30370 ( .A(n31532), .B(n31535), .Z(n31533) );
  IV U30371 ( .A(n31514), .Z(n31518) );
  XOR U30372 ( .A(n31514), .B(n31496), .Z(n31516) );
  XOR U30373 ( .A(n31536), .B(n31537), .Z(n31496) );
  AND U30374 ( .A(n1890), .B(n31538), .Z(n31536) );
  XOR U30375 ( .A(n31539), .B(n31537), .Z(n31538) );
  NANDN U30376 ( .A(n31498), .B(n31500), .Z(n31514) );
  XOR U30377 ( .A(n31540), .B(n31541), .Z(n31500) );
  AND U30378 ( .A(n1890), .B(n31542), .Z(n31540) );
  XOR U30379 ( .A(n31541), .B(n31543), .Z(n31542) );
  XOR U30380 ( .A(n31544), .B(n31545), .Z(n1890) );
  AND U30381 ( .A(n31546), .B(n31547), .Z(n31544) );
  XNOR U30382 ( .A(n31545), .B(n31511), .Z(n31547) );
  XNOR U30383 ( .A(n31548), .B(n31549), .Z(n31511) );
  ANDN U30384 ( .B(n31550), .A(n31551), .Z(n31548) );
  XOR U30385 ( .A(n31549), .B(n31552), .Z(n31550) );
  XOR U30386 ( .A(n31545), .B(n31513), .Z(n31546) );
  XOR U30387 ( .A(n31553), .B(n31554), .Z(n31513) );
  AND U30388 ( .A(n1894), .B(n31555), .Z(n31553) );
  XOR U30389 ( .A(n31556), .B(n31554), .Z(n31555) );
  XNOR U30390 ( .A(n31557), .B(n31558), .Z(n31545) );
  NAND U30391 ( .A(n31559), .B(n31560), .Z(n31558) );
  XOR U30392 ( .A(n31561), .B(n31537), .Z(n31560) );
  XOR U30393 ( .A(n31551), .B(n31552), .Z(n31537) );
  XOR U30394 ( .A(n31562), .B(n31563), .Z(n31552) );
  ANDN U30395 ( .B(n31564), .A(n31565), .Z(n31562) );
  XOR U30396 ( .A(n31563), .B(n31566), .Z(n31564) );
  XOR U30397 ( .A(n31567), .B(n31568), .Z(n31551) );
  XOR U30398 ( .A(n31569), .B(n31570), .Z(n31568) );
  ANDN U30399 ( .B(n31571), .A(n31572), .Z(n31569) );
  XOR U30400 ( .A(n31573), .B(n31570), .Z(n31571) );
  IV U30401 ( .A(n31549), .Z(n31567) );
  XOR U30402 ( .A(n31574), .B(n31575), .Z(n31549) );
  ANDN U30403 ( .B(n31576), .A(n31577), .Z(n31574) );
  XOR U30404 ( .A(n31575), .B(n31578), .Z(n31576) );
  IV U30405 ( .A(n31557), .Z(n31561) );
  XOR U30406 ( .A(n31557), .B(n31539), .Z(n31559) );
  XOR U30407 ( .A(n31579), .B(n31580), .Z(n31539) );
  AND U30408 ( .A(n1894), .B(n31581), .Z(n31579) );
  XOR U30409 ( .A(n31582), .B(n31580), .Z(n31581) );
  NANDN U30410 ( .A(n31541), .B(n31543), .Z(n31557) );
  XOR U30411 ( .A(n31583), .B(n31584), .Z(n31543) );
  AND U30412 ( .A(n1894), .B(n31585), .Z(n31583) );
  XOR U30413 ( .A(n31584), .B(n31586), .Z(n31585) );
  XOR U30414 ( .A(n31587), .B(n31588), .Z(n1894) );
  AND U30415 ( .A(n31589), .B(n31590), .Z(n31587) );
  XNOR U30416 ( .A(n31588), .B(n31554), .Z(n31590) );
  XNOR U30417 ( .A(n31591), .B(n31592), .Z(n31554) );
  ANDN U30418 ( .B(n31593), .A(n31594), .Z(n31591) );
  XOR U30419 ( .A(n31592), .B(n31595), .Z(n31593) );
  XOR U30420 ( .A(n31588), .B(n31556), .Z(n31589) );
  XOR U30421 ( .A(n31596), .B(n31597), .Z(n31556) );
  AND U30422 ( .A(n1898), .B(n31598), .Z(n31596) );
  XOR U30423 ( .A(n31599), .B(n31597), .Z(n31598) );
  XNOR U30424 ( .A(n31600), .B(n31601), .Z(n31588) );
  NAND U30425 ( .A(n31602), .B(n31603), .Z(n31601) );
  XOR U30426 ( .A(n31604), .B(n31580), .Z(n31603) );
  XOR U30427 ( .A(n31594), .B(n31595), .Z(n31580) );
  XOR U30428 ( .A(n31605), .B(n31606), .Z(n31595) );
  ANDN U30429 ( .B(n31607), .A(n31608), .Z(n31605) );
  XOR U30430 ( .A(n31606), .B(n31609), .Z(n31607) );
  XOR U30431 ( .A(n31610), .B(n31611), .Z(n31594) );
  XOR U30432 ( .A(n31612), .B(n31613), .Z(n31611) );
  ANDN U30433 ( .B(n31614), .A(n31615), .Z(n31612) );
  XOR U30434 ( .A(n31616), .B(n31613), .Z(n31614) );
  IV U30435 ( .A(n31592), .Z(n31610) );
  XOR U30436 ( .A(n31617), .B(n31618), .Z(n31592) );
  ANDN U30437 ( .B(n31619), .A(n31620), .Z(n31617) );
  XOR U30438 ( .A(n31618), .B(n31621), .Z(n31619) );
  IV U30439 ( .A(n31600), .Z(n31604) );
  XOR U30440 ( .A(n31600), .B(n31582), .Z(n31602) );
  XOR U30441 ( .A(n31622), .B(n31623), .Z(n31582) );
  AND U30442 ( .A(n1898), .B(n31624), .Z(n31622) );
  XOR U30443 ( .A(n31625), .B(n31623), .Z(n31624) );
  NANDN U30444 ( .A(n31584), .B(n31586), .Z(n31600) );
  XOR U30445 ( .A(n31626), .B(n31627), .Z(n31586) );
  AND U30446 ( .A(n1898), .B(n31628), .Z(n31626) );
  XOR U30447 ( .A(n31627), .B(n31629), .Z(n31628) );
  XOR U30448 ( .A(n31630), .B(n31631), .Z(n1898) );
  AND U30449 ( .A(n31632), .B(n31633), .Z(n31630) );
  XNOR U30450 ( .A(n31631), .B(n31597), .Z(n31633) );
  XNOR U30451 ( .A(n31634), .B(n31635), .Z(n31597) );
  ANDN U30452 ( .B(n31636), .A(n31637), .Z(n31634) );
  XOR U30453 ( .A(n31635), .B(n31638), .Z(n31636) );
  XOR U30454 ( .A(n31631), .B(n31599), .Z(n31632) );
  XOR U30455 ( .A(n31639), .B(n31640), .Z(n31599) );
  AND U30456 ( .A(n1902), .B(n31641), .Z(n31639) );
  XOR U30457 ( .A(n31642), .B(n31640), .Z(n31641) );
  XNOR U30458 ( .A(n31643), .B(n31644), .Z(n31631) );
  NAND U30459 ( .A(n31645), .B(n31646), .Z(n31644) );
  XOR U30460 ( .A(n31647), .B(n31623), .Z(n31646) );
  XOR U30461 ( .A(n31637), .B(n31638), .Z(n31623) );
  XOR U30462 ( .A(n31648), .B(n31649), .Z(n31638) );
  ANDN U30463 ( .B(n31650), .A(n31651), .Z(n31648) );
  XOR U30464 ( .A(n31649), .B(n31652), .Z(n31650) );
  XOR U30465 ( .A(n31653), .B(n31654), .Z(n31637) );
  XOR U30466 ( .A(n31655), .B(n31656), .Z(n31654) );
  ANDN U30467 ( .B(n31657), .A(n31658), .Z(n31655) );
  XOR U30468 ( .A(n31659), .B(n31656), .Z(n31657) );
  IV U30469 ( .A(n31635), .Z(n31653) );
  XOR U30470 ( .A(n31660), .B(n31661), .Z(n31635) );
  ANDN U30471 ( .B(n31662), .A(n31663), .Z(n31660) );
  XOR U30472 ( .A(n31661), .B(n31664), .Z(n31662) );
  IV U30473 ( .A(n31643), .Z(n31647) );
  XOR U30474 ( .A(n31643), .B(n31625), .Z(n31645) );
  XOR U30475 ( .A(n31665), .B(n31666), .Z(n31625) );
  AND U30476 ( .A(n1902), .B(n31667), .Z(n31665) );
  XOR U30477 ( .A(n31668), .B(n31666), .Z(n31667) );
  NANDN U30478 ( .A(n31627), .B(n31629), .Z(n31643) );
  XOR U30479 ( .A(n31669), .B(n31670), .Z(n31629) );
  AND U30480 ( .A(n1902), .B(n31671), .Z(n31669) );
  XOR U30481 ( .A(n31670), .B(n31672), .Z(n31671) );
  XOR U30482 ( .A(n31673), .B(n31674), .Z(n1902) );
  AND U30483 ( .A(n31675), .B(n31676), .Z(n31673) );
  XNOR U30484 ( .A(n31674), .B(n31640), .Z(n31676) );
  XNOR U30485 ( .A(n31677), .B(n31678), .Z(n31640) );
  ANDN U30486 ( .B(n31679), .A(n31680), .Z(n31677) );
  XOR U30487 ( .A(n31678), .B(n31681), .Z(n31679) );
  XOR U30488 ( .A(n31674), .B(n31642), .Z(n31675) );
  XOR U30489 ( .A(n31682), .B(n31683), .Z(n31642) );
  AND U30490 ( .A(n1906), .B(n31684), .Z(n31682) );
  XOR U30491 ( .A(n31685), .B(n31683), .Z(n31684) );
  XNOR U30492 ( .A(n31686), .B(n31687), .Z(n31674) );
  NAND U30493 ( .A(n31688), .B(n31689), .Z(n31687) );
  XOR U30494 ( .A(n31690), .B(n31666), .Z(n31689) );
  XOR U30495 ( .A(n31680), .B(n31681), .Z(n31666) );
  XOR U30496 ( .A(n31691), .B(n31692), .Z(n31681) );
  ANDN U30497 ( .B(n31693), .A(n31694), .Z(n31691) );
  XOR U30498 ( .A(n31692), .B(n31695), .Z(n31693) );
  XOR U30499 ( .A(n31696), .B(n31697), .Z(n31680) );
  XOR U30500 ( .A(n31698), .B(n31699), .Z(n31697) );
  ANDN U30501 ( .B(n31700), .A(n31701), .Z(n31698) );
  XOR U30502 ( .A(n31702), .B(n31699), .Z(n31700) );
  IV U30503 ( .A(n31678), .Z(n31696) );
  XOR U30504 ( .A(n31703), .B(n31704), .Z(n31678) );
  ANDN U30505 ( .B(n31705), .A(n31706), .Z(n31703) );
  XOR U30506 ( .A(n31704), .B(n31707), .Z(n31705) );
  IV U30507 ( .A(n31686), .Z(n31690) );
  XOR U30508 ( .A(n31686), .B(n31668), .Z(n31688) );
  XOR U30509 ( .A(n31708), .B(n31709), .Z(n31668) );
  AND U30510 ( .A(n1906), .B(n31710), .Z(n31708) );
  XOR U30511 ( .A(n31711), .B(n31709), .Z(n31710) );
  NANDN U30512 ( .A(n31670), .B(n31672), .Z(n31686) );
  XOR U30513 ( .A(n31712), .B(n31713), .Z(n31672) );
  AND U30514 ( .A(n1906), .B(n31714), .Z(n31712) );
  XOR U30515 ( .A(n31713), .B(n31715), .Z(n31714) );
  XOR U30516 ( .A(n31716), .B(n31717), .Z(n1906) );
  AND U30517 ( .A(n31718), .B(n31719), .Z(n31716) );
  XNOR U30518 ( .A(n31717), .B(n31683), .Z(n31719) );
  XNOR U30519 ( .A(n31720), .B(n31721), .Z(n31683) );
  ANDN U30520 ( .B(n31722), .A(n31723), .Z(n31720) );
  XOR U30521 ( .A(n31721), .B(n31724), .Z(n31722) );
  XOR U30522 ( .A(n31717), .B(n31685), .Z(n31718) );
  XOR U30523 ( .A(n31725), .B(n31726), .Z(n31685) );
  AND U30524 ( .A(n1910), .B(n31727), .Z(n31725) );
  XOR U30525 ( .A(n31728), .B(n31726), .Z(n31727) );
  XNOR U30526 ( .A(n31729), .B(n31730), .Z(n31717) );
  NAND U30527 ( .A(n31731), .B(n31732), .Z(n31730) );
  XOR U30528 ( .A(n31733), .B(n31709), .Z(n31732) );
  XOR U30529 ( .A(n31723), .B(n31724), .Z(n31709) );
  XOR U30530 ( .A(n31734), .B(n31735), .Z(n31724) );
  ANDN U30531 ( .B(n31736), .A(n31737), .Z(n31734) );
  XOR U30532 ( .A(n31735), .B(n31738), .Z(n31736) );
  XOR U30533 ( .A(n31739), .B(n31740), .Z(n31723) );
  XOR U30534 ( .A(n31741), .B(n31742), .Z(n31740) );
  ANDN U30535 ( .B(n31743), .A(n31744), .Z(n31741) );
  XOR U30536 ( .A(n31745), .B(n31742), .Z(n31743) );
  IV U30537 ( .A(n31721), .Z(n31739) );
  XOR U30538 ( .A(n31746), .B(n31747), .Z(n31721) );
  ANDN U30539 ( .B(n31748), .A(n31749), .Z(n31746) );
  XOR U30540 ( .A(n31747), .B(n31750), .Z(n31748) );
  IV U30541 ( .A(n31729), .Z(n31733) );
  XOR U30542 ( .A(n31729), .B(n31711), .Z(n31731) );
  XOR U30543 ( .A(n31751), .B(n31752), .Z(n31711) );
  AND U30544 ( .A(n1910), .B(n31753), .Z(n31751) );
  XOR U30545 ( .A(n31754), .B(n31752), .Z(n31753) );
  NANDN U30546 ( .A(n31713), .B(n31715), .Z(n31729) );
  XOR U30547 ( .A(n31755), .B(n31756), .Z(n31715) );
  AND U30548 ( .A(n1910), .B(n31757), .Z(n31755) );
  XOR U30549 ( .A(n31756), .B(n31758), .Z(n31757) );
  XOR U30550 ( .A(n31759), .B(n31760), .Z(n1910) );
  AND U30551 ( .A(n31761), .B(n31762), .Z(n31759) );
  XNOR U30552 ( .A(n31760), .B(n31726), .Z(n31762) );
  XNOR U30553 ( .A(n31763), .B(n31764), .Z(n31726) );
  ANDN U30554 ( .B(n31765), .A(n31766), .Z(n31763) );
  XOR U30555 ( .A(n31764), .B(n31767), .Z(n31765) );
  XOR U30556 ( .A(n31760), .B(n31728), .Z(n31761) );
  XOR U30557 ( .A(n31768), .B(n31769), .Z(n31728) );
  AND U30558 ( .A(n1914), .B(n31770), .Z(n31768) );
  XOR U30559 ( .A(n31771), .B(n31769), .Z(n31770) );
  XNOR U30560 ( .A(n31772), .B(n31773), .Z(n31760) );
  NAND U30561 ( .A(n31774), .B(n31775), .Z(n31773) );
  XOR U30562 ( .A(n31776), .B(n31752), .Z(n31775) );
  XOR U30563 ( .A(n31766), .B(n31767), .Z(n31752) );
  XOR U30564 ( .A(n31777), .B(n31778), .Z(n31767) );
  ANDN U30565 ( .B(n31779), .A(n31780), .Z(n31777) );
  XOR U30566 ( .A(n31778), .B(n31781), .Z(n31779) );
  XOR U30567 ( .A(n31782), .B(n31783), .Z(n31766) );
  XOR U30568 ( .A(n31784), .B(n31785), .Z(n31783) );
  ANDN U30569 ( .B(n31786), .A(n31787), .Z(n31784) );
  XOR U30570 ( .A(n31788), .B(n31785), .Z(n31786) );
  IV U30571 ( .A(n31764), .Z(n31782) );
  XOR U30572 ( .A(n31789), .B(n31790), .Z(n31764) );
  ANDN U30573 ( .B(n31791), .A(n31792), .Z(n31789) );
  XOR U30574 ( .A(n31790), .B(n31793), .Z(n31791) );
  IV U30575 ( .A(n31772), .Z(n31776) );
  XOR U30576 ( .A(n31772), .B(n31754), .Z(n31774) );
  XOR U30577 ( .A(n31794), .B(n31795), .Z(n31754) );
  AND U30578 ( .A(n1914), .B(n31796), .Z(n31794) );
  XOR U30579 ( .A(n31797), .B(n31795), .Z(n31796) );
  NANDN U30580 ( .A(n31756), .B(n31758), .Z(n31772) );
  XOR U30581 ( .A(n31798), .B(n31799), .Z(n31758) );
  AND U30582 ( .A(n1914), .B(n31800), .Z(n31798) );
  XOR U30583 ( .A(n31799), .B(n31801), .Z(n31800) );
  XOR U30584 ( .A(n31802), .B(n31803), .Z(n1914) );
  AND U30585 ( .A(n31804), .B(n31805), .Z(n31802) );
  XNOR U30586 ( .A(n31803), .B(n31769), .Z(n31805) );
  XNOR U30587 ( .A(n31806), .B(n31807), .Z(n31769) );
  ANDN U30588 ( .B(n31808), .A(n31809), .Z(n31806) );
  XOR U30589 ( .A(n31807), .B(n31810), .Z(n31808) );
  XOR U30590 ( .A(n31803), .B(n31771), .Z(n31804) );
  XOR U30591 ( .A(n31811), .B(n31812), .Z(n31771) );
  AND U30592 ( .A(n1918), .B(n31813), .Z(n31811) );
  XOR U30593 ( .A(n31814), .B(n31812), .Z(n31813) );
  XNOR U30594 ( .A(n31815), .B(n31816), .Z(n31803) );
  NAND U30595 ( .A(n31817), .B(n31818), .Z(n31816) );
  XOR U30596 ( .A(n31819), .B(n31795), .Z(n31818) );
  XOR U30597 ( .A(n31809), .B(n31810), .Z(n31795) );
  XOR U30598 ( .A(n31820), .B(n31821), .Z(n31810) );
  ANDN U30599 ( .B(n31822), .A(n31823), .Z(n31820) );
  XOR U30600 ( .A(n31821), .B(n31824), .Z(n31822) );
  XOR U30601 ( .A(n31825), .B(n31826), .Z(n31809) );
  XOR U30602 ( .A(n31827), .B(n31828), .Z(n31826) );
  ANDN U30603 ( .B(n31829), .A(n31830), .Z(n31827) );
  XOR U30604 ( .A(n31831), .B(n31828), .Z(n31829) );
  IV U30605 ( .A(n31807), .Z(n31825) );
  XOR U30606 ( .A(n31832), .B(n31833), .Z(n31807) );
  ANDN U30607 ( .B(n31834), .A(n31835), .Z(n31832) );
  XOR U30608 ( .A(n31833), .B(n31836), .Z(n31834) );
  IV U30609 ( .A(n31815), .Z(n31819) );
  XOR U30610 ( .A(n31815), .B(n31797), .Z(n31817) );
  XOR U30611 ( .A(n31837), .B(n31838), .Z(n31797) );
  AND U30612 ( .A(n1918), .B(n31839), .Z(n31837) );
  XOR U30613 ( .A(n31840), .B(n31838), .Z(n31839) );
  NANDN U30614 ( .A(n31799), .B(n31801), .Z(n31815) );
  XOR U30615 ( .A(n31841), .B(n31842), .Z(n31801) );
  AND U30616 ( .A(n1918), .B(n31843), .Z(n31841) );
  XOR U30617 ( .A(n31842), .B(n31844), .Z(n31843) );
  XOR U30618 ( .A(n31845), .B(n31846), .Z(n1918) );
  AND U30619 ( .A(n31847), .B(n31848), .Z(n31845) );
  XNOR U30620 ( .A(n31846), .B(n31812), .Z(n31848) );
  XNOR U30621 ( .A(n31849), .B(n31850), .Z(n31812) );
  ANDN U30622 ( .B(n31851), .A(n31852), .Z(n31849) );
  XOR U30623 ( .A(n31850), .B(n31853), .Z(n31851) );
  XOR U30624 ( .A(n31846), .B(n31814), .Z(n31847) );
  XOR U30625 ( .A(n31854), .B(n31855), .Z(n31814) );
  AND U30626 ( .A(n1922), .B(n31856), .Z(n31854) );
  XOR U30627 ( .A(n31857), .B(n31855), .Z(n31856) );
  XNOR U30628 ( .A(n31858), .B(n31859), .Z(n31846) );
  NAND U30629 ( .A(n31860), .B(n31861), .Z(n31859) );
  XOR U30630 ( .A(n31862), .B(n31838), .Z(n31861) );
  XOR U30631 ( .A(n31852), .B(n31853), .Z(n31838) );
  XOR U30632 ( .A(n31863), .B(n31864), .Z(n31853) );
  ANDN U30633 ( .B(n31865), .A(n31866), .Z(n31863) );
  XOR U30634 ( .A(n31864), .B(n31867), .Z(n31865) );
  XOR U30635 ( .A(n31868), .B(n31869), .Z(n31852) );
  XOR U30636 ( .A(n31870), .B(n31871), .Z(n31869) );
  ANDN U30637 ( .B(n31872), .A(n31873), .Z(n31870) );
  XOR U30638 ( .A(n31874), .B(n31871), .Z(n31872) );
  IV U30639 ( .A(n31850), .Z(n31868) );
  XOR U30640 ( .A(n31875), .B(n31876), .Z(n31850) );
  ANDN U30641 ( .B(n31877), .A(n31878), .Z(n31875) );
  XOR U30642 ( .A(n31876), .B(n31879), .Z(n31877) );
  IV U30643 ( .A(n31858), .Z(n31862) );
  XOR U30644 ( .A(n31858), .B(n31840), .Z(n31860) );
  XOR U30645 ( .A(n31880), .B(n31881), .Z(n31840) );
  AND U30646 ( .A(n1922), .B(n31882), .Z(n31880) );
  XOR U30647 ( .A(n31883), .B(n31881), .Z(n31882) );
  NANDN U30648 ( .A(n31842), .B(n31844), .Z(n31858) );
  XOR U30649 ( .A(n31884), .B(n31885), .Z(n31844) );
  AND U30650 ( .A(n1922), .B(n31886), .Z(n31884) );
  XOR U30651 ( .A(n31885), .B(n31887), .Z(n31886) );
  XOR U30652 ( .A(n31888), .B(n31889), .Z(n1922) );
  AND U30653 ( .A(n31890), .B(n31891), .Z(n31888) );
  XNOR U30654 ( .A(n31889), .B(n31855), .Z(n31891) );
  XNOR U30655 ( .A(n31892), .B(n31893), .Z(n31855) );
  ANDN U30656 ( .B(n31894), .A(n31895), .Z(n31892) );
  XOR U30657 ( .A(n31893), .B(n31896), .Z(n31894) );
  XOR U30658 ( .A(n31889), .B(n31857), .Z(n31890) );
  XOR U30659 ( .A(n31897), .B(n31898), .Z(n31857) );
  AND U30660 ( .A(n1926), .B(n31899), .Z(n31897) );
  XOR U30661 ( .A(n31900), .B(n31898), .Z(n31899) );
  XNOR U30662 ( .A(n31901), .B(n31902), .Z(n31889) );
  NAND U30663 ( .A(n31903), .B(n31904), .Z(n31902) );
  XOR U30664 ( .A(n31905), .B(n31881), .Z(n31904) );
  XOR U30665 ( .A(n31895), .B(n31896), .Z(n31881) );
  XOR U30666 ( .A(n31906), .B(n31907), .Z(n31896) );
  ANDN U30667 ( .B(n31908), .A(n31909), .Z(n31906) );
  XOR U30668 ( .A(n31907), .B(n31910), .Z(n31908) );
  XOR U30669 ( .A(n31911), .B(n31912), .Z(n31895) );
  XOR U30670 ( .A(n31913), .B(n31914), .Z(n31912) );
  ANDN U30671 ( .B(n31915), .A(n31916), .Z(n31913) );
  XOR U30672 ( .A(n31917), .B(n31914), .Z(n31915) );
  IV U30673 ( .A(n31893), .Z(n31911) );
  XOR U30674 ( .A(n31918), .B(n31919), .Z(n31893) );
  ANDN U30675 ( .B(n31920), .A(n31921), .Z(n31918) );
  XOR U30676 ( .A(n31919), .B(n31922), .Z(n31920) );
  IV U30677 ( .A(n31901), .Z(n31905) );
  XOR U30678 ( .A(n31901), .B(n31883), .Z(n31903) );
  XOR U30679 ( .A(n31923), .B(n31924), .Z(n31883) );
  AND U30680 ( .A(n1926), .B(n31925), .Z(n31923) );
  XOR U30681 ( .A(n31926), .B(n31924), .Z(n31925) );
  NANDN U30682 ( .A(n31885), .B(n31887), .Z(n31901) );
  XOR U30683 ( .A(n31927), .B(n31928), .Z(n31887) );
  AND U30684 ( .A(n1926), .B(n31929), .Z(n31927) );
  XOR U30685 ( .A(n31928), .B(n31930), .Z(n31929) );
  XOR U30686 ( .A(n31931), .B(n31932), .Z(n1926) );
  AND U30687 ( .A(n31933), .B(n31934), .Z(n31931) );
  XNOR U30688 ( .A(n31932), .B(n31898), .Z(n31934) );
  XNOR U30689 ( .A(n31935), .B(n31936), .Z(n31898) );
  ANDN U30690 ( .B(n31937), .A(n31938), .Z(n31935) );
  XOR U30691 ( .A(n31936), .B(n31939), .Z(n31937) );
  XOR U30692 ( .A(n31932), .B(n31900), .Z(n31933) );
  XOR U30693 ( .A(n31940), .B(n31941), .Z(n31900) );
  AND U30694 ( .A(n1930), .B(n31942), .Z(n31940) );
  XOR U30695 ( .A(n31943), .B(n31941), .Z(n31942) );
  XNOR U30696 ( .A(n31944), .B(n31945), .Z(n31932) );
  NAND U30697 ( .A(n31946), .B(n31947), .Z(n31945) );
  XOR U30698 ( .A(n31948), .B(n31924), .Z(n31947) );
  XOR U30699 ( .A(n31938), .B(n31939), .Z(n31924) );
  XOR U30700 ( .A(n31949), .B(n31950), .Z(n31939) );
  ANDN U30701 ( .B(n31951), .A(n31952), .Z(n31949) );
  XOR U30702 ( .A(n31950), .B(n31953), .Z(n31951) );
  XOR U30703 ( .A(n31954), .B(n31955), .Z(n31938) );
  XOR U30704 ( .A(n31956), .B(n31957), .Z(n31955) );
  ANDN U30705 ( .B(n31958), .A(n31959), .Z(n31956) );
  XOR U30706 ( .A(n31960), .B(n31957), .Z(n31958) );
  IV U30707 ( .A(n31936), .Z(n31954) );
  XOR U30708 ( .A(n31961), .B(n31962), .Z(n31936) );
  ANDN U30709 ( .B(n31963), .A(n31964), .Z(n31961) );
  XOR U30710 ( .A(n31962), .B(n31965), .Z(n31963) );
  IV U30711 ( .A(n31944), .Z(n31948) );
  XOR U30712 ( .A(n31944), .B(n31926), .Z(n31946) );
  XOR U30713 ( .A(n31966), .B(n31967), .Z(n31926) );
  AND U30714 ( .A(n1930), .B(n31968), .Z(n31966) );
  XOR U30715 ( .A(n31969), .B(n31967), .Z(n31968) );
  NANDN U30716 ( .A(n31928), .B(n31930), .Z(n31944) );
  XOR U30717 ( .A(n31970), .B(n31971), .Z(n31930) );
  AND U30718 ( .A(n1930), .B(n31972), .Z(n31970) );
  XOR U30719 ( .A(n31971), .B(n31973), .Z(n31972) );
  XOR U30720 ( .A(n31974), .B(n31975), .Z(n1930) );
  AND U30721 ( .A(n31976), .B(n31977), .Z(n31974) );
  XNOR U30722 ( .A(n31975), .B(n31941), .Z(n31977) );
  XNOR U30723 ( .A(n31978), .B(n31979), .Z(n31941) );
  ANDN U30724 ( .B(n31980), .A(n31981), .Z(n31978) );
  XOR U30725 ( .A(n31979), .B(n31982), .Z(n31980) );
  XOR U30726 ( .A(n31975), .B(n31943), .Z(n31976) );
  XOR U30727 ( .A(n31983), .B(n31984), .Z(n31943) );
  AND U30728 ( .A(n1934), .B(n31985), .Z(n31983) );
  XOR U30729 ( .A(n31986), .B(n31984), .Z(n31985) );
  XNOR U30730 ( .A(n31987), .B(n31988), .Z(n31975) );
  NAND U30731 ( .A(n31989), .B(n31990), .Z(n31988) );
  XOR U30732 ( .A(n31991), .B(n31967), .Z(n31990) );
  XOR U30733 ( .A(n31981), .B(n31982), .Z(n31967) );
  XOR U30734 ( .A(n31992), .B(n31993), .Z(n31982) );
  ANDN U30735 ( .B(n31994), .A(n31995), .Z(n31992) );
  XOR U30736 ( .A(n31993), .B(n31996), .Z(n31994) );
  XOR U30737 ( .A(n31997), .B(n31998), .Z(n31981) );
  XOR U30738 ( .A(n31999), .B(n32000), .Z(n31998) );
  ANDN U30739 ( .B(n32001), .A(n32002), .Z(n31999) );
  XOR U30740 ( .A(n32003), .B(n32000), .Z(n32001) );
  IV U30741 ( .A(n31979), .Z(n31997) );
  XOR U30742 ( .A(n32004), .B(n32005), .Z(n31979) );
  ANDN U30743 ( .B(n32006), .A(n32007), .Z(n32004) );
  XOR U30744 ( .A(n32005), .B(n32008), .Z(n32006) );
  IV U30745 ( .A(n31987), .Z(n31991) );
  XOR U30746 ( .A(n31987), .B(n31969), .Z(n31989) );
  XOR U30747 ( .A(n32009), .B(n32010), .Z(n31969) );
  AND U30748 ( .A(n1934), .B(n32011), .Z(n32009) );
  XOR U30749 ( .A(n32012), .B(n32010), .Z(n32011) );
  NANDN U30750 ( .A(n31971), .B(n31973), .Z(n31987) );
  XOR U30751 ( .A(n32013), .B(n32014), .Z(n31973) );
  AND U30752 ( .A(n1934), .B(n32015), .Z(n32013) );
  XOR U30753 ( .A(n32014), .B(n32016), .Z(n32015) );
  XOR U30754 ( .A(n32017), .B(n32018), .Z(n1934) );
  AND U30755 ( .A(n32019), .B(n32020), .Z(n32017) );
  XNOR U30756 ( .A(n32018), .B(n31984), .Z(n32020) );
  XNOR U30757 ( .A(n32021), .B(n32022), .Z(n31984) );
  ANDN U30758 ( .B(n32023), .A(n32024), .Z(n32021) );
  XOR U30759 ( .A(n32022), .B(n32025), .Z(n32023) );
  XOR U30760 ( .A(n32018), .B(n31986), .Z(n32019) );
  XOR U30761 ( .A(n32026), .B(n32027), .Z(n31986) );
  AND U30762 ( .A(n1938), .B(n32028), .Z(n32026) );
  XOR U30763 ( .A(n32029), .B(n32027), .Z(n32028) );
  XNOR U30764 ( .A(n32030), .B(n32031), .Z(n32018) );
  NAND U30765 ( .A(n32032), .B(n32033), .Z(n32031) );
  XOR U30766 ( .A(n32034), .B(n32010), .Z(n32033) );
  XOR U30767 ( .A(n32024), .B(n32025), .Z(n32010) );
  XOR U30768 ( .A(n32035), .B(n32036), .Z(n32025) );
  ANDN U30769 ( .B(n32037), .A(n32038), .Z(n32035) );
  XOR U30770 ( .A(n32036), .B(n32039), .Z(n32037) );
  XOR U30771 ( .A(n32040), .B(n32041), .Z(n32024) );
  XOR U30772 ( .A(n32042), .B(n32043), .Z(n32041) );
  ANDN U30773 ( .B(n32044), .A(n32045), .Z(n32042) );
  XOR U30774 ( .A(n32046), .B(n32043), .Z(n32044) );
  IV U30775 ( .A(n32022), .Z(n32040) );
  XOR U30776 ( .A(n32047), .B(n32048), .Z(n32022) );
  ANDN U30777 ( .B(n32049), .A(n32050), .Z(n32047) );
  XOR U30778 ( .A(n32048), .B(n32051), .Z(n32049) );
  IV U30779 ( .A(n32030), .Z(n32034) );
  XOR U30780 ( .A(n32030), .B(n32012), .Z(n32032) );
  XOR U30781 ( .A(n32052), .B(n32053), .Z(n32012) );
  AND U30782 ( .A(n1938), .B(n32054), .Z(n32052) );
  XOR U30783 ( .A(n32055), .B(n32053), .Z(n32054) );
  NANDN U30784 ( .A(n32014), .B(n32016), .Z(n32030) );
  XOR U30785 ( .A(n32056), .B(n32057), .Z(n32016) );
  AND U30786 ( .A(n1938), .B(n32058), .Z(n32056) );
  XOR U30787 ( .A(n32057), .B(n32059), .Z(n32058) );
  XOR U30788 ( .A(n32060), .B(n32061), .Z(n1938) );
  AND U30789 ( .A(n32062), .B(n32063), .Z(n32060) );
  XNOR U30790 ( .A(n32061), .B(n32027), .Z(n32063) );
  XNOR U30791 ( .A(n32064), .B(n32065), .Z(n32027) );
  ANDN U30792 ( .B(n32066), .A(n32067), .Z(n32064) );
  XOR U30793 ( .A(n32065), .B(n32068), .Z(n32066) );
  XOR U30794 ( .A(n32061), .B(n32029), .Z(n32062) );
  XOR U30795 ( .A(n32069), .B(n32070), .Z(n32029) );
  AND U30796 ( .A(n1942), .B(n32071), .Z(n32069) );
  XOR U30797 ( .A(n32072), .B(n32070), .Z(n32071) );
  XNOR U30798 ( .A(n32073), .B(n32074), .Z(n32061) );
  NAND U30799 ( .A(n32075), .B(n32076), .Z(n32074) );
  XOR U30800 ( .A(n32077), .B(n32053), .Z(n32076) );
  XOR U30801 ( .A(n32067), .B(n32068), .Z(n32053) );
  XOR U30802 ( .A(n32078), .B(n32079), .Z(n32068) );
  ANDN U30803 ( .B(n32080), .A(n32081), .Z(n32078) );
  XOR U30804 ( .A(n32079), .B(n32082), .Z(n32080) );
  XOR U30805 ( .A(n32083), .B(n32084), .Z(n32067) );
  XOR U30806 ( .A(n32085), .B(n32086), .Z(n32084) );
  ANDN U30807 ( .B(n32087), .A(n32088), .Z(n32085) );
  XOR U30808 ( .A(n32089), .B(n32086), .Z(n32087) );
  IV U30809 ( .A(n32065), .Z(n32083) );
  XOR U30810 ( .A(n32090), .B(n32091), .Z(n32065) );
  ANDN U30811 ( .B(n32092), .A(n32093), .Z(n32090) );
  XOR U30812 ( .A(n32091), .B(n32094), .Z(n32092) );
  IV U30813 ( .A(n32073), .Z(n32077) );
  XOR U30814 ( .A(n32073), .B(n32055), .Z(n32075) );
  XOR U30815 ( .A(n32095), .B(n32096), .Z(n32055) );
  AND U30816 ( .A(n1942), .B(n32097), .Z(n32095) );
  XOR U30817 ( .A(n32098), .B(n32096), .Z(n32097) );
  NANDN U30818 ( .A(n32057), .B(n32059), .Z(n32073) );
  XOR U30819 ( .A(n32099), .B(n32100), .Z(n32059) );
  AND U30820 ( .A(n1942), .B(n32101), .Z(n32099) );
  XOR U30821 ( .A(n32100), .B(n32102), .Z(n32101) );
  XOR U30822 ( .A(n32103), .B(n32104), .Z(n1942) );
  AND U30823 ( .A(n32105), .B(n32106), .Z(n32103) );
  XNOR U30824 ( .A(n32104), .B(n32070), .Z(n32106) );
  XNOR U30825 ( .A(n32107), .B(n32108), .Z(n32070) );
  ANDN U30826 ( .B(n32109), .A(n32110), .Z(n32107) );
  XOR U30827 ( .A(n32108), .B(n32111), .Z(n32109) );
  XOR U30828 ( .A(n32104), .B(n32072), .Z(n32105) );
  XOR U30829 ( .A(n32112), .B(n32113), .Z(n32072) );
  AND U30830 ( .A(n1946), .B(n32114), .Z(n32112) );
  XOR U30831 ( .A(n32115), .B(n32113), .Z(n32114) );
  XNOR U30832 ( .A(n32116), .B(n32117), .Z(n32104) );
  NAND U30833 ( .A(n32118), .B(n32119), .Z(n32117) );
  XOR U30834 ( .A(n32120), .B(n32096), .Z(n32119) );
  XOR U30835 ( .A(n32110), .B(n32111), .Z(n32096) );
  XOR U30836 ( .A(n32121), .B(n32122), .Z(n32111) );
  ANDN U30837 ( .B(n32123), .A(n32124), .Z(n32121) );
  XOR U30838 ( .A(n32122), .B(n32125), .Z(n32123) );
  XOR U30839 ( .A(n32126), .B(n32127), .Z(n32110) );
  XOR U30840 ( .A(n32128), .B(n32129), .Z(n32127) );
  ANDN U30841 ( .B(n32130), .A(n32131), .Z(n32128) );
  XOR U30842 ( .A(n32132), .B(n32129), .Z(n32130) );
  IV U30843 ( .A(n32108), .Z(n32126) );
  XOR U30844 ( .A(n32133), .B(n32134), .Z(n32108) );
  ANDN U30845 ( .B(n32135), .A(n32136), .Z(n32133) );
  XOR U30846 ( .A(n32134), .B(n32137), .Z(n32135) );
  IV U30847 ( .A(n32116), .Z(n32120) );
  XOR U30848 ( .A(n32116), .B(n32098), .Z(n32118) );
  XOR U30849 ( .A(n32138), .B(n32139), .Z(n32098) );
  AND U30850 ( .A(n1946), .B(n32140), .Z(n32138) );
  XOR U30851 ( .A(n32141), .B(n32139), .Z(n32140) );
  NANDN U30852 ( .A(n32100), .B(n32102), .Z(n32116) );
  XOR U30853 ( .A(n32142), .B(n32143), .Z(n32102) );
  AND U30854 ( .A(n1946), .B(n32144), .Z(n32142) );
  XOR U30855 ( .A(n32143), .B(n32145), .Z(n32144) );
  XOR U30856 ( .A(n32146), .B(n32147), .Z(n1946) );
  AND U30857 ( .A(n32148), .B(n32149), .Z(n32146) );
  XNOR U30858 ( .A(n32147), .B(n32113), .Z(n32149) );
  XNOR U30859 ( .A(n32150), .B(n32151), .Z(n32113) );
  ANDN U30860 ( .B(n32152), .A(n32153), .Z(n32150) );
  XOR U30861 ( .A(n32151), .B(n32154), .Z(n32152) );
  XOR U30862 ( .A(n32147), .B(n32115), .Z(n32148) );
  XOR U30863 ( .A(n32155), .B(n32156), .Z(n32115) );
  AND U30864 ( .A(n1950), .B(n32157), .Z(n32155) );
  XOR U30865 ( .A(n32158), .B(n32156), .Z(n32157) );
  XNOR U30866 ( .A(n32159), .B(n32160), .Z(n32147) );
  NAND U30867 ( .A(n32161), .B(n32162), .Z(n32160) );
  XOR U30868 ( .A(n32163), .B(n32139), .Z(n32162) );
  XOR U30869 ( .A(n32153), .B(n32154), .Z(n32139) );
  XOR U30870 ( .A(n32164), .B(n32165), .Z(n32154) );
  ANDN U30871 ( .B(n32166), .A(n32167), .Z(n32164) );
  XOR U30872 ( .A(n32165), .B(n32168), .Z(n32166) );
  XOR U30873 ( .A(n32169), .B(n32170), .Z(n32153) );
  XOR U30874 ( .A(n32171), .B(n32172), .Z(n32170) );
  ANDN U30875 ( .B(n32173), .A(n32174), .Z(n32171) );
  XOR U30876 ( .A(n32175), .B(n32172), .Z(n32173) );
  IV U30877 ( .A(n32151), .Z(n32169) );
  XOR U30878 ( .A(n32176), .B(n32177), .Z(n32151) );
  ANDN U30879 ( .B(n32178), .A(n32179), .Z(n32176) );
  XOR U30880 ( .A(n32177), .B(n32180), .Z(n32178) );
  IV U30881 ( .A(n32159), .Z(n32163) );
  XOR U30882 ( .A(n32159), .B(n32141), .Z(n32161) );
  XOR U30883 ( .A(n32181), .B(n32182), .Z(n32141) );
  AND U30884 ( .A(n1950), .B(n32183), .Z(n32181) );
  XOR U30885 ( .A(n32184), .B(n32182), .Z(n32183) );
  NANDN U30886 ( .A(n32143), .B(n32145), .Z(n32159) );
  XOR U30887 ( .A(n32185), .B(n32186), .Z(n32145) );
  AND U30888 ( .A(n1950), .B(n32187), .Z(n32185) );
  XOR U30889 ( .A(n32186), .B(n32188), .Z(n32187) );
  XOR U30890 ( .A(n32189), .B(n32190), .Z(n1950) );
  AND U30891 ( .A(n32191), .B(n32192), .Z(n32189) );
  XNOR U30892 ( .A(n32190), .B(n32156), .Z(n32192) );
  XNOR U30893 ( .A(n32193), .B(n32194), .Z(n32156) );
  ANDN U30894 ( .B(n32195), .A(n32196), .Z(n32193) );
  XOR U30895 ( .A(n32194), .B(n32197), .Z(n32195) );
  XOR U30896 ( .A(n32190), .B(n32158), .Z(n32191) );
  XOR U30897 ( .A(n32198), .B(n32199), .Z(n32158) );
  AND U30898 ( .A(n1954), .B(n32200), .Z(n32198) );
  XOR U30899 ( .A(n32201), .B(n32199), .Z(n32200) );
  XNOR U30900 ( .A(n32202), .B(n32203), .Z(n32190) );
  NAND U30901 ( .A(n32204), .B(n32205), .Z(n32203) );
  XOR U30902 ( .A(n32206), .B(n32182), .Z(n32205) );
  XOR U30903 ( .A(n32196), .B(n32197), .Z(n32182) );
  XOR U30904 ( .A(n32207), .B(n32208), .Z(n32197) );
  ANDN U30905 ( .B(n32209), .A(n32210), .Z(n32207) );
  XOR U30906 ( .A(n32208), .B(n32211), .Z(n32209) );
  XOR U30907 ( .A(n32212), .B(n32213), .Z(n32196) );
  XOR U30908 ( .A(n32214), .B(n32215), .Z(n32213) );
  ANDN U30909 ( .B(n32216), .A(n32217), .Z(n32214) );
  XOR U30910 ( .A(n32218), .B(n32215), .Z(n32216) );
  IV U30911 ( .A(n32194), .Z(n32212) );
  XOR U30912 ( .A(n32219), .B(n32220), .Z(n32194) );
  ANDN U30913 ( .B(n32221), .A(n32222), .Z(n32219) );
  XOR U30914 ( .A(n32220), .B(n32223), .Z(n32221) );
  IV U30915 ( .A(n32202), .Z(n32206) );
  XOR U30916 ( .A(n32202), .B(n32184), .Z(n32204) );
  XOR U30917 ( .A(n32224), .B(n32225), .Z(n32184) );
  AND U30918 ( .A(n1954), .B(n32226), .Z(n32224) );
  XOR U30919 ( .A(n32227), .B(n32225), .Z(n32226) );
  NANDN U30920 ( .A(n32186), .B(n32188), .Z(n32202) );
  XOR U30921 ( .A(n32228), .B(n32229), .Z(n32188) );
  AND U30922 ( .A(n1954), .B(n32230), .Z(n32228) );
  XOR U30923 ( .A(n32229), .B(n32231), .Z(n32230) );
  XOR U30924 ( .A(n32232), .B(n32233), .Z(n1954) );
  AND U30925 ( .A(n32234), .B(n32235), .Z(n32232) );
  XNOR U30926 ( .A(n32233), .B(n32199), .Z(n32235) );
  XNOR U30927 ( .A(n32236), .B(n32237), .Z(n32199) );
  ANDN U30928 ( .B(n32238), .A(n32239), .Z(n32236) );
  XOR U30929 ( .A(n32237), .B(n32240), .Z(n32238) );
  XOR U30930 ( .A(n32233), .B(n32201), .Z(n32234) );
  XOR U30931 ( .A(n32241), .B(n32242), .Z(n32201) );
  AND U30932 ( .A(n1958), .B(n32243), .Z(n32241) );
  XOR U30933 ( .A(n32244), .B(n32242), .Z(n32243) );
  XNOR U30934 ( .A(n32245), .B(n32246), .Z(n32233) );
  NAND U30935 ( .A(n32247), .B(n32248), .Z(n32246) );
  XOR U30936 ( .A(n32249), .B(n32225), .Z(n32248) );
  XOR U30937 ( .A(n32239), .B(n32240), .Z(n32225) );
  XOR U30938 ( .A(n32250), .B(n32251), .Z(n32240) );
  ANDN U30939 ( .B(n32252), .A(n32253), .Z(n32250) );
  XOR U30940 ( .A(n32251), .B(n32254), .Z(n32252) );
  XOR U30941 ( .A(n32255), .B(n32256), .Z(n32239) );
  XOR U30942 ( .A(n32257), .B(n32258), .Z(n32256) );
  ANDN U30943 ( .B(n32259), .A(n32260), .Z(n32257) );
  XOR U30944 ( .A(n32261), .B(n32258), .Z(n32259) );
  IV U30945 ( .A(n32237), .Z(n32255) );
  XOR U30946 ( .A(n32262), .B(n32263), .Z(n32237) );
  ANDN U30947 ( .B(n32264), .A(n32265), .Z(n32262) );
  XOR U30948 ( .A(n32263), .B(n32266), .Z(n32264) );
  IV U30949 ( .A(n32245), .Z(n32249) );
  XOR U30950 ( .A(n32245), .B(n32227), .Z(n32247) );
  XOR U30951 ( .A(n32267), .B(n32268), .Z(n32227) );
  AND U30952 ( .A(n1958), .B(n32269), .Z(n32267) );
  XOR U30953 ( .A(n32270), .B(n32268), .Z(n32269) );
  NANDN U30954 ( .A(n32229), .B(n32231), .Z(n32245) );
  XOR U30955 ( .A(n32271), .B(n32272), .Z(n32231) );
  AND U30956 ( .A(n1958), .B(n32273), .Z(n32271) );
  XOR U30957 ( .A(n32272), .B(n32274), .Z(n32273) );
  XOR U30958 ( .A(n32275), .B(n32276), .Z(n1958) );
  AND U30959 ( .A(n32277), .B(n32278), .Z(n32275) );
  XNOR U30960 ( .A(n32276), .B(n32242), .Z(n32278) );
  XNOR U30961 ( .A(n32279), .B(n32280), .Z(n32242) );
  ANDN U30962 ( .B(n32281), .A(n32282), .Z(n32279) );
  XOR U30963 ( .A(n32280), .B(n32283), .Z(n32281) );
  XOR U30964 ( .A(n32276), .B(n32244), .Z(n32277) );
  XOR U30965 ( .A(n32284), .B(n32285), .Z(n32244) );
  AND U30966 ( .A(n1962), .B(n32286), .Z(n32284) );
  XOR U30967 ( .A(n32287), .B(n32285), .Z(n32286) );
  XNOR U30968 ( .A(n32288), .B(n32289), .Z(n32276) );
  NAND U30969 ( .A(n32290), .B(n32291), .Z(n32289) );
  XOR U30970 ( .A(n32292), .B(n32268), .Z(n32291) );
  XOR U30971 ( .A(n32282), .B(n32283), .Z(n32268) );
  XOR U30972 ( .A(n32293), .B(n32294), .Z(n32283) );
  ANDN U30973 ( .B(n32295), .A(n32296), .Z(n32293) );
  XOR U30974 ( .A(n32294), .B(n32297), .Z(n32295) );
  XOR U30975 ( .A(n32298), .B(n32299), .Z(n32282) );
  XOR U30976 ( .A(n32300), .B(n32301), .Z(n32299) );
  ANDN U30977 ( .B(n32302), .A(n32303), .Z(n32300) );
  XOR U30978 ( .A(n32304), .B(n32301), .Z(n32302) );
  IV U30979 ( .A(n32280), .Z(n32298) );
  XOR U30980 ( .A(n32305), .B(n32306), .Z(n32280) );
  ANDN U30981 ( .B(n32307), .A(n32308), .Z(n32305) );
  XOR U30982 ( .A(n32306), .B(n32309), .Z(n32307) );
  IV U30983 ( .A(n32288), .Z(n32292) );
  XOR U30984 ( .A(n32288), .B(n32270), .Z(n32290) );
  XOR U30985 ( .A(n32310), .B(n32311), .Z(n32270) );
  AND U30986 ( .A(n1962), .B(n32312), .Z(n32310) );
  XOR U30987 ( .A(n32313), .B(n32311), .Z(n32312) );
  NANDN U30988 ( .A(n32272), .B(n32274), .Z(n32288) );
  XOR U30989 ( .A(n32314), .B(n32315), .Z(n32274) );
  AND U30990 ( .A(n1962), .B(n32316), .Z(n32314) );
  XOR U30991 ( .A(n32315), .B(n32317), .Z(n32316) );
  XOR U30992 ( .A(n32318), .B(n32319), .Z(n1962) );
  AND U30993 ( .A(n32320), .B(n32321), .Z(n32318) );
  XNOR U30994 ( .A(n32319), .B(n32285), .Z(n32321) );
  XNOR U30995 ( .A(n32322), .B(n32323), .Z(n32285) );
  ANDN U30996 ( .B(n32324), .A(n32325), .Z(n32322) );
  XOR U30997 ( .A(n32323), .B(n32326), .Z(n32324) );
  XOR U30998 ( .A(n32319), .B(n32287), .Z(n32320) );
  XOR U30999 ( .A(n32327), .B(n32328), .Z(n32287) );
  AND U31000 ( .A(n1966), .B(n32329), .Z(n32327) );
  XOR U31001 ( .A(n32330), .B(n32328), .Z(n32329) );
  XNOR U31002 ( .A(n32331), .B(n32332), .Z(n32319) );
  NAND U31003 ( .A(n32333), .B(n32334), .Z(n32332) );
  XOR U31004 ( .A(n32335), .B(n32311), .Z(n32334) );
  XOR U31005 ( .A(n32325), .B(n32326), .Z(n32311) );
  XOR U31006 ( .A(n32336), .B(n32337), .Z(n32326) );
  ANDN U31007 ( .B(n32338), .A(n32339), .Z(n32336) );
  XOR U31008 ( .A(n32337), .B(n32340), .Z(n32338) );
  XOR U31009 ( .A(n32341), .B(n32342), .Z(n32325) );
  XOR U31010 ( .A(n32343), .B(n32344), .Z(n32342) );
  ANDN U31011 ( .B(n32345), .A(n32346), .Z(n32343) );
  XOR U31012 ( .A(n32347), .B(n32344), .Z(n32345) );
  IV U31013 ( .A(n32323), .Z(n32341) );
  XOR U31014 ( .A(n32348), .B(n32349), .Z(n32323) );
  ANDN U31015 ( .B(n32350), .A(n32351), .Z(n32348) );
  XOR U31016 ( .A(n32349), .B(n32352), .Z(n32350) );
  IV U31017 ( .A(n32331), .Z(n32335) );
  XOR U31018 ( .A(n32331), .B(n32313), .Z(n32333) );
  XOR U31019 ( .A(n32353), .B(n32354), .Z(n32313) );
  AND U31020 ( .A(n1966), .B(n32355), .Z(n32353) );
  XOR U31021 ( .A(n32356), .B(n32354), .Z(n32355) );
  NANDN U31022 ( .A(n32315), .B(n32317), .Z(n32331) );
  XOR U31023 ( .A(n32357), .B(n32358), .Z(n32317) );
  AND U31024 ( .A(n1966), .B(n32359), .Z(n32357) );
  XOR U31025 ( .A(n32358), .B(n32360), .Z(n32359) );
  XOR U31026 ( .A(n32361), .B(n32362), .Z(n1966) );
  AND U31027 ( .A(n32363), .B(n32364), .Z(n32361) );
  XNOR U31028 ( .A(n32362), .B(n32328), .Z(n32364) );
  XNOR U31029 ( .A(n32365), .B(n32366), .Z(n32328) );
  ANDN U31030 ( .B(n32367), .A(n32368), .Z(n32365) );
  XOR U31031 ( .A(n32366), .B(n32369), .Z(n32367) );
  XOR U31032 ( .A(n32362), .B(n32330), .Z(n32363) );
  XOR U31033 ( .A(n32370), .B(n32371), .Z(n32330) );
  AND U31034 ( .A(n1970), .B(n32372), .Z(n32370) );
  XOR U31035 ( .A(n32373), .B(n32371), .Z(n32372) );
  XNOR U31036 ( .A(n32374), .B(n32375), .Z(n32362) );
  NAND U31037 ( .A(n32376), .B(n32377), .Z(n32375) );
  XOR U31038 ( .A(n32378), .B(n32354), .Z(n32377) );
  XOR U31039 ( .A(n32368), .B(n32369), .Z(n32354) );
  XOR U31040 ( .A(n32379), .B(n32380), .Z(n32369) );
  ANDN U31041 ( .B(n32381), .A(n32382), .Z(n32379) );
  XOR U31042 ( .A(n32380), .B(n32383), .Z(n32381) );
  XOR U31043 ( .A(n32384), .B(n32385), .Z(n32368) );
  XOR U31044 ( .A(n32386), .B(n32387), .Z(n32385) );
  ANDN U31045 ( .B(n32388), .A(n32389), .Z(n32386) );
  XOR U31046 ( .A(n32390), .B(n32387), .Z(n32388) );
  IV U31047 ( .A(n32366), .Z(n32384) );
  XOR U31048 ( .A(n32391), .B(n32392), .Z(n32366) );
  ANDN U31049 ( .B(n32393), .A(n32394), .Z(n32391) );
  XOR U31050 ( .A(n32392), .B(n32395), .Z(n32393) );
  IV U31051 ( .A(n32374), .Z(n32378) );
  XOR U31052 ( .A(n32374), .B(n32356), .Z(n32376) );
  XOR U31053 ( .A(n32396), .B(n32397), .Z(n32356) );
  AND U31054 ( .A(n1970), .B(n32398), .Z(n32396) );
  XOR U31055 ( .A(n32399), .B(n32397), .Z(n32398) );
  NANDN U31056 ( .A(n32358), .B(n32360), .Z(n32374) );
  XOR U31057 ( .A(n32400), .B(n32401), .Z(n32360) );
  AND U31058 ( .A(n1970), .B(n32402), .Z(n32400) );
  XOR U31059 ( .A(n32401), .B(n32403), .Z(n32402) );
  XOR U31060 ( .A(n32404), .B(n32405), .Z(n1970) );
  AND U31061 ( .A(n32406), .B(n32407), .Z(n32404) );
  XNOR U31062 ( .A(n32405), .B(n32371), .Z(n32407) );
  XNOR U31063 ( .A(n32408), .B(n32409), .Z(n32371) );
  ANDN U31064 ( .B(n32410), .A(n32411), .Z(n32408) );
  XOR U31065 ( .A(n32409), .B(n32412), .Z(n32410) );
  XOR U31066 ( .A(n32405), .B(n32373), .Z(n32406) );
  XOR U31067 ( .A(n32413), .B(n32414), .Z(n32373) );
  AND U31068 ( .A(n1974), .B(n32415), .Z(n32413) );
  XOR U31069 ( .A(n32416), .B(n32414), .Z(n32415) );
  XNOR U31070 ( .A(n32417), .B(n32418), .Z(n32405) );
  NAND U31071 ( .A(n32419), .B(n32420), .Z(n32418) );
  XOR U31072 ( .A(n32421), .B(n32397), .Z(n32420) );
  XOR U31073 ( .A(n32411), .B(n32412), .Z(n32397) );
  XOR U31074 ( .A(n32422), .B(n32423), .Z(n32412) );
  ANDN U31075 ( .B(n32424), .A(n32425), .Z(n32422) );
  XOR U31076 ( .A(n32423), .B(n32426), .Z(n32424) );
  XOR U31077 ( .A(n32427), .B(n32428), .Z(n32411) );
  XOR U31078 ( .A(n32429), .B(n32430), .Z(n32428) );
  ANDN U31079 ( .B(n32431), .A(n32432), .Z(n32429) );
  XOR U31080 ( .A(n32433), .B(n32430), .Z(n32431) );
  IV U31081 ( .A(n32409), .Z(n32427) );
  XOR U31082 ( .A(n32434), .B(n32435), .Z(n32409) );
  ANDN U31083 ( .B(n32436), .A(n32437), .Z(n32434) );
  XOR U31084 ( .A(n32435), .B(n32438), .Z(n32436) );
  IV U31085 ( .A(n32417), .Z(n32421) );
  XOR U31086 ( .A(n32417), .B(n32399), .Z(n32419) );
  XOR U31087 ( .A(n32439), .B(n32440), .Z(n32399) );
  AND U31088 ( .A(n1974), .B(n32441), .Z(n32439) );
  XOR U31089 ( .A(n32442), .B(n32440), .Z(n32441) );
  NANDN U31090 ( .A(n32401), .B(n32403), .Z(n32417) );
  XOR U31091 ( .A(n32443), .B(n32444), .Z(n32403) );
  AND U31092 ( .A(n1974), .B(n32445), .Z(n32443) );
  XOR U31093 ( .A(n32444), .B(n32446), .Z(n32445) );
  XOR U31094 ( .A(n32447), .B(n32448), .Z(n1974) );
  AND U31095 ( .A(n32449), .B(n32450), .Z(n32447) );
  XNOR U31096 ( .A(n32448), .B(n32414), .Z(n32450) );
  XNOR U31097 ( .A(n32451), .B(n32452), .Z(n32414) );
  ANDN U31098 ( .B(n32453), .A(n32454), .Z(n32451) );
  XOR U31099 ( .A(n32452), .B(n32455), .Z(n32453) );
  XOR U31100 ( .A(n32448), .B(n32416), .Z(n32449) );
  XOR U31101 ( .A(n32456), .B(n32457), .Z(n32416) );
  AND U31102 ( .A(n1978), .B(n32458), .Z(n32456) );
  XOR U31103 ( .A(n32459), .B(n32457), .Z(n32458) );
  XNOR U31104 ( .A(n32460), .B(n32461), .Z(n32448) );
  NAND U31105 ( .A(n32462), .B(n32463), .Z(n32461) );
  XOR U31106 ( .A(n32464), .B(n32440), .Z(n32463) );
  XOR U31107 ( .A(n32454), .B(n32455), .Z(n32440) );
  XOR U31108 ( .A(n32465), .B(n32466), .Z(n32455) );
  ANDN U31109 ( .B(n32467), .A(n32468), .Z(n32465) );
  XOR U31110 ( .A(n32466), .B(n32469), .Z(n32467) );
  XOR U31111 ( .A(n32470), .B(n32471), .Z(n32454) );
  XOR U31112 ( .A(n32472), .B(n32473), .Z(n32471) );
  ANDN U31113 ( .B(n32474), .A(n32475), .Z(n32472) );
  XOR U31114 ( .A(n32476), .B(n32473), .Z(n32474) );
  IV U31115 ( .A(n32452), .Z(n32470) );
  XOR U31116 ( .A(n32477), .B(n32478), .Z(n32452) );
  ANDN U31117 ( .B(n32479), .A(n32480), .Z(n32477) );
  XOR U31118 ( .A(n32478), .B(n32481), .Z(n32479) );
  IV U31119 ( .A(n32460), .Z(n32464) );
  XOR U31120 ( .A(n32460), .B(n32442), .Z(n32462) );
  XOR U31121 ( .A(n32482), .B(n32483), .Z(n32442) );
  AND U31122 ( .A(n1978), .B(n32484), .Z(n32482) );
  XOR U31123 ( .A(n32485), .B(n32483), .Z(n32484) );
  NANDN U31124 ( .A(n32444), .B(n32446), .Z(n32460) );
  XOR U31125 ( .A(n32486), .B(n32487), .Z(n32446) );
  AND U31126 ( .A(n1978), .B(n32488), .Z(n32486) );
  XOR U31127 ( .A(n32487), .B(n32489), .Z(n32488) );
  XOR U31128 ( .A(n32490), .B(n32491), .Z(n1978) );
  AND U31129 ( .A(n32492), .B(n32493), .Z(n32490) );
  XNOR U31130 ( .A(n32491), .B(n32457), .Z(n32493) );
  XNOR U31131 ( .A(n32494), .B(n32495), .Z(n32457) );
  ANDN U31132 ( .B(n32496), .A(n32497), .Z(n32494) );
  XOR U31133 ( .A(n32495), .B(n32498), .Z(n32496) );
  XOR U31134 ( .A(n32491), .B(n32459), .Z(n32492) );
  XOR U31135 ( .A(n32499), .B(n32500), .Z(n32459) );
  AND U31136 ( .A(n1982), .B(n32501), .Z(n32499) );
  XOR U31137 ( .A(n32502), .B(n32500), .Z(n32501) );
  XNOR U31138 ( .A(n32503), .B(n32504), .Z(n32491) );
  NAND U31139 ( .A(n32505), .B(n32506), .Z(n32504) );
  XOR U31140 ( .A(n32507), .B(n32483), .Z(n32506) );
  XOR U31141 ( .A(n32497), .B(n32498), .Z(n32483) );
  XOR U31142 ( .A(n32508), .B(n32509), .Z(n32498) );
  ANDN U31143 ( .B(n32510), .A(n32511), .Z(n32508) );
  XOR U31144 ( .A(n32509), .B(n32512), .Z(n32510) );
  XOR U31145 ( .A(n32513), .B(n32514), .Z(n32497) );
  XOR U31146 ( .A(n32515), .B(n32516), .Z(n32514) );
  ANDN U31147 ( .B(n32517), .A(n32518), .Z(n32515) );
  XOR U31148 ( .A(n32519), .B(n32516), .Z(n32517) );
  IV U31149 ( .A(n32495), .Z(n32513) );
  XOR U31150 ( .A(n32520), .B(n32521), .Z(n32495) );
  ANDN U31151 ( .B(n32522), .A(n32523), .Z(n32520) );
  XOR U31152 ( .A(n32521), .B(n32524), .Z(n32522) );
  IV U31153 ( .A(n32503), .Z(n32507) );
  XOR U31154 ( .A(n32503), .B(n32485), .Z(n32505) );
  XOR U31155 ( .A(n32525), .B(n32526), .Z(n32485) );
  AND U31156 ( .A(n1982), .B(n32527), .Z(n32525) );
  XOR U31157 ( .A(n32528), .B(n32526), .Z(n32527) );
  NANDN U31158 ( .A(n32487), .B(n32489), .Z(n32503) );
  XOR U31159 ( .A(n32529), .B(n32530), .Z(n32489) );
  AND U31160 ( .A(n1982), .B(n32531), .Z(n32529) );
  XOR U31161 ( .A(n32530), .B(n32532), .Z(n32531) );
  XOR U31162 ( .A(n32533), .B(n32534), .Z(n1982) );
  AND U31163 ( .A(n32535), .B(n32536), .Z(n32533) );
  XNOR U31164 ( .A(n32534), .B(n32500), .Z(n32536) );
  XNOR U31165 ( .A(n32537), .B(n32538), .Z(n32500) );
  ANDN U31166 ( .B(n32539), .A(n32540), .Z(n32537) );
  XOR U31167 ( .A(n32538), .B(n32541), .Z(n32539) );
  XOR U31168 ( .A(n32534), .B(n32502), .Z(n32535) );
  XOR U31169 ( .A(n32542), .B(n32543), .Z(n32502) );
  AND U31170 ( .A(n1986), .B(n32544), .Z(n32542) );
  XOR U31171 ( .A(n32545), .B(n32543), .Z(n32544) );
  XNOR U31172 ( .A(n32546), .B(n32547), .Z(n32534) );
  NAND U31173 ( .A(n32548), .B(n32549), .Z(n32547) );
  XOR U31174 ( .A(n32550), .B(n32526), .Z(n32549) );
  XOR U31175 ( .A(n32540), .B(n32541), .Z(n32526) );
  XOR U31176 ( .A(n32551), .B(n32552), .Z(n32541) );
  ANDN U31177 ( .B(n32553), .A(n32554), .Z(n32551) );
  XOR U31178 ( .A(n32552), .B(n32555), .Z(n32553) );
  XOR U31179 ( .A(n32556), .B(n32557), .Z(n32540) );
  XOR U31180 ( .A(n32558), .B(n32559), .Z(n32557) );
  ANDN U31181 ( .B(n32560), .A(n32561), .Z(n32558) );
  XOR U31182 ( .A(n32562), .B(n32559), .Z(n32560) );
  IV U31183 ( .A(n32538), .Z(n32556) );
  XOR U31184 ( .A(n32563), .B(n32564), .Z(n32538) );
  ANDN U31185 ( .B(n32565), .A(n32566), .Z(n32563) );
  XOR U31186 ( .A(n32564), .B(n32567), .Z(n32565) );
  IV U31187 ( .A(n32546), .Z(n32550) );
  XOR U31188 ( .A(n32546), .B(n32528), .Z(n32548) );
  XOR U31189 ( .A(n32568), .B(n32569), .Z(n32528) );
  AND U31190 ( .A(n1986), .B(n32570), .Z(n32568) );
  XOR U31191 ( .A(n32571), .B(n32569), .Z(n32570) );
  NANDN U31192 ( .A(n32530), .B(n32532), .Z(n32546) );
  XOR U31193 ( .A(n32572), .B(n32573), .Z(n32532) );
  AND U31194 ( .A(n1986), .B(n32574), .Z(n32572) );
  XOR U31195 ( .A(n32573), .B(n32575), .Z(n32574) );
  XOR U31196 ( .A(n32576), .B(n32577), .Z(n1986) );
  AND U31197 ( .A(n32578), .B(n32579), .Z(n32576) );
  XNOR U31198 ( .A(n32577), .B(n32543), .Z(n32579) );
  XNOR U31199 ( .A(n32580), .B(n32581), .Z(n32543) );
  ANDN U31200 ( .B(n32582), .A(n32583), .Z(n32580) );
  XOR U31201 ( .A(n32581), .B(n32584), .Z(n32582) );
  XOR U31202 ( .A(n32577), .B(n32545), .Z(n32578) );
  XOR U31203 ( .A(n32585), .B(n32586), .Z(n32545) );
  AND U31204 ( .A(n1990), .B(n32587), .Z(n32585) );
  XOR U31205 ( .A(n32588), .B(n32586), .Z(n32587) );
  XNOR U31206 ( .A(n32589), .B(n32590), .Z(n32577) );
  NAND U31207 ( .A(n32591), .B(n32592), .Z(n32590) );
  XOR U31208 ( .A(n32593), .B(n32569), .Z(n32592) );
  XOR U31209 ( .A(n32583), .B(n32584), .Z(n32569) );
  XOR U31210 ( .A(n32594), .B(n32595), .Z(n32584) );
  ANDN U31211 ( .B(n32596), .A(n32597), .Z(n32594) );
  XOR U31212 ( .A(n32595), .B(n32598), .Z(n32596) );
  XOR U31213 ( .A(n32599), .B(n32600), .Z(n32583) );
  XOR U31214 ( .A(n32601), .B(n32602), .Z(n32600) );
  ANDN U31215 ( .B(n32603), .A(n32604), .Z(n32601) );
  XOR U31216 ( .A(n32605), .B(n32602), .Z(n32603) );
  IV U31217 ( .A(n32581), .Z(n32599) );
  XOR U31218 ( .A(n32606), .B(n32607), .Z(n32581) );
  ANDN U31219 ( .B(n32608), .A(n32609), .Z(n32606) );
  XOR U31220 ( .A(n32607), .B(n32610), .Z(n32608) );
  IV U31221 ( .A(n32589), .Z(n32593) );
  XOR U31222 ( .A(n32589), .B(n32571), .Z(n32591) );
  XOR U31223 ( .A(n32611), .B(n32612), .Z(n32571) );
  AND U31224 ( .A(n1990), .B(n32613), .Z(n32611) );
  XOR U31225 ( .A(n32614), .B(n32612), .Z(n32613) );
  NANDN U31226 ( .A(n32573), .B(n32575), .Z(n32589) );
  XOR U31227 ( .A(n32615), .B(n32616), .Z(n32575) );
  AND U31228 ( .A(n1990), .B(n32617), .Z(n32615) );
  XOR U31229 ( .A(n32616), .B(n32618), .Z(n32617) );
  XOR U31230 ( .A(n32619), .B(n32620), .Z(n1990) );
  AND U31231 ( .A(n32621), .B(n32622), .Z(n32619) );
  XNOR U31232 ( .A(n32620), .B(n32586), .Z(n32622) );
  XNOR U31233 ( .A(n32623), .B(n32624), .Z(n32586) );
  ANDN U31234 ( .B(n32625), .A(n32626), .Z(n32623) );
  XOR U31235 ( .A(n32624), .B(n32627), .Z(n32625) );
  XOR U31236 ( .A(n32620), .B(n32588), .Z(n32621) );
  XOR U31237 ( .A(n32628), .B(n32629), .Z(n32588) );
  AND U31238 ( .A(n1994), .B(n32630), .Z(n32628) );
  XOR U31239 ( .A(n32631), .B(n32629), .Z(n32630) );
  XNOR U31240 ( .A(n32632), .B(n32633), .Z(n32620) );
  NAND U31241 ( .A(n32634), .B(n32635), .Z(n32633) );
  XOR U31242 ( .A(n32636), .B(n32612), .Z(n32635) );
  XOR U31243 ( .A(n32626), .B(n32627), .Z(n32612) );
  XOR U31244 ( .A(n32637), .B(n32638), .Z(n32627) );
  ANDN U31245 ( .B(n32639), .A(n32640), .Z(n32637) );
  XOR U31246 ( .A(n32638), .B(n32641), .Z(n32639) );
  XOR U31247 ( .A(n32642), .B(n32643), .Z(n32626) );
  XOR U31248 ( .A(n32644), .B(n32645), .Z(n32643) );
  ANDN U31249 ( .B(n32646), .A(n32647), .Z(n32644) );
  XOR U31250 ( .A(n32648), .B(n32645), .Z(n32646) );
  IV U31251 ( .A(n32624), .Z(n32642) );
  XOR U31252 ( .A(n32649), .B(n32650), .Z(n32624) );
  ANDN U31253 ( .B(n32651), .A(n32652), .Z(n32649) );
  XOR U31254 ( .A(n32650), .B(n32653), .Z(n32651) );
  IV U31255 ( .A(n32632), .Z(n32636) );
  XOR U31256 ( .A(n32632), .B(n32614), .Z(n32634) );
  XOR U31257 ( .A(n32654), .B(n32655), .Z(n32614) );
  AND U31258 ( .A(n1994), .B(n32656), .Z(n32654) );
  XOR U31259 ( .A(n32657), .B(n32655), .Z(n32656) );
  NANDN U31260 ( .A(n32616), .B(n32618), .Z(n32632) );
  XOR U31261 ( .A(n32658), .B(n32659), .Z(n32618) );
  AND U31262 ( .A(n1994), .B(n32660), .Z(n32658) );
  XOR U31263 ( .A(n32659), .B(n32661), .Z(n32660) );
  XOR U31264 ( .A(n32662), .B(n32663), .Z(n1994) );
  AND U31265 ( .A(n32664), .B(n32665), .Z(n32662) );
  XNOR U31266 ( .A(n32663), .B(n32629), .Z(n32665) );
  XNOR U31267 ( .A(n32666), .B(n32667), .Z(n32629) );
  ANDN U31268 ( .B(n32668), .A(n32669), .Z(n32666) );
  XOR U31269 ( .A(n32667), .B(n32670), .Z(n32668) );
  XOR U31270 ( .A(n32663), .B(n32631), .Z(n32664) );
  XOR U31271 ( .A(n32671), .B(n32672), .Z(n32631) );
  AND U31272 ( .A(n1998), .B(n32673), .Z(n32671) );
  XOR U31273 ( .A(n32674), .B(n32672), .Z(n32673) );
  XNOR U31274 ( .A(n32675), .B(n32676), .Z(n32663) );
  NAND U31275 ( .A(n32677), .B(n32678), .Z(n32676) );
  XOR U31276 ( .A(n32679), .B(n32655), .Z(n32678) );
  XOR U31277 ( .A(n32669), .B(n32670), .Z(n32655) );
  XOR U31278 ( .A(n32680), .B(n32681), .Z(n32670) );
  ANDN U31279 ( .B(n32682), .A(n32683), .Z(n32680) );
  XOR U31280 ( .A(n32681), .B(n32684), .Z(n32682) );
  XOR U31281 ( .A(n32685), .B(n32686), .Z(n32669) );
  XOR U31282 ( .A(n32687), .B(n32688), .Z(n32686) );
  ANDN U31283 ( .B(n32689), .A(n32690), .Z(n32687) );
  XOR U31284 ( .A(n32691), .B(n32688), .Z(n32689) );
  IV U31285 ( .A(n32667), .Z(n32685) );
  XOR U31286 ( .A(n32692), .B(n32693), .Z(n32667) );
  ANDN U31287 ( .B(n32694), .A(n32695), .Z(n32692) );
  XOR U31288 ( .A(n32693), .B(n32696), .Z(n32694) );
  IV U31289 ( .A(n32675), .Z(n32679) );
  XOR U31290 ( .A(n32675), .B(n32657), .Z(n32677) );
  XOR U31291 ( .A(n32697), .B(n32698), .Z(n32657) );
  AND U31292 ( .A(n1998), .B(n32699), .Z(n32697) );
  XOR U31293 ( .A(n32700), .B(n32698), .Z(n32699) );
  NANDN U31294 ( .A(n32659), .B(n32661), .Z(n32675) );
  XOR U31295 ( .A(n32701), .B(n32702), .Z(n32661) );
  AND U31296 ( .A(n1998), .B(n32703), .Z(n32701) );
  XOR U31297 ( .A(n32702), .B(n32704), .Z(n32703) );
  XOR U31298 ( .A(n32705), .B(n32706), .Z(n1998) );
  AND U31299 ( .A(n32707), .B(n32708), .Z(n32705) );
  XNOR U31300 ( .A(n32706), .B(n32672), .Z(n32708) );
  XNOR U31301 ( .A(n32709), .B(n32710), .Z(n32672) );
  ANDN U31302 ( .B(n32711), .A(n32712), .Z(n32709) );
  XOR U31303 ( .A(n32710), .B(n32713), .Z(n32711) );
  XOR U31304 ( .A(n32706), .B(n32674), .Z(n32707) );
  XOR U31305 ( .A(n32714), .B(n32715), .Z(n32674) );
  AND U31306 ( .A(n2002), .B(n32716), .Z(n32714) );
  XOR U31307 ( .A(n32717), .B(n32715), .Z(n32716) );
  XNOR U31308 ( .A(n32718), .B(n32719), .Z(n32706) );
  NAND U31309 ( .A(n32720), .B(n32721), .Z(n32719) );
  XOR U31310 ( .A(n32722), .B(n32698), .Z(n32721) );
  XOR U31311 ( .A(n32712), .B(n32713), .Z(n32698) );
  XOR U31312 ( .A(n32723), .B(n32724), .Z(n32713) );
  ANDN U31313 ( .B(n32725), .A(n32726), .Z(n32723) );
  XOR U31314 ( .A(n32724), .B(n32727), .Z(n32725) );
  XOR U31315 ( .A(n32728), .B(n32729), .Z(n32712) );
  XOR U31316 ( .A(n32730), .B(n32731), .Z(n32729) );
  ANDN U31317 ( .B(n32732), .A(n32733), .Z(n32730) );
  XOR U31318 ( .A(n32734), .B(n32731), .Z(n32732) );
  IV U31319 ( .A(n32710), .Z(n32728) );
  XOR U31320 ( .A(n32735), .B(n32736), .Z(n32710) );
  ANDN U31321 ( .B(n32737), .A(n32738), .Z(n32735) );
  XOR U31322 ( .A(n32736), .B(n32739), .Z(n32737) );
  IV U31323 ( .A(n32718), .Z(n32722) );
  XOR U31324 ( .A(n32718), .B(n32700), .Z(n32720) );
  XOR U31325 ( .A(n32740), .B(n32741), .Z(n32700) );
  AND U31326 ( .A(n2002), .B(n32742), .Z(n32740) );
  XOR U31327 ( .A(n32743), .B(n32741), .Z(n32742) );
  NANDN U31328 ( .A(n32702), .B(n32704), .Z(n32718) );
  XOR U31329 ( .A(n32744), .B(n32745), .Z(n32704) );
  AND U31330 ( .A(n2002), .B(n32746), .Z(n32744) );
  XOR U31331 ( .A(n32745), .B(n32747), .Z(n32746) );
  XOR U31332 ( .A(n32748), .B(n32749), .Z(n2002) );
  AND U31333 ( .A(n32750), .B(n32751), .Z(n32748) );
  XNOR U31334 ( .A(n32749), .B(n32715), .Z(n32751) );
  XNOR U31335 ( .A(n32752), .B(n32753), .Z(n32715) );
  ANDN U31336 ( .B(n32754), .A(n32755), .Z(n32752) );
  XOR U31337 ( .A(n32753), .B(n32756), .Z(n32754) );
  XOR U31338 ( .A(n32749), .B(n32717), .Z(n32750) );
  XOR U31339 ( .A(n32757), .B(n32758), .Z(n32717) );
  AND U31340 ( .A(n2006), .B(n32759), .Z(n32757) );
  XOR U31341 ( .A(n32760), .B(n32758), .Z(n32759) );
  XNOR U31342 ( .A(n32761), .B(n32762), .Z(n32749) );
  NAND U31343 ( .A(n32763), .B(n32764), .Z(n32762) );
  XOR U31344 ( .A(n32765), .B(n32741), .Z(n32764) );
  XOR U31345 ( .A(n32755), .B(n32756), .Z(n32741) );
  XOR U31346 ( .A(n32766), .B(n32767), .Z(n32756) );
  ANDN U31347 ( .B(n32768), .A(n32769), .Z(n32766) );
  XOR U31348 ( .A(n32767), .B(n32770), .Z(n32768) );
  XOR U31349 ( .A(n32771), .B(n32772), .Z(n32755) );
  XOR U31350 ( .A(n32773), .B(n32774), .Z(n32772) );
  ANDN U31351 ( .B(n32775), .A(n32776), .Z(n32773) );
  XOR U31352 ( .A(n32777), .B(n32774), .Z(n32775) );
  IV U31353 ( .A(n32753), .Z(n32771) );
  XOR U31354 ( .A(n32778), .B(n32779), .Z(n32753) );
  ANDN U31355 ( .B(n32780), .A(n32781), .Z(n32778) );
  XOR U31356 ( .A(n32779), .B(n32782), .Z(n32780) );
  IV U31357 ( .A(n32761), .Z(n32765) );
  XOR U31358 ( .A(n32761), .B(n32743), .Z(n32763) );
  XOR U31359 ( .A(n32783), .B(n32784), .Z(n32743) );
  AND U31360 ( .A(n2006), .B(n32785), .Z(n32783) );
  XOR U31361 ( .A(n32786), .B(n32784), .Z(n32785) );
  NANDN U31362 ( .A(n32745), .B(n32747), .Z(n32761) );
  XOR U31363 ( .A(n32787), .B(n32788), .Z(n32747) );
  AND U31364 ( .A(n2006), .B(n32789), .Z(n32787) );
  XOR U31365 ( .A(n32788), .B(n32790), .Z(n32789) );
  XOR U31366 ( .A(n32791), .B(n32792), .Z(n2006) );
  AND U31367 ( .A(n32793), .B(n32794), .Z(n32791) );
  XNOR U31368 ( .A(n32792), .B(n32758), .Z(n32794) );
  XNOR U31369 ( .A(n32795), .B(n32796), .Z(n32758) );
  ANDN U31370 ( .B(n32797), .A(n32798), .Z(n32795) );
  XOR U31371 ( .A(n32796), .B(n32799), .Z(n32797) );
  XOR U31372 ( .A(n32792), .B(n32760), .Z(n32793) );
  XOR U31373 ( .A(n32800), .B(n32801), .Z(n32760) );
  AND U31374 ( .A(n2010), .B(n32802), .Z(n32800) );
  XOR U31375 ( .A(n32803), .B(n32801), .Z(n32802) );
  XNOR U31376 ( .A(n32804), .B(n32805), .Z(n32792) );
  NAND U31377 ( .A(n32806), .B(n32807), .Z(n32805) );
  XOR U31378 ( .A(n32808), .B(n32784), .Z(n32807) );
  XOR U31379 ( .A(n32798), .B(n32799), .Z(n32784) );
  XOR U31380 ( .A(n32809), .B(n32810), .Z(n32799) );
  ANDN U31381 ( .B(n32811), .A(n32812), .Z(n32809) );
  XOR U31382 ( .A(n32810), .B(n32813), .Z(n32811) );
  XOR U31383 ( .A(n32814), .B(n32815), .Z(n32798) );
  XOR U31384 ( .A(n32816), .B(n32817), .Z(n32815) );
  ANDN U31385 ( .B(n32818), .A(n32819), .Z(n32816) );
  XOR U31386 ( .A(n32820), .B(n32817), .Z(n32818) );
  IV U31387 ( .A(n32796), .Z(n32814) );
  XOR U31388 ( .A(n32821), .B(n32822), .Z(n32796) );
  ANDN U31389 ( .B(n32823), .A(n32824), .Z(n32821) );
  XOR U31390 ( .A(n32822), .B(n32825), .Z(n32823) );
  IV U31391 ( .A(n32804), .Z(n32808) );
  XOR U31392 ( .A(n32804), .B(n32786), .Z(n32806) );
  XOR U31393 ( .A(n32826), .B(n32827), .Z(n32786) );
  AND U31394 ( .A(n2010), .B(n32828), .Z(n32826) );
  XOR U31395 ( .A(n32829), .B(n32827), .Z(n32828) );
  NANDN U31396 ( .A(n32788), .B(n32790), .Z(n32804) );
  XOR U31397 ( .A(n32830), .B(n32831), .Z(n32790) );
  AND U31398 ( .A(n2010), .B(n32832), .Z(n32830) );
  XOR U31399 ( .A(n32831), .B(n32833), .Z(n32832) );
  XOR U31400 ( .A(n32834), .B(n32835), .Z(n2010) );
  AND U31401 ( .A(n32836), .B(n32837), .Z(n32834) );
  XNOR U31402 ( .A(n32835), .B(n32801), .Z(n32837) );
  XNOR U31403 ( .A(n32838), .B(n32839), .Z(n32801) );
  ANDN U31404 ( .B(n32840), .A(n32841), .Z(n32838) );
  XOR U31405 ( .A(n32839), .B(n32842), .Z(n32840) );
  XOR U31406 ( .A(n32835), .B(n32803), .Z(n32836) );
  XOR U31407 ( .A(n32843), .B(n32844), .Z(n32803) );
  AND U31408 ( .A(n2014), .B(n32845), .Z(n32843) );
  XOR U31409 ( .A(n32846), .B(n32844), .Z(n32845) );
  XNOR U31410 ( .A(n32847), .B(n32848), .Z(n32835) );
  NAND U31411 ( .A(n32849), .B(n32850), .Z(n32848) );
  XOR U31412 ( .A(n32851), .B(n32827), .Z(n32850) );
  XOR U31413 ( .A(n32841), .B(n32842), .Z(n32827) );
  XOR U31414 ( .A(n32852), .B(n32853), .Z(n32842) );
  ANDN U31415 ( .B(n32854), .A(n32855), .Z(n32852) );
  XOR U31416 ( .A(n32853), .B(n32856), .Z(n32854) );
  XOR U31417 ( .A(n32857), .B(n32858), .Z(n32841) );
  XOR U31418 ( .A(n32859), .B(n32860), .Z(n32858) );
  ANDN U31419 ( .B(n32861), .A(n32862), .Z(n32859) );
  XOR U31420 ( .A(n32863), .B(n32860), .Z(n32861) );
  IV U31421 ( .A(n32839), .Z(n32857) );
  XOR U31422 ( .A(n32864), .B(n32865), .Z(n32839) );
  ANDN U31423 ( .B(n32866), .A(n32867), .Z(n32864) );
  XOR U31424 ( .A(n32865), .B(n32868), .Z(n32866) );
  IV U31425 ( .A(n32847), .Z(n32851) );
  XOR U31426 ( .A(n32847), .B(n32829), .Z(n32849) );
  XOR U31427 ( .A(n32869), .B(n32870), .Z(n32829) );
  AND U31428 ( .A(n2014), .B(n32871), .Z(n32869) );
  XOR U31429 ( .A(n32872), .B(n32870), .Z(n32871) );
  NANDN U31430 ( .A(n32831), .B(n32833), .Z(n32847) );
  XOR U31431 ( .A(n32873), .B(n32874), .Z(n32833) );
  AND U31432 ( .A(n2014), .B(n32875), .Z(n32873) );
  XOR U31433 ( .A(n32874), .B(n32876), .Z(n32875) );
  XOR U31434 ( .A(n32877), .B(n32878), .Z(n2014) );
  AND U31435 ( .A(n32879), .B(n32880), .Z(n32877) );
  XNOR U31436 ( .A(n32878), .B(n32844), .Z(n32880) );
  XNOR U31437 ( .A(n32881), .B(n32882), .Z(n32844) );
  ANDN U31438 ( .B(n32883), .A(n32884), .Z(n32881) );
  XOR U31439 ( .A(n32882), .B(n32885), .Z(n32883) );
  XOR U31440 ( .A(n32878), .B(n32846), .Z(n32879) );
  XOR U31441 ( .A(n32886), .B(n32887), .Z(n32846) );
  AND U31442 ( .A(n2018), .B(n32888), .Z(n32886) );
  XOR U31443 ( .A(n32889), .B(n32887), .Z(n32888) );
  XNOR U31444 ( .A(n32890), .B(n32891), .Z(n32878) );
  NAND U31445 ( .A(n32892), .B(n32893), .Z(n32891) );
  XOR U31446 ( .A(n32894), .B(n32870), .Z(n32893) );
  XOR U31447 ( .A(n32884), .B(n32885), .Z(n32870) );
  XOR U31448 ( .A(n32895), .B(n32896), .Z(n32885) );
  ANDN U31449 ( .B(n32897), .A(n32898), .Z(n32895) );
  XOR U31450 ( .A(n32896), .B(n32899), .Z(n32897) );
  XOR U31451 ( .A(n32900), .B(n32901), .Z(n32884) );
  XOR U31452 ( .A(n32902), .B(n32903), .Z(n32901) );
  ANDN U31453 ( .B(n32904), .A(n32905), .Z(n32902) );
  XOR U31454 ( .A(n32906), .B(n32903), .Z(n32904) );
  IV U31455 ( .A(n32882), .Z(n32900) );
  XOR U31456 ( .A(n32907), .B(n32908), .Z(n32882) );
  ANDN U31457 ( .B(n32909), .A(n32910), .Z(n32907) );
  XOR U31458 ( .A(n32908), .B(n32911), .Z(n32909) );
  IV U31459 ( .A(n32890), .Z(n32894) );
  XOR U31460 ( .A(n32890), .B(n32872), .Z(n32892) );
  XOR U31461 ( .A(n32912), .B(n32913), .Z(n32872) );
  AND U31462 ( .A(n2018), .B(n32914), .Z(n32912) );
  XOR U31463 ( .A(n32915), .B(n32913), .Z(n32914) );
  NANDN U31464 ( .A(n32874), .B(n32876), .Z(n32890) );
  XOR U31465 ( .A(n32916), .B(n32917), .Z(n32876) );
  AND U31466 ( .A(n2018), .B(n32918), .Z(n32916) );
  XOR U31467 ( .A(n32917), .B(n32919), .Z(n32918) );
  XOR U31468 ( .A(n32920), .B(n32921), .Z(n2018) );
  AND U31469 ( .A(n32922), .B(n32923), .Z(n32920) );
  XNOR U31470 ( .A(n32921), .B(n32887), .Z(n32923) );
  XNOR U31471 ( .A(n32924), .B(n32925), .Z(n32887) );
  ANDN U31472 ( .B(n32926), .A(n32927), .Z(n32924) );
  XOR U31473 ( .A(n32925), .B(n32928), .Z(n32926) );
  XOR U31474 ( .A(n32921), .B(n32889), .Z(n32922) );
  XOR U31475 ( .A(n32929), .B(n32930), .Z(n32889) );
  AND U31476 ( .A(n2022), .B(n32931), .Z(n32929) );
  XOR U31477 ( .A(n32932), .B(n32930), .Z(n32931) );
  XNOR U31478 ( .A(n32933), .B(n32934), .Z(n32921) );
  NAND U31479 ( .A(n32935), .B(n32936), .Z(n32934) );
  XOR U31480 ( .A(n32937), .B(n32913), .Z(n32936) );
  XOR U31481 ( .A(n32927), .B(n32928), .Z(n32913) );
  XOR U31482 ( .A(n32938), .B(n32939), .Z(n32928) );
  ANDN U31483 ( .B(n32940), .A(n32941), .Z(n32938) );
  XOR U31484 ( .A(n32939), .B(n32942), .Z(n32940) );
  XOR U31485 ( .A(n32943), .B(n32944), .Z(n32927) );
  XOR U31486 ( .A(n32945), .B(n32946), .Z(n32944) );
  ANDN U31487 ( .B(n32947), .A(n32948), .Z(n32945) );
  XOR U31488 ( .A(n32949), .B(n32946), .Z(n32947) );
  IV U31489 ( .A(n32925), .Z(n32943) );
  XOR U31490 ( .A(n32950), .B(n32951), .Z(n32925) );
  ANDN U31491 ( .B(n32952), .A(n32953), .Z(n32950) );
  XOR U31492 ( .A(n32951), .B(n32954), .Z(n32952) );
  IV U31493 ( .A(n32933), .Z(n32937) );
  XOR U31494 ( .A(n32933), .B(n32915), .Z(n32935) );
  XOR U31495 ( .A(n32955), .B(n32956), .Z(n32915) );
  AND U31496 ( .A(n2022), .B(n32957), .Z(n32955) );
  XOR U31497 ( .A(n32958), .B(n32956), .Z(n32957) );
  NANDN U31498 ( .A(n32917), .B(n32919), .Z(n32933) );
  XOR U31499 ( .A(n32959), .B(n32960), .Z(n32919) );
  AND U31500 ( .A(n2022), .B(n32961), .Z(n32959) );
  XOR U31501 ( .A(n32960), .B(n32962), .Z(n32961) );
  XOR U31502 ( .A(n32963), .B(n32964), .Z(n2022) );
  AND U31503 ( .A(n32965), .B(n32966), .Z(n32963) );
  XNOR U31504 ( .A(n32964), .B(n32930), .Z(n32966) );
  XNOR U31505 ( .A(n32967), .B(n32968), .Z(n32930) );
  ANDN U31506 ( .B(n32969), .A(n32970), .Z(n32967) );
  XOR U31507 ( .A(n32968), .B(n32971), .Z(n32969) );
  XOR U31508 ( .A(n32964), .B(n32932), .Z(n32965) );
  XOR U31509 ( .A(n32972), .B(n32973), .Z(n32932) );
  AND U31510 ( .A(n2026), .B(n32974), .Z(n32972) );
  XOR U31511 ( .A(n32975), .B(n32973), .Z(n32974) );
  XNOR U31512 ( .A(n32976), .B(n32977), .Z(n32964) );
  NAND U31513 ( .A(n32978), .B(n32979), .Z(n32977) );
  XOR U31514 ( .A(n32980), .B(n32956), .Z(n32979) );
  XOR U31515 ( .A(n32970), .B(n32971), .Z(n32956) );
  XOR U31516 ( .A(n32981), .B(n32982), .Z(n32971) );
  ANDN U31517 ( .B(n32983), .A(n32984), .Z(n32981) );
  XOR U31518 ( .A(n32982), .B(n32985), .Z(n32983) );
  XOR U31519 ( .A(n32986), .B(n32987), .Z(n32970) );
  XOR U31520 ( .A(n32988), .B(n32989), .Z(n32987) );
  ANDN U31521 ( .B(n32990), .A(n32991), .Z(n32988) );
  XOR U31522 ( .A(n32992), .B(n32989), .Z(n32990) );
  IV U31523 ( .A(n32968), .Z(n32986) );
  XOR U31524 ( .A(n32993), .B(n32994), .Z(n32968) );
  ANDN U31525 ( .B(n32995), .A(n32996), .Z(n32993) );
  XOR U31526 ( .A(n32994), .B(n32997), .Z(n32995) );
  IV U31527 ( .A(n32976), .Z(n32980) );
  XOR U31528 ( .A(n32976), .B(n32958), .Z(n32978) );
  XOR U31529 ( .A(n32998), .B(n32999), .Z(n32958) );
  AND U31530 ( .A(n2026), .B(n33000), .Z(n32998) );
  XOR U31531 ( .A(n33001), .B(n32999), .Z(n33000) );
  NANDN U31532 ( .A(n32960), .B(n32962), .Z(n32976) );
  XOR U31533 ( .A(n33002), .B(n33003), .Z(n32962) );
  AND U31534 ( .A(n2026), .B(n33004), .Z(n33002) );
  XOR U31535 ( .A(n33003), .B(n33005), .Z(n33004) );
  XOR U31536 ( .A(n33006), .B(n33007), .Z(n2026) );
  AND U31537 ( .A(n33008), .B(n33009), .Z(n33006) );
  XNOR U31538 ( .A(n33007), .B(n32973), .Z(n33009) );
  XNOR U31539 ( .A(n33010), .B(n33011), .Z(n32973) );
  ANDN U31540 ( .B(n33012), .A(n33013), .Z(n33010) );
  XOR U31541 ( .A(n33011), .B(n33014), .Z(n33012) );
  XOR U31542 ( .A(n33007), .B(n32975), .Z(n33008) );
  XOR U31543 ( .A(n33015), .B(n33016), .Z(n32975) );
  AND U31544 ( .A(n2030), .B(n33017), .Z(n33015) );
  XOR U31545 ( .A(n33018), .B(n33016), .Z(n33017) );
  XNOR U31546 ( .A(n33019), .B(n33020), .Z(n33007) );
  NAND U31547 ( .A(n33021), .B(n33022), .Z(n33020) );
  XOR U31548 ( .A(n33023), .B(n32999), .Z(n33022) );
  XOR U31549 ( .A(n33013), .B(n33014), .Z(n32999) );
  XOR U31550 ( .A(n33024), .B(n33025), .Z(n33014) );
  ANDN U31551 ( .B(n33026), .A(n33027), .Z(n33024) );
  XOR U31552 ( .A(n33025), .B(n33028), .Z(n33026) );
  XOR U31553 ( .A(n33029), .B(n33030), .Z(n33013) );
  XOR U31554 ( .A(n33031), .B(n33032), .Z(n33030) );
  ANDN U31555 ( .B(n33033), .A(n33034), .Z(n33031) );
  XOR U31556 ( .A(n33035), .B(n33032), .Z(n33033) );
  IV U31557 ( .A(n33011), .Z(n33029) );
  XOR U31558 ( .A(n33036), .B(n33037), .Z(n33011) );
  ANDN U31559 ( .B(n33038), .A(n33039), .Z(n33036) );
  XOR U31560 ( .A(n33037), .B(n33040), .Z(n33038) );
  IV U31561 ( .A(n33019), .Z(n33023) );
  XOR U31562 ( .A(n33019), .B(n33001), .Z(n33021) );
  XOR U31563 ( .A(n33041), .B(n33042), .Z(n33001) );
  AND U31564 ( .A(n2030), .B(n33043), .Z(n33041) );
  XOR U31565 ( .A(n33044), .B(n33042), .Z(n33043) );
  NANDN U31566 ( .A(n33003), .B(n33005), .Z(n33019) );
  XOR U31567 ( .A(n33045), .B(n33046), .Z(n33005) );
  AND U31568 ( .A(n2030), .B(n33047), .Z(n33045) );
  XOR U31569 ( .A(n33046), .B(n33048), .Z(n33047) );
  XOR U31570 ( .A(n33049), .B(n33050), .Z(n2030) );
  AND U31571 ( .A(n33051), .B(n33052), .Z(n33049) );
  XNOR U31572 ( .A(n33050), .B(n33016), .Z(n33052) );
  XNOR U31573 ( .A(n33053), .B(n33054), .Z(n33016) );
  ANDN U31574 ( .B(n33055), .A(n33056), .Z(n33053) );
  XOR U31575 ( .A(n33054), .B(n33057), .Z(n33055) );
  XOR U31576 ( .A(n33050), .B(n33018), .Z(n33051) );
  XOR U31577 ( .A(n33058), .B(n33059), .Z(n33018) );
  AND U31578 ( .A(n2034), .B(n33060), .Z(n33058) );
  XOR U31579 ( .A(n33061), .B(n33059), .Z(n33060) );
  XNOR U31580 ( .A(n33062), .B(n33063), .Z(n33050) );
  NAND U31581 ( .A(n33064), .B(n33065), .Z(n33063) );
  XOR U31582 ( .A(n33066), .B(n33042), .Z(n33065) );
  XOR U31583 ( .A(n33056), .B(n33057), .Z(n33042) );
  XOR U31584 ( .A(n33067), .B(n33068), .Z(n33057) );
  ANDN U31585 ( .B(n33069), .A(n33070), .Z(n33067) );
  XOR U31586 ( .A(n33068), .B(n33071), .Z(n33069) );
  XOR U31587 ( .A(n33072), .B(n33073), .Z(n33056) );
  XOR U31588 ( .A(n33074), .B(n33075), .Z(n33073) );
  ANDN U31589 ( .B(n33076), .A(n33077), .Z(n33074) );
  XOR U31590 ( .A(n33078), .B(n33075), .Z(n33076) );
  IV U31591 ( .A(n33054), .Z(n33072) );
  XOR U31592 ( .A(n33079), .B(n33080), .Z(n33054) );
  ANDN U31593 ( .B(n33081), .A(n33082), .Z(n33079) );
  XOR U31594 ( .A(n33080), .B(n33083), .Z(n33081) );
  IV U31595 ( .A(n33062), .Z(n33066) );
  XOR U31596 ( .A(n33062), .B(n33044), .Z(n33064) );
  XOR U31597 ( .A(n33084), .B(n33085), .Z(n33044) );
  AND U31598 ( .A(n2034), .B(n33086), .Z(n33084) );
  XOR U31599 ( .A(n33087), .B(n33085), .Z(n33086) );
  NANDN U31600 ( .A(n33046), .B(n33048), .Z(n33062) );
  XOR U31601 ( .A(n33088), .B(n33089), .Z(n33048) );
  AND U31602 ( .A(n2034), .B(n33090), .Z(n33088) );
  XOR U31603 ( .A(n33089), .B(n33091), .Z(n33090) );
  XOR U31604 ( .A(n33092), .B(n33093), .Z(n2034) );
  AND U31605 ( .A(n33094), .B(n33095), .Z(n33092) );
  XNOR U31606 ( .A(n33093), .B(n33059), .Z(n33095) );
  XNOR U31607 ( .A(n33096), .B(n33097), .Z(n33059) );
  ANDN U31608 ( .B(n33098), .A(n33099), .Z(n33096) );
  XOR U31609 ( .A(n33097), .B(n33100), .Z(n33098) );
  XOR U31610 ( .A(n33093), .B(n33061), .Z(n33094) );
  XOR U31611 ( .A(n33101), .B(n33102), .Z(n33061) );
  AND U31612 ( .A(n2038), .B(n33103), .Z(n33101) );
  XOR U31613 ( .A(n33104), .B(n33102), .Z(n33103) );
  XNOR U31614 ( .A(n33105), .B(n33106), .Z(n33093) );
  NAND U31615 ( .A(n33107), .B(n33108), .Z(n33106) );
  XOR U31616 ( .A(n33109), .B(n33085), .Z(n33108) );
  XOR U31617 ( .A(n33099), .B(n33100), .Z(n33085) );
  XOR U31618 ( .A(n33110), .B(n33111), .Z(n33100) );
  ANDN U31619 ( .B(n33112), .A(n33113), .Z(n33110) );
  XOR U31620 ( .A(n33111), .B(n33114), .Z(n33112) );
  XOR U31621 ( .A(n33115), .B(n33116), .Z(n33099) );
  XOR U31622 ( .A(n33117), .B(n33118), .Z(n33116) );
  ANDN U31623 ( .B(n33119), .A(n33120), .Z(n33117) );
  XOR U31624 ( .A(n33121), .B(n33118), .Z(n33119) );
  IV U31625 ( .A(n33097), .Z(n33115) );
  XOR U31626 ( .A(n33122), .B(n33123), .Z(n33097) );
  ANDN U31627 ( .B(n33124), .A(n33125), .Z(n33122) );
  XOR U31628 ( .A(n33123), .B(n33126), .Z(n33124) );
  IV U31629 ( .A(n33105), .Z(n33109) );
  XOR U31630 ( .A(n33105), .B(n33087), .Z(n33107) );
  XOR U31631 ( .A(n33127), .B(n33128), .Z(n33087) );
  AND U31632 ( .A(n2038), .B(n33129), .Z(n33127) );
  XOR U31633 ( .A(n33130), .B(n33128), .Z(n33129) );
  NANDN U31634 ( .A(n33089), .B(n33091), .Z(n33105) );
  XOR U31635 ( .A(n33131), .B(n33132), .Z(n33091) );
  AND U31636 ( .A(n2038), .B(n33133), .Z(n33131) );
  XOR U31637 ( .A(n33132), .B(n33134), .Z(n33133) );
  XOR U31638 ( .A(n33135), .B(n33136), .Z(n2038) );
  AND U31639 ( .A(n33137), .B(n33138), .Z(n33135) );
  XNOR U31640 ( .A(n33136), .B(n33102), .Z(n33138) );
  XNOR U31641 ( .A(n33139), .B(n33140), .Z(n33102) );
  ANDN U31642 ( .B(n33141), .A(n33142), .Z(n33139) );
  XOR U31643 ( .A(n33140), .B(n33143), .Z(n33141) );
  XOR U31644 ( .A(n33136), .B(n33104), .Z(n33137) );
  XOR U31645 ( .A(n33144), .B(n33145), .Z(n33104) );
  AND U31646 ( .A(n2042), .B(n33146), .Z(n33144) );
  XOR U31647 ( .A(n33147), .B(n33145), .Z(n33146) );
  XNOR U31648 ( .A(n33148), .B(n33149), .Z(n33136) );
  NAND U31649 ( .A(n33150), .B(n33151), .Z(n33149) );
  XOR U31650 ( .A(n33152), .B(n33128), .Z(n33151) );
  XOR U31651 ( .A(n33142), .B(n33143), .Z(n33128) );
  XOR U31652 ( .A(n33153), .B(n33154), .Z(n33143) );
  ANDN U31653 ( .B(n33155), .A(n33156), .Z(n33153) );
  XOR U31654 ( .A(n33154), .B(n33157), .Z(n33155) );
  XOR U31655 ( .A(n33158), .B(n33159), .Z(n33142) );
  XOR U31656 ( .A(n33160), .B(n33161), .Z(n33159) );
  ANDN U31657 ( .B(n33162), .A(n33163), .Z(n33160) );
  XOR U31658 ( .A(n33164), .B(n33161), .Z(n33162) );
  IV U31659 ( .A(n33140), .Z(n33158) );
  XOR U31660 ( .A(n33165), .B(n33166), .Z(n33140) );
  ANDN U31661 ( .B(n33167), .A(n33168), .Z(n33165) );
  XOR U31662 ( .A(n33166), .B(n33169), .Z(n33167) );
  IV U31663 ( .A(n33148), .Z(n33152) );
  XOR U31664 ( .A(n33148), .B(n33130), .Z(n33150) );
  XOR U31665 ( .A(n33170), .B(n33171), .Z(n33130) );
  AND U31666 ( .A(n2042), .B(n33172), .Z(n33170) );
  XNOR U31667 ( .A(n33173), .B(n33171), .Z(n33172) );
  NANDN U31668 ( .A(n33132), .B(n33134), .Z(n33148) );
  XOR U31669 ( .A(n33174), .B(n33175), .Z(n33134) );
  AND U31670 ( .A(n2042), .B(n33176), .Z(n33174) );
  XOR U31671 ( .A(n33175), .B(n33177), .Z(n33176) );
  XOR U31672 ( .A(n33178), .B(n33179), .Z(n2042) );
  AND U31673 ( .A(n33180), .B(n33181), .Z(n33178) );
  XNOR U31674 ( .A(n33179), .B(n33145), .Z(n33181) );
  XNOR U31675 ( .A(n33182), .B(n33183), .Z(n33145) );
  ANDN U31676 ( .B(n33184), .A(n33185), .Z(n33182) );
  XOR U31677 ( .A(n33183), .B(n33186), .Z(n33184) );
  XOR U31678 ( .A(n33179), .B(n33147), .Z(n33180) );
  XNOR U31679 ( .A(n33187), .B(n33188), .Z(n33147) );
  ANDN U31680 ( .B(n33189), .A(n33190), .Z(n33187) );
  XOR U31681 ( .A(n33188), .B(n33191), .Z(n33189) );
  XNOR U31682 ( .A(n33192), .B(n33193), .Z(n33179) );
  NAND U31683 ( .A(n33194), .B(n33195), .Z(n33193) );
  XOR U31684 ( .A(n33196), .B(n33171), .Z(n33195) );
  XOR U31685 ( .A(n33185), .B(n33186), .Z(n33171) );
  XOR U31686 ( .A(n33197), .B(n33198), .Z(n33186) );
  ANDN U31687 ( .B(n33199), .A(n33200), .Z(n33197) );
  XOR U31688 ( .A(n33198), .B(n33201), .Z(n33199) );
  XOR U31689 ( .A(n33202), .B(n33203), .Z(n33185) );
  XOR U31690 ( .A(n33204), .B(n33205), .Z(n33203) );
  ANDN U31691 ( .B(n33206), .A(n33207), .Z(n33204) );
  XOR U31692 ( .A(n33208), .B(n33205), .Z(n33206) );
  IV U31693 ( .A(n33183), .Z(n33202) );
  XOR U31694 ( .A(n33209), .B(n33210), .Z(n33183) );
  ANDN U31695 ( .B(n33211), .A(n33212), .Z(n33209) );
  XOR U31696 ( .A(n33210), .B(n33213), .Z(n33211) );
  IV U31697 ( .A(n33192), .Z(n33196) );
  XNOR U31698 ( .A(n33192), .B(n33173), .Z(n33194) );
  XOR U31699 ( .A(n33214), .B(n33191), .Z(n33173) );
  XOR U31700 ( .A(n33215), .B(n33216), .Z(n33191) );
  ANDN U31701 ( .B(n33217), .A(n33218), .Z(n33215) );
  XOR U31702 ( .A(n33216), .B(n33219), .Z(n33217) );
  IV U31703 ( .A(n33190), .Z(n33214) );
  XOR U31704 ( .A(n33220), .B(n33221), .Z(n33190) );
  XOR U31705 ( .A(n33222), .B(n33223), .Z(n33221) );
  ANDN U31706 ( .B(n33224), .A(n33225), .Z(n33222) );
  XOR U31707 ( .A(n33226), .B(n33223), .Z(n33224) );
  IV U31708 ( .A(n33188), .Z(n33220) );
  XNOR U31709 ( .A(n33227), .B(n33228), .Z(n33188) );
  ANDN U31710 ( .B(n33229), .A(n33230), .Z(n33227) );
  XNOR U31711 ( .A(n33228), .B(n33231), .Z(n33229) );
  NANDN U31712 ( .A(n33175), .B(n33177), .Z(n33192) );
  XOR U31713 ( .A(n33232), .B(n33231), .Z(n33177) );
  XOR U31714 ( .A(n33233), .B(n33219), .Z(n33231) );
  XNOR U31715 ( .A(q[6]), .B(DB[6]), .Z(n33219) );
  IV U31716 ( .A(n33218), .Z(n33233) );
  XNOR U31717 ( .A(n33216), .B(n33234), .Z(n33218) );
  XNOR U31718 ( .A(q[5]), .B(DB[5]), .Z(n33234) );
  XNOR U31719 ( .A(q[4]), .B(DB[4]), .Z(n33216) );
  IV U31720 ( .A(n33230), .Z(n33232) );
  XOR U31721 ( .A(n33235), .B(n33236), .Z(n33230) );
  XOR U31722 ( .A(n33228), .B(n33226), .Z(n33236) );
  XNOR U31723 ( .A(q[3]), .B(DB[3]), .Z(n33226) );
  XOR U31724 ( .A(q[0]), .B(DB[0]), .Z(n33228) );
  IV U31725 ( .A(n33225), .Z(n33235) );
  XNOR U31726 ( .A(n33223), .B(n33237), .Z(n33225) );
  XNOR U31727 ( .A(q[2]), .B(DB[2]), .Z(n33237) );
  XNOR U31728 ( .A(q[1]), .B(DB[1]), .Z(n33223) );
  XOR U31729 ( .A(n33238), .B(n33213), .Z(n33175) );
  XOR U31730 ( .A(n33239), .B(n33201), .Z(n33213) );
  XNOR U31731 ( .A(q[6]), .B(DB[13]), .Z(n33201) );
  IV U31732 ( .A(n33200), .Z(n33239) );
  XNOR U31733 ( .A(n33198), .B(n33240), .Z(n33200) );
  XNOR U31734 ( .A(q[5]), .B(DB[12]), .Z(n33240) );
  XNOR U31735 ( .A(q[4]), .B(DB[11]), .Z(n33198) );
  IV U31736 ( .A(n33212), .Z(n33238) );
  XOR U31737 ( .A(n33241), .B(n33242), .Z(n33212) );
  XNOR U31738 ( .A(n33208), .B(n33210), .Z(n33242) );
  XNOR U31739 ( .A(q[0]), .B(DB[7]), .Z(n33210) );
  XNOR U31740 ( .A(q[3]), .B(DB[10]), .Z(n33208) );
  IV U31741 ( .A(n33207), .Z(n33241) );
  XNOR U31742 ( .A(n33205), .B(n33243), .Z(n33207) );
  XNOR U31743 ( .A(q[2]), .B(DB[9]), .Z(n33243) );
  XNOR U31744 ( .A(q[1]), .B(DB[8]), .Z(n33205) );
  XOR U31745 ( .A(n33244), .B(n33169), .Z(n33132) );
  XOR U31746 ( .A(n33245), .B(n33157), .Z(n33169) );
  XNOR U31747 ( .A(q[6]), .B(DB[20]), .Z(n33157) );
  IV U31748 ( .A(n33156), .Z(n33245) );
  XNOR U31749 ( .A(n33154), .B(n33246), .Z(n33156) );
  XNOR U31750 ( .A(q[5]), .B(DB[19]), .Z(n33246) );
  XNOR U31751 ( .A(q[4]), .B(DB[18]), .Z(n33154) );
  IV U31752 ( .A(n33168), .Z(n33244) );
  XOR U31753 ( .A(n33247), .B(n33248), .Z(n33168) );
  XNOR U31754 ( .A(n33164), .B(n33166), .Z(n33248) );
  XNOR U31755 ( .A(q[0]), .B(DB[14]), .Z(n33166) );
  XNOR U31756 ( .A(q[3]), .B(DB[17]), .Z(n33164) );
  IV U31757 ( .A(n33163), .Z(n33247) );
  XNOR U31758 ( .A(n33161), .B(n33249), .Z(n33163) );
  XNOR U31759 ( .A(q[2]), .B(DB[16]), .Z(n33249) );
  XNOR U31760 ( .A(q[1]), .B(DB[15]), .Z(n33161) );
  XOR U31761 ( .A(n33250), .B(n33126), .Z(n33089) );
  XOR U31762 ( .A(n33251), .B(n33114), .Z(n33126) );
  XNOR U31763 ( .A(q[6]), .B(DB[27]), .Z(n33114) );
  IV U31764 ( .A(n33113), .Z(n33251) );
  XNOR U31765 ( .A(n33111), .B(n33252), .Z(n33113) );
  XNOR U31766 ( .A(q[5]), .B(DB[26]), .Z(n33252) );
  XNOR U31767 ( .A(q[4]), .B(DB[25]), .Z(n33111) );
  IV U31768 ( .A(n33125), .Z(n33250) );
  XOR U31769 ( .A(n33253), .B(n33254), .Z(n33125) );
  XNOR U31770 ( .A(n33121), .B(n33123), .Z(n33254) );
  XNOR U31771 ( .A(q[0]), .B(DB[21]), .Z(n33123) );
  XNOR U31772 ( .A(q[3]), .B(DB[24]), .Z(n33121) );
  IV U31773 ( .A(n33120), .Z(n33253) );
  XNOR U31774 ( .A(n33118), .B(n33255), .Z(n33120) );
  XNOR U31775 ( .A(q[2]), .B(DB[23]), .Z(n33255) );
  XNOR U31776 ( .A(q[1]), .B(DB[22]), .Z(n33118) );
  XOR U31777 ( .A(n33256), .B(n33083), .Z(n33046) );
  XOR U31778 ( .A(n33257), .B(n33071), .Z(n33083) );
  XNOR U31779 ( .A(q[6]), .B(DB[34]), .Z(n33071) );
  IV U31780 ( .A(n33070), .Z(n33257) );
  XNOR U31781 ( .A(n33068), .B(n33258), .Z(n33070) );
  XNOR U31782 ( .A(q[5]), .B(DB[33]), .Z(n33258) );
  XNOR U31783 ( .A(q[4]), .B(DB[32]), .Z(n33068) );
  IV U31784 ( .A(n33082), .Z(n33256) );
  XOR U31785 ( .A(n33259), .B(n33260), .Z(n33082) );
  XNOR U31786 ( .A(n33078), .B(n33080), .Z(n33260) );
  XNOR U31787 ( .A(q[0]), .B(DB[28]), .Z(n33080) );
  XNOR U31788 ( .A(q[3]), .B(DB[31]), .Z(n33078) );
  IV U31789 ( .A(n33077), .Z(n33259) );
  XNOR U31790 ( .A(n33075), .B(n33261), .Z(n33077) );
  XNOR U31791 ( .A(q[2]), .B(DB[30]), .Z(n33261) );
  XNOR U31792 ( .A(q[1]), .B(DB[29]), .Z(n33075) );
  XOR U31793 ( .A(n33262), .B(n33040), .Z(n33003) );
  XOR U31794 ( .A(n33263), .B(n33028), .Z(n33040) );
  XNOR U31795 ( .A(q[6]), .B(DB[41]), .Z(n33028) );
  IV U31796 ( .A(n33027), .Z(n33263) );
  XNOR U31797 ( .A(n33025), .B(n33264), .Z(n33027) );
  XNOR U31798 ( .A(q[5]), .B(DB[40]), .Z(n33264) );
  XNOR U31799 ( .A(q[4]), .B(DB[39]), .Z(n33025) );
  IV U31800 ( .A(n33039), .Z(n33262) );
  XOR U31801 ( .A(n33265), .B(n33266), .Z(n33039) );
  XNOR U31802 ( .A(n33035), .B(n33037), .Z(n33266) );
  XNOR U31803 ( .A(q[0]), .B(DB[35]), .Z(n33037) );
  XNOR U31804 ( .A(q[3]), .B(DB[38]), .Z(n33035) );
  IV U31805 ( .A(n33034), .Z(n33265) );
  XNOR U31806 ( .A(n33032), .B(n33267), .Z(n33034) );
  XNOR U31807 ( .A(q[2]), .B(DB[37]), .Z(n33267) );
  XNOR U31808 ( .A(q[1]), .B(DB[36]), .Z(n33032) );
  XOR U31809 ( .A(n33268), .B(n32997), .Z(n32960) );
  XOR U31810 ( .A(n33269), .B(n32985), .Z(n32997) );
  XNOR U31811 ( .A(q[6]), .B(DB[48]), .Z(n32985) );
  IV U31812 ( .A(n32984), .Z(n33269) );
  XNOR U31813 ( .A(n32982), .B(n33270), .Z(n32984) );
  XNOR U31814 ( .A(q[5]), .B(DB[47]), .Z(n33270) );
  XNOR U31815 ( .A(q[4]), .B(DB[46]), .Z(n32982) );
  IV U31816 ( .A(n32996), .Z(n33268) );
  XOR U31817 ( .A(n33271), .B(n33272), .Z(n32996) );
  XNOR U31818 ( .A(n32992), .B(n32994), .Z(n33272) );
  XNOR U31819 ( .A(q[0]), .B(DB[42]), .Z(n32994) );
  XNOR U31820 ( .A(q[3]), .B(DB[45]), .Z(n32992) );
  IV U31821 ( .A(n32991), .Z(n33271) );
  XNOR U31822 ( .A(n32989), .B(n33273), .Z(n32991) );
  XNOR U31823 ( .A(q[2]), .B(DB[44]), .Z(n33273) );
  XNOR U31824 ( .A(q[1]), .B(DB[43]), .Z(n32989) );
  XOR U31825 ( .A(n33274), .B(n32954), .Z(n32917) );
  XOR U31826 ( .A(n33275), .B(n32942), .Z(n32954) );
  XNOR U31827 ( .A(q[6]), .B(DB[55]), .Z(n32942) );
  IV U31828 ( .A(n32941), .Z(n33275) );
  XNOR U31829 ( .A(n32939), .B(n33276), .Z(n32941) );
  XNOR U31830 ( .A(q[5]), .B(DB[54]), .Z(n33276) );
  XNOR U31831 ( .A(q[4]), .B(DB[53]), .Z(n32939) );
  IV U31832 ( .A(n32953), .Z(n33274) );
  XOR U31833 ( .A(n33277), .B(n33278), .Z(n32953) );
  XNOR U31834 ( .A(n32949), .B(n32951), .Z(n33278) );
  XNOR U31835 ( .A(q[0]), .B(DB[49]), .Z(n32951) );
  XNOR U31836 ( .A(q[3]), .B(DB[52]), .Z(n32949) );
  IV U31837 ( .A(n32948), .Z(n33277) );
  XNOR U31838 ( .A(n32946), .B(n33279), .Z(n32948) );
  XNOR U31839 ( .A(q[2]), .B(DB[51]), .Z(n33279) );
  XNOR U31840 ( .A(q[1]), .B(DB[50]), .Z(n32946) );
  XOR U31841 ( .A(n33280), .B(n32911), .Z(n32874) );
  XOR U31842 ( .A(n33281), .B(n32899), .Z(n32911) );
  XNOR U31843 ( .A(q[6]), .B(DB[62]), .Z(n32899) );
  IV U31844 ( .A(n32898), .Z(n33281) );
  XNOR U31845 ( .A(n32896), .B(n33282), .Z(n32898) );
  XNOR U31846 ( .A(q[5]), .B(DB[61]), .Z(n33282) );
  XNOR U31847 ( .A(q[4]), .B(DB[60]), .Z(n32896) );
  IV U31848 ( .A(n32910), .Z(n33280) );
  XOR U31849 ( .A(n33283), .B(n33284), .Z(n32910) );
  XNOR U31850 ( .A(n32906), .B(n32908), .Z(n33284) );
  XNOR U31851 ( .A(q[0]), .B(DB[56]), .Z(n32908) );
  XNOR U31852 ( .A(q[3]), .B(DB[59]), .Z(n32906) );
  IV U31853 ( .A(n32905), .Z(n33283) );
  XNOR U31854 ( .A(n32903), .B(n33285), .Z(n32905) );
  XNOR U31855 ( .A(q[2]), .B(DB[58]), .Z(n33285) );
  XNOR U31856 ( .A(q[1]), .B(DB[57]), .Z(n32903) );
  XOR U31857 ( .A(n33286), .B(n32868), .Z(n32831) );
  XOR U31858 ( .A(n33287), .B(n32856), .Z(n32868) );
  XNOR U31859 ( .A(q[6]), .B(DB[69]), .Z(n32856) );
  IV U31860 ( .A(n32855), .Z(n33287) );
  XNOR U31861 ( .A(n32853), .B(n33288), .Z(n32855) );
  XNOR U31862 ( .A(q[5]), .B(DB[68]), .Z(n33288) );
  XNOR U31863 ( .A(q[4]), .B(DB[67]), .Z(n32853) );
  IV U31864 ( .A(n32867), .Z(n33286) );
  XOR U31865 ( .A(n33289), .B(n33290), .Z(n32867) );
  XNOR U31866 ( .A(n32863), .B(n32865), .Z(n33290) );
  XNOR U31867 ( .A(q[0]), .B(DB[63]), .Z(n32865) );
  XNOR U31868 ( .A(q[3]), .B(DB[66]), .Z(n32863) );
  IV U31869 ( .A(n32862), .Z(n33289) );
  XNOR U31870 ( .A(n32860), .B(n33291), .Z(n32862) );
  XNOR U31871 ( .A(q[2]), .B(DB[65]), .Z(n33291) );
  XNOR U31872 ( .A(q[1]), .B(DB[64]), .Z(n32860) );
  XOR U31873 ( .A(n33292), .B(n32825), .Z(n32788) );
  XOR U31874 ( .A(n33293), .B(n32813), .Z(n32825) );
  XNOR U31875 ( .A(q[6]), .B(DB[76]), .Z(n32813) );
  IV U31876 ( .A(n32812), .Z(n33293) );
  XNOR U31877 ( .A(n32810), .B(n33294), .Z(n32812) );
  XNOR U31878 ( .A(q[5]), .B(DB[75]), .Z(n33294) );
  XNOR U31879 ( .A(q[4]), .B(DB[74]), .Z(n32810) );
  IV U31880 ( .A(n32824), .Z(n33292) );
  XOR U31881 ( .A(n33295), .B(n33296), .Z(n32824) );
  XNOR U31882 ( .A(n32820), .B(n32822), .Z(n33296) );
  XNOR U31883 ( .A(q[0]), .B(DB[70]), .Z(n32822) );
  XNOR U31884 ( .A(q[3]), .B(DB[73]), .Z(n32820) );
  IV U31885 ( .A(n32819), .Z(n33295) );
  XNOR U31886 ( .A(n32817), .B(n33297), .Z(n32819) );
  XNOR U31887 ( .A(q[2]), .B(DB[72]), .Z(n33297) );
  XNOR U31888 ( .A(q[1]), .B(DB[71]), .Z(n32817) );
  XOR U31889 ( .A(n33298), .B(n32782), .Z(n32745) );
  XOR U31890 ( .A(n33299), .B(n32770), .Z(n32782) );
  XNOR U31891 ( .A(q[6]), .B(DB[83]), .Z(n32770) );
  IV U31892 ( .A(n32769), .Z(n33299) );
  XNOR U31893 ( .A(n32767), .B(n33300), .Z(n32769) );
  XNOR U31894 ( .A(q[5]), .B(DB[82]), .Z(n33300) );
  XNOR U31895 ( .A(q[4]), .B(DB[81]), .Z(n32767) );
  IV U31896 ( .A(n32781), .Z(n33298) );
  XOR U31897 ( .A(n33301), .B(n33302), .Z(n32781) );
  XNOR U31898 ( .A(n32777), .B(n32779), .Z(n33302) );
  XNOR U31899 ( .A(q[0]), .B(DB[77]), .Z(n32779) );
  XNOR U31900 ( .A(q[3]), .B(DB[80]), .Z(n32777) );
  IV U31901 ( .A(n32776), .Z(n33301) );
  XNOR U31902 ( .A(n32774), .B(n33303), .Z(n32776) );
  XNOR U31903 ( .A(q[2]), .B(DB[79]), .Z(n33303) );
  XNOR U31904 ( .A(q[1]), .B(DB[78]), .Z(n32774) );
  XOR U31905 ( .A(n33304), .B(n32739), .Z(n32702) );
  XOR U31906 ( .A(n33305), .B(n32727), .Z(n32739) );
  XNOR U31907 ( .A(q[6]), .B(DB[90]), .Z(n32727) );
  IV U31908 ( .A(n32726), .Z(n33305) );
  XNOR U31909 ( .A(n32724), .B(n33306), .Z(n32726) );
  XNOR U31910 ( .A(q[5]), .B(DB[89]), .Z(n33306) );
  XNOR U31911 ( .A(q[4]), .B(DB[88]), .Z(n32724) );
  IV U31912 ( .A(n32738), .Z(n33304) );
  XOR U31913 ( .A(n33307), .B(n33308), .Z(n32738) );
  XNOR U31914 ( .A(n32734), .B(n32736), .Z(n33308) );
  XNOR U31915 ( .A(q[0]), .B(DB[84]), .Z(n32736) );
  XNOR U31916 ( .A(q[3]), .B(DB[87]), .Z(n32734) );
  IV U31917 ( .A(n32733), .Z(n33307) );
  XNOR U31918 ( .A(n32731), .B(n33309), .Z(n32733) );
  XNOR U31919 ( .A(q[2]), .B(DB[86]), .Z(n33309) );
  XNOR U31920 ( .A(q[1]), .B(DB[85]), .Z(n32731) );
  XOR U31921 ( .A(n33310), .B(n32696), .Z(n32659) );
  XOR U31922 ( .A(n33311), .B(n32684), .Z(n32696) );
  XNOR U31923 ( .A(q[6]), .B(DB[97]), .Z(n32684) );
  IV U31924 ( .A(n32683), .Z(n33311) );
  XNOR U31925 ( .A(n32681), .B(n33312), .Z(n32683) );
  XNOR U31926 ( .A(q[5]), .B(DB[96]), .Z(n33312) );
  XNOR U31927 ( .A(q[4]), .B(DB[95]), .Z(n32681) );
  IV U31928 ( .A(n32695), .Z(n33310) );
  XOR U31929 ( .A(n33313), .B(n33314), .Z(n32695) );
  XNOR U31930 ( .A(n32691), .B(n32693), .Z(n33314) );
  XNOR U31931 ( .A(q[0]), .B(DB[91]), .Z(n32693) );
  XNOR U31932 ( .A(q[3]), .B(DB[94]), .Z(n32691) );
  IV U31933 ( .A(n32690), .Z(n33313) );
  XNOR U31934 ( .A(n32688), .B(n33315), .Z(n32690) );
  XNOR U31935 ( .A(q[2]), .B(DB[93]), .Z(n33315) );
  XNOR U31936 ( .A(q[1]), .B(DB[92]), .Z(n32688) );
  XOR U31937 ( .A(n33316), .B(n32653), .Z(n32616) );
  XOR U31938 ( .A(n33317), .B(n32641), .Z(n32653) );
  XNOR U31939 ( .A(q[6]), .B(DB[104]), .Z(n32641) );
  IV U31940 ( .A(n32640), .Z(n33317) );
  XNOR U31941 ( .A(n32638), .B(n33318), .Z(n32640) );
  XNOR U31942 ( .A(q[5]), .B(DB[103]), .Z(n33318) );
  XNOR U31943 ( .A(q[4]), .B(DB[102]), .Z(n32638) );
  IV U31944 ( .A(n32652), .Z(n33316) );
  XOR U31945 ( .A(n33319), .B(n33320), .Z(n32652) );
  XNOR U31946 ( .A(n32648), .B(n32650), .Z(n33320) );
  XNOR U31947 ( .A(q[0]), .B(DB[98]), .Z(n32650) );
  XNOR U31948 ( .A(q[3]), .B(DB[101]), .Z(n32648) );
  IV U31949 ( .A(n32647), .Z(n33319) );
  XNOR U31950 ( .A(n32645), .B(n33321), .Z(n32647) );
  XNOR U31951 ( .A(q[2]), .B(DB[100]), .Z(n33321) );
  XNOR U31952 ( .A(q[1]), .B(DB[99]), .Z(n32645) );
  XOR U31953 ( .A(n33322), .B(n32610), .Z(n32573) );
  XOR U31954 ( .A(n33323), .B(n32598), .Z(n32610) );
  XNOR U31955 ( .A(q[6]), .B(DB[111]), .Z(n32598) );
  IV U31956 ( .A(n32597), .Z(n33323) );
  XNOR U31957 ( .A(n32595), .B(n33324), .Z(n32597) );
  XNOR U31958 ( .A(q[5]), .B(DB[110]), .Z(n33324) );
  XNOR U31959 ( .A(q[4]), .B(DB[109]), .Z(n32595) );
  IV U31960 ( .A(n32609), .Z(n33322) );
  XOR U31961 ( .A(n33325), .B(n33326), .Z(n32609) );
  XNOR U31962 ( .A(n32605), .B(n32607), .Z(n33326) );
  XNOR U31963 ( .A(q[0]), .B(DB[105]), .Z(n32607) );
  XNOR U31964 ( .A(q[3]), .B(DB[108]), .Z(n32605) );
  IV U31965 ( .A(n32604), .Z(n33325) );
  XNOR U31966 ( .A(n32602), .B(n33327), .Z(n32604) );
  XNOR U31967 ( .A(q[2]), .B(DB[107]), .Z(n33327) );
  XNOR U31968 ( .A(q[1]), .B(DB[106]), .Z(n32602) );
  XOR U31969 ( .A(n33328), .B(n32567), .Z(n32530) );
  XOR U31970 ( .A(n33329), .B(n32555), .Z(n32567) );
  XNOR U31971 ( .A(q[6]), .B(DB[118]), .Z(n32555) );
  IV U31972 ( .A(n32554), .Z(n33329) );
  XNOR U31973 ( .A(n32552), .B(n33330), .Z(n32554) );
  XNOR U31974 ( .A(q[5]), .B(DB[117]), .Z(n33330) );
  XNOR U31975 ( .A(q[4]), .B(DB[116]), .Z(n32552) );
  IV U31976 ( .A(n32566), .Z(n33328) );
  XOR U31977 ( .A(n33331), .B(n33332), .Z(n32566) );
  XNOR U31978 ( .A(n32562), .B(n32564), .Z(n33332) );
  XNOR U31979 ( .A(q[0]), .B(DB[112]), .Z(n32564) );
  XNOR U31980 ( .A(q[3]), .B(DB[115]), .Z(n32562) );
  IV U31981 ( .A(n32561), .Z(n33331) );
  XNOR U31982 ( .A(n32559), .B(n33333), .Z(n32561) );
  XNOR U31983 ( .A(q[2]), .B(DB[114]), .Z(n33333) );
  XNOR U31984 ( .A(q[1]), .B(DB[113]), .Z(n32559) );
  XOR U31985 ( .A(n33334), .B(n32524), .Z(n32487) );
  XOR U31986 ( .A(n33335), .B(n32512), .Z(n32524) );
  XNOR U31987 ( .A(q[6]), .B(DB[125]), .Z(n32512) );
  IV U31988 ( .A(n32511), .Z(n33335) );
  XNOR U31989 ( .A(n32509), .B(n33336), .Z(n32511) );
  XNOR U31990 ( .A(q[5]), .B(DB[124]), .Z(n33336) );
  XNOR U31991 ( .A(q[4]), .B(DB[123]), .Z(n32509) );
  IV U31992 ( .A(n32523), .Z(n33334) );
  XOR U31993 ( .A(n33337), .B(n33338), .Z(n32523) );
  XNOR U31994 ( .A(n32519), .B(n32521), .Z(n33338) );
  XNOR U31995 ( .A(q[0]), .B(DB[119]), .Z(n32521) );
  XNOR U31996 ( .A(q[3]), .B(DB[122]), .Z(n32519) );
  IV U31997 ( .A(n32518), .Z(n33337) );
  XNOR U31998 ( .A(n32516), .B(n33339), .Z(n32518) );
  XNOR U31999 ( .A(q[2]), .B(DB[121]), .Z(n33339) );
  XNOR U32000 ( .A(q[1]), .B(DB[120]), .Z(n32516) );
  XOR U32001 ( .A(n33340), .B(n32481), .Z(n32444) );
  XOR U32002 ( .A(n33341), .B(n32469), .Z(n32481) );
  XNOR U32003 ( .A(q[6]), .B(DB[132]), .Z(n32469) );
  IV U32004 ( .A(n32468), .Z(n33341) );
  XNOR U32005 ( .A(n32466), .B(n33342), .Z(n32468) );
  XNOR U32006 ( .A(q[5]), .B(DB[131]), .Z(n33342) );
  XNOR U32007 ( .A(q[4]), .B(DB[130]), .Z(n32466) );
  IV U32008 ( .A(n32480), .Z(n33340) );
  XOR U32009 ( .A(n33343), .B(n33344), .Z(n32480) );
  XNOR U32010 ( .A(n32476), .B(n32478), .Z(n33344) );
  XNOR U32011 ( .A(q[0]), .B(DB[126]), .Z(n32478) );
  XNOR U32012 ( .A(q[3]), .B(DB[129]), .Z(n32476) );
  IV U32013 ( .A(n32475), .Z(n33343) );
  XNOR U32014 ( .A(n32473), .B(n33345), .Z(n32475) );
  XNOR U32015 ( .A(q[2]), .B(DB[128]), .Z(n33345) );
  XNOR U32016 ( .A(q[1]), .B(DB[127]), .Z(n32473) );
  XOR U32017 ( .A(n33346), .B(n32438), .Z(n32401) );
  XOR U32018 ( .A(n33347), .B(n32426), .Z(n32438) );
  XNOR U32019 ( .A(q[6]), .B(DB[139]), .Z(n32426) );
  IV U32020 ( .A(n32425), .Z(n33347) );
  XNOR U32021 ( .A(n32423), .B(n33348), .Z(n32425) );
  XNOR U32022 ( .A(q[5]), .B(DB[138]), .Z(n33348) );
  XNOR U32023 ( .A(q[4]), .B(DB[137]), .Z(n32423) );
  IV U32024 ( .A(n32437), .Z(n33346) );
  XOR U32025 ( .A(n33349), .B(n33350), .Z(n32437) );
  XNOR U32026 ( .A(n32433), .B(n32435), .Z(n33350) );
  XNOR U32027 ( .A(q[0]), .B(DB[133]), .Z(n32435) );
  XNOR U32028 ( .A(q[3]), .B(DB[136]), .Z(n32433) );
  IV U32029 ( .A(n32432), .Z(n33349) );
  XNOR U32030 ( .A(n32430), .B(n33351), .Z(n32432) );
  XNOR U32031 ( .A(q[2]), .B(DB[135]), .Z(n33351) );
  XNOR U32032 ( .A(q[1]), .B(DB[134]), .Z(n32430) );
  XOR U32033 ( .A(n33352), .B(n32395), .Z(n32358) );
  XOR U32034 ( .A(n33353), .B(n32383), .Z(n32395) );
  XNOR U32035 ( .A(q[6]), .B(DB[146]), .Z(n32383) );
  IV U32036 ( .A(n32382), .Z(n33353) );
  XNOR U32037 ( .A(n32380), .B(n33354), .Z(n32382) );
  XNOR U32038 ( .A(q[5]), .B(DB[145]), .Z(n33354) );
  XNOR U32039 ( .A(q[4]), .B(DB[144]), .Z(n32380) );
  IV U32040 ( .A(n32394), .Z(n33352) );
  XOR U32041 ( .A(n33355), .B(n33356), .Z(n32394) );
  XNOR U32042 ( .A(n32390), .B(n32392), .Z(n33356) );
  XNOR U32043 ( .A(q[0]), .B(DB[140]), .Z(n32392) );
  XNOR U32044 ( .A(q[3]), .B(DB[143]), .Z(n32390) );
  IV U32045 ( .A(n32389), .Z(n33355) );
  XNOR U32046 ( .A(n32387), .B(n33357), .Z(n32389) );
  XNOR U32047 ( .A(q[2]), .B(DB[142]), .Z(n33357) );
  XNOR U32048 ( .A(q[1]), .B(DB[141]), .Z(n32387) );
  XOR U32049 ( .A(n33358), .B(n32352), .Z(n32315) );
  XOR U32050 ( .A(n33359), .B(n32340), .Z(n32352) );
  XNOR U32051 ( .A(q[6]), .B(DB[153]), .Z(n32340) );
  IV U32052 ( .A(n32339), .Z(n33359) );
  XNOR U32053 ( .A(n32337), .B(n33360), .Z(n32339) );
  XNOR U32054 ( .A(q[5]), .B(DB[152]), .Z(n33360) );
  XNOR U32055 ( .A(q[4]), .B(DB[151]), .Z(n32337) );
  IV U32056 ( .A(n32351), .Z(n33358) );
  XOR U32057 ( .A(n33361), .B(n33362), .Z(n32351) );
  XNOR U32058 ( .A(n32347), .B(n32349), .Z(n33362) );
  XNOR U32059 ( .A(q[0]), .B(DB[147]), .Z(n32349) );
  XNOR U32060 ( .A(q[3]), .B(DB[150]), .Z(n32347) );
  IV U32061 ( .A(n32346), .Z(n33361) );
  XNOR U32062 ( .A(n32344), .B(n33363), .Z(n32346) );
  XNOR U32063 ( .A(q[2]), .B(DB[149]), .Z(n33363) );
  XNOR U32064 ( .A(q[1]), .B(DB[148]), .Z(n32344) );
  XOR U32065 ( .A(n33364), .B(n32309), .Z(n32272) );
  XOR U32066 ( .A(n33365), .B(n32297), .Z(n32309) );
  XNOR U32067 ( .A(q[6]), .B(DB[160]), .Z(n32297) );
  IV U32068 ( .A(n32296), .Z(n33365) );
  XNOR U32069 ( .A(n32294), .B(n33366), .Z(n32296) );
  XNOR U32070 ( .A(q[5]), .B(DB[159]), .Z(n33366) );
  XNOR U32071 ( .A(q[4]), .B(DB[158]), .Z(n32294) );
  IV U32072 ( .A(n32308), .Z(n33364) );
  XOR U32073 ( .A(n33367), .B(n33368), .Z(n32308) );
  XNOR U32074 ( .A(n32304), .B(n32306), .Z(n33368) );
  XNOR U32075 ( .A(q[0]), .B(DB[154]), .Z(n32306) );
  XNOR U32076 ( .A(q[3]), .B(DB[157]), .Z(n32304) );
  IV U32077 ( .A(n32303), .Z(n33367) );
  XNOR U32078 ( .A(n32301), .B(n33369), .Z(n32303) );
  XNOR U32079 ( .A(q[2]), .B(DB[156]), .Z(n33369) );
  XNOR U32080 ( .A(q[1]), .B(DB[155]), .Z(n32301) );
  XOR U32081 ( .A(n33370), .B(n32266), .Z(n32229) );
  XOR U32082 ( .A(n33371), .B(n32254), .Z(n32266) );
  XNOR U32083 ( .A(q[6]), .B(DB[167]), .Z(n32254) );
  IV U32084 ( .A(n32253), .Z(n33371) );
  XNOR U32085 ( .A(n32251), .B(n33372), .Z(n32253) );
  XNOR U32086 ( .A(q[5]), .B(DB[166]), .Z(n33372) );
  XNOR U32087 ( .A(q[4]), .B(DB[165]), .Z(n32251) );
  IV U32088 ( .A(n32265), .Z(n33370) );
  XOR U32089 ( .A(n33373), .B(n33374), .Z(n32265) );
  XNOR U32090 ( .A(n32261), .B(n32263), .Z(n33374) );
  XNOR U32091 ( .A(q[0]), .B(DB[161]), .Z(n32263) );
  XNOR U32092 ( .A(q[3]), .B(DB[164]), .Z(n32261) );
  IV U32093 ( .A(n32260), .Z(n33373) );
  XNOR U32094 ( .A(n32258), .B(n33375), .Z(n32260) );
  XNOR U32095 ( .A(q[2]), .B(DB[163]), .Z(n33375) );
  XNOR U32096 ( .A(q[1]), .B(DB[162]), .Z(n32258) );
  XOR U32097 ( .A(n33376), .B(n32223), .Z(n32186) );
  XOR U32098 ( .A(n33377), .B(n32211), .Z(n32223) );
  XNOR U32099 ( .A(q[6]), .B(DB[174]), .Z(n32211) );
  IV U32100 ( .A(n32210), .Z(n33377) );
  XNOR U32101 ( .A(n32208), .B(n33378), .Z(n32210) );
  XNOR U32102 ( .A(q[5]), .B(DB[173]), .Z(n33378) );
  XNOR U32103 ( .A(q[4]), .B(DB[172]), .Z(n32208) );
  IV U32104 ( .A(n32222), .Z(n33376) );
  XOR U32105 ( .A(n33379), .B(n33380), .Z(n32222) );
  XNOR U32106 ( .A(n32218), .B(n32220), .Z(n33380) );
  XNOR U32107 ( .A(q[0]), .B(DB[168]), .Z(n32220) );
  XNOR U32108 ( .A(q[3]), .B(DB[171]), .Z(n32218) );
  IV U32109 ( .A(n32217), .Z(n33379) );
  XNOR U32110 ( .A(n32215), .B(n33381), .Z(n32217) );
  XNOR U32111 ( .A(q[2]), .B(DB[170]), .Z(n33381) );
  XNOR U32112 ( .A(q[1]), .B(DB[169]), .Z(n32215) );
  XOR U32113 ( .A(n33382), .B(n32180), .Z(n32143) );
  XOR U32114 ( .A(n33383), .B(n32168), .Z(n32180) );
  XNOR U32115 ( .A(q[6]), .B(DB[181]), .Z(n32168) );
  IV U32116 ( .A(n32167), .Z(n33383) );
  XNOR U32117 ( .A(n32165), .B(n33384), .Z(n32167) );
  XNOR U32118 ( .A(q[5]), .B(DB[180]), .Z(n33384) );
  XNOR U32119 ( .A(q[4]), .B(DB[179]), .Z(n32165) );
  IV U32120 ( .A(n32179), .Z(n33382) );
  XOR U32121 ( .A(n33385), .B(n33386), .Z(n32179) );
  XNOR U32122 ( .A(n32175), .B(n32177), .Z(n33386) );
  XNOR U32123 ( .A(q[0]), .B(DB[175]), .Z(n32177) );
  XNOR U32124 ( .A(q[3]), .B(DB[178]), .Z(n32175) );
  IV U32125 ( .A(n32174), .Z(n33385) );
  XNOR U32126 ( .A(n32172), .B(n33387), .Z(n32174) );
  XNOR U32127 ( .A(q[2]), .B(DB[177]), .Z(n33387) );
  XNOR U32128 ( .A(q[1]), .B(DB[176]), .Z(n32172) );
  XOR U32129 ( .A(n33388), .B(n32137), .Z(n32100) );
  XOR U32130 ( .A(n33389), .B(n32125), .Z(n32137) );
  XNOR U32131 ( .A(q[6]), .B(DB[188]), .Z(n32125) );
  IV U32132 ( .A(n32124), .Z(n33389) );
  XNOR U32133 ( .A(n32122), .B(n33390), .Z(n32124) );
  XNOR U32134 ( .A(q[5]), .B(DB[187]), .Z(n33390) );
  XNOR U32135 ( .A(q[4]), .B(DB[186]), .Z(n32122) );
  IV U32136 ( .A(n32136), .Z(n33388) );
  XOR U32137 ( .A(n33391), .B(n33392), .Z(n32136) );
  XNOR U32138 ( .A(n32132), .B(n32134), .Z(n33392) );
  XNOR U32139 ( .A(q[0]), .B(DB[182]), .Z(n32134) );
  XNOR U32140 ( .A(q[3]), .B(DB[185]), .Z(n32132) );
  IV U32141 ( .A(n32131), .Z(n33391) );
  XNOR U32142 ( .A(n32129), .B(n33393), .Z(n32131) );
  XNOR U32143 ( .A(q[2]), .B(DB[184]), .Z(n33393) );
  XNOR U32144 ( .A(q[1]), .B(DB[183]), .Z(n32129) );
  XOR U32145 ( .A(n33394), .B(n32094), .Z(n32057) );
  XOR U32146 ( .A(n33395), .B(n32082), .Z(n32094) );
  XNOR U32147 ( .A(q[6]), .B(DB[195]), .Z(n32082) );
  IV U32148 ( .A(n32081), .Z(n33395) );
  XNOR U32149 ( .A(n32079), .B(n33396), .Z(n32081) );
  XNOR U32150 ( .A(q[5]), .B(DB[194]), .Z(n33396) );
  XNOR U32151 ( .A(q[4]), .B(DB[193]), .Z(n32079) );
  IV U32152 ( .A(n32093), .Z(n33394) );
  XOR U32153 ( .A(n33397), .B(n33398), .Z(n32093) );
  XNOR U32154 ( .A(n32089), .B(n32091), .Z(n33398) );
  XNOR U32155 ( .A(q[0]), .B(DB[189]), .Z(n32091) );
  XNOR U32156 ( .A(q[3]), .B(DB[192]), .Z(n32089) );
  IV U32157 ( .A(n32088), .Z(n33397) );
  XNOR U32158 ( .A(n32086), .B(n33399), .Z(n32088) );
  XNOR U32159 ( .A(q[2]), .B(DB[191]), .Z(n33399) );
  XNOR U32160 ( .A(q[1]), .B(DB[190]), .Z(n32086) );
  XOR U32161 ( .A(n33400), .B(n32051), .Z(n32014) );
  XOR U32162 ( .A(n33401), .B(n32039), .Z(n32051) );
  XNOR U32163 ( .A(q[6]), .B(DB[202]), .Z(n32039) );
  IV U32164 ( .A(n32038), .Z(n33401) );
  XNOR U32165 ( .A(n32036), .B(n33402), .Z(n32038) );
  XNOR U32166 ( .A(q[5]), .B(DB[201]), .Z(n33402) );
  XNOR U32167 ( .A(q[4]), .B(DB[200]), .Z(n32036) );
  IV U32168 ( .A(n32050), .Z(n33400) );
  XOR U32169 ( .A(n33403), .B(n33404), .Z(n32050) );
  XNOR U32170 ( .A(n32046), .B(n32048), .Z(n33404) );
  XNOR U32171 ( .A(q[0]), .B(DB[196]), .Z(n32048) );
  XNOR U32172 ( .A(q[3]), .B(DB[199]), .Z(n32046) );
  IV U32173 ( .A(n32045), .Z(n33403) );
  XNOR U32174 ( .A(n32043), .B(n33405), .Z(n32045) );
  XNOR U32175 ( .A(q[2]), .B(DB[198]), .Z(n33405) );
  XNOR U32176 ( .A(q[1]), .B(DB[197]), .Z(n32043) );
  XOR U32177 ( .A(n33406), .B(n32008), .Z(n31971) );
  XOR U32178 ( .A(n33407), .B(n31996), .Z(n32008) );
  XNOR U32179 ( .A(q[6]), .B(DB[209]), .Z(n31996) );
  IV U32180 ( .A(n31995), .Z(n33407) );
  XNOR U32181 ( .A(n31993), .B(n33408), .Z(n31995) );
  XNOR U32182 ( .A(q[5]), .B(DB[208]), .Z(n33408) );
  XNOR U32183 ( .A(q[4]), .B(DB[207]), .Z(n31993) );
  IV U32184 ( .A(n32007), .Z(n33406) );
  XOR U32185 ( .A(n33409), .B(n33410), .Z(n32007) );
  XNOR U32186 ( .A(n32003), .B(n32005), .Z(n33410) );
  XNOR U32187 ( .A(q[0]), .B(DB[203]), .Z(n32005) );
  XNOR U32188 ( .A(q[3]), .B(DB[206]), .Z(n32003) );
  IV U32189 ( .A(n32002), .Z(n33409) );
  XNOR U32190 ( .A(n32000), .B(n33411), .Z(n32002) );
  XNOR U32191 ( .A(q[2]), .B(DB[205]), .Z(n33411) );
  XNOR U32192 ( .A(q[1]), .B(DB[204]), .Z(n32000) );
  XOR U32193 ( .A(n33412), .B(n31965), .Z(n31928) );
  XOR U32194 ( .A(n33413), .B(n31953), .Z(n31965) );
  XNOR U32195 ( .A(q[6]), .B(DB[216]), .Z(n31953) );
  IV U32196 ( .A(n31952), .Z(n33413) );
  XNOR U32197 ( .A(n31950), .B(n33414), .Z(n31952) );
  XNOR U32198 ( .A(q[5]), .B(DB[215]), .Z(n33414) );
  XNOR U32199 ( .A(q[4]), .B(DB[214]), .Z(n31950) );
  IV U32200 ( .A(n31964), .Z(n33412) );
  XOR U32201 ( .A(n33415), .B(n33416), .Z(n31964) );
  XNOR U32202 ( .A(n31960), .B(n31962), .Z(n33416) );
  XNOR U32203 ( .A(q[0]), .B(DB[210]), .Z(n31962) );
  XNOR U32204 ( .A(q[3]), .B(DB[213]), .Z(n31960) );
  IV U32205 ( .A(n31959), .Z(n33415) );
  XNOR U32206 ( .A(n31957), .B(n33417), .Z(n31959) );
  XNOR U32207 ( .A(q[2]), .B(DB[212]), .Z(n33417) );
  XNOR U32208 ( .A(q[1]), .B(DB[211]), .Z(n31957) );
  XOR U32209 ( .A(n33418), .B(n31922), .Z(n31885) );
  XOR U32210 ( .A(n33419), .B(n31910), .Z(n31922) );
  XNOR U32211 ( .A(q[6]), .B(DB[223]), .Z(n31910) );
  IV U32212 ( .A(n31909), .Z(n33419) );
  XNOR U32213 ( .A(n31907), .B(n33420), .Z(n31909) );
  XNOR U32214 ( .A(q[5]), .B(DB[222]), .Z(n33420) );
  XNOR U32215 ( .A(q[4]), .B(DB[221]), .Z(n31907) );
  IV U32216 ( .A(n31921), .Z(n33418) );
  XOR U32217 ( .A(n33421), .B(n33422), .Z(n31921) );
  XNOR U32218 ( .A(n31917), .B(n31919), .Z(n33422) );
  XNOR U32219 ( .A(q[0]), .B(DB[217]), .Z(n31919) );
  XNOR U32220 ( .A(q[3]), .B(DB[220]), .Z(n31917) );
  IV U32221 ( .A(n31916), .Z(n33421) );
  XNOR U32222 ( .A(n31914), .B(n33423), .Z(n31916) );
  XNOR U32223 ( .A(q[2]), .B(DB[219]), .Z(n33423) );
  XNOR U32224 ( .A(q[1]), .B(DB[218]), .Z(n31914) );
  XOR U32225 ( .A(n33424), .B(n31879), .Z(n31842) );
  XOR U32226 ( .A(n33425), .B(n31867), .Z(n31879) );
  XNOR U32227 ( .A(q[6]), .B(DB[230]), .Z(n31867) );
  IV U32228 ( .A(n31866), .Z(n33425) );
  XNOR U32229 ( .A(n31864), .B(n33426), .Z(n31866) );
  XNOR U32230 ( .A(q[5]), .B(DB[229]), .Z(n33426) );
  XNOR U32231 ( .A(q[4]), .B(DB[228]), .Z(n31864) );
  IV U32232 ( .A(n31878), .Z(n33424) );
  XOR U32233 ( .A(n33427), .B(n33428), .Z(n31878) );
  XNOR U32234 ( .A(n31874), .B(n31876), .Z(n33428) );
  XNOR U32235 ( .A(q[0]), .B(DB[224]), .Z(n31876) );
  XNOR U32236 ( .A(q[3]), .B(DB[227]), .Z(n31874) );
  IV U32237 ( .A(n31873), .Z(n33427) );
  XNOR U32238 ( .A(n31871), .B(n33429), .Z(n31873) );
  XNOR U32239 ( .A(q[2]), .B(DB[226]), .Z(n33429) );
  XNOR U32240 ( .A(q[1]), .B(DB[225]), .Z(n31871) );
  XOR U32241 ( .A(n33430), .B(n31836), .Z(n31799) );
  XOR U32242 ( .A(n33431), .B(n31824), .Z(n31836) );
  XNOR U32243 ( .A(q[6]), .B(DB[237]), .Z(n31824) );
  IV U32244 ( .A(n31823), .Z(n33431) );
  XNOR U32245 ( .A(n31821), .B(n33432), .Z(n31823) );
  XNOR U32246 ( .A(q[5]), .B(DB[236]), .Z(n33432) );
  XNOR U32247 ( .A(q[4]), .B(DB[235]), .Z(n31821) );
  IV U32248 ( .A(n31835), .Z(n33430) );
  XOR U32249 ( .A(n33433), .B(n33434), .Z(n31835) );
  XNOR U32250 ( .A(n31831), .B(n31833), .Z(n33434) );
  XNOR U32251 ( .A(q[0]), .B(DB[231]), .Z(n31833) );
  XNOR U32252 ( .A(q[3]), .B(DB[234]), .Z(n31831) );
  IV U32253 ( .A(n31830), .Z(n33433) );
  XNOR U32254 ( .A(n31828), .B(n33435), .Z(n31830) );
  XNOR U32255 ( .A(q[2]), .B(DB[233]), .Z(n33435) );
  XNOR U32256 ( .A(q[1]), .B(DB[232]), .Z(n31828) );
  XOR U32257 ( .A(n33436), .B(n31793), .Z(n31756) );
  XOR U32258 ( .A(n33437), .B(n31781), .Z(n31793) );
  XNOR U32259 ( .A(q[6]), .B(DB[244]), .Z(n31781) );
  IV U32260 ( .A(n31780), .Z(n33437) );
  XNOR U32261 ( .A(n31778), .B(n33438), .Z(n31780) );
  XNOR U32262 ( .A(q[5]), .B(DB[243]), .Z(n33438) );
  XNOR U32263 ( .A(q[4]), .B(DB[242]), .Z(n31778) );
  IV U32264 ( .A(n31792), .Z(n33436) );
  XOR U32265 ( .A(n33439), .B(n33440), .Z(n31792) );
  XNOR U32266 ( .A(n31788), .B(n31790), .Z(n33440) );
  XNOR U32267 ( .A(q[0]), .B(DB[238]), .Z(n31790) );
  XNOR U32268 ( .A(q[3]), .B(DB[241]), .Z(n31788) );
  IV U32269 ( .A(n31787), .Z(n33439) );
  XNOR U32270 ( .A(n31785), .B(n33441), .Z(n31787) );
  XNOR U32271 ( .A(q[2]), .B(DB[240]), .Z(n33441) );
  XNOR U32272 ( .A(q[1]), .B(DB[239]), .Z(n31785) );
  XOR U32273 ( .A(n33442), .B(n31750), .Z(n31713) );
  XOR U32274 ( .A(n33443), .B(n31738), .Z(n31750) );
  XNOR U32275 ( .A(q[6]), .B(DB[251]), .Z(n31738) );
  IV U32276 ( .A(n31737), .Z(n33443) );
  XNOR U32277 ( .A(n31735), .B(n33444), .Z(n31737) );
  XNOR U32278 ( .A(q[5]), .B(DB[250]), .Z(n33444) );
  XNOR U32279 ( .A(q[4]), .B(DB[249]), .Z(n31735) );
  IV U32280 ( .A(n31749), .Z(n33442) );
  XOR U32281 ( .A(n33445), .B(n33446), .Z(n31749) );
  XNOR U32282 ( .A(n31745), .B(n31747), .Z(n33446) );
  XNOR U32283 ( .A(q[0]), .B(DB[245]), .Z(n31747) );
  XNOR U32284 ( .A(q[3]), .B(DB[248]), .Z(n31745) );
  IV U32285 ( .A(n31744), .Z(n33445) );
  XNOR U32286 ( .A(n31742), .B(n33447), .Z(n31744) );
  XNOR U32287 ( .A(q[2]), .B(DB[247]), .Z(n33447) );
  XNOR U32288 ( .A(q[1]), .B(DB[246]), .Z(n31742) );
  XOR U32289 ( .A(n33448), .B(n31707), .Z(n31670) );
  XOR U32290 ( .A(n33449), .B(n31695), .Z(n31707) );
  XNOR U32291 ( .A(q[6]), .B(DB[258]), .Z(n31695) );
  IV U32292 ( .A(n31694), .Z(n33449) );
  XNOR U32293 ( .A(n31692), .B(n33450), .Z(n31694) );
  XNOR U32294 ( .A(q[5]), .B(DB[257]), .Z(n33450) );
  XNOR U32295 ( .A(q[4]), .B(DB[256]), .Z(n31692) );
  IV U32296 ( .A(n31706), .Z(n33448) );
  XOR U32297 ( .A(n33451), .B(n33452), .Z(n31706) );
  XNOR U32298 ( .A(n31702), .B(n31704), .Z(n33452) );
  XNOR U32299 ( .A(q[0]), .B(DB[252]), .Z(n31704) );
  XNOR U32300 ( .A(q[3]), .B(DB[255]), .Z(n31702) );
  IV U32301 ( .A(n31701), .Z(n33451) );
  XNOR U32302 ( .A(n31699), .B(n33453), .Z(n31701) );
  XNOR U32303 ( .A(q[2]), .B(DB[254]), .Z(n33453) );
  XNOR U32304 ( .A(q[1]), .B(DB[253]), .Z(n31699) );
  XOR U32305 ( .A(n33454), .B(n31664), .Z(n31627) );
  XOR U32306 ( .A(n33455), .B(n31652), .Z(n31664) );
  XNOR U32307 ( .A(q[6]), .B(DB[265]), .Z(n31652) );
  IV U32308 ( .A(n31651), .Z(n33455) );
  XNOR U32309 ( .A(n31649), .B(n33456), .Z(n31651) );
  XNOR U32310 ( .A(q[5]), .B(DB[264]), .Z(n33456) );
  XNOR U32311 ( .A(q[4]), .B(DB[263]), .Z(n31649) );
  IV U32312 ( .A(n31663), .Z(n33454) );
  XOR U32313 ( .A(n33457), .B(n33458), .Z(n31663) );
  XNOR U32314 ( .A(n31659), .B(n31661), .Z(n33458) );
  XNOR U32315 ( .A(q[0]), .B(DB[259]), .Z(n31661) );
  XNOR U32316 ( .A(q[3]), .B(DB[262]), .Z(n31659) );
  IV U32317 ( .A(n31658), .Z(n33457) );
  XNOR U32318 ( .A(n31656), .B(n33459), .Z(n31658) );
  XNOR U32319 ( .A(q[2]), .B(DB[261]), .Z(n33459) );
  XNOR U32320 ( .A(q[1]), .B(DB[260]), .Z(n31656) );
  XOR U32321 ( .A(n33460), .B(n31621), .Z(n31584) );
  XOR U32322 ( .A(n33461), .B(n31609), .Z(n31621) );
  XNOR U32323 ( .A(q[6]), .B(DB[272]), .Z(n31609) );
  IV U32324 ( .A(n31608), .Z(n33461) );
  XNOR U32325 ( .A(n31606), .B(n33462), .Z(n31608) );
  XNOR U32326 ( .A(q[5]), .B(DB[271]), .Z(n33462) );
  XNOR U32327 ( .A(q[4]), .B(DB[270]), .Z(n31606) );
  IV U32328 ( .A(n31620), .Z(n33460) );
  XOR U32329 ( .A(n33463), .B(n33464), .Z(n31620) );
  XNOR U32330 ( .A(n31616), .B(n31618), .Z(n33464) );
  XNOR U32331 ( .A(q[0]), .B(DB[266]), .Z(n31618) );
  XNOR U32332 ( .A(q[3]), .B(DB[269]), .Z(n31616) );
  IV U32333 ( .A(n31615), .Z(n33463) );
  XNOR U32334 ( .A(n31613), .B(n33465), .Z(n31615) );
  XNOR U32335 ( .A(q[2]), .B(DB[268]), .Z(n33465) );
  XNOR U32336 ( .A(q[1]), .B(DB[267]), .Z(n31613) );
  XOR U32337 ( .A(n33466), .B(n31578), .Z(n31541) );
  XOR U32338 ( .A(n33467), .B(n31566), .Z(n31578) );
  XNOR U32339 ( .A(q[6]), .B(DB[279]), .Z(n31566) );
  IV U32340 ( .A(n31565), .Z(n33467) );
  XNOR U32341 ( .A(n31563), .B(n33468), .Z(n31565) );
  XNOR U32342 ( .A(q[5]), .B(DB[278]), .Z(n33468) );
  XNOR U32343 ( .A(q[4]), .B(DB[277]), .Z(n31563) );
  IV U32344 ( .A(n31577), .Z(n33466) );
  XOR U32345 ( .A(n33469), .B(n33470), .Z(n31577) );
  XNOR U32346 ( .A(n31573), .B(n31575), .Z(n33470) );
  XNOR U32347 ( .A(q[0]), .B(DB[273]), .Z(n31575) );
  XNOR U32348 ( .A(q[3]), .B(DB[276]), .Z(n31573) );
  IV U32349 ( .A(n31572), .Z(n33469) );
  XNOR U32350 ( .A(n31570), .B(n33471), .Z(n31572) );
  XNOR U32351 ( .A(q[2]), .B(DB[275]), .Z(n33471) );
  XNOR U32352 ( .A(q[1]), .B(DB[274]), .Z(n31570) );
  XOR U32353 ( .A(n33472), .B(n31535), .Z(n31498) );
  XOR U32354 ( .A(n33473), .B(n31523), .Z(n31535) );
  XNOR U32355 ( .A(q[6]), .B(DB[286]), .Z(n31523) );
  IV U32356 ( .A(n31522), .Z(n33473) );
  XNOR U32357 ( .A(n31520), .B(n33474), .Z(n31522) );
  XNOR U32358 ( .A(q[5]), .B(DB[285]), .Z(n33474) );
  XNOR U32359 ( .A(q[4]), .B(DB[284]), .Z(n31520) );
  IV U32360 ( .A(n31534), .Z(n33472) );
  XOR U32361 ( .A(n33475), .B(n33476), .Z(n31534) );
  XNOR U32362 ( .A(n31530), .B(n31532), .Z(n33476) );
  XNOR U32363 ( .A(q[0]), .B(DB[280]), .Z(n31532) );
  XNOR U32364 ( .A(q[3]), .B(DB[283]), .Z(n31530) );
  IV U32365 ( .A(n31529), .Z(n33475) );
  XNOR U32366 ( .A(n31527), .B(n33477), .Z(n31529) );
  XNOR U32367 ( .A(q[2]), .B(DB[282]), .Z(n33477) );
  XNOR U32368 ( .A(q[1]), .B(DB[281]), .Z(n31527) );
  XOR U32369 ( .A(n33478), .B(n31492), .Z(n31455) );
  XOR U32370 ( .A(n33479), .B(n31480), .Z(n31492) );
  XNOR U32371 ( .A(q[6]), .B(DB[293]), .Z(n31480) );
  IV U32372 ( .A(n31479), .Z(n33479) );
  XNOR U32373 ( .A(n31477), .B(n33480), .Z(n31479) );
  XNOR U32374 ( .A(q[5]), .B(DB[292]), .Z(n33480) );
  XNOR U32375 ( .A(q[4]), .B(DB[291]), .Z(n31477) );
  IV U32376 ( .A(n31491), .Z(n33478) );
  XOR U32377 ( .A(n33481), .B(n33482), .Z(n31491) );
  XNOR U32378 ( .A(n31487), .B(n31489), .Z(n33482) );
  XNOR U32379 ( .A(q[0]), .B(DB[287]), .Z(n31489) );
  XNOR U32380 ( .A(q[3]), .B(DB[290]), .Z(n31487) );
  IV U32381 ( .A(n31486), .Z(n33481) );
  XNOR U32382 ( .A(n31484), .B(n33483), .Z(n31486) );
  XNOR U32383 ( .A(q[2]), .B(DB[289]), .Z(n33483) );
  XNOR U32384 ( .A(q[1]), .B(DB[288]), .Z(n31484) );
  XOR U32385 ( .A(n33484), .B(n31449), .Z(n31412) );
  XOR U32386 ( .A(n33485), .B(n31437), .Z(n31449) );
  XNOR U32387 ( .A(q[6]), .B(DB[300]), .Z(n31437) );
  IV U32388 ( .A(n31436), .Z(n33485) );
  XNOR U32389 ( .A(n31434), .B(n33486), .Z(n31436) );
  XNOR U32390 ( .A(q[5]), .B(DB[299]), .Z(n33486) );
  XNOR U32391 ( .A(q[4]), .B(DB[298]), .Z(n31434) );
  IV U32392 ( .A(n31448), .Z(n33484) );
  XOR U32393 ( .A(n33487), .B(n33488), .Z(n31448) );
  XNOR U32394 ( .A(n31444), .B(n31446), .Z(n33488) );
  XNOR U32395 ( .A(q[0]), .B(DB[294]), .Z(n31446) );
  XNOR U32396 ( .A(q[3]), .B(DB[297]), .Z(n31444) );
  IV U32397 ( .A(n31443), .Z(n33487) );
  XNOR U32398 ( .A(n31441), .B(n33489), .Z(n31443) );
  XNOR U32399 ( .A(q[2]), .B(DB[296]), .Z(n33489) );
  XNOR U32400 ( .A(q[1]), .B(DB[295]), .Z(n31441) );
  XOR U32401 ( .A(n33490), .B(n31406), .Z(n31369) );
  XOR U32402 ( .A(n33491), .B(n31394), .Z(n31406) );
  XNOR U32403 ( .A(q[6]), .B(DB[307]), .Z(n31394) );
  IV U32404 ( .A(n31393), .Z(n33491) );
  XNOR U32405 ( .A(n31391), .B(n33492), .Z(n31393) );
  XNOR U32406 ( .A(q[5]), .B(DB[306]), .Z(n33492) );
  XNOR U32407 ( .A(q[4]), .B(DB[305]), .Z(n31391) );
  IV U32408 ( .A(n31405), .Z(n33490) );
  XOR U32409 ( .A(n33493), .B(n33494), .Z(n31405) );
  XNOR U32410 ( .A(n31401), .B(n31403), .Z(n33494) );
  XNOR U32411 ( .A(q[0]), .B(DB[301]), .Z(n31403) );
  XNOR U32412 ( .A(q[3]), .B(DB[304]), .Z(n31401) );
  IV U32413 ( .A(n31400), .Z(n33493) );
  XNOR U32414 ( .A(n31398), .B(n33495), .Z(n31400) );
  XNOR U32415 ( .A(q[2]), .B(DB[303]), .Z(n33495) );
  XNOR U32416 ( .A(q[1]), .B(DB[302]), .Z(n31398) );
  XOR U32417 ( .A(n33496), .B(n31363), .Z(n31326) );
  XOR U32418 ( .A(n33497), .B(n31351), .Z(n31363) );
  XNOR U32419 ( .A(q[6]), .B(DB[314]), .Z(n31351) );
  IV U32420 ( .A(n31350), .Z(n33497) );
  XNOR U32421 ( .A(n31348), .B(n33498), .Z(n31350) );
  XNOR U32422 ( .A(q[5]), .B(DB[313]), .Z(n33498) );
  XNOR U32423 ( .A(q[4]), .B(DB[312]), .Z(n31348) );
  IV U32424 ( .A(n31362), .Z(n33496) );
  XOR U32425 ( .A(n33499), .B(n33500), .Z(n31362) );
  XNOR U32426 ( .A(n31358), .B(n31360), .Z(n33500) );
  XNOR U32427 ( .A(q[0]), .B(DB[308]), .Z(n31360) );
  XNOR U32428 ( .A(q[3]), .B(DB[311]), .Z(n31358) );
  IV U32429 ( .A(n31357), .Z(n33499) );
  XNOR U32430 ( .A(n31355), .B(n33501), .Z(n31357) );
  XNOR U32431 ( .A(q[2]), .B(DB[310]), .Z(n33501) );
  XNOR U32432 ( .A(q[1]), .B(DB[309]), .Z(n31355) );
  XOR U32433 ( .A(n33502), .B(n31320), .Z(n31283) );
  XOR U32434 ( .A(n33503), .B(n31308), .Z(n31320) );
  XNOR U32435 ( .A(q[6]), .B(DB[321]), .Z(n31308) );
  IV U32436 ( .A(n31307), .Z(n33503) );
  XNOR U32437 ( .A(n31305), .B(n33504), .Z(n31307) );
  XNOR U32438 ( .A(q[5]), .B(DB[320]), .Z(n33504) );
  XNOR U32439 ( .A(q[4]), .B(DB[319]), .Z(n31305) );
  IV U32440 ( .A(n31319), .Z(n33502) );
  XOR U32441 ( .A(n33505), .B(n33506), .Z(n31319) );
  XNOR U32442 ( .A(n31315), .B(n31317), .Z(n33506) );
  XNOR U32443 ( .A(q[0]), .B(DB[315]), .Z(n31317) );
  XNOR U32444 ( .A(q[3]), .B(DB[318]), .Z(n31315) );
  IV U32445 ( .A(n31314), .Z(n33505) );
  XNOR U32446 ( .A(n31312), .B(n33507), .Z(n31314) );
  XNOR U32447 ( .A(q[2]), .B(DB[317]), .Z(n33507) );
  XNOR U32448 ( .A(q[1]), .B(DB[316]), .Z(n31312) );
  XOR U32449 ( .A(n33508), .B(n31277), .Z(n31240) );
  XOR U32450 ( .A(n33509), .B(n31265), .Z(n31277) );
  XNOR U32451 ( .A(q[6]), .B(DB[328]), .Z(n31265) );
  IV U32452 ( .A(n31264), .Z(n33509) );
  XNOR U32453 ( .A(n31262), .B(n33510), .Z(n31264) );
  XNOR U32454 ( .A(q[5]), .B(DB[327]), .Z(n33510) );
  XNOR U32455 ( .A(q[4]), .B(DB[326]), .Z(n31262) );
  IV U32456 ( .A(n31276), .Z(n33508) );
  XOR U32457 ( .A(n33511), .B(n33512), .Z(n31276) );
  XNOR U32458 ( .A(n31272), .B(n31274), .Z(n33512) );
  XNOR U32459 ( .A(q[0]), .B(DB[322]), .Z(n31274) );
  XNOR U32460 ( .A(q[3]), .B(DB[325]), .Z(n31272) );
  IV U32461 ( .A(n31271), .Z(n33511) );
  XNOR U32462 ( .A(n31269), .B(n33513), .Z(n31271) );
  XNOR U32463 ( .A(q[2]), .B(DB[324]), .Z(n33513) );
  XNOR U32464 ( .A(q[1]), .B(DB[323]), .Z(n31269) );
  XOR U32465 ( .A(n33514), .B(n31234), .Z(n31197) );
  XOR U32466 ( .A(n33515), .B(n31222), .Z(n31234) );
  XNOR U32467 ( .A(q[6]), .B(DB[335]), .Z(n31222) );
  IV U32468 ( .A(n31221), .Z(n33515) );
  XNOR U32469 ( .A(n31219), .B(n33516), .Z(n31221) );
  XNOR U32470 ( .A(q[5]), .B(DB[334]), .Z(n33516) );
  XNOR U32471 ( .A(q[4]), .B(DB[333]), .Z(n31219) );
  IV U32472 ( .A(n31233), .Z(n33514) );
  XOR U32473 ( .A(n33517), .B(n33518), .Z(n31233) );
  XNOR U32474 ( .A(n31229), .B(n31231), .Z(n33518) );
  XNOR U32475 ( .A(q[0]), .B(DB[329]), .Z(n31231) );
  XNOR U32476 ( .A(q[3]), .B(DB[332]), .Z(n31229) );
  IV U32477 ( .A(n31228), .Z(n33517) );
  XNOR U32478 ( .A(n31226), .B(n33519), .Z(n31228) );
  XNOR U32479 ( .A(q[2]), .B(DB[331]), .Z(n33519) );
  XNOR U32480 ( .A(q[1]), .B(DB[330]), .Z(n31226) );
  XOR U32481 ( .A(n33520), .B(n31191), .Z(n31154) );
  XOR U32482 ( .A(n33521), .B(n31179), .Z(n31191) );
  XNOR U32483 ( .A(q[6]), .B(DB[342]), .Z(n31179) );
  IV U32484 ( .A(n31178), .Z(n33521) );
  XNOR U32485 ( .A(n31176), .B(n33522), .Z(n31178) );
  XNOR U32486 ( .A(q[5]), .B(DB[341]), .Z(n33522) );
  XNOR U32487 ( .A(q[4]), .B(DB[340]), .Z(n31176) );
  IV U32488 ( .A(n31190), .Z(n33520) );
  XOR U32489 ( .A(n33523), .B(n33524), .Z(n31190) );
  XNOR U32490 ( .A(n31186), .B(n31188), .Z(n33524) );
  XNOR U32491 ( .A(q[0]), .B(DB[336]), .Z(n31188) );
  XNOR U32492 ( .A(q[3]), .B(DB[339]), .Z(n31186) );
  IV U32493 ( .A(n31185), .Z(n33523) );
  XNOR U32494 ( .A(n31183), .B(n33525), .Z(n31185) );
  XNOR U32495 ( .A(q[2]), .B(DB[338]), .Z(n33525) );
  XNOR U32496 ( .A(q[1]), .B(DB[337]), .Z(n31183) );
  XOR U32497 ( .A(n33526), .B(n31148), .Z(n31111) );
  XOR U32498 ( .A(n33527), .B(n31136), .Z(n31148) );
  XNOR U32499 ( .A(q[6]), .B(DB[349]), .Z(n31136) );
  IV U32500 ( .A(n31135), .Z(n33527) );
  XNOR U32501 ( .A(n31133), .B(n33528), .Z(n31135) );
  XNOR U32502 ( .A(q[5]), .B(DB[348]), .Z(n33528) );
  XNOR U32503 ( .A(q[4]), .B(DB[347]), .Z(n31133) );
  IV U32504 ( .A(n31147), .Z(n33526) );
  XOR U32505 ( .A(n33529), .B(n33530), .Z(n31147) );
  XNOR U32506 ( .A(n31143), .B(n31145), .Z(n33530) );
  XNOR U32507 ( .A(q[0]), .B(DB[343]), .Z(n31145) );
  XNOR U32508 ( .A(q[3]), .B(DB[346]), .Z(n31143) );
  IV U32509 ( .A(n31142), .Z(n33529) );
  XNOR U32510 ( .A(n31140), .B(n33531), .Z(n31142) );
  XNOR U32511 ( .A(q[2]), .B(DB[345]), .Z(n33531) );
  XNOR U32512 ( .A(q[1]), .B(DB[344]), .Z(n31140) );
  XOR U32513 ( .A(n33532), .B(n31105), .Z(n31068) );
  XOR U32514 ( .A(n33533), .B(n31093), .Z(n31105) );
  XNOR U32515 ( .A(q[6]), .B(DB[356]), .Z(n31093) );
  IV U32516 ( .A(n31092), .Z(n33533) );
  XNOR U32517 ( .A(n31090), .B(n33534), .Z(n31092) );
  XNOR U32518 ( .A(q[5]), .B(DB[355]), .Z(n33534) );
  XNOR U32519 ( .A(q[4]), .B(DB[354]), .Z(n31090) );
  IV U32520 ( .A(n31104), .Z(n33532) );
  XOR U32521 ( .A(n33535), .B(n33536), .Z(n31104) );
  XNOR U32522 ( .A(n31100), .B(n31102), .Z(n33536) );
  XNOR U32523 ( .A(q[0]), .B(DB[350]), .Z(n31102) );
  XNOR U32524 ( .A(q[3]), .B(DB[353]), .Z(n31100) );
  IV U32525 ( .A(n31099), .Z(n33535) );
  XNOR U32526 ( .A(n31097), .B(n33537), .Z(n31099) );
  XNOR U32527 ( .A(q[2]), .B(DB[352]), .Z(n33537) );
  XNOR U32528 ( .A(q[1]), .B(DB[351]), .Z(n31097) );
  XOR U32529 ( .A(n33538), .B(n31062), .Z(n31025) );
  XOR U32530 ( .A(n33539), .B(n31050), .Z(n31062) );
  XNOR U32531 ( .A(q[6]), .B(DB[363]), .Z(n31050) );
  IV U32532 ( .A(n31049), .Z(n33539) );
  XNOR U32533 ( .A(n31047), .B(n33540), .Z(n31049) );
  XNOR U32534 ( .A(q[5]), .B(DB[362]), .Z(n33540) );
  XNOR U32535 ( .A(q[4]), .B(DB[361]), .Z(n31047) );
  IV U32536 ( .A(n31061), .Z(n33538) );
  XOR U32537 ( .A(n33541), .B(n33542), .Z(n31061) );
  XNOR U32538 ( .A(n31057), .B(n31059), .Z(n33542) );
  XNOR U32539 ( .A(q[0]), .B(DB[357]), .Z(n31059) );
  XNOR U32540 ( .A(q[3]), .B(DB[360]), .Z(n31057) );
  IV U32541 ( .A(n31056), .Z(n33541) );
  XNOR U32542 ( .A(n31054), .B(n33543), .Z(n31056) );
  XNOR U32543 ( .A(q[2]), .B(DB[359]), .Z(n33543) );
  XNOR U32544 ( .A(q[1]), .B(DB[358]), .Z(n31054) );
  XOR U32545 ( .A(n33544), .B(n31019), .Z(n30982) );
  XOR U32546 ( .A(n33545), .B(n31007), .Z(n31019) );
  XNOR U32547 ( .A(q[6]), .B(DB[370]), .Z(n31007) );
  IV U32548 ( .A(n31006), .Z(n33545) );
  XNOR U32549 ( .A(n31004), .B(n33546), .Z(n31006) );
  XNOR U32550 ( .A(q[5]), .B(DB[369]), .Z(n33546) );
  XNOR U32551 ( .A(q[4]), .B(DB[368]), .Z(n31004) );
  IV U32552 ( .A(n31018), .Z(n33544) );
  XOR U32553 ( .A(n33547), .B(n33548), .Z(n31018) );
  XNOR U32554 ( .A(n31014), .B(n31016), .Z(n33548) );
  XNOR U32555 ( .A(q[0]), .B(DB[364]), .Z(n31016) );
  XNOR U32556 ( .A(q[3]), .B(DB[367]), .Z(n31014) );
  IV U32557 ( .A(n31013), .Z(n33547) );
  XNOR U32558 ( .A(n31011), .B(n33549), .Z(n31013) );
  XNOR U32559 ( .A(q[2]), .B(DB[366]), .Z(n33549) );
  XNOR U32560 ( .A(q[1]), .B(DB[365]), .Z(n31011) );
  XOR U32561 ( .A(n33550), .B(n30976), .Z(n30939) );
  XOR U32562 ( .A(n33551), .B(n30964), .Z(n30976) );
  XNOR U32563 ( .A(q[6]), .B(DB[377]), .Z(n30964) );
  IV U32564 ( .A(n30963), .Z(n33551) );
  XNOR U32565 ( .A(n30961), .B(n33552), .Z(n30963) );
  XNOR U32566 ( .A(q[5]), .B(DB[376]), .Z(n33552) );
  XNOR U32567 ( .A(q[4]), .B(DB[375]), .Z(n30961) );
  IV U32568 ( .A(n30975), .Z(n33550) );
  XOR U32569 ( .A(n33553), .B(n33554), .Z(n30975) );
  XNOR U32570 ( .A(n30971), .B(n30973), .Z(n33554) );
  XNOR U32571 ( .A(q[0]), .B(DB[371]), .Z(n30973) );
  XNOR U32572 ( .A(q[3]), .B(DB[374]), .Z(n30971) );
  IV U32573 ( .A(n30970), .Z(n33553) );
  XNOR U32574 ( .A(n30968), .B(n33555), .Z(n30970) );
  XNOR U32575 ( .A(q[2]), .B(DB[373]), .Z(n33555) );
  XNOR U32576 ( .A(q[1]), .B(DB[372]), .Z(n30968) );
  XOR U32577 ( .A(n33556), .B(n30933), .Z(n30896) );
  XOR U32578 ( .A(n33557), .B(n30921), .Z(n30933) );
  XNOR U32579 ( .A(q[6]), .B(DB[384]), .Z(n30921) );
  IV U32580 ( .A(n30920), .Z(n33557) );
  XNOR U32581 ( .A(n30918), .B(n33558), .Z(n30920) );
  XNOR U32582 ( .A(q[5]), .B(DB[383]), .Z(n33558) );
  XNOR U32583 ( .A(q[4]), .B(DB[382]), .Z(n30918) );
  IV U32584 ( .A(n30932), .Z(n33556) );
  XOR U32585 ( .A(n33559), .B(n33560), .Z(n30932) );
  XNOR U32586 ( .A(n30928), .B(n30930), .Z(n33560) );
  XNOR U32587 ( .A(q[0]), .B(DB[378]), .Z(n30930) );
  XNOR U32588 ( .A(q[3]), .B(DB[381]), .Z(n30928) );
  IV U32589 ( .A(n30927), .Z(n33559) );
  XNOR U32590 ( .A(n30925), .B(n33561), .Z(n30927) );
  XNOR U32591 ( .A(q[2]), .B(DB[380]), .Z(n33561) );
  XNOR U32592 ( .A(q[1]), .B(DB[379]), .Z(n30925) );
  XOR U32593 ( .A(n33562), .B(n30890), .Z(n30853) );
  XOR U32594 ( .A(n33563), .B(n30878), .Z(n30890) );
  XNOR U32595 ( .A(q[6]), .B(DB[391]), .Z(n30878) );
  IV U32596 ( .A(n30877), .Z(n33563) );
  XNOR U32597 ( .A(n30875), .B(n33564), .Z(n30877) );
  XNOR U32598 ( .A(q[5]), .B(DB[390]), .Z(n33564) );
  XNOR U32599 ( .A(q[4]), .B(DB[389]), .Z(n30875) );
  IV U32600 ( .A(n30889), .Z(n33562) );
  XOR U32601 ( .A(n33565), .B(n33566), .Z(n30889) );
  XNOR U32602 ( .A(n30885), .B(n30887), .Z(n33566) );
  XNOR U32603 ( .A(q[0]), .B(DB[385]), .Z(n30887) );
  XNOR U32604 ( .A(q[3]), .B(DB[388]), .Z(n30885) );
  IV U32605 ( .A(n30884), .Z(n33565) );
  XNOR U32606 ( .A(n30882), .B(n33567), .Z(n30884) );
  XNOR U32607 ( .A(q[2]), .B(DB[387]), .Z(n33567) );
  XNOR U32608 ( .A(q[1]), .B(DB[386]), .Z(n30882) );
  XOR U32609 ( .A(n33568), .B(n30847), .Z(n30810) );
  XOR U32610 ( .A(n33569), .B(n30835), .Z(n30847) );
  XNOR U32611 ( .A(q[6]), .B(DB[398]), .Z(n30835) );
  IV U32612 ( .A(n30834), .Z(n33569) );
  XNOR U32613 ( .A(n30832), .B(n33570), .Z(n30834) );
  XNOR U32614 ( .A(q[5]), .B(DB[397]), .Z(n33570) );
  XNOR U32615 ( .A(q[4]), .B(DB[396]), .Z(n30832) );
  IV U32616 ( .A(n30846), .Z(n33568) );
  XOR U32617 ( .A(n33571), .B(n33572), .Z(n30846) );
  XNOR U32618 ( .A(n30842), .B(n30844), .Z(n33572) );
  XNOR U32619 ( .A(q[0]), .B(DB[392]), .Z(n30844) );
  XNOR U32620 ( .A(q[3]), .B(DB[395]), .Z(n30842) );
  IV U32621 ( .A(n30841), .Z(n33571) );
  XNOR U32622 ( .A(n30839), .B(n33573), .Z(n30841) );
  XNOR U32623 ( .A(q[2]), .B(DB[394]), .Z(n33573) );
  XNOR U32624 ( .A(q[1]), .B(DB[393]), .Z(n30839) );
  XOR U32625 ( .A(n33574), .B(n30804), .Z(n30767) );
  XOR U32626 ( .A(n33575), .B(n30792), .Z(n30804) );
  XNOR U32627 ( .A(q[6]), .B(DB[405]), .Z(n30792) );
  IV U32628 ( .A(n30791), .Z(n33575) );
  XNOR U32629 ( .A(n30789), .B(n33576), .Z(n30791) );
  XNOR U32630 ( .A(q[5]), .B(DB[404]), .Z(n33576) );
  XNOR U32631 ( .A(q[4]), .B(DB[403]), .Z(n30789) );
  IV U32632 ( .A(n30803), .Z(n33574) );
  XOR U32633 ( .A(n33577), .B(n33578), .Z(n30803) );
  XNOR U32634 ( .A(n30799), .B(n30801), .Z(n33578) );
  XNOR U32635 ( .A(q[0]), .B(DB[399]), .Z(n30801) );
  XNOR U32636 ( .A(q[3]), .B(DB[402]), .Z(n30799) );
  IV U32637 ( .A(n30798), .Z(n33577) );
  XNOR U32638 ( .A(n30796), .B(n33579), .Z(n30798) );
  XNOR U32639 ( .A(q[2]), .B(DB[401]), .Z(n33579) );
  XNOR U32640 ( .A(q[1]), .B(DB[400]), .Z(n30796) );
  XOR U32641 ( .A(n33580), .B(n30761), .Z(n30724) );
  XOR U32642 ( .A(n33581), .B(n30749), .Z(n30761) );
  XNOR U32643 ( .A(q[6]), .B(DB[412]), .Z(n30749) );
  IV U32644 ( .A(n30748), .Z(n33581) );
  XNOR U32645 ( .A(n30746), .B(n33582), .Z(n30748) );
  XNOR U32646 ( .A(q[5]), .B(DB[411]), .Z(n33582) );
  XNOR U32647 ( .A(q[4]), .B(DB[410]), .Z(n30746) );
  IV U32648 ( .A(n30760), .Z(n33580) );
  XOR U32649 ( .A(n33583), .B(n33584), .Z(n30760) );
  XNOR U32650 ( .A(n30756), .B(n30758), .Z(n33584) );
  XNOR U32651 ( .A(q[0]), .B(DB[406]), .Z(n30758) );
  XNOR U32652 ( .A(q[3]), .B(DB[409]), .Z(n30756) );
  IV U32653 ( .A(n30755), .Z(n33583) );
  XNOR U32654 ( .A(n30753), .B(n33585), .Z(n30755) );
  XNOR U32655 ( .A(q[2]), .B(DB[408]), .Z(n33585) );
  XNOR U32656 ( .A(q[1]), .B(DB[407]), .Z(n30753) );
  XOR U32657 ( .A(n33586), .B(n30718), .Z(n30681) );
  XOR U32658 ( .A(n33587), .B(n30706), .Z(n30718) );
  XNOR U32659 ( .A(q[6]), .B(DB[419]), .Z(n30706) );
  IV U32660 ( .A(n30705), .Z(n33587) );
  XNOR U32661 ( .A(n30703), .B(n33588), .Z(n30705) );
  XNOR U32662 ( .A(q[5]), .B(DB[418]), .Z(n33588) );
  XNOR U32663 ( .A(q[4]), .B(DB[417]), .Z(n30703) );
  IV U32664 ( .A(n30717), .Z(n33586) );
  XOR U32665 ( .A(n33589), .B(n33590), .Z(n30717) );
  XNOR U32666 ( .A(n30713), .B(n30715), .Z(n33590) );
  XNOR U32667 ( .A(q[0]), .B(DB[413]), .Z(n30715) );
  XNOR U32668 ( .A(q[3]), .B(DB[416]), .Z(n30713) );
  IV U32669 ( .A(n30712), .Z(n33589) );
  XNOR U32670 ( .A(n30710), .B(n33591), .Z(n30712) );
  XNOR U32671 ( .A(q[2]), .B(DB[415]), .Z(n33591) );
  XNOR U32672 ( .A(q[1]), .B(DB[414]), .Z(n30710) );
  XOR U32673 ( .A(n33592), .B(n30675), .Z(n30638) );
  XOR U32674 ( .A(n33593), .B(n30663), .Z(n30675) );
  XNOR U32675 ( .A(q[6]), .B(DB[426]), .Z(n30663) );
  IV U32676 ( .A(n30662), .Z(n33593) );
  XNOR U32677 ( .A(n30660), .B(n33594), .Z(n30662) );
  XNOR U32678 ( .A(q[5]), .B(DB[425]), .Z(n33594) );
  XNOR U32679 ( .A(q[4]), .B(DB[424]), .Z(n30660) );
  IV U32680 ( .A(n30674), .Z(n33592) );
  XOR U32681 ( .A(n33595), .B(n33596), .Z(n30674) );
  XNOR U32682 ( .A(n30670), .B(n30672), .Z(n33596) );
  XNOR U32683 ( .A(q[0]), .B(DB[420]), .Z(n30672) );
  XNOR U32684 ( .A(q[3]), .B(DB[423]), .Z(n30670) );
  IV U32685 ( .A(n30669), .Z(n33595) );
  XNOR U32686 ( .A(n30667), .B(n33597), .Z(n30669) );
  XNOR U32687 ( .A(q[2]), .B(DB[422]), .Z(n33597) );
  XNOR U32688 ( .A(q[1]), .B(DB[421]), .Z(n30667) );
  XOR U32689 ( .A(n33598), .B(n30632), .Z(n30595) );
  XOR U32690 ( .A(n33599), .B(n30620), .Z(n30632) );
  XNOR U32691 ( .A(q[6]), .B(DB[433]), .Z(n30620) );
  IV U32692 ( .A(n30619), .Z(n33599) );
  XNOR U32693 ( .A(n30617), .B(n33600), .Z(n30619) );
  XNOR U32694 ( .A(q[5]), .B(DB[432]), .Z(n33600) );
  XNOR U32695 ( .A(q[4]), .B(DB[431]), .Z(n30617) );
  IV U32696 ( .A(n30631), .Z(n33598) );
  XOR U32697 ( .A(n33601), .B(n33602), .Z(n30631) );
  XNOR U32698 ( .A(n30627), .B(n30629), .Z(n33602) );
  XNOR U32699 ( .A(q[0]), .B(DB[427]), .Z(n30629) );
  XNOR U32700 ( .A(q[3]), .B(DB[430]), .Z(n30627) );
  IV U32701 ( .A(n30626), .Z(n33601) );
  XNOR U32702 ( .A(n30624), .B(n33603), .Z(n30626) );
  XNOR U32703 ( .A(q[2]), .B(DB[429]), .Z(n33603) );
  XNOR U32704 ( .A(q[1]), .B(DB[428]), .Z(n30624) );
  XOR U32705 ( .A(n33604), .B(n30589), .Z(n30552) );
  XOR U32706 ( .A(n33605), .B(n30577), .Z(n30589) );
  XNOR U32707 ( .A(q[6]), .B(DB[440]), .Z(n30577) );
  IV U32708 ( .A(n30576), .Z(n33605) );
  XNOR U32709 ( .A(n30574), .B(n33606), .Z(n30576) );
  XNOR U32710 ( .A(q[5]), .B(DB[439]), .Z(n33606) );
  XNOR U32711 ( .A(q[4]), .B(DB[438]), .Z(n30574) );
  IV U32712 ( .A(n30588), .Z(n33604) );
  XOR U32713 ( .A(n33607), .B(n33608), .Z(n30588) );
  XNOR U32714 ( .A(n30584), .B(n30586), .Z(n33608) );
  XNOR U32715 ( .A(q[0]), .B(DB[434]), .Z(n30586) );
  XNOR U32716 ( .A(q[3]), .B(DB[437]), .Z(n30584) );
  IV U32717 ( .A(n30583), .Z(n33607) );
  XNOR U32718 ( .A(n30581), .B(n33609), .Z(n30583) );
  XNOR U32719 ( .A(q[2]), .B(DB[436]), .Z(n33609) );
  XNOR U32720 ( .A(q[1]), .B(DB[435]), .Z(n30581) );
  XOR U32721 ( .A(n33610), .B(n30546), .Z(n30509) );
  XOR U32722 ( .A(n33611), .B(n30534), .Z(n30546) );
  XNOR U32723 ( .A(q[6]), .B(DB[447]), .Z(n30534) );
  IV U32724 ( .A(n30533), .Z(n33611) );
  XNOR U32725 ( .A(n30531), .B(n33612), .Z(n30533) );
  XNOR U32726 ( .A(q[5]), .B(DB[446]), .Z(n33612) );
  XNOR U32727 ( .A(q[4]), .B(DB[445]), .Z(n30531) );
  IV U32728 ( .A(n30545), .Z(n33610) );
  XOR U32729 ( .A(n33613), .B(n33614), .Z(n30545) );
  XNOR U32730 ( .A(n30541), .B(n30543), .Z(n33614) );
  XNOR U32731 ( .A(q[0]), .B(DB[441]), .Z(n30543) );
  XNOR U32732 ( .A(q[3]), .B(DB[444]), .Z(n30541) );
  IV U32733 ( .A(n30540), .Z(n33613) );
  XNOR U32734 ( .A(n30538), .B(n33615), .Z(n30540) );
  XNOR U32735 ( .A(q[2]), .B(DB[443]), .Z(n33615) );
  XNOR U32736 ( .A(q[1]), .B(DB[442]), .Z(n30538) );
  XOR U32737 ( .A(n33616), .B(n30503), .Z(n30466) );
  XOR U32738 ( .A(n33617), .B(n30491), .Z(n30503) );
  XNOR U32739 ( .A(q[6]), .B(DB[454]), .Z(n30491) );
  IV U32740 ( .A(n30490), .Z(n33617) );
  XNOR U32741 ( .A(n30488), .B(n33618), .Z(n30490) );
  XNOR U32742 ( .A(q[5]), .B(DB[453]), .Z(n33618) );
  XNOR U32743 ( .A(q[4]), .B(DB[452]), .Z(n30488) );
  IV U32744 ( .A(n30502), .Z(n33616) );
  XOR U32745 ( .A(n33619), .B(n33620), .Z(n30502) );
  XNOR U32746 ( .A(n30498), .B(n30500), .Z(n33620) );
  XNOR U32747 ( .A(q[0]), .B(DB[448]), .Z(n30500) );
  XNOR U32748 ( .A(q[3]), .B(DB[451]), .Z(n30498) );
  IV U32749 ( .A(n30497), .Z(n33619) );
  XNOR U32750 ( .A(n30495), .B(n33621), .Z(n30497) );
  XNOR U32751 ( .A(q[2]), .B(DB[450]), .Z(n33621) );
  XNOR U32752 ( .A(q[1]), .B(DB[449]), .Z(n30495) );
  XOR U32753 ( .A(n33622), .B(n30460), .Z(n30423) );
  XOR U32754 ( .A(n33623), .B(n30448), .Z(n30460) );
  XNOR U32755 ( .A(q[6]), .B(DB[461]), .Z(n30448) );
  IV U32756 ( .A(n30447), .Z(n33623) );
  XNOR U32757 ( .A(n30445), .B(n33624), .Z(n30447) );
  XNOR U32758 ( .A(q[5]), .B(DB[460]), .Z(n33624) );
  XNOR U32759 ( .A(q[4]), .B(DB[459]), .Z(n30445) );
  IV U32760 ( .A(n30459), .Z(n33622) );
  XOR U32761 ( .A(n33625), .B(n33626), .Z(n30459) );
  XNOR U32762 ( .A(n30455), .B(n30457), .Z(n33626) );
  XNOR U32763 ( .A(q[0]), .B(DB[455]), .Z(n30457) );
  XNOR U32764 ( .A(q[3]), .B(DB[458]), .Z(n30455) );
  IV U32765 ( .A(n30454), .Z(n33625) );
  XNOR U32766 ( .A(n30452), .B(n33627), .Z(n30454) );
  XNOR U32767 ( .A(q[2]), .B(DB[457]), .Z(n33627) );
  XNOR U32768 ( .A(q[1]), .B(DB[456]), .Z(n30452) );
  XOR U32769 ( .A(n33628), .B(n30417), .Z(n30380) );
  XOR U32770 ( .A(n33629), .B(n30405), .Z(n30417) );
  XNOR U32771 ( .A(q[6]), .B(DB[468]), .Z(n30405) );
  IV U32772 ( .A(n30404), .Z(n33629) );
  XNOR U32773 ( .A(n30402), .B(n33630), .Z(n30404) );
  XNOR U32774 ( .A(q[5]), .B(DB[467]), .Z(n33630) );
  XNOR U32775 ( .A(q[4]), .B(DB[466]), .Z(n30402) );
  IV U32776 ( .A(n30416), .Z(n33628) );
  XOR U32777 ( .A(n33631), .B(n33632), .Z(n30416) );
  XNOR U32778 ( .A(n30412), .B(n30414), .Z(n33632) );
  XNOR U32779 ( .A(q[0]), .B(DB[462]), .Z(n30414) );
  XNOR U32780 ( .A(q[3]), .B(DB[465]), .Z(n30412) );
  IV U32781 ( .A(n30411), .Z(n33631) );
  XNOR U32782 ( .A(n30409), .B(n33633), .Z(n30411) );
  XNOR U32783 ( .A(q[2]), .B(DB[464]), .Z(n33633) );
  XNOR U32784 ( .A(q[1]), .B(DB[463]), .Z(n30409) );
  XOR U32785 ( .A(n33634), .B(n30374), .Z(n30337) );
  XOR U32786 ( .A(n33635), .B(n30362), .Z(n30374) );
  XNOR U32787 ( .A(q[6]), .B(DB[475]), .Z(n30362) );
  IV U32788 ( .A(n30361), .Z(n33635) );
  XNOR U32789 ( .A(n30359), .B(n33636), .Z(n30361) );
  XNOR U32790 ( .A(q[5]), .B(DB[474]), .Z(n33636) );
  XNOR U32791 ( .A(q[4]), .B(DB[473]), .Z(n30359) );
  IV U32792 ( .A(n30373), .Z(n33634) );
  XOR U32793 ( .A(n33637), .B(n33638), .Z(n30373) );
  XNOR U32794 ( .A(n30369), .B(n30371), .Z(n33638) );
  XNOR U32795 ( .A(q[0]), .B(DB[469]), .Z(n30371) );
  XNOR U32796 ( .A(q[3]), .B(DB[472]), .Z(n30369) );
  IV U32797 ( .A(n30368), .Z(n33637) );
  XNOR U32798 ( .A(n30366), .B(n33639), .Z(n30368) );
  XNOR U32799 ( .A(q[2]), .B(DB[471]), .Z(n33639) );
  XNOR U32800 ( .A(q[1]), .B(DB[470]), .Z(n30366) );
  XOR U32801 ( .A(n33640), .B(n30331), .Z(n30294) );
  XOR U32802 ( .A(n33641), .B(n30319), .Z(n30331) );
  XNOR U32803 ( .A(q[6]), .B(DB[482]), .Z(n30319) );
  IV U32804 ( .A(n30318), .Z(n33641) );
  XNOR U32805 ( .A(n30316), .B(n33642), .Z(n30318) );
  XNOR U32806 ( .A(q[5]), .B(DB[481]), .Z(n33642) );
  XNOR U32807 ( .A(q[4]), .B(DB[480]), .Z(n30316) );
  IV U32808 ( .A(n30330), .Z(n33640) );
  XOR U32809 ( .A(n33643), .B(n33644), .Z(n30330) );
  XNOR U32810 ( .A(n30326), .B(n30328), .Z(n33644) );
  XNOR U32811 ( .A(q[0]), .B(DB[476]), .Z(n30328) );
  XNOR U32812 ( .A(q[3]), .B(DB[479]), .Z(n30326) );
  IV U32813 ( .A(n30325), .Z(n33643) );
  XNOR U32814 ( .A(n30323), .B(n33645), .Z(n30325) );
  XNOR U32815 ( .A(q[2]), .B(DB[478]), .Z(n33645) );
  XNOR U32816 ( .A(q[1]), .B(DB[477]), .Z(n30323) );
  XOR U32817 ( .A(n33646), .B(n30288), .Z(n30251) );
  XOR U32818 ( .A(n33647), .B(n30276), .Z(n30288) );
  XNOR U32819 ( .A(q[6]), .B(DB[489]), .Z(n30276) );
  IV U32820 ( .A(n30275), .Z(n33647) );
  XNOR U32821 ( .A(n30273), .B(n33648), .Z(n30275) );
  XNOR U32822 ( .A(q[5]), .B(DB[488]), .Z(n33648) );
  XNOR U32823 ( .A(q[4]), .B(DB[487]), .Z(n30273) );
  IV U32824 ( .A(n30287), .Z(n33646) );
  XOR U32825 ( .A(n33649), .B(n33650), .Z(n30287) );
  XNOR U32826 ( .A(n30283), .B(n30285), .Z(n33650) );
  XNOR U32827 ( .A(q[0]), .B(DB[483]), .Z(n30285) );
  XNOR U32828 ( .A(q[3]), .B(DB[486]), .Z(n30283) );
  IV U32829 ( .A(n30282), .Z(n33649) );
  XNOR U32830 ( .A(n30280), .B(n33651), .Z(n30282) );
  XNOR U32831 ( .A(q[2]), .B(DB[485]), .Z(n33651) );
  XNOR U32832 ( .A(q[1]), .B(DB[484]), .Z(n30280) );
  XOR U32833 ( .A(n33652), .B(n30245), .Z(n30208) );
  XOR U32834 ( .A(n33653), .B(n30233), .Z(n30245) );
  XNOR U32835 ( .A(q[6]), .B(DB[496]), .Z(n30233) );
  IV U32836 ( .A(n30232), .Z(n33653) );
  XNOR U32837 ( .A(n30230), .B(n33654), .Z(n30232) );
  XNOR U32838 ( .A(q[5]), .B(DB[495]), .Z(n33654) );
  XNOR U32839 ( .A(q[4]), .B(DB[494]), .Z(n30230) );
  IV U32840 ( .A(n30244), .Z(n33652) );
  XOR U32841 ( .A(n33655), .B(n33656), .Z(n30244) );
  XNOR U32842 ( .A(n30240), .B(n30242), .Z(n33656) );
  XNOR U32843 ( .A(q[0]), .B(DB[490]), .Z(n30242) );
  XNOR U32844 ( .A(q[3]), .B(DB[493]), .Z(n30240) );
  IV U32845 ( .A(n30239), .Z(n33655) );
  XNOR U32846 ( .A(n30237), .B(n33657), .Z(n30239) );
  XNOR U32847 ( .A(q[2]), .B(DB[492]), .Z(n33657) );
  XNOR U32848 ( .A(q[1]), .B(DB[491]), .Z(n30237) );
  XOR U32849 ( .A(n33658), .B(n30202), .Z(n30165) );
  XOR U32850 ( .A(n33659), .B(n30190), .Z(n30202) );
  XNOR U32851 ( .A(q[6]), .B(DB[503]), .Z(n30190) );
  IV U32852 ( .A(n30189), .Z(n33659) );
  XNOR U32853 ( .A(n30187), .B(n33660), .Z(n30189) );
  XNOR U32854 ( .A(q[5]), .B(DB[502]), .Z(n33660) );
  XNOR U32855 ( .A(q[4]), .B(DB[501]), .Z(n30187) );
  IV U32856 ( .A(n30201), .Z(n33658) );
  XOR U32857 ( .A(n33661), .B(n33662), .Z(n30201) );
  XNOR U32858 ( .A(n30197), .B(n30199), .Z(n33662) );
  XNOR U32859 ( .A(q[0]), .B(DB[497]), .Z(n30199) );
  XNOR U32860 ( .A(q[3]), .B(DB[500]), .Z(n30197) );
  IV U32861 ( .A(n30196), .Z(n33661) );
  XNOR U32862 ( .A(n30194), .B(n33663), .Z(n30196) );
  XNOR U32863 ( .A(q[2]), .B(DB[499]), .Z(n33663) );
  XNOR U32864 ( .A(q[1]), .B(DB[498]), .Z(n30194) );
  XOR U32865 ( .A(n33664), .B(n30159), .Z(n30122) );
  XOR U32866 ( .A(n33665), .B(n30147), .Z(n30159) );
  XNOR U32867 ( .A(q[6]), .B(DB[510]), .Z(n30147) );
  IV U32868 ( .A(n30146), .Z(n33665) );
  XNOR U32869 ( .A(n30144), .B(n33666), .Z(n30146) );
  XNOR U32870 ( .A(q[5]), .B(DB[509]), .Z(n33666) );
  XNOR U32871 ( .A(q[4]), .B(DB[508]), .Z(n30144) );
  IV U32872 ( .A(n30158), .Z(n33664) );
  XOR U32873 ( .A(n33667), .B(n33668), .Z(n30158) );
  XNOR U32874 ( .A(n30154), .B(n30156), .Z(n33668) );
  XNOR U32875 ( .A(q[0]), .B(DB[504]), .Z(n30156) );
  XNOR U32876 ( .A(q[3]), .B(DB[507]), .Z(n30154) );
  IV U32877 ( .A(n30153), .Z(n33667) );
  XNOR U32878 ( .A(n30151), .B(n33669), .Z(n30153) );
  XNOR U32879 ( .A(q[2]), .B(DB[506]), .Z(n33669) );
  XNOR U32880 ( .A(q[1]), .B(DB[505]), .Z(n30151) );
  XOR U32881 ( .A(n33670), .B(n30116), .Z(n30079) );
  XOR U32882 ( .A(n33671), .B(n30104), .Z(n30116) );
  XNOR U32883 ( .A(q[6]), .B(DB[517]), .Z(n30104) );
  IV U32884 ( .A(n30103), .Z(n33671) );
  XNOR U32885 ( .A(n30101), .B(n33672), .Z(n30103) );
  XNOR U32886 ( .A(q[5]), .B(DB[516]), .Z(n33672) );
  XNOR U32887 ( .A(q[4]), .B(DB[515]), .Z(n30101) );
  IV U32888 ( .A(n30115), .Z(n33670) );
  XOR U32889 ( .A(n33673), .B(n33674), .Z(n30115) );
  XNOR U32890 ( .A(n30111), .B(n30113), .Z(n33674) );
  XNOR U32891 ( .A(q[0]), .B(DB[511]), .Z(n30113) );
  XNOR U32892 ( .A(q[3]), .B(DB[514]), .Z(n30111) );
  IV U32893 ( .A(n30110), .Z(n33673) );
  XNOR U32894 ( .A(n30108), .B(n33675), .Z(n30110) );
  XNOR U32895 ( .A(q[2]), .B(DB[513]), .Z(n33675) );
  XNOR U32896 ( .A(q[1]), .B(DB[512]), .Z(n30108) );
  XOR U32897 ( .A(n33676), .B(n30073), .Z(n30036) );
  XOR U32898 ( .A(n33677), .B(n30061), .Z(n30073) );
  XNOR U32899 ( .A(q[6]), .B(DB[524]), .Z(n30061) );
  IV U32900 ( .A(n30060), .Z(n33677) );
  XNOR U32901 ( .A(n30058), .B(n33678), .Z(n30060) );
  XNOR U32902 ( .A(q[5]), .B(DB[523]), .Z(n33678) );
  XNOR U32903 ( .A(q[4]), .B(DB[522]), .Z(n30058) );
  IV U32904 ( .A(n30072), .Z(n33676) );
  XOR U32905 ( .A(n33679), .B(n33680), .Z(n30072) );
  XNOR U32906 ( .A(n30068), .B(n30070), .Z(n33680) );
  XNOR U32907 ( .A(q[0]), .B(DB[518]), .Z(n30070) );
  XNOR U32908 ( .A(q[3]), .B(DB[521]), .Z(n30068) );
  IV U32909 ( .A(n30067), .Z(n33679) );
  XNOR U32910 ( .A(n30065), .B(n33681), .Z(n30067) );
  XNOR U32911 ( .A(q[2]), .B(DB[520]), .Z(n33681) );
  XNOR U32912 ( .A(q[1]), .B(DB[519]), .Z(n30065) );
  XOR U32913 ( .A(n33682), .B(n30030), .Z(n29993) );
  XOR U32914 ( .A(n33683), .B(n30018), .Z(n30030) );
  XNOR U32915 ( .A(q[6]), .B(DB[531]), .Z(n30018) );
  IV U32916 ( .A(n30017), .Z(n33683) );
  XNOR U32917 ( .A(n30015), .B(n33684), .Z(n30017) );
  XNOR U32918 ( .A(q[5]), .B(DB[530]), .Z(n33684) );
  XNOR U32919 ( .A(q[4]), .B(DB[529]), .Z(n30015) );
  IV U32920 ( .A(n30029), .Z(n33682) );
  XOR U32921 ( .A(n33685), .B(n33686), .Z(n30029) );
  XNOR U32922 ( .A(n30025), .B(n30027), .Z(n33686) );
  XNOR U32923 ( .A(q[0]), .B(DB[525]), .Z(n30027) );
  XNOR U32924 ( .A(q[3]), .B(DB[528]), .Z(n30025) );
  IV U32925 ( .A(n30024), .Z(n33685) );
  XNOR U32926 ( .A(n30022), .B(n33687), .Z(n30024) );
  XNOR U32927 ( .A(q[2]), .B(DB[527]), .Z(n33687) );
  XNOR U32928 ( .A(q[1]), .B(DB[526]), .Z(n30022) );
  XOR U32929 ( .A(n33688), .B(n29987), .Z(n29950) );
  XOR U32930 ( .A(n33689), .B(n29975), .Z(n29987) );
  XNOR U32931 ( .A(q[6]), .B(DB[538]), .Z(n29975) );
  IV U32932 ( .A(n29974), .Z(n33689) );
  XNOR U32933 ( .A(n29972), .B(n33690), .Z(n29974) );
  XNOR U32934 ( .A(q[5]), .B(DB[537]), .Z(n33690) );
  XNOR U32935 ( .A(q[4]), .B(DB[536]), .Z(n29972) );
  IV U32936 ( .A(n29986), .Z(n33688) );
  XOR U32937 ( .A(n33691), .B(n33692), .Z(n29986) );
  XNOR U32938 ( .A(n29982), .B(n29984), .Z(n33692) );
  XNOR U32939 ( .A(q[0]), .B(DB[532]), .Z(n29984) );
  XNOR U32940 ( .A(q[3]), .B(DB[535]), .Z(n29982) );
  IV U32941 ( .A(n29981), .Z(n33691) );
  XNOR U32942 ( .A(n29979), .B(n33693), .Z(n29981) );
  XNOR U32943 ( .A(q[2]), .B(DB[534]), .Z(n33693) );
  XNOR U32944 ( .A(q[1]), .B(DB[533]), .Z(n29979) );
  XOR U32945 ( .A(n33694), .B(n29944), .Z(n29907) );
  XOR U32946 ( .A(n33695), .B(n29932), .Z(n29944) );
  XNOR U32947 ( .A(q[6]), .B(DB[545]), .Z(n29932) );
  IV U32948 ( .A(n29931), .Z(n33695) );
  XNOR U32949 ( .A(n29929), .B(n33696), .Z(n29931) );
  XNOR U32950 ( .A(q[5]), .B(DB[544]), .Z(n33696) );
  XNOR U32951 ( .A(q[4]), .B(DB[543]), .Z(n29929) );
  IV U32952 ( .A(n29943), .Z(n33694) );
  XOR U32953 ( .A(n33697), .B(n33698), .Z(n29943) );
  XNOR U32954 ( .A(n29939), .B(n29941), .Z(n33698) );
  XNOR U32955 ( .A(q[0]), .B(DB[539]), .Z(n29941) );
  XNOR U32956 ( .A(q[3]), .B(DB[542]), .Z(n29939) );
  IV U32957 ( .A(n29938), .Z(n33697) );
  XNOR U32958 ( .A(n29936), .B(n33699), .Z(n29938) );
  XNOR U32959 ( .A(q[2]), .B(DB[541]), .Z(n33699) );
  XNOR U32960 ( .A(q[1]), .B(DB[540]), .Z(n29936) );
  XOR U32961 ( .A(n33700), .B(n29901), .Z(n29864) );
  XOR U32962 ( .A(n33701), .B(n29889), .Z(n29901) );
  XNOR U32963 ( .A(q[6]), .B(DB[552]), .Z(n29889) );
  IV U32964 ( .A(n29888), .Z(n33701) );
  XNOR U32965 ( .A(n29886), .B(n33702), .Z(n29888) );
  XNOR U32966 ( .A(q[5]), .B(DB[551]), .Z(n33702) );
  XNOR U32967 ( .A(q[4]), .B(DB[550]), .Z(n29886) );
  IV U32968 ( .A(n29900), .Z(n33700) );
  XOR U32969 ( .A(n33703), .B(n33704), .Z(n29900) );
  XNOR U32970 ( .A(n29896), .B(n29898), .Z(n33704) );
  XNOR U32971 ( .A(q[0]), .B(DB[546]), .Z(n29898) );
  XNOR U32972 ( .A(q[3]), .B(DB[549]), .Z(n29896) );
  IV U32973 ( .A(n29895), .Z(n33703) );
  XNOR U32974 ( .A(n29893), .B(n33705), .Z(n29895) );
  XNOR U32975 ( .A(q[2]), .B(DB[548]), .Z(n33705) );
  XNOR U32976 ( .A(q[1]), .B(DB[547]), .Z(n29893) );
  XOR U32977 ( .A(n33706), .B(n29858), .Z(n29821) );
  XOR U32978 ( .A(n33707), .B(n29846), .Z(n29858) );
  XNOR U32979 ( .A(q[6]), .B(DB[559]), .Z(n29846) );
  IV U32980 ( .A(n29845), .Z(n33707) );
  XNOR U32981 ( .A(n29843), .B(n33708), .Z(n29845) );
  XNOR U32982 ( .A(q[5]), .B(DB[558]), .Z(n33708) );
  XNOR U32983 ( .A(q[4]), .B(DB[557]), .Z(n29843) );
  IV U32984 ( .A(n29857), .Z(n33706) );
  XOR U32985 ( .A(n33709), .B(n33710), .Z(n29857) );
  XNOR U32986 ( .A(n29853), .B(n29855), .Z(n33710) );
  XNOR U32987 ( .A(q[0]), .B(DB[553]), .Z(n29855) );
  XNOR U32988 ( .A(q[3]), .B(DB[556]), .Z(n29853) );
  IV U32989 ( .A(n29852), .Z(n33709) );
  XNOR U32990 ( .A(n29850), .B(n33711), .Z(n29852) );
  XNOR U32991 ( .A(q[2]), .B(DB[555]), .Z(n33711) );
  XNOR U32992 ( .A(q[1]), .B(DB[554]), .Z(n29850) );
  XOR U32993 ( .A(n33712), .B(n29815), .Z(n29778) );
  XOR U32994 ( .A(n33713), .B(n29803), .Z(n29815) );
  XNOR U32995 ( .A(q[6]), .B(DB[566]), .Z(n29803) );
  IV U32996 ( .A(n29802), .Z(n33713) );
  XNOR U32997 ( .A(n29800), .B(n33714), .Z(n29802) );
  XNOR U32998 ( .A(q[5]), .B(DB[565]), .Z(n33714) );
  XNOR U32999 ( .A(q[4]), .B(DB[564]), .Z(n29800) );
  IV U33000 ( .A(n29814), .Z(n33712) );
  XOR U33001 ( .A(n33715), .B(n33716), .Z(n29814) );
  XNOR U33002 ( .A(n29810), .B(n29812), .Z(n33716) );
  XNOR U33003 ( .A(q[0]), .B(DB[560]), .Z(n29812) );
  XNOR U33004 ( .A(q[3]), .B(DB[563]), .Z(n29810) );
  IV U33005 ( .A(n29809), .Z(n33715) );
  XNOR U33006 ( .A(n29807), .B(n33717), .Z(n29809) );
  XNOR U33007 ( .A(q[2]), .B(DB[562]), .Z(n33717) );
  XNOR U33008 ( .A(q[1]), .B(DB[561]), .Z(n29807) );
  XOR U33009 ( .A(n33718), .B(n29772), .Z(n29735) );
  XOR U33010 ( .A(n33719), .B(n29760), .Z(n29772) );
  XNOR U33011 ( .A(q[6]), .B(DB[573]), .Z(n29760) );
  IV U33012 ( .A(n29759), .Z(n33719) );
  XNOR U33013 ( .A(n29757), .B(n33720), .Z(n29759) );
  XNOR U33014 ( .A(q[5]), .B(DB[572]), .Z(n33720) );
  XNOR U33015 ( .A(q[4]), .B(DB[571]), .Z(n29757) );
  IV U33016 ( .A(n29771), .Z(n33718) );
  XOR U33017 ( .A(n33721), .B(n33722), .Z(n29771) );
  XNOR U33018 ( .A(n29767), .B(n29769), .Z(n33722) );
  XNOR U33019 ( .A(q[0]), .B(DB[567]), .Z(n29769) );
  XNOR U33020 ( .A(q[3]), .B(DB[570]), .Z(n29767) );
  IV U33021 ( .A(n29766), .Z(n33721) );
  XNOR U33022 ( .A(n29764), .B(n33723), .Z(n29766) );
  XNOR U33023 ( .A(q[2]), .B(DB[569]), .Z(n33723) );
  XNOR U33024 ( .A(q[1]), .B(DB[568]), .Z(n29764) );
  XOR U33025 ( .A(n33724), .B(n29729), .Z(n29692) );
  XOR U33026 ( .A(n33725), .B(n29717), .Z(n29729) );
  XNOR U33027 ( .A(q[6]), .B(DB[580]), .Z(n29717) );
  IV U33028 ( .A(n29716), .Z(n33725) );
  XNOR U33029 ( .A(n29714), .B(n33726), .Z(n29716) );
  XNOR U33030 ( .A(q[5]), .B(DB[579]), .Z(n33726) );
  XNOR U33031 ( .A(q[4]), .B(DB[578]), .Z(n29714) );
  IV U33032 ( .A(n29728), .Z(n33724) );
  XOR U33033 ( .A(n33727), .B(n33728), .Z(n29728) );
  XNOR U33034 ( .A(n29724), .B(n29726), .Z(n33728) );
  XNOR U33035 ( .A(q[0]), .B(DB[574]), .Z(n29726) );
  XNOR U33036 ( .A(q[3]), .B(DB[577]), .Z(n29724) );
  IV U33037 ( .A(n29723), .Z(n33727) );
  XNOR U33038 ( .A(n29721), .B(n33729), .Z(n29723) );
  XNOR U33039 ( .A(q[2]), .B(DB[576]), .Z(n33729) );
  XNOR U33040 ( .A(q[1]), .B(DB[575]), .Z(n29721) );
  XOR U33041 ( .A(n33730), .B(n29686), .Z(n29649) );
  XOR U33042 ( .A(n33731), .B(n29674), .Z(n29686) );
  XNOR U33043 ( .A(q[6]), .B(DB[587]), .Z(n29674) );
  IV U33044 ( .A(n29673), .Z(n33731) );
  XNOR U33045 ( .A(n29671), .B(n33732), .Z(n29673) );
  XNOR U33046 ( .A(q[5]), .B(DB[586]), .Z(n33732) );
  XNOR U33047 ( .A(q[4]), .B(DB[585]), .Z(n29671) );
  IV U33048 ( .A(n29685), .Z(n33730) );
  XOR U33049 ( .A(n33733), .B(n33734), .Z(n29685) );
  XNOR U33050 ( .A(n29681), .B(n29683), .Z(n33734) );
  XNOR U33051 ( .A(q[0]), .B(DB[581]), .Z(n29683) );
  XNOR U33052 ( .A(q[3]), .B(DB[584]), .Z(n29681) );
  IV U33053 ( .A(n29680), .Z(n33733) );
  XNOR U33054 ( .A(n29678), .B(n33735), .Z(n29680) );
  XNOR U33055 ( .A(q[2]), .B(DB[583]), .Z(n33735) );
  XNOR U33056 ( .A(q[1]), .B(DB[582]), .Z(n29678) );
  XOR U33057 ( .A(n33736), .B(n29643), .Z(n29606) );
  XOR U33058 ( .A(n33737), .B(n29631), .Z(n29643) );
  XNOR U33059 ( .A(q[6]), .B(DB[594]), .Z(n29631) );
  IV U33060 ( .A(n29630), .Z(n33737) );
  XNOR U33061 ( .A(n29628), .B(n33738), .Z(n29630) );
  XNOR U33062 ( .A(q[5]), .B(DB[593]), .Z(n33738) );
  XNOR U33063 ( .A(q[4]), .B(DB[592]), .Z(n29628) );
  IV U33064 ( .A(n29642), .Z(n33736) );
  XOR U33065 ( .A(n33739), .B(n33740), .Z(n29642) );
  XNOR U33066 ( .A(n29638), .B(n29640), .Z(n33740) );
  XNOR U33067 ( .A(q[0]), .B(DB[588]), .Z(n29640) );
  XNOR U33068 ( .A(q[3]), .B(DB[591]), .Z(n29638) );
  IV U33069 ( .A(n29637), .Z(n33739) );
  XNOR U33070 ( .A(n29635), .B(n33741), .Z(n29637) );
  XNOR U33071 ( .A(q[2]), .B(DB[590]), .Z(n33741) );
  XNOR U33072 ( .A(q[1]), .B(DB[589]), .Z(n29635) );
  XOR U33073 ( .A(n33742), .B(n29600), .Z(n29563) );
  XOR U33074 ( .A(n33743), .B(n29588), .Z(n29600) );
  XNOR U33075 ( .A(q[6]), .B(DB[601]), .Z(n29588) );
  IV U33076 ( .A(n29587), .Z(n33743) );
  XNOR U33077 ( .A(n29585), .B(n33744), .Z(n29587) );
  XNOR U33078 ( .A(q[5]), .B(DB[600]), .Z(n33744) );
  XNOR U33079 ( .A(q[4]), .B(DB[599]), .Z(n29585) );
  IV U33080 ( .A(n29599), .Z(n33742) );
  XOR U33081 ( .A(n33745), .B(n33746), .Z(n29599) );
  XNOR U33082 ( .A(n29595), .B(n29597), .Z(n33746) );
  XNOR U33083 ( .A(q[0]), .B(DB[595]), .Z(n29597) );
  XNOR U33084 ( .A(q[3]), .B(DB[598]), .Z(n29595) );
  IV U33085 ( .A(n29594), .Z(n33745) );
  XNOR U33086 ( .A(n29592), .B(n33747), .Z(n29594) );
  XNOR U33087 ( .A(q[2]), .B(DB[597]), .Z(n33747) );
  XNOR U33088 ( .A(q[1]), .B(DB[596]), .Z(n29592) );
  XOR U33089 ( .A(n33748), .B(n29557), .Z(n29520) );
  XOR U33090 ( .A(n33749), .B(n29545), .Z(n29557) );
  XNOR U33091 ( .A(q[6]), .B(DB[608]), .Z(n29545) );
  IV U33092 ( .A(n29544), .Z(n33749) );
  XNOR U33093 ( .A(n29542), .B(n33750), .Z(n29544) );
  XNOR U33094 ( .A(q[5]), .B(DB[607]), .Z(n33750) );
  XNOR U33095 ( .A(q[4]), .B(DB[606]), .Z(n29542) );
  IV U33096 ( .A(n29556), .Z(n33748) );
  XOR U33097 ( .A(n33751), .B(n33752), .Z(n29556) );
  XNOR U33098 ( .A(n29552), .B(n29554), .Z(n33752) );
  XNOR U33099 ( .A(q[0]), .B(DB[602]), .Z(n29554) );
  XNOR U33100 ( .A(q[3]), .B(DB[605]), .Z(n29552) );
  IV U33101 ( .A(n29551), .Z(n33751) );
  XNOR U33102 ( .A(n29549), .B(n33753), .Z(n29551) );
  XNOR U33103 ( .A(q[2]), .B(DB[604]), .Z(n33753) );
  XNOR U33104 ( .A(q[1]), .B(DB[603]), .Z(n29549) );
  XOR U33105 ( .A(n33754), .B(n29514), .Z(n29477) );
  XOR U33106 ( .A(n33755), .B(n29502), .Z(n29514) );
  XNOR U33107 ( .A(q[6]), .B(DB[615]), .Z(n29502) );
  IV U33108 ( .A(n29501), .Z(n33755) );
  XNOR U33109 ( .A(n29499), .B(n33756), .Z(n29501) );
  XNOR U33110 ( .A(q[5]), .B(DB[614]), .Z(n33756) );
  XNOR U33111 ( .A(q[4]), .B(DB[613]), .Z(n29499) );
  IV U33112 ( .A(n29513), .Z(n33754) );
  XOR U33113 ( .A(n33757), .B(n33758), .Z(n29513) );
  XNOR U33114 ( .A(n29509), .B(n29511), .Z(n33758) );
  XNOR U33115 ( .A(q[0]), .B(DB[609]), .Z(n29511) );
  XNOR U33116 ( .A(q[3]), .B(DB[612]), .Z(n29509) );
  IV U33117 ( .A(n29508), .Z(n33757) );
  XNOR U33118 ( .A(n29506), .B(n33759), .Z(n29508) );
  XNOR U33119 ( .A(q[2]), .B(DB[611]), .Z(n33759) );
  XNOR U33120 ( .A(q[1]), .B(DB[610]), .Z(n29506) );
  XOR U33121 ( .A(n33760), .B(n29471), .Z(n29434) );
  XOR U33122 ( .A(n33761), .B(n29459), .Z(n29471) );
  XNOR U33123 ( .A(q[6]), .B(DB[622]), .Z(n29459) );
  IV U33124 ( .A(n29458), .Z(n33761) );
  XNOR U33125 ( .A(n29456), .B(n33762), .Z(n29458) );
  XNOR U33126 ( .A(q[5]), .B(DB[621]), .Z(n33762) );
  XNOR U33127 ( .A(q[4]), .B(DB[620]), .Z(n29456) );
  IV U33128 ( .A(n29470), .Z(n33760) );
  XOR U33129 ( .A(n33763), .B(n33764), .Z(n29470) );
  XNOR U33130 ( .A(n29466), .B(n29468), .Z(n33764) );
  XNOR U33131 ( .A(q[0]), .B(DB[616]), .Z(n29468) );
  XNOR U33132 ( .A(q[3]), .B(DB[619]), .Z(n29466) );
  IV U33133 ( .A(n29465), .Z(n33763) );
  XNOR U33134 ( .A(n29463), .B(n33765), .Z(n29465) );
  XNOR U33135 ( .A(q[2]), .B(DB[618]), .Z(n33765) );
  XNOR U33136 ( .A(q[1]), .B(DB[617]), .Z(n29463) );
  XOR U33137 ( .A(n33766), .B(n29428), .Z(n29391) );
  XOR U33138 ( .A(n33767), .B(n29416), .Z(n29428) );
  XNOR U33139 ( .A(q[6]), .B(DB[629]), .Z(n29416) );
  IV U33140 ( .A(n29415), .Z(n33767) );
  XNOR U33141 ( .A(n29413), .B(n33768), .Z(n29415) );
  XNOR U33142 ( .A(q[5]), .B(DB[628]), .Z(n33768) );
  XNOR U33143 ( .A(q[4]), .B(DB[627]), .Z(n29413) );
  IV U33144 ( .A(n29427), .Z(n33766) );
  XOR U33145 ( .A(n33769), .B(n33770), .Z(n29427) );
  XNOR U33146 ( .A(n29423), .B(n29425), .Z(n33770) );
  XNOR U33147 ( .A(q[0]), .B(DB[623]), .Z(n29425) );
  XNOR U33148 ( .A(q[3]), .B(DB[626]), .Z(n29423) );
  IV U33149 ( .A(n29422), .Z(n33769) );
  XNOR U33150 ( .A(n29420), .B(n33771), .Z(n29422) );
  XNOR U33151 ( .A(q[2]), .B(DB[625]), .Z(n33771) );
  XNOR U33152 ( .A(q[1]), .B(DB[624]), .Z(n29420) );
  XOR U33153 ( .A(n33772), .B(n29385), .Z(n29348) );
  XOR U33154 ( .A(n33773), .B(n29373), .Z(n29385) );
  XNOR U33155 ( .A(q[6]), .B(DB[636]), .Z(n29373) );
  IV U33156 ( .A(n29372), .Z(n33773) );
  XNOR U33157 ( .A(n29370), .B(n33774), .Z(n29372) );
  XNOR U33158 ( .A(q[5]), .B(DB[635]), .Z(n33774) );
  XNOR U33159 ( .A(q[4]), .B(DB[634]), .Z(n29370) );
  IV U33160 ( .A(n29384), .Z(n33772) );
  XOR U33161 ( .A(n33775), .B(n33776), .Z(n29384) );
  XNOR U33162 ( .A(n29380), .B(n29382), .Z(n33776) );
  XNOR U33163 ( .A(q[0]), .B(DB[630]), .Z(n29382) );
  XNOR U33164 ( .A(q[3]), .B(DB[633]), .Z(n29380) );
  IV U33165 ( .A(n29379), .Z(n33775) );
  XNOR U33166 ( .A(n29377), .B(n33777), .Z(n29379) );
  XNOR U33167 ( .A(q[2]), .B(DB[632]), .Z(n33777) );
  XNOR U33168 ( .A(q[1]), .B(DB[631]), .Z(n29377) );
  XOR U33169 ( .A(n33778), .B(n29342), .Z(n29305) );
  XOR U33170 ( .A(n33779), .B(n29330), .Z(n29342) );
  XNOR U33171 ( .A(q[6]), .B(DB[643]), .Z(n29330) );
  IV U33172 ( .A(n29329), .Z(n33779) );
  XNOR U33173 ( .A(n29327), .B(n33780), .Z(n29329) );
  XNOR U33174 ( .A(q[5]), .B(DB[642]), .Z(n33780) );
  XNOR U33175 ( .A(q[4]), .B(DB[641]), .Z(n29327) );
  IV U33176 ( .A(n29341), .Z(n33778) );
  XOR U33177 ( .A(n33781), .B(n33782), .Z(n29341) );
  XNOR U33178 ( .A(n29337), .B(n29339), .Z(n33782) );
  XNOR U33179 ( .A(q[0]), .B(DB[637]), .Z(n29339) );
  XNOR U33180 ( .A(q[3]), .B(DB[640]), .Z(n29337) );
  IV U33181 ( .A(n29336), .Z(n33781) );
  XNOR U33182 ( .A(n29334), .B(n33783), .Z(n29336) );
  XNOR U33183 ( .A(q[2]), .B(DB[639]), .Z(n33783) );
  XNOR U33184 ( .A(q[1]), .B(DB[638]), .Z(n29334) );
  XOR U33185 ( .A(n33784), .B(n29299), .Z(n29262) );
  XOR U33186 ( .A(n33785), .B(n29287), .Z(n29299) );
  XNOR U33187 ( .A(q[6]), .B(DB[650]), .Z(n29287) );
  IV U33188 ( .A(n29286), .Z(n33785) );
  XNOR U33189 ( .A(n29284), .B(n33786), .Z(n29286) );
  XNOR U33190 ( .A(q[5]), .B(DB[649]), .Z(n33786) );
  XNOR U33191 ( .A(q[4]), .B(DB[648]), .Z(n29284) );
  IV U33192 ( .A(n29298), .Z(n33784) );
  XOR U33193 ( .A(n33787), .B(n33788), .Z(n29298) );
  XNOR U33194 ( .A(n29294), .B(n29296), .Z(n33788) );
  XNOR U33195 ( .A(q[0]), .B(DB[644]), .Z(n29296) );
  XNOR U33196 ( .A(q[3]), .B(DB[647]), .Z(n29294) );
  IV U33197 ( .A(n29293), .Z(n33787) );
  XNOR U33198 ( .A(n29291), .B(n33789), .Z(n29293) );
  XNOR U33199 ( .A(q[2]), .B(DB[646]), .Z(n33789) );
  XNOR U33200 ( .A(q[1]), .B(DB[645]), .Z(n29291) );
  XOR U33201 ( .A(n33790), .B(n29256), .Z(n29219) );
  XOR U33202 ( .A(n33791), .B(n29244), .Z(n29256) );
  XNOR U33203 ( .A(q[6]), .B(DB[657]), .Z(n29244) );
  IV U33204 ( .A(n29243), .Z(n33791) );
  XNOR U33205 ( .A(n29241), .B(n33792), .Z(n29243) );
  XNOR U33206 ( .A(q[5]), .B(DB[656]), .Z(n33792) );
  XNOR U33207 ( .A(q[4]), .B(DB[655]), .Z(n29241) );
  IV U33208 ( .A(n29255), .Z(n33790) );
  XOR U33209 ( .A(n33793), .B(n33794), .Z(n29255) );
  XNOR U33210 ( .A(n29251), .B(n29253), .Z(n33794) );
  XNOR U33211 ( .A(q[0]), .B(DB[651]), .Z(n29253) );
  XNOR U33212 ( .A(q[3]), .B(DB[654]), .Z(n29251) );
  IV U33213 ( .A(n29250), .Z(n33793) );
  XNOR U33214 ( .A(n29248), .B(n33795), .Z(n29250) );
  XNOR U33215 ( .A(q[2]), .B(DB[653]), .Z(n33795) );
  XNOR U33216 ( .A(q[1]), .B(DB[652]), .Z(n29248) );
  XOR U33217 ( .A(n33796), .B(n29213), .Z(n29176) );
  XOR U33218 ( .A(n33797), .B(n29201), .Z(n29213) );
  XNOR U33219 ( .A(q[6]), .B(DB[664]), .Z(n29201) );
  IV U33220 ( .A(n29200), .Z(n33797) );
  XNOR U33221 ( .A(n29198), .B(n33798), .Z(n29200) );
  XNOR U33222 ( .A(q[5]), .B(DB[663]), .Z(n33798) );
  XNOR U33223 ( .A(q[4]), .B(DB[662]), .Z(n29198) );
  IV U33224 ( .A(n29212), .Z(n33796) );
  XOR U33225 ( .A(n33799), .B(n33800), .Z(n29212) );
  XNOR U33226 ( .A(n29208), .B(n29210), .Z(n33800) );
  XNOR U33227 ( .A(q[0]), .B(DB[658]), .Z(n29210) );
  XNOR U33228 ( .A(q[3]), .B(DB[661]), .Z(n29208) );
  IV U33229 ( .A(n29207), .Z(n33799) );
  XNOR U33230 ( .A(n29205), .B(n33801), .Z(n29207) );
  XNOR U33231 ( .A(q[2]), .B(DB[660]), .Z(n33801) );
  XNOR U33232 ( .A(q[1]), .B(DB[659]), .Z(n29205) );
  XOR U33233 ( .A(n33802), .B(n29170), .Z(n29133) );
  XOR U33234 ( .A(n33803), .B(n29158), .Z(n29170) );
  XNOR U33235 ( .A(q[6]), .B(DB[671]), .Z(n29158) );
  IV U33236 ( .A(n29157), .Z(n33803) );
  XNOR U33237 ( .A(n29155), .B(n33804), .Z(n29157) );
  XNOR U33238 ( .A(q[5]), .B(DB[670]), .Z(n33804) );
  XNOR U33239 ( .A(q[4]), .B(DB[669]), .Z(n29155) );
  IV U33240 ( .A(n29169), .Z(n33802) );
  XOR U33241 ( .A(n33805), .B(n33806), .Z(n29169) );
  XNOR U33242 ( .A(n29165), .B(n29167), .Z(n33806) );
  XNOR U33243 ( .A(q[0]), .B(DB[665]), .Z(n29167) );
  XNOR U33244 ( .A(q[3]), .B(DB[668]), .Z(n29165) );
  IV U33245 ( .A(n29164), .Z(n33805) );
  XNOR U33246 ( .A(n29162), .B(n33807), .Z(n29164) );
  XNOR U33247 ( .A(q[2]), .B(DB[667]), .Z(n33807) );
  XNOR U33248 ( .A(q[1]), .B(DB[666]), .Z(n29162) );
  XOR U33249 ( .A(n33808), .B(n29127), .Z(n29090) );
  XOR U33250 ( .A(n33809), .B(n29115), .Z(n29127) );
  XNOR U33251 ( .A(q[6]), .B(DB[678]), .Z(n29115) );
  IV U33252 ( .A(n29114), .Z(n33809) );
  XNOR U33253 ( .A(n29112), .B(n33810), .Z(n29114) );
  XNOR U33254 ( .A(q[5]), .B(DB[677]), .Z(n33810) );
  XNOR U33255 ( .A(q[4]), .B(DB[676]), .Z(n29112) );
  IV U33256 ( .A(n29126), .Z(n33808) );
  XOR U33257 ( .A(n33811), .B(n33812), .Z(n29126) );
  XNOR U33258 ( .A(n29122), .B(n29124), .Z(n33812) );
  XNOR U33259 ( .A(q[0]), .B(DB[672]), .Z(n29124) );
  XNOR U33260 ( .A(q[3]), .B(DB[675]), .Z(n29122) );
  IV U33261 ( .A(n29121), .Z(n33811) );
  XNOR U33262 ( .A(n29119), .B(n33813), .Z(n29121) );
  XNOR U33263 ( .A(q[2]), .B(DB[674]), .Z(n33813) );
  XNOR U33264 ( .A(q[1]), .B(DB[673]), .Z(n29119) );
  XOR U33265 ( .A(n33814), .B(n29084), .Z(n29047) );
  XOR U33266 ( .A(n33815), .B(n29072), .Z(n29084) );
  XNOR U33267 ( .A(q[6]), .B(DB[685]), .Z(n29072) );
  IV U33268 ( .A(n29071), .Z(n33815) );
  XNOR U33269 ( .A(n29069), .B(n33816), .Z(n29071) );
  XNOR U33270 ( .A(q[5]), .B(DB[684]), .Z(n33816) );
  XNOR U33271 ( .A(q[4]), .B(DB[683]), .Z(n29069) );
  IV U33272 ( .A(n29083), .Z(n33814) );
  XOR U33273 ( .A(n33817), .B(n33818), .Z(n29083) );
  XNOR U33274 ( .A(n29079), .B(n29081), .Z(n33818) );
  XNOR U33275 ( .A(q[0]), .B(DB[679]), .Z(n29081) );
  XNOR U33276 ( .A(q[3]), .B(DB[682]), .Z(n29079) );
  IV U33277 ( .A(n29078), .Z(n33817) );
  XNOR U33278 ( .A(n29076), .B(n33819), .Z(n29078) );
  XNOR U33279 ( .A(q[2]), .B(DB[681]), .Z(n33819) );
  XNOR U33280 ( .A(q[1]), .B(DB[680]), .Z(n29076) );
  XOR U33281 ( .A(n33820), .B(n29041), .Z(n29004) );
  XOR U33282 ( .A(n33821), .B(n29029), .Z(n29041) );
  XNOR U33283 ( .A(q[6]), .B(DB[692]), .Z(n29029) );
  IV U33284 ( .A(n29028), .Z(n33821) );
  XNOR U33285 ( .A(n29026), .B(n33822), .Z(n29028) );
  XNOR U33286 ( .A(q[5]), .B(DB[691]), .Z(n33822) );
  XNOR U33287 ( .A(q[4]), .B(DB[690]), .Z(n29026) );
  IV U33288 ( .A(n29040), .Z(n33820) );
  XOR U33289 ( .A(n33823), .B(n33824), .Z(n29040) );
  XNOR U33290 ( .A(n29036), .B(n29038), .Z(n33824) );
  XNOR U33291 ( .A(q[0]), .B(DB[686]), .Z(n29038) );
  XNOR U33292 ( .A(q[3]), .B(DB[689]), .Z(n29036) );
  IV U33293 ( .A(n29035), .Z(n33823) );
  XNOR U33294 ( .A(n29033), .B(n33825), .Z(n29035) );
  XNOR U33295 ( .A(q[2]), .B(DB[688]), .Z(n33825) );
  XNOR U33296 ( .A(q[1]), .B(DB[687]), .Z(n29033) );
  XOR U33297 ( .A(n33826), .B(n28998), .Z(n28961) );
  XOR U33298 ( .A(n33827), .B(n28986), .Z(n28998) );
  XNOR U33299 ( .A(q[6]), .B(DB[699]), .Z(n28986) );
  IV U33300 ( .A(n28985), .Z(n33827) );
  XNOR U33301 ( .A(n28983), .B(n33828), .Z(n28985) );
  XNOR U33302 ( .A(q[5]), .B(DB[698]), .Z(n33828) );
  XNOR U33303 ( .A(q[4]), .B(DB[697]), .Z(n28983) );
  IV U33304 ( .A(n28997), .Z(n33826) );
  XOR U33305 ( .A(n33829), .B(n33830), .Z(n28997) );
  XNOR U33306 ( .A(n28993), .B(n28995), .Z(n33830) );
  XNOR U33307 ( .A(q[0]), .B(DB[693]), .Z(n28995) );
  XNOR U33308 ( .A(q[3]), .B(DB[696]), .Z(n28993) );
  IV U33309 ( .A(n28992), .Z(n33829) );
  XNOR U33310 ( .A(n28990), .B(n33831), .Z(n28992) );
  XNOR U33311 ( .A(q[2]), .B(DB[695]), .Z(n33831) );
  XNOR U33312 ( .A(q[1]), .B(DB[694]), .Z(n28990) );
  XOR U33313 ( .A(n33832), .B(n28955), .Z(n28918) );
  XOR U33314 ( .A(n33833), .B(n28943), .Z(n28955) );
  XNOR U33315 ( .A(q[6]), .B(DB[706]), .Z(n28943) );
  IV U33316 ( .A(n28942), .Z(n33833) );
  XNOR U33317 ( .A(n28940), .B(n33834), .Z(n28942) );
  XNOR U33318 ( .A(q[5]), .B(DB[705]), .Z(n33834) );
  XNOR U33319 ( .A(q[4]), .B(DB[704]), .Z(n28940) );
  IV U33320 ( .A(n28954), .Z(n33832) );
  XOR U33321 ( .A(n33835), .B(n33836), .Z(n28954) );
  XNOR U33322 ( .A(n28950), .B(n28952), .Z(n33836) );
  XNOR U33323 ( .A(q[0]), .B(DB[700]), .Z(n28952) );
  XNOR U33324 ( .A(q[3]), .B(DB[703]), .Z(n28950) );
  IV U33325 ( .A(n28949), .Z(n33835) );
  XNOR U33326 ( .A(n28947), .B(n33837), .Z(n28949) );
  XNOR U33327 ( .A(q[2]), .B(DB[702]), .Z(n33837) );
  XNOR U33328 ( .A(q[1]), .B(DB[701]), .Z(n28947) );
  XOR U33329 ( .A(n33838), .B(n28912), .Z(n28875) );
  XOR U33330 ( .A(n33839), .B(n28900), .Z(n28912) );
  XNOR U33331 ( .A(q[6]), .B(DB[713]), .Z(n28900) );
  IV U33332 ( .A(n28899), .Z(n33839) );
  XNOR U33333 ( .A(n28897), .B(n33840), .Z(n28899) );
  XNOR U33334 ( .A(q[5]), .B(DB[712]), .Z(n33840) );
  XNOR U33335 ( .A(q[4]), .B(DB[711]), .Z(n28897) );
  IV U33336 ( .A(n28911), .Z(n33838) );
  XOR U33337 ( .A(n33841), .B(n33842), .Z(n28911) );
  XNOR U33338 ( .A(n28907), .B(n28909), .Z(n33842) );
  XNOR U33339 ( .A(q[0]), .B(DB[707]), .Z(n28909) );
  XNOR U33340 ( .A(q[3]), .B(DB[710]), .Z(n28907) );
  IV U33341 ( .A(n28906), .Z(n33841) );
  XNOR U33342 ( .A(n28904), .B(n33843), .Z(n28906) );
  XNOR U33343 ( .A(q[2]), .B(DB[709]), .Z(n33843) );
  XNOR U33344 ( .A(q[1]), .B(DB[708]), .Z(n28904) );
  XOR U33345 ( .A(n33844), .B(n28869), .Z(n28832) );
  XOR U33346 ( .A(n33845), .B(n28857), .Z(n28869) );
  XNOR U33347 ( .A(q[6]), .B(DB[720]), .Z(n28857) );
  IV U33348 ( .A(n28856), .Z(n33845) );
  XNOR U33349 ( .A(n28854), .B(n33846), .Z(n28856) );
  XNOR U33350 ( .A(q[5]), .B(DB[719]), .Z(n33846) );
  XNOR U33351 ( .A(q[4]), .B(DB[718]), .Z(n28854) );
  IV U33352 ( .A(n28868), .Z(n33844) );
  XOR U33353 ( .A(n33847), .B(n33848), .Z(n28868) );
  XNOR U33354 ( .A(n28864), .B(n28866), .Z(n33848) );
  XNOR U33355 ( .A(q[0]), .B(DB[714]), .Z(n28866) );
  XNOR U33356 ( .A(q[3]), .B(DB[717]), .Z(n28864) );
  IV U33357 ( .A(n28863), .Z(n33847) );
  XNOR U33358 ( .A(n28861), .B(n33849), .Z(n28863) );
  XNOR U33359 ( .A(q[2]), .B(DB[716]), .Z(n33849) );
  XNOR U33360 ( .A(q[1]), .B(DB[715]), .Z(n28861) );
  XOR U33361 ( .A(n33850), .B(n28826), .Z(n28789) );
  XOR U33362 ( .A(n33851), .B(n28814), .Z(n28826) );
  XNOR U33363 ( .A(q[6]), .B(DB[727]), .Z(n28814) );
  IV U33364 ( .A(n28813), .Z(n33851) );
  XNOR U33365 ( .A(n28811), .B(n33852), .Z(n28813) );
  XNOR U33366 ( .A(q[5]), .B(DB[726]), .Z(n33852) );
  XNOR U33367 ( .A(q[4]), .B(DB[725]), .Z(n28811) );
  IV U33368 ( .A(n28825), .Z(n33850) );
  XOR U33369 ( .A(n33853), .B(n33854), .Z(n28825) );
  XNOR U33370 ( .A(n28821), .B(n28823), .Z(n33854) );
  XNOR U33371 ( .A(q[0]), .B(DB[721]), .Z(n28823) );
  XNOR U33372 ( .A(q[3]), .B(DB[724]), .Z(n28821) );
  IV U33373 ( .A(n28820), .Z(n33853) );
  XNOR U33374 ( .A(n28818), .B(n33855), .Z(n28820) );
  XNOR U33375 ( .A(q[2]), .B(DB[723]), .Z(n33855) );
  XNOR U33376 ( .A(q[1]), .B(DB[722]), .Z(n28818) );
  XOR U33377 ( .A(n33856), .B(n28783), .Z(n28746) );
  XOR U33378 ( .A(n33857), .B(n28771), .Z(n28783) );
  XNOR U33379 ( .A(q[6]), .B(DB[734]), .Z(n28771) );
  IV U33380 ( .A(n28770), .Z(n33857) );
  XNOR U33381 ( .A(n28768), .B(n33858), .Z(n28770) );
  XNOR U33382 ( .A(q[5]), .B(DB[733]), .Z(n33858) );
  XNOR U33383 ( .A(q[4]), .B(DB[732]), .Z(n28768) );
  IV U33384 ( .A(n28782), .Z(n33856) );
  XOR U33385 ( .A(n33859), .B(n33860), .Z(n28782) );
  XNOR U33386 ( .A(n28778), .B(n28780), .Z(n33860) );
  XNOR U33387 ( .A(q[0]), .B(DB[728]), .Z(n28780) );
  XNOR U33388 ( .A(q[3]), .B(DB[731]), .Z(n28778) );
  IV U33389 ( .A(n28777), .Z(n33859) );
  XNOR U33390 ( .A(n28775), .B(n33861), .Z(n28777) );
  XNOR U33391 ( .A(q[2]), .B(DB[730]), .Z(n33861) );
  XNOR U33392 ( .A(q[1]), .B(DB[729]), .Z(n28775) );
  XOR U33393 ( .A(n33862), .B(n28740), .Z(n28703) );
  XOR U33394 ( .A(n33863), .B(n28728), .Z(n28740) );
  XNOR U33395 ( .A(q[6]), .B(DB[741]), .Z(n28728) );
  IV U33396 ( .A(n28727), .Z(n33863) );
  XNOR U33397 ( .A(n28725), .B(n33864), .Z(n28727) );
  XNOR U33398 ( .A(q[5]), .B(DB[740]), .Z(n33864) );
  XNOR U33399 ( .A(q[4]), .B(DB[739]), .Z(n28725) );
  IV U33400 ( .A(n28739), .Z(n33862) );
  XOR U33401 ( .A(n33865), .B(n33866), .Z(n28739) );
  XNOR U33402 ( .A(n28735), .B(n28737), .Z(n33866) );
  XNOR U33403 ( .A(q[0]), .B(DB[735]), .Z(n28737) );
  XNOR U33404 ( .A(q[3]), .B(DB[738]), .Z(n28735) );
  IV U33405 ( .A(n28734), .Z(n33865) );
  XNOR U33406 ( .A(n28732), .B(n33867), .Z(n28734) );
  XNOR U33407 ( .A(q[2]), .B(DB[737]), .Z(n33867) );
  XNOR U33408 ( .A(q[1]), .B(DB[736]), .Z(n28732) );
  XOR U33409 ( .A(n33868), .B(n28697), .Z(n28660) );
  XOR U33410 ( .A(n33869), .B(n28685), .Z(n28697) );
  XNOR U33411 ( .A(q[6]), .B(DB[748]), .Z(n28685) );
  IV U33412 ( .A(n28684), .Z(n33869) );
  XNOR U33413 ( .A(n28682), .B(n33870), .Z(n28684) );
  XNOR U33414 ( .A(q[5]), .B(DB[747]), .Z(n33870) );
  XNOR U33415 ( .A(q[4]), .B(DB[746]), .Z(n28682) );
  IV U33416 ( .A(n28696), .Z(n33868) );
  XOR U33417 ( .A(n33871), .B(n33872), .Z(n28696) );
  XNOR U33418 ( .A(n28692), .B(n28694), .Z(n33872) );
  XNOR U33419 ( .A(q[0]), .B(DB[742]), .Z(n28694) );
  XNOR U33420 ( .A(q[3]), .B(DB[745]), .Z(n28692) );
  IV U33421 ( .A(n28691), .Z(n33871) );
  XNOR U33422 ( .A(n28689), .B(n33873), .Z(n28691) );
  XNOR U33423 ( .A(q[2]), .B(DB[744]), .Z(n33873) );
  XNOR U33424 ( .A(q[1]), .B(DB[743]), .Z(n28689) );
  XOR U33425 ( .A(n33874), .B(n28654), .Z(n28617) );
  XOR U33426 ( .A(n33875), .B(n28642), .Z(n28654) );
  XNOR U33427 ( .A(q[6]), .B(DB[755]), .Z(n28642) );
  IV U33428 ( .A(n28641), .Z(n33875) );
  XNOR U33429 ( .A(n28639), .B(n33876), .Z(n28641) );
  XNOR U33430 ( .A(q[5]), .B(DB[754]), .Z(n33876) );
  XNOR U33431 ( .A(q[4]), .B(DB[753]), .Z(n28639) );
  IV U33432 ( .A(n28653), .Z(n33874) );
  XOR U33433 ( .A(n33877), .B(n33878), .Z(n28653) );
  XNOR U33434 ( .A(n28649), .B(n28651), .Z(n33878) );
  XNOR U33435 ( .A(q[0]), .B(DB[749]), .Z(n28651) );
  XNOR U33436 ( .A(q[3]), .B(DB[752]), .Z(n28649) );
  IV U33437 ( .A(n28648), .Z(n33877) );
  XNOR U33438 ( .A(n28646), .B(n33879), .Z(n28648) );
  XNOR U33439 ( .A(q[2]), .B(DB[751]), .Z(n33879) );
  XNOR U33440 ( .A(q[1]), .B(DB[750]), .Z(n28646) );
  XOR U33441 ( .A(n33880), .B(n28611), .Z(n28574) );
  XOR U33442 ( .A(n33881), .B(n28599), .Z(n28611) );
  XNOR U33443 ( .A(q[6]), .B(DB[762]), .Z(n28599) );
  IV U33444 ( .A(n28598), .Z(n33881) );
  XNOR U33445 ( .A(n28596), .B(n33882), .Z(n28598) );
  XNOR U33446 ( .A(q[5]), .B(DB[761]), .Z(n33882) );
  XNOR U33447 ( .A(q[4]), .B(DB[760]), .Z(n28596) );
  IV U33448 ( .A(n28610), .Z(n33880) );
  XOR U33449 ( .A(n33883), .B(n33884), .Z(n28610) );
  XNOR U33450 ( .A(n28606), .B(n28608), .Z(n33884) );
  XNOR U33451 ( .A(q[0]), .B(DB[756]), .Z(n28608) );
  XNOR U33452 ( .A(q[3]), .B(DB[759]), .Z(n28606) );
  IV U33453 ( .A(n28605), .Z(n33883) );
  XNOR U33454 ( .A(n28603), .B(n33885), .Z(n28605) );
  XNOR U33455 ( .A(q[2]), .B(DB[758]), .Z(n33885) );
  XNOR U33456 ( .A(q[1]), .B(DB[757]), .Z(n28603) );
  XOR U33457 ( .A(n33886), .B(n28568), .Z(n28531) );
  XOR U33458 ( .A(n33887), .B(n28556), .Z(n28568) );
  XNOR U33459 ( .A(q[6]), .B(DB[769]), .Z(n28556) );
  IV U33460 ( .A(n28555), .Z(n33887) );
  XNOR U33461 ( .A(n28553), .B(n33888), .Z(n28555) );
  XNOR U33462 ( .A(q[5]), .B(DB[768]), .Z(n33888) );
  XNOR U33463 ( .A(q[4]), .B(DB[767]), .Z(n28553) );
  IV U33464 ( .A(n28567), .Z(n33886) );
  XOR U33465 ( .A(n33889), .B(n33890), .Z(n28567) );
  XNOR U33466 ( .A(n28563), .B(n28565), .Z(n33890) );
  XNOR U33467 ( .A(q[0]), .B(DB[763]), .Z(n28565) );
  XNOR U33468 ( .A(q[3]), .B(DB[766]), .Z(n28563) );
  IV U33469 ( .A(n28562), .Z(n33889) );
  XNOR U33470 ( .A(n28560), .B(n33891), .Z(n28562) );
  XNOR U33471 ( .A(q[2]), .B(DB[765]), .Z(n33891) );
  XNOR U33472 ( .A(q[1]), .B(DB[764]), .Z(n28560) );
  XOR U33473 ( .A(n33892), .B(n28525), .Z(n28488) );
  XOR U33474 ( .A(n33893), .B(n28513), .Z(n28525) );
  XNOR U33475 ( .A(q[6]), .B(DB[776]), .Z(n28513) );
  IV U33476 ( .A(n28512), .Z(n33893) );
  XNOR U33477 ( .A(n28510), .B(n33894), .Z(n28512) );
  XNOR U33478 ( .A(q[5]), .B(DB[775]), .Z(n33894) );
  XNOR U33479 ( .A(q[4]), .B(DB[774]), .Z(n28510) );
  IV U33480 ( .A(n28524), .Z(n33892) );
  XOR U33481 ( .A(n33895), .B(n33896), .Z(n28524) );
  XNOR U33482 ( .A(n28520), .B(n28522), .Z(n33896) );
  XNOR U33483 ( .A(q[0]), .B(DB[770]), .Z(n28522) );
  XNOR U33484 ( .A(q[3]), .B(DB[773]), .Z(n28520) );
  IV U33485 ( .A(n28519), .Z(n33895) );
  XNOR U33486 ( .A(n28517), .B(n33897), .Z(n28519) );
  XNOR U33487 ( .A(q[2]), .B(DB[772]), .Z(n33897) );
  XNOR U33488 ( .A(q[1]), .B(DB[771]), .Z(n28517) );
  XOR U33489 ( .A(n33898), .B(n28482), .Z(n28445) );
  XOR U33490 ( .A(n33899), .B(n28470), .Z(n28482) );
  XNOR U33491 ( .A(q[6]), .B(DB[783]), .Z(n28470) );
  IV U33492 ( .A(n28469), .Z(n33899) );
  XNOR U33493 ( .A(n28467), .B(n33900), .Z(n28469) );
  XNOR U33494 ( .A(q[5]), .B(DB[782]), .Z(n33900) );
  XNOR U33495 ( .A(q[4]), .B(DB[781]), .Z(n28467) );
  IV U33496 ( .A(n28481), .Z(n33898) );
  XOR U33497 ( .A(n33901), .B(n33902), .Z(n28481) );
  XNOR U33498 ( .A(n28477), .B(n28479), .Z(n33902) );
  XNOR U33499 ( .A(q[0]), .B(DB[777]), .Z(n28479) );
  XNOR U33500 ( .A(q[3]), .B(DB[780]), .Z(n28477) );
  IV U33501 ( .A(n28476), .Z(n33901) );
  XNOR U33502 ( .A(n28474), .B(n33903), .Z(n28476) );
  XNOR U33503 ( .A(q[2]), .B(DB[779]), .Z(n33903) );
  XNOR U33504 ( .A(q[1]), .B(DB[778]), .Z(n28474) );
  XOR U33505 ( .A(n33904), .B(n28439), .Z(n28402) );
  XOR U33506 ( .A(n33905), .B(n28427), .Z(n28439) );
  XNOR U33507 ( .A(q[6]), .B(DB[790]), .Z(n28427) );
  IV U33508 ( .A(n28426), .Z(n33905) );
  XNOR U33509 ( .A(n28424), .B(n33906), .Z(n28426) );
  XNOR U33510 ( .A(q[5]), .B(DB[789]), .Z(n33906) );
  XNOR U33511 ( .A(q[4]), .B(DB[788]), .Z(n28424) );
  IV U33512 ( .A(n28438), .Z(n33904) );
  XOR U33513 ( .A(n33907), .B(n33908), .Z(n28438) );
  XNOR U33514 ( .A(n28434), .B(n28436), .Z(n33908) );
  XNOR U33515 ( .A(q[0]), .B(DB[784]), .Z(n28436) );
  XNOR U33516 ( .A(q[3]), .B(DB[787]), .Z(n28434) );
  IV U33517 ( .A(n28433), .Z(n33907) );
  XNOR U33518 ( .A(n28431), .B(n33909), .Z(n28433) );
  XNOR U33519 ( .A(q[2]), .B(DB[786]), .Z(n33909) );
  XNOR U33520 ( .A(q[1]), .B(DB[785]), .Z(n28431) );
  XOR U33521 ( .A(n33910), .B(n28396), .Z(n28359) );
  XOR U33522 ( .A(n33911), .B(n28384), .Z(n28396) );
  XNOR U33523 ( .A(q[6]), .B(DB[797]), .Z(n28384) );
  IV U33524 ( .A(n28383), .Z(n33911) );
  XNOR U33525 ( .A(n28381), .B(n33912), .Z(n28383) );
  XNOR U33526 ( .A(q[5]), .B(DB[796]), .Z(n33912) );
  XNOR U33527 ( .A(q[4]), .B(DB[795]), .Z(n28381) );
  IV U33528 ( .A(n28395), .Z(n33910) );
  XOR U33529 ( .A(n33913), .B(n33914), .Z(n28395) );
  XNOR U33530 ( .A(n28391), .B(n28393), .Z(n33914) );
  XNOR U33531 ( .A(q[0]), .B(DB[791]), .Z(n28393) );
  XNOR U33532 ( .A(q[3]), .B(DB[794]), .Z(n28391) );
  IV U33533 ( .A(n28390), .Z(n33913) );
  XNOR U33534 ( .A(n28388), .B(n33915), .Z(n28390) );
  XNOR U33535 ( .A(q[2]), .B(DB[793]), .Z(n33915) );
  XNOR U33536 ( .A(q[1]), .B(DB[792]), .Z(n28388) );
  XOR U33537 ( .A(n33916), .B(n28353), .Z(n28316) );
  XOR U33538 ( .A(n33917), .B(n28341), .Z(n28353) );
  XNOR U33539 ( .A(q[6]), .B(DB[804]), .Z(n28341) );
  IV U33540 ( .A(n28340), .Z(n33917) );
  XNOR U33541 ( .A(n28338), .B(n33918), .Z(n28340) );
  XNOR U33542 ( .A(q[5]), .B(DB[803]), .Z(n33918) );
  XNOR U33543 ( .A(q[4]), .B(DB[802]), .Z(n28338) );
  IV U33544 ( .A(n28352), .Z(n33916) );
  XOR U33545 ( .A(n33919), .B(n33920), .Z(n28352) );
  XNOR U33546 ( .A(n28348), .B(n28350), .Z(n33920) );
  XNOR U33547 ( .A(q[0]), .B(DB[798]), .Z(n28350) );
  XNOR U33548 ( .A(q[3]), .B(DB[801]), .Z(n28348) );
  IV U33549 ( .A(n28347), .Z(n33919) );
  XNOR U33550 ( .A(n28345), .B(n33921), .Z(n28347) );
  XNOR U33551 ( .A(q[2]), .B(DB[800]), .Z(n33921) );
  XNOR U33552 ( .A(q[1]), .B(DB[799]), .Z(n28345) );
  XOR U33553 ( .A(n33922), .B(n28310), .Z(n28273) );
  XOR U33554 ( .A(n33923), .B(n28298), .Z(n28310) );
  XNOR U33555 ( .A(q[6]), .B(DB[811]), .Z(n28298) );
  IV U33556 ( .A(n28297), .Z(n33923) );
  XNOR U33557 ( .A(n28295), .B(n33924), .Z(n28297) );
  XNOR U33558 ( .A(q[5]), .B(DB[810]), .Z(n33924) );
  XNOR U33559 ( .A(q[4]), .B(DB[809]), .Z(n28295) );
  IV U33560 ( .A(n28309), .Z(n33922) );
  XOR U33561 ( .A(n33925), .B(n33926), .Z(n28309) );
  XNOR U33562 ( .A(n28305), .B(n28307), .Z(n33926) );
  XNOR U33563 ( .A(q[0]), .B(DB[805]), .Z(n28307) );
  XNOR U33564 ( .A(q[3]), .B(DB[808]), .Z(n28305) );
  IV U33565 ( .A(n28304), .Z(n33925) );
  XNOR U33566 ( .A(n28302), .B(n33927), .Z(n28304) );
  XNOR U33567 ( .A(q[2]), .B(DB[807]), .Z(n33927) );
  XNOR U33568 ( .A(q[1]), .B(DB[806]), .Z(n28302) );
  XOR U33569 ( .A(n33928), .B(n28267), .Z(n28230) );
  XOR U33570 ( .A(n33929), .B(n28255), .Z(n28267) );
  XNOR U33571 ( .A(q[6]), .B(DB[818]), .Z(n28255) );
  IV U33572 ( .A(n28254), .Z(n33929) );
  XNOR U33573 ( .A(n28252), .B(n33930), .Z(n28254) );
  XNOR U33574 ( .A(q[5]), .B(DB[817]), .Z(n33930) );
  XNOR U33575 ( .A(q[4]), .B(DB[816]), .Z(n28252) );
  IV U33576 ( .A(n28266), .Z(n33928) );
  XOR U33577 ( .A(n33931), .B(n33932), .Z(n28266) );
  XNOR U33578 ( .A(n28262), .B(n28264), .Z(n33932) );
  XNOR U33579 ( .A(q[0]), .B(DB[812]), .Z(n28264) );
  XNOR U33580 ( .A(q[3]), .B(DB[815]), .Z(n28262) );
  IV U33581 ( .A(n28261), .Z(n33931) );
  XNOR U33582 ( .A(n28259), .B(n33933), .Z(n28261) );
  XNOR U33583 ( .A(q[2]), .B(DB[814]), .Z(n33933) );
  XNOR U33584 ( .A(q[1]), .B(DB[813]), .Z(n28259) );
  XOR U33585 ( .A(n33934), .B(n28224), .Z(n28187) );
  XOR U33586 ( .A(n33935), .B(n28212), .Z(n28224) );
  XNOR U33587 ( .A(q[6]), .B(DB[825]), .Z(n28212) );
  IV U33588 ( .A(n28211), .Z(n33935) );
  XNOR U33589 ( .A(n28209), .B(n33936), .Z(n28211) );
  XNOR U33590 ( .A(q[5]), .B(DB[824]), .Z(n33936) );
  XNOR U33591 ( .A(q[4]), .B(DB[823]), .Z(n28209) );
  IV U33592 ( .A(n28223), .Z(n33934) );
  XOR U33593 ( .A(n33937), .B(n33938), .Z(n28223) );
  XNOR U33594 ( .A(n28219), .B(n28221), .Z(n33938) );
  XNOR U33595 ( .A(q[0]), .B(DB[819]), .Z(n28221) );
  XNOR U33596 ( .A(q[3]), .B(DB[822]), .Z(n28219) );
  IV U33597 ( .A(n28218), .Z(n33937) );
  XNOR U33598 ( .A(n28216), .B(n33939), .Z(n28218) );
  XNOR U33599 ( .A(q[2]), .B(DB[821]), .Z(n33939) );
  XNOR U33600 ( .A(q[1]), .B(DB[820]), .Z(n28216) );
  XOR U33601 ( .A(n33940), .B(n28181), .Z(n28144) );
  XOR U33602 ( .A(n33941), .B(n28169), .Z(n28181) );
  XNOR U33603 ( .A(q[6]), .B(DB[832]), .Z(n28169) );
  IV U33604 ( .A(n28168), .Z(n33941) );
  XNOR U33605 ( .A(n28166), .B(n33942), .Z(n28168) );
  XNOR U33606 ( .A(q[5]), .B(DB[831]), .Z(n33942) );
  XNOR U33607 ( .A(q[4]), .B(DB[830]), .Z(n28166) );
  IV U33608 ( .A(n28180), .Z(n33940) );
  XOR U33609 ( .A(n33943), .B(n33944), .Z(n28180) );
  XNOR U33610 ( .A(n28176), .B(n28178), .Z(n33944) );
  XNOR U33611 ( .A(q[0]), .B(DB[826]), .Z(n28178) );
  XNOR U33612 ( .A(q[3]), .B(DB[829]), .Z(n28176) );
  IV U33613 ( .A(n28175), .Z(n33943) );
  XNOR U33614 ( .A(n28173), .B(n33945), .Z(n28175) );
  XNOR U33615 ( .A(q[2]), .B(DB[828]), .Z(n33945) );
  XNOR U33616 ( .A(q[1]), .B(DB[827]), .Z(n28173) );
  XOR U33617 ( .A(n33946), .B(n28138), .Z(n28101) );
  XOR U33618 ( .A(n33947), .B(n28126), .Z(n28138) );
  XNOR U33619 ( .A(q[6]), .B(DB[839]), .Z(n28126) );
  IV U33620 ( .A(n28125), .Z(n33947) );
  XNOR U33621 ( .A(n28123), .B(n33948), .Z(n28125) );
  XNOR U33622 ( .A(q[5]), .B(DB[838]), .Z(n33948) );
  XNOR U33623 ( .A(q[4]), .B(DB[837]), .Z(n28123) );
  IV U33624 ( .A(n28137), .Z(n33946) );
  XOR U33625 ( .A(n33949), .B(n33950), .Z(n28137) );
  XNOR U33626 ( .A(n28133), .B(n28135), .Z(n33950) );
  XNOR U33627 ( .A(q[0]), .B(DB[833]), .Z(n28135) );
  XNOR U33628 ( .A(q[3]), .B(DB[836]), .Z(n28133) );
  IV U33629 ( .A(n28132), .Z(n33949) );
  XNOR U33630 ( .A(n28130), .B(n33951), .Z(n28132) );
  XNOR U33631 ( .A(q[2]), .B(DB[835]), .Z(n33951) );
  XNOR U33632 ( .A(q[1]), .B(DB[834]), .Z(n28130) );
  XOR U33633 ( .A(n33952), .B(n28095), .Z(n28058) );
  XOR U33634 ( .A(n33953), .B(n28083), .Z(n28095) );
  XNOR U33635 ( .A(q[6]), .B(DB[846]), .Z(n28083) );
  IV U33636 ( .A(n28082), .Z(n33953) );
  XNOR U33637 ( .A(n28080), .B(n33954), .Z(n28082) );
  XNOR U33638 ( .A(q[5]), .B(DB[845]), .Z(n33954) );
  XNOR U33639 ( .A(q[4]), .B(DB[844]), .Z(n28080) );
  IV U33640 ( .A(n28094), .Z(n33952) );
  XOR U33641 ( .A(n33955), .B(n33956), .Z(n28094) );
  XNOR U33642 ( .A(n28090), .B(n28092), .Z(n33956) );
  XNOR U33643 ( .A(q[0]), .B(DB[840]), .Z(n28092) );
  XNOR U33644 ( .A(q[3]), .B(DB[843]), .Z(n28090) );
  IV U33645 ( .A(n28089), .Z(n33955) );
  XNOR U33646 ( .A(n28087), .B(n33957), .Z(n28089) );
  XNOR U33647 ( .A(q[2]), .B(DB[842]), .Z(n33957) );
  XNOR U33648 ( .A(q[1]), .B(DB[841]), .Z(n28087) );
  XOR U33649 ( .A(n33958), .B(n28052), .Z(n28015) );
  XOR U33650 ( .A(n33959), .B(n28040), .Z(n28052) );
  XNOR U33651 ( .A(q[6]), .B(DB[853]), .Z(n28040) );
  IV U33652 ( .A(n28039), .Z(n33959) );
  XNOR U33653 ( .A(n28037), .B(n33960), .Z(n28039) );
  XNOR U33654 ( .A(q[5]), .B(DB[852]), .Z(n33960) );
  XNOR U33655 ( .A(q[4]), .B(DB[851]), .Z(n28037) );
  IV U33656 ( .A(n28051), .Z(n33958) );
  XOR U33657 ( .A(n33961), .B(n33962), .Z(n28051) );
  XNOR U33658 ( .A(n28047), .B(n28049), .Z(n33962) );
  XNOR U33659 ( .A(q[0]), .B(DB[847]), .Z(n28049) );
  XNOR U33660 ( .A(q[3]), .B(DB[850]), .Z(n28047) );
  IV U33661 ( .A(n28046), .Z(n33961) );
  XNOR U33662 ( .A(n28044), .B(n33963), .Z(n28046) );
  XNOR U33663 ( .A(q[2]), .B(DB[849]), .Z(n33963) );
  XNOR U33664 ( .A(q[1]), .B(DB[848]), .Z(n28044) );
  XOR U33665 ( .A(n33964), .B(n28009), .Z(n27972) );
  XOR U33666 ( .A(n33965), .B(n27997), .Z(n28009) );
  XNOR U33667 ( .A(q[6]), .B(DB[860]), .Z(n27997) );
  IV U33668 ( .A(n27996), .Z(n33965) );
  XNOR U33669 ( .A(n27994), .B(n33966), .Z(n27996) );
  XNOR U33670 ( .A(q[5]), .B(DB[859]), .Z(n33966) );
  XNOR U33671 ( .A(q[4]), .B(DB[858]), .Z(n27994) );
  IV U33672 ( .A(n28008), .Z(n33964) );
  XOR U33673 ( .A(n33967), .B(n33968), .Z(n28008) );
  XNOR U33674 ( .A(n28004), .B(n28006), .Z(n33968) );
  XNOR U33675 ( .A(q[0]), .B(DB[854]), .Z(n28006) );
  XNOR U33676 ( .A(q[3]), .B(DB[857]), .Z(n28004) );
  IV U33677 ( .A(n28003), .Z(n33967) );
  XNOR U33678 ( .A(n28001), .B(n33969), .Z(n28003) );
  XNOR U33679 ( .A(q[2]), .B(DB[856]), .Z(n33969) );
  XNOR U33680 ( .A(q[1]), .B(DB[855]), .Z(n28001) );
  XOR U33681 ( .A(n33970), .B(n27966), .Z(n27929) );
  XOR U33682 ( .A(n33971), .B(n27954), .Z(n27966) );
  XNOR U33683 ( .A(q[6]), .B(DB[867]), .Z(n27954) );
  IV U33684 ( .A(n27953), .Z(n33971) );
  XNOR U33685 ( .A(n27951), .B(n33972), .Z(n27953) );
  XNOR U33686 ( .A(q[5]), .B(DB[866]), .Z(n33972) );
  XNOR U33687 ( .A(q[4]), .B(DB[865]), .Z(n27951) );
  IV U33688 ( .A(n27965), .Z(n33970) );
  XOR U33689 ( .A(n33973), .B(n33974), .Z(n27965) );
  XNOR U33690 ( .A(n27961), .B(n27963), .Z(n33974) );
  XNOR U33691 ( .A(q[0]), .B(DB[861]), .Z(n27963) );
  XNOR U33692 ( .A(q[3]), .B(DB[864]), .Z(n27961) );
  IV U33693 ( .A(n27960), .Z(n33973) );
  XNOR U33694 ( .A(n27958), .B(n33975), .Z(n27960) );
  XNOR U33695 ( .A(q[2]), .B(DB[863]), .Z(n33975) );
  XNOR U33696 ( .A(q[1]), .B(DB[862]), .Z(n27958) );
  XOR U33697 ( .A(n33976), .B(n27923), .Z(n27886) );
  XOR U33698 ( .A(n33977), .B(n27911), .Z(n27923) );
  XNOR U33699 ( .A(q[6]), .B(DB[874]), .Z(n27911) );
  IV U33700 ( .A(n27910), .Z(n33977) );
  XNOR U33701 ( .A(n27908), .B(n33978), .Z(n27910) );
  XNOR U33702 ( .A(q[5]), .B(DB[873]), .Z(n33978) );
  XNOR U33703 ( .A(q[4]), .B(DB[872]), .Z(n27908) );
  IV U33704 ( .A(n27922), .Z(n33976) );
  XOR U33705 ( .A(n33979), .B(n33980), .Z(n27922) );
  XNOR U33706 ( .A(n27918), .B(n27920), .Z(n33980) );
  XNOR U33707 ( .A(q[0]), .B(DB[868]), .Z(n27920) );
  XNOR U33708 ( .A(q[3]), .B(DB[871]), .Z(n27918) );
  IV U33709 ( .A(n27917), .Z(n33979) );
  XNOR U33710 ( .A(n27915), .B(n33981), .Z(n27917) );
  XNOR U33711 ( .A(q[2]), .B(DB[870]), .Z(n33981) );
  XNOR U33712 ( .A(q[1]), .B(DB[869]), .Z(n27915) );
  XOR U33713 ( .A(n33982), .B(n27880), .Z(n27843) );
  XOR U33714 ( .A(n33983), .B(n27868), .Z(n27880) );
  XNOR U33715 ( .A(q[6]), .B(DB[881]), .Z(n27868) );
  IV U33716 ( .A(n27867), .Z(n33983) );
  XNOR U33717 ( .A(n27865), .B(n33984), .Z(n27867) );
  XNOR U33718 ( .A(q[5]), .B(DB[880]), .Z(n33984) );
  XNOR U33719 ( .A(q[4]), .B(DB[879]), .Z(n27865) );
  IV U33720 ( .A(n27879), .Z(n33982) );
  XOR U33721 ( .A(n33985), .B(n33986), .Z(n27879) );
  XNOR U33722 ( .A(n27875), .B(n27877), .Z(n33986) );
  XNOR U33723 ( .A(q[0]), .B(DB[875]), .Z(n27877) );
  XNOR U33724 ( .A(q[3]), .B(DB[878]), .Z(n27875) );
  IV U33725 ( .A(n27874), .Z(n33985) );
  XNOR U33726 ( .A(n27872), .B(n33987), .Z(n27874) );
  XNOR U33727 ( .A(q[2]), .B(DB[877]), .Z(n33987) );
  XNOR U33728 ( .A(q[1]), .B(DB[876]), .Z(n27872) );
  XOR U33729 ( .A(n33988), .B(n27837), .Z(n27800) );
  XOR U33730 ( .A(n33989), .B(n27825), .Z(n27837) );
  XNOR U33731 ( .A(q[6]), .B(DB[888]), .Z(n27825) );
  IV U33732 ( .A(n27824), .Z(n33989) );
  XNOR U33733 ( .A(n27822), .B(n33990), .Z(n27824) );
  XNOR U33734 ( .A(q[5]), .B(DB[887]), .Z(n33990) );
  XNOR U33735 ( .A(q[4]), .B(DB[886]), .Z(n27822) );
  IV U33736 ( .A(n27836), .Z(n33988) );
  XOR U33737 ( .A(n33991), .B(n33992), .Z(n27836) );
  XNOR U33738 ( .A(n27832), .B(n27834), .Z(n33992) );
  XNOR U33739 ( .A(q[0]), .B(DB[882]), .Z(n27834) );
  XNOR U33740 ( .A(q[3]), .B(DB[885]), .Z(n27832) );
  IV U33741 ( .A(n27831), .Z(n33991) );
  XNOR U33742 ( .A(n27829), .B(n33993), .Z(n27831) );
  XNOR U33743 ( .A(q[2]), .B(DB[884]), .Z(n33993) );
  XNOR U33744 ( .A(q[1]), .B(DB[883]), .Z(n27829) );
  XOR U33745 ( .A(n33994), .B(n27794), .Z(n27757) );
  XOR U33746 ( .A(n33995), .B(n27782), .Z(n27794) );
  XNOR U33747 ( .A(q[6]), .B(DB[895]), .Z(n27782) );
  IV U33748 ( .A(n27781), .Z(n33995) );
  XNOR U33749 ( .A(n27779), .B(n33996), .Z(n27781) );
  XNOR U33750 ( .A(q[5]), .B(DB[894]), .Z(n33996) );
  XNOR U33751 ( .A(q[4]), .B(DB[893]), .Z(n27779) );
  IV U33752 ( .A(n27793), .Z(n33994) );
  XOR U33753 ( .A(n33997), .B(n33998), .Z(n27793) );
  XNOR U33754 ( .A(n27789), .B(n27791), .Z(n33998) );
  XNOR U33755 ( .A(q[0]), .B(DB[889]), .Z(n27791) );
  XNOR U33756 ( .A(q[3]), .B(DB[892]), .Z(n27789) );
  IV U33757 ( .A(n27788), .Z(n33997) );
  XNOR U33758 ( .A(n27786), .B(n33999), .Z(n27788) );
  XNOR U33759 ( .A(q[2]), .B(DB[891]), .Z(n33999) );
  XNOR U33760 ( .A(q[1]), .B(DB[890]), .Z(n27786) );
  XOR U33761 ( .A(n34000), .B(n27751), .Z(n27714) );
  XOR U33762 ( .A(n34001), .B(n27739), .Z(n27751) );
  XNOR U33763 ( .A(q[6]), .B(DB[902]), .Z(n27739) );
  IV U33764 ( .A(n27738), .Z(n34001) );
  XNOR U33765 ( .A(n27736), .B(n34002), .Z(n27738) );
  XNOR U33766 ( .A(q[5]), .B(DB[901]), .Z(n34002) );
  XNOR U33767 ( .A(q[4]), .B(DB[900]), .Z(n27736) );
  IV U33768 ( .A(n27750), .Z(n34000) );
  XOR U33769 ( .A(n34003), .B(n34004), .Z(n27750) );
  XNOR U33770 ( .A(n27746), .B(n27748), .Z(n34004) );
  XNOR U33771 ( .A(q[0]), .B(DB[896]), .Z(n27748) );
  XNOR U33772 ( .A(q[3]), .B(DB[899]), .Z(n27746) );
  IV U33773 ( .A(n27745), .Z(n34003) );
  XNOR U33774 ( .A(n27743), .B(n34005), .Z(n27745) );
  XNOR U33775 ( .A(q[2]), .B(DB[898]), .Z(n34005) );
  XNOR U33776 ( .A(q[1]), .B(DB[897]), .Z(n27743) );
  XOR U33777 ( .A(n34006), .B(n27708), .Z(n27671) );
  XOR U33778 ( .A(n34007), .B(n27696), .Z(n27708) );
  XNOR U33779 ( .A(q[6]), .B(DB[909]), .Z(n27696) );
  IV U33780 ( .A(n27695), .Z(n34007) );
  XNOR U33781 ( .A(n27693), .B(n34008), .Z(n27695) );
  XNOR U33782 ( .A(q[5]), .B(DB[908]), .Z(n34008) );
  XNOR U33783 ( .A(q[4]), .B(DB[907]), .Z(n27693) );
  IV U33784 ( .A(n27707), .Z(n34006) );
  XOR U33785 ( .A(n34009), .B(n34010), .Z(n27707) );
  XNOR U33786 ( .A(n27703), .B(n27705), .Z(n34010) );
  XNOR U33787 ( .A(q[0]), .B(DB[903]), .Z(n27705) );
  XNOR U33788 ( .A(q[3]), .B(DB[906]), .Z(n27703) );
  IV U33789 ( .A(n27702), .Z(n34009) );
  XNOR U33790 ( .A(n27700), .B(n34011), .Z(n27702) );
  XNOR U33791 ( .A(q[2]), .B(DB[905]), .Z(n34011) );
  XNOR U33792 ( .A(q[1]), .B(DB[904]), .Z(n27700) );
  XOR U33793 ( .A(n34012), .B(n27665), .Z(n27628) );
  XOR U33794 ( .A(n34013), .B(n27653), .Z(n27665) );
  XNOR U33795 ( .A(q[6]), .B(DB[916]), .Z(n27653) );
  IV U33796 ( .A(n27652), .Z(n34013) );
  XNOR U33797 ( .A(n27650), .B(n34014), .Z(n27652) );
  XNOR U33798 ( .A(q[5]), .B(DB[915]), .Z(n34014) );
  XNOR U33799 ( .A(q[4]), .B(DB[914]), .Z(n27650) );
  IV U33800 ( .A(n27664), .Z(n34012) );
  XOR U33801 ( .A(n34015), .B(n34016), .Z(n27664) );
  XNOR U33802 ( .A(n27660), .B(n27662), .Z(n34016) );
  XNOR U33803 ( .A(q[0]), .B(DB[910]), .Z(n27662) );
  XNOR U33804 ( .A(q[3]), .B(DB[913]), .Z(n27660) );
  IV U33805 ( .A(n27659), .Z(n34015) );
  XNOR U33806 ( .A(n27657), .B(n34017), .Z(n27659) );
  XNOR U33807 ( .A(q[2]), .B(DB[912]), .Z(n34017) );
  XNOR U33808 ( .A(q[1]), .B(DB[911]), .Z(n27657) );
  XOR U33809 ( .A(n34018), .B(n27622), .Z(n27585) );
  XOR U33810 ( .A(n34019), .B(n27610), .Z(n27622) );
  XNOR U33811 ( .A(q[6]), .B(DB[923]), .Z(n27610) );
  IV U33812 ( .A(n27609), .Z(n34019) );
  XNOR U33813 ( .A(n27607), .B(n34020), .Z(n27609) );
  XNOR U33814 ( .A(q[5]), .B(DB[922]), .Z(n34020) );
  XNOR U33815 ( .A(q[4]), .B(DB[921]), .Z(n27607) );
  IV U33816 ( .A(n27621), .Z(n34018) );
  XOR U33817 ( .A(n34021), .B(n34022), .Z(n27621) );
  XNOR U33818 ( .A(n27617), .B(n27619), .Z(n34022) );
  XNOR U33819 ( .A(q[0]), .B(DB[917]), .Z(n27619) );
  XNOR U33820 ( .A(q[3]), .B(DB[920]), .Z(n27617) );
  IV U33821 ( .A(n27616), .Z(n34021) );
  XNOR U33822 ( .A(n27614), .B(n34023), .Z(n27616) );
  XNOR U33823 ( .A(q[2]), .B(DB[919]), .Z(n34023) );
  XNOR U33824 ( .A(q[1]), .B(DB[918]), .Z(n27614) );
  XOR U33825 ( .A(n34024), .B(n27579), .Z(n27542) );
  XOR U33826 ( .A(n34025), .B(n27567), .Z(n27579) );
  XNOR U33827 ( .A(q[6]), .B(DB[930]), .Z(n27567) );
  IV U33828 ( .A(n27566), .Z(n34025) );
  XNOR U33829 ( .A(n27564), .B(n34026), .Z(n27566) );
  XNOR U33830 ( .A(q[5]), .B(DB[929]), .Z(n34026) );
  XNOR U33831 ( .A(q[4]), .B(DB[928]), .Z(n27564) );
  IV U33832 ( .A(n27578), .Z(n34024) );
  XOR U33833 ( .A(n34027), .B(n34028), .Z(n27578) );
  XNOR U33834 ( .A(n27574), .B(n27576), .Z(n34028) );
  XNOR U33835 ( .A(q[0]), .B(DB[924]), .Z(n27576) );
  XNOR U33836 ( .A(q[3]), .B(DB[927]), .Z(n27574) );
  IV U33837 ( .A(n27573), .Z(n34027) );
  XNOR U33838 ( .A(n27571), .B(n34029), .Z(n27573) );
  XNOR U33839 ( .A(q[2]), .B(DB[926]), .Z(n34029) );
  XNOR U33840 ( .A(q[1]), .B(DB[925]), .Z(n27571) );
  XOR U33841 ( .A(n34030), .B(n27536), .Z(n27499) );
  XOR U33842 ( .A(n34031), .B(n27524), .Z(n27536) );
  XNOR U33843 ( .A(q[6]), .B(DB[937]), .Z(n27524) );
  IV U33844 ( .A(n27523), .Z(n34031) );
  XNOR U33845 ( .A(n27521), .B(n34032), .Z(n27523) );
  XNOR U33846 ( .A(q[5]), .B(DB[936]), .Z(n34032) );
  XNOR U33847 ( .A(q[4]), .B(DB[935]), .Z(n27521) );
  IV U33848 ( .A(n27535), .Z(n34030) );
  XOR U33849 ( .A(n34033), .B(n34034), .Z(n27535) );
  XNOR U33850 ( .A(n27531), .B(n27533), .Z(n34034) );
  XNOR U33851 ( .A(q[0]), .B(DB[931]), .Z(n27533) );
  XNOR U33852 ( .A(q[3]), .B(DB[934]), .Z(n27531) );
  IV U33853 ( .A(n27530), .Z(n34033) );
  XNOR U33854 ( .A(n27528), .B(n34035), .Z(n27530) );
  XNOR U33855 ( .A(q[2]), .B(DB[933]), .Z(n34035) );
  XNOR U33856 ( .A(q[1]), .B(DB[932]), .Z(n27528) );
  XOR U33857 ( .A(n34036), .B(n27493), .Z(n27456) );
  XOR U33858 ( .A(n34037), .B(n27481), .Z(n27493) );
  XNOR U33859 ( .A(q[6]), .B(DB[944]), .Z(n27481) );
  IV U33860 ( .A(n27480), .Z(n34037) );
  XNOR U33861 ( .A(n27478), .B(n34038), .Z(n27480) );
  XNOR U33862 ( .A(q[5]), .B(DB[943]), .Z(n34038) );
  XNOR U33863 ( .A(q[4]), .B(DB[942]), .Z(n27478) );
  IV U33864 ( .A(n27492), .Z(n34036) );
  XOR U33865 ( .A(n34039), .B(n34040), .Z(n27492) );
  XNOR U33866 ( .A(n27488), .B(n27490), .Z(n34040) );
  XNOR U33867 ( .A(q[0]), .B(DB[938]), .Z(n27490) );
  XNOR U33868 ( .A(q[3]), .B(DB[941]), .Z(n27488) );
  IV U33869 ( .A(n27487), .Z(n34039) );
  XNOR U33870 ( .A(n27485), .B(n34041), .Z(n27487) );
  XNOR U33871 ( .A(q[2]), .B(DB[940]), .Z(n34041) );
  XNOR U33872 ( .A(q[1]), .B(DB[939]), .Z(n27485) );
  XOR U33873 ( .A(n34042), .B(n27450), .Z(n27413) );
  XOR U33874 ( .A(n34043), .B(n27438), .Z(n27450) );
  XNOR U33875 ( .A(q[6]), .B(DB[951]), .Z(n27438) );
  IV U33876 ( .A(n27437), .Z(n34043) );
  XNOR U33877 ( .A(n27435), .B(n34044), .Z(n27437) );
  XNOR U33878 ( .A(q[5]), .B(DB[950]), .Z(n34044) );
  XNOR U33879 ( .A(q[4]), .B(DB[949]), .Z(n27435) );
  IV U33880 ( .A(n27449), .Z(n34042) );
  XOR U33881 ( .A(n34045), .B(n34046), .Z(n27449) );
  XNOR U33882 ( .A(n27445), .B(n27447), .Z(n34046) );
  XNOR U33883 ( .A(q[0]), .B(DB[945]), .Z(n27447) );
  XNOR U33884 ( .A(q[3]), .B(DB[948]), .Z(n27445) );
  IV U33885 ( .A(n27444), .Z(n34045) );
  XNOR U33886 ( .A(n27442), .B(n34047), .Z(n27444) );
  XNOR U33887 ( .A(q[2]), .B(DB[947]), .Z(n34047) );
  XNOR U33888 ( .A(q[1]), .B(DB[946]), .Z(n27442) );
  XOR U33889 ( .A(n34048), .B(n27407), .Z(n27370) );
  XOR U33890 ( .A(n34049), .B(n27395), .Z(n27407) );
  XNOR U33891 ( .A(q[6]), .B(DB[958]), .Z(n27395) );
  IV U33892 ( .A(n27394), .Z(n34049) );
  XNOR U33893 ( .A(n27392), .B(n34050), .Z(n27394) );
  XNOR U33894 ( .A(q[5]), .B(DB[957]), .Z(n34050) );
  XNOR U33895 ( .A(q[4]), .B(DB[956]), .Z(n27392) );
  IV U33896 ( .A(n27406), .Z(n34048) );
  XOR U33897 ( .A(n34051), .B(n34052), .Z(n27406) );
  XNOR U33898 ( .A(n27402), .B(n27404), .Z(n34052) );
  XNOR U33899 ( .A(q[0]), .B(DB[952]), .Z(n27404) );
  XNOR U33900 ( .A(q[3]), .B(DB[955]), .Z(n27402) );
  IV U33901 ( .A(n27401), .Z(n34051) );
  XNOR U33902 ( .A(n27399), .B(n34053), .Z(n27401) );
  XNOR U33903 ( .A(q[2]), .B(DB[954]), .Z(n34053) );
  XNOR U33904 ( .A(q[1]), .B(DB[953]), .Z(n27399) );
  XOR U33905 ( .A(n34054), .B(n27364), .Z(n27327) );
  XOR U33906 ( .A(n34055), .B(n27352), .Z(n27364) );
  XNOR U33907 ( .A(q[6]), .B(DB[965]), .Z(n27352) );
  IV U33908 ( .A(n27351), .Z(n34055) );
  XNOR U33909 ( .A(n27349), .B(n34056), .Z(n27351) );
  XNOR U33910 ( .A(q[5]), .B(DB[964]), .Z(n34056) );
  XNOR U33911 ( .A(q[4]), .B(DB[963]), .Z(n27349) );
  IV U33912 ( .A(n27363), .Z(n34054) );
  XOR U33913 ( .A(n34057), .B(n34058), .Z(n27363) );
  XNOR U33914 ( .A(n27359), .B(n27361), .Z(n34058) );
  XNOR U33915 ( .A(q[0]), .B(DB[959]), .Z(n27361) );
  XNOR U33916 ( .A(q[3]), .B(DB[962]), .Z(n27359) );
  IV U33917 ( .A(n27358), .Z(n34057) );
  XNOR U33918 ( .A(n27356), .B(n34059), .Z(n27358) );
  XNOR U33919 ( .A(q[2]), .B(DB[961]), .Z(n34059) );
  XNOR U33920 ( .A(q[1]), .B(DB[960]), .Z(n27356) );
  XOR U33921 ( .A(n34060), .B(n27321), .Z(n27284) );
  XOR U33922 ( .A(n34061), .B(n27309), .Z(n27321) );
  XNOR U33923 ( .A(q[6]), .B(DB[972]), .Z(n27309) );
  IV U33924 ( .A(n27308), .Z(n34061) );
  XNOR U33925 ( .A(n27306), .B(n34062), .Z(n27308) );
  XNOR U33926 ( .A(q[5]), .B(DB[971]), .Z(n34062) );
  XNOR U33927 ( .A(q[4]), .B(DB[970]), .Z(n27306) );
  IV U33928 ( .A(n27320), .Z(n34060) );
  XOR U33929 ( .A(n34063), .B(n34064), .Z(n27320) );
  XNOR U33930 ( .A(n27316), .B(n27318), .Z(n34064) );
  XNOR U33931 ( .A(q[0]), .B(DB[966]), .Z(n27318) );
  XNOR U33932 ( .A(q[3]), .B(DB[969]), .Z(n27316) );
  IV U33933 ( .A(n27315), .Z(n34063) );
  XNOR U33934 ( .A(n27313), .B(n34065), .Z(n27315) );
  XNOR U33935 ( .A(q[2]), .B(DB[968]), .Z(n34065) );
  XNOR U33936 ( .A(q[1]), .B(DB[967]), .Z(n27313) );
  XOR U33937 ( .A(n34066), .B(n27278), .Z(n27241) );
  XOR U33938 ( .A(n34067), .B(n27266), .Z(n27278) );
  XNOR U33939 ( .A(q[6]), .B(DB[979]), .Z(n27266) );
  IV U33940 ( .A(n27265), .Z(n34067) );
  XNOR U33941 ( .A(n27263), .B(n34068), .Z(n27265) );
  XNOR U33942 ( .A(q[5]), .B(DB[978]), .Z(n34068) );
  XNOR U33943 ( .A(q[4]), .B(DB[977]), .Z(n27263) );
  IV U33944 ( .A(n27277), .Z(n34066) );
  XOR U33945 ( .A(n34069), .B(n34070), .Z(n27277) );
  XNOR U33946 ( .A(n27273), .B(n27275), .Z(n34070) );
  XNOR U33947 ( .A(q[0]), .B(DB[973]), .Z(n27275) );
  XNOR U33948 ( .A(q[3]), .B(DB[976]), .Z(n27273) );
  IV U33949 ( .A(n27272), .Z(n34069) );
  XNOR U33950 ( .A(n27270), .B(n34071), .Z(n27272) );
  XNOR U33951 ( .A(q[2]), .B(DB[975]), .Z(n34071) );
  XNOR U33952 ( .A(q[1]), .B(DB[974]), .Z(n27270) );
  XOR U33953 ( .A(n34072), .B(n27235), .Z(n27198) );
  XOR U33954 ( .A(n34073), .B(n27223), .Z(n27235) );
  XNOR U33955 ( .A(q[6]), .B(DB[986]), .Z(n27223) );
  IV U33956 ( .A(n27222), .Z(n34073) );
  XNOR U33957 ( .A(n27220), .B(n34074), .Z(n27222) );
  XNOR U33958 ( .A(q[5]), .B(DB[985]), .Z(n34074) );
  XNOR U33959 ( .A(q[4]), .B(DB[984]), .Z(n27220) );
  IV U33960 ( .A(n27234), .Z(n34072) );
  XOR U33961 ( .A(n34075), .B(n34076), .Z(n27234) );
  XNOR U33962 ( .A(n27230), .B(n27232), .Z(n34076) );
  XNOR U33963 ( .A(q[0]), .B(DB[980]), .Z(n27232) );
  XNOR U33964 ( .A(q[3]), .B(DB[983]), .Z(n27230) );
  IV U33965 ( .A(n27229), .Z(n34075) );
  XNOR U33966 ( .A(n27227), .B(n34077), .Z(n27229) );
  XNOR U33967 ( .A(q[2]), .B(DB[982]), .Z(n34077) );
  XNOR U33968 ( .A(q[1]), .B(DB[981]), .Z(n27227) );
  XOR U33969 ( .A(n34078), .B(n27192), .Z(n27155) );
  XOR U33970 ( .A(n34079), .B(n27180), .Z(n27192) );
  XNOR U33971 ( .A(q[6]), .B(DB[993]), .Z(n27180) );
  IV U33972 ( .A(n27179), .Z(n34079) );
  XNOR U33973 ( .A(n27177), .B(n34080), .Z(n27179) );
  XNOR U33974 ( .A(q[5]), .B(DB[992]), .Z(n34080) );
  XNOR U33975 ( .A(q[4]), .B(DB[991]), .Z(n27177) );
  IV U33976 ( .A(n27191), .Z(n34078) );
  XOR U33977 ( .A(n34081), .B(n34082), .Z(n27191) );
  XNOR U33978 ( .A(n27187), .B(n27189), .Z(n34082) );
  XNOR U33979 ( .A(q[0]), .B(DB[987]), .Z(n27189) );
  XNOR U33980 ( .A(q[3]), .B(DB[990]), .Z(n27187) );
  IV U33981 ( .A(n27186), .Z(n34081) );
  XNOR U33982 ( .A(n27184), .B(n34083), .Z(n27186) );
  XNOR U33983 ( .A(q[2]), .B(DB[989]), .Z(n34083) );
  XNOR U33984 ( .A(q[1]), .B(DB[988]), .Z(n27184) );
  XOR U33985 ( .A(n34084), .B(n27149), .Z(n27112) );
  XOR U33986 ( .A(n34085), .B(n27137), .Z(n27149) );
  XNOR U33987 ( .A(q[6]), .B(DB[1000]), .Z(n27137) );
  IV U33988 ( .A(n27136), .Z(n34085) );
  XNOR U33989 ( .A(n27134), .B(n34086), .Z(n27136) );
  XNOR U33990 ( .A(q[5]), .B(DB[999]), .Z(n34086) );
  XNOR U33991 ( .A(q[4]), .B(DB[998]), .Z(n27134) );
  IV U33992 ( .A(n27148), .Z(n34084) );
  XOR U33993 ( .A(n34087), .B(n34088), .Z(n27148) );
  XNOR U33994 ( .A(n27144), .B(n27146), .Z(n34088) );
  XNOR U33995 ( .A(q[0]), .B(DB[994]), .Z(n27146) );
  XNOR U33996 ( .A(q[3]), .B(DB[997]), .Z(n27144) );
  IV U33997 ( .A(n27143), .Z(n34087) );
  XNOR U33998 ( .A(n27141), .B(n34089), .Z(n27143) );
  XNOR U33999 ( .A(q[2]), .B(DB[996]), .Z(n34089) );
  XNOR U34000 ( .A(q[1]), .B(DB[995]), .Z(n27141) );
  XOR U34001 ( .A(n34090), .B(n27106), .Z(n27069) );
  XOR U34002 ( .A(n34091), .B(n27094), .Z(n27106) );
  XNOR U34003 ( .A(q[6]), .B(DB[1007]), .Z(n27094) );
  IV U34004 ( .A(n27093), .Z(n34091) );
  XNOR U34005 ( .A(n27091), .B(n34092), .Z(n27093) );
  XNOR U34006 ( .A(q[5]), .B(DB[1006]), .Z(n34092) );
  XNOR U34007 ( .A(q[4]), .B(DB[1005]), .Z(n27091) );
  IV U34008 ( .A(n27105), .Z(n34090) );
  XOR U34009 ( .A(n34093), .B(n34094), .Z(n27105) );
  XNOR U34010 ( .A(n27101), .B(n27103), .Z(n34094) );
  XNOR U34011 ( .A(q[0]), .B(DB[1001]), .Z(n27103) );
  XNOR U34012 ( .A(q[3]), .B(DB[1004]), .Z(n27101) );
  IV U34013 ( .A(n27100), .Z(n34093) );
  XNOR U34014 ( .A(n27098), .B(n34095), .Z(n27100) );
  XNOR U34015 ( .A(q[2]), .B(DB[1003]), .Z(n34095) );
  XNOR U34016 ( .A(q[1]), .B(DB[1002]), .Z(n27098) );
  XOR U34017 ( .A(n34096), .B(n27063), .Z(n27026) );
  XOR U34018 ( .A(n34097), .B(n27051), .Z(n27063) );
  XNOR U34019 ( .A(q[6]), .B(DB[1014]), .Z(n27051) );
  IV U34020 ( .A(n27050), .Z(n34097) );
  XNOR U34021 ( .A(n27048), .B(n34098), .Z(n27050) );
  XNOR U34022 ( .A(q[5]), .B(DB[1013]), .Z(n34098) );
  XNOR U34023 ( .A(q[4]), .B(DB[1012]), .Z(n27048) );
  IV U34024 ( .A(n27062), .Z(n34096) );
  XOR U34025 ( .A(n34099), .B(n34100), .Z(n27062) );
  XNOR U34026 ( .A(n27058), .B(n27060), .Z(n34100) );
  XNOR U34027 ( .A(q[0]), .B(DB[1008]), .Z(n27060) );
  XNOR U34028 ( .A(q[3]), .B(DB[1011]), .Z(n27058) );
  IV U34029 ( .A(n27057), .Z(n34099) );
  XNOR U34030 ( .A(n27055), .B(n34101), .Z(n27057) );
  XNOR U34031 ( .A(q[2]), .B(DB[1010]), .Z(n34101) );
  XNOR U34032 ( .A(q[1]), .B(DB[1009]), .Z(n27055) );
  XOR U34033 ( .A(n34102), .B(n27020), .Z(n26983) );
  XOR U34034 ( .A(n34103), .B(n27008), .Z(n27020) );
  XNOR U34035 ( .A(q[6]), .B(DB[1021]), .Z(n27008) );
  IV U34036 ( .A(n27007), .Z(n34103) );
  XNOR U34037 ( .A(n27005), .B(n34104), .Z(n27007) );
  XNOR U34038 ( .A(q[5]), .B(DB[1020]), .Z(n34104) );
  XNOR U34039 ( .A(q[4]), .B(DB[1019]), .Z(n27005) );
  IV U34040 ( .A(n27019), .Z(n34102) );
  XOR U34041 ( .A(n34105), .B(n34106), .Z(n27019) );
  XNOR U34042 ( .A(n27015), .B(n27017), .Z(n34106) );
  XNOR U34043 ( .A(q[0]), .B(DB[1015]), .Z(n27017) );
  XNOR U34044 ( .A(q[3]), .B(DB[1018]), .Z(n27015) );
  IV U34045 ( .A(n27014), .Z(n34105) );
  XNOR U34046 ( .A(n27012), .B(n34107), .Z(n27014) );
  XNOR U34047 ( .A(q[2]), .B(DB[1017]), .Z(n34107) );
  XNOR U34048 ( .A(q[1]), .B(DB[1016]), .Z(n27012) );
  XOR U34049 ( .A(n34108), .B(n26977), .Z(n26940) );
  XOR U34050 ( .A(n34109), .B(n26965), .Z(n26977) );
  XNOR U34051 ( .A(q[6]), .B(DB[1028]), .Z(n26965) );
  IV U34052 ( .A(n26964), .Z(n34109) );
  XNOR U34053 ( .A(n26962), .B(n34110), .Z(n26964) );
  XNOR U34054 ( .A(q[5]), .B(DB[1027]), .Z(n34110) );
  XNOR U34055 ( .A(q[4]), .B(DB[1026]), .Z(n26962) );
  IV U34056 ( .A(n26976), .Z(n34108) );
  XOR U34057 ( .A(n34111), .B(n34112), .Z(n26976) );
  XNOR U34058 ( .A(n26972), .B(n26974), .Z(n34112) );
  XNOR U34059 ( .A(q[0]), .B(DB[1022]), .Z(n26974) );
  XNOR U34060 ( .A(q[3]), .B(DB[1025]), .Z(n26972) );
  IV U34061 ( .A(n26971), .Z(n34111) );
  XNOR U34062 ( .A(n26969), .B(n34113), .Z(n26971) );
  XNOR U34063 ( .A(q[2]), .B(DB[1024]), .Z(n34113) );
  XNOR U34064 ( .A(q[1]), .B(DB[1023]), .Z(n26969) );
  XOR U34065 ( .A(n34114), .B(n26934), .Z(n26897) );
  XOR U34066 ( .A(n34115), .B(n26922), .Z(n26934) );
  XNOR U34067 ( .A(q[6]), .B(DB[1035]), .Z(n26922) );
  IV U34068 ( .A(n26921), .Z(n34115) );
  XNOR U34069 ( .A(n26919), .B(n34116), .Z(n26921) );
  XNOR U34070 ( .A(q[5]), .B(DB[1034]), .Z(n34116) );
  XNOR U34071 ( .A(q[4]), .B(DB[1033]), .Z(n26919) );
  IV U34072 ( .A(n26933), .Z(n34114) );
  XOR U34073 ( .A(n34117), .B(n34118), .Z(n26933) );
  XNOR U34074 ( .A(n26929), .B(n26931), .Z(n34118) );
  XNOR U34075 ( .A(q[0]), .B(DB[1029]), .Z(n26931) );
  XNOR U34076 ( .A(q[3]), .B(DB[1032]), .Z(n26929) );
  IV U34077 ( .A(n26928), .Z(n34117) );
  XNOR U34078 ( .A(n26926), .B(n34119), .Z(n26928) );
  XNOR U34079 ( .A(q[2]), .B(DB[1031]), .Z(n34119) );
  XNOR U34080 ( .A(q[1]), .B(DB[1030]), .Z(n26926) );
  XOR U34081 ( .A(n34120), .B(n26891), .Z(n26854) );
  XOR U34082 ( .A(n34121), .B(n26879), .Z(n26891) );
  XNOR U34083 ( .A(q[6]), .B(DB[1042]), .Z(n26879) );
  IV U34084 ( .A(n26878), .Z(n34121) );
  XNOR U34085 ( .A(n26876), .B(n34122), .Z(n26878) );
  XNOR U34086 ( .A(q[5]), .B(DB[1041]), .Z(n34122) );
  XNOR U34087 ( .A(q[4]), .B(DB[1040]), .Z(n26876) );
  IV U34088 ( .A(n26890), .Z(n34120) );
  XOR U34089 ( .A(n34123), .B(n34124), .Z(n26890) );
  XNOR U34090 ( .A(n26886), .B(n26888), .Z(n34124) );
  XNOR U34091 ( .A(q[0]), .B(DB[1036]), .Z(n26888) );
  XNOR U34092 ( .A(q[3]), .B(DB[1039]), .Z(n26886) );
  IV U34093 ( .A(n26885), .Z(n34123) );
  XNOR U34094 ( .A(n26883), .B(n34125), .Z(n26885) );
  XNOR U34095 ( .A(q[2]), .B(DB[1038]), .Z(n34125) );
  XNOR U34096 ( .A(q[1]), .B(DB[1037]), .Z(n26883) );
  XOR U34097 ( .A(n34126), .B(n26848), .Z(n26811) );
  XOR U34098 ( .A(n34127), .B(n26836), .Z(n26848) );
  XNOR U34099 ( .A(q[6]), .B(DB[1049]), .Z(n26836) );
  IV U34100 ( .A(n26835), .Z(n34127) );
  XNOR U34101 ( .A(n26833), .B(n34128), .Z(n26835) );
  XNOR U34102 ( .A(q[5]), .B(DB[1048]), .Z(n34128) );
  XNOR U34103 ( .A(q[4]), .B(DB[1047]), .Z(n26833) );
  IV U34104 ( .A(n26847), .Z(n34126) );
  XOR U34105 ( .A(n34129), .B(n34130), .Z(n26847) );
  XNOR U34106 ( .A(n26843), .B(n26845), .Z(n34130) );
  XNOR U34107 ( .A(q[0]), .B(DB[1043]), .Z(n26845) );
  XNOR U34108 ( .A(q[3]), .B(DB[1046]), .Z(n26843) );
  IV U34109 ( .A(n26842), .Z(n34129) );
  XNOR U34110 ( .A(n26840), .B(n34131), .Z(n26842) );
  XNOR U34111 ( .A(q[2]), .B(DB[1045]), .Z(n34131) );
  XNOR U34112 ( .A(q[1]), .B(DB[1044]), .Z(n26840) );
  XOR U34113 ( .A(n34132), .B(n26805), .Z(n26768) );
  XOR U34114 ( .A(n34133), .B(n26793), .Z(n26805) );
  XNOR U34115 ( .A(q[6]), .B(DB[1056]), .Z(n26793) );
  IV U34116 ( .A(n26792), .Z(n34133) );
  XNOR U34117 ( .A(n26790), .B(n34134), .Z(n26792) );
  XNOR U34118 ( .A(q[5]), .B(DB[1055]), .Z(n34134) );
  XNOR U34119 ( .A(q[4]), .B(DB[1054]), .Z(n26790) );
  IV U34120 ( .A(n26804), .Z(n34132) );
  XOR U34121 ( .A(n34135), .B(n34136), .Z(n26804) );
  XNOR U34122 ( .A(n26800), .B(n26802), .Z(n34136) );
  XNOR U34123 ( .A(q[0]), .B(DB[1050]), .Z(n26802) );
  XNOR U34124 ( .A(q[3]), .B(DB[1053]), .Z(n26800) );
  IV U34125 ( .A(n26799), .Z(n34135) );
  XNOR U34126 ( .A(n26797), .B(n34137), .Z(n26799) );
  XNOR U34127 ( .A(q[2]), .B(DB[1052]), .Z(n34137) );
  XNOR U34128 ( .A(q[1]), .B(DB[1051]), .Z(n26797) );
  XOR U34129 ( .A(n34138), .B(n26762), .Z(n26725) );
  XOR U34130 ( .A(n34139), .B(n26750), .Z(n26762) );
  XNOR U34131 ( .A(q[6]), .B(DB[1063]), .Z(n26750) );
  IV U34132 ( .A(n26749), .Z(n34139) );
  XNOR U34133 ( .A(n26747), .B(n34140), .Z(n26749) );
  XNOR U34134 ( .A(q[5]), .B(DB[1062]), .Z(n34140) );
  XNOR U34135 ( .A(q[4]), .B(DB[1061]), .Z(n26747) );
  IV U34136 ( .A(n26761), .Z(n34138) );
  XOR U34137 ( .A(n34141), .B(n34142), .Z(n26761) );
  XNOR U34138 ( .A(n26757), .B(n26759), .Z(n34142) );
  XNOR U34139 ( .A(q[0]), .B(DB[1057]), .Z(n26759) );
  XNOR U34140 ( .A(q[3]), .B(DB[1060]), .Z(n26757) );
  IV U34141 ( .A(n26756), .Z(n34141) );
  XNOR U34142 ( .A(n26754), .B(n34143), .Z(n26756) );
  XNOR U34143 ( .A(q[2]), .B(DB[1059]), .Z(n34143) );
  XNOR U34144 ( .A(q[1]), .B(DB[1058]), .Z(n26754) );
  XOR U34145 ( .A(n34144), .B(n26719), .Z(n26682) );
  XOR U34146 ( .A(n34145), .B(n26707), .Z(n26719) );
  XNOR U34147 ( .A(q[6]), .B(DB[1070]), .Z(n26707) );
  IV U34148 ( .A(n26706), .Z(n34145) );
  XNOR U34149 ( .A(n26704), .B(n34146), .Z(n26706) );
  XNOR U34150 ( .A(q[5]), .B(DB[1069]), .Z(n34146) );
  XNOR U34151 ( .A(q[4]), .B(DB[1068]), .Z(n26704) );
  IV U34152 ( .A(n26718), .Z(n34144) );
  XOR U34153 ( .A(n34147), .B(n34148), .Z(n26718) );
  XNOR U34154 ( .A(n26714), .B(n26716), .Z(n34148) );
  XNOR U34155 ( .A(q[0]), .B(DB[1064]), .Z(n26716) );
  XNOR U34156 ( .A(q[3]), .B(DB[1067]), .Z(n26714) );
  IV U34157 ( .A(n26713), .Z(n34147) );
  XNOR U34158 ( .A(n26711), .B(n34149), .Z(n26713) );
  XNOR U34159 ( .A(q[2]), .B(DB[1066]), .Z(n34149) );
  XNOR U34160 ( .A(q[1]), .B(DB[1065]), .Z(n26711) );
  XOR U34161 ( .A(n34150), .B(n26676), .Z(n26639) );
  XOR U34162 ( .A(n34151), .B(n26664), .Z(n26676) );
  XNOR U34163 ( .A(q[6]), .B(DB[1077]), .Z(n26664) );
  IV U34164 ( .A(n26663), .Z(n34151) );
  XNOR U34165 ( .A(n26661), .B(n34152), .Z(n26663) );
  XNOR U34166 ( .A(q[5]), .B(DB[1076]), .Z(n34152) );
  XNOR U34167 ( .A(q[4]), .B(DB[1075]), .Z(n26661) );
  IV U34168 ( .A(n26675), .Z(n34150) );
  XOR U34169 ( .A(n34153), .B(n34154), .Z(n26675) );
  XNOR U34170 ( .A(n26671), .B(n26673), .Z(n34154) );
  XNOR U34171 ( .A(q[0]), .B(DB[1071]), .Z(n26673) );
  XNOR U34172 ( .A(q[3]), .B(DB[1074]), .Z(n26671) );
  IV U34173 ( .A(n26670), .Z(n34153) );
  XNOR U34174 ( .A(n26668), .B(n34155), .Z(n26670) );
  XNOR U34175 ( .A(q[2]), .B(DB[1073]), .Z(n34155) );
  XNOR U34176 ( .A(q[1]), .B(DB[1072]), .Z(n26668) );
  XOR U34177 ( .A(n34156), .B(n26633), .Z(n26596) );
  XOR U34178 ( .A(n34157), .B(n26621), .Z(n26633) );
  XNOR U34179 ( .A(q[6]), .B(DB[1084]), .Z(n26621) );
  IV U34180 ( .A(n26620), .Z(n34157) );
  XNOR U34181 ( .A(n26618), .B(n34158), .Z(n26620) );
  XNOR U34182 ( .A(q[5]), .B(DB[1083]), .Z(n34158) );
  XNOR U34183 ( .A(q[4]), .B(DB[1082]), .Z(n26618) );
  IV U34184 ( .A(n26632), .Z(n34156) );
  XOR U34185 ( .A(n34159), .B(n34160), .Z(n26632) );
  XNOR U34186 ( .A(n26628), .B(n26630), .Z(n34160) );
  XNOR U34187 ( .A(q[0]), .B(DB[1078]), .Z(n26630) );
  XNOR U34188 ( .A(q[3]), .B(DB[1081]), .Z(n26628) );
  IV U34189 ( .A(n26627), .Z(n34159) );
  XNOR U34190 ( .A(n26625), .B(n34161), .Z(n26627) );
  XNOR U34191 ( .A(q[2]), .B(DB[1080]), .Z(n34161) );
  XNOR U34192 ( .A(q[1]), .B(DB[1079]), .Z(n26625) );
  XOR U34193 ( .A(n34162), .B(n26590), .Z(n26553) );
  XOR U34194 ( .A(n34163), .B(n26578), .Z(n26590) );
  XNOR U34195 ( .A(q[6]), .B(DB[1091]), .Z(n26578) );
  IV U34196 ( .A(n26577), .Z(n34163) );
  XNOR U34197 ( .A(n26575), .B(n34164), .Z(n26577) );
  XNOR U34198 ( .A(q[5]), .B(DB[1090]), .Z(n34164) );
  XNOR U34199 ( .A(q[4]), .B(DB[1089]), .Z(n26575) );
  IV U34200 ( .A(n26589), .Z(n34162) );
  XOR U34201 ( .A(n34165), .B(n34166), .Z(n26589) );
  XNOR U34202 ( .A(n26585), .B(n26587), .Z(n34166) );
  XNOR U34203 ( .A(q[0]), .B(DB[1085]), .Z(n26587) );
  XNOR U34204 ( .A(q[3]), .B(DB[1088]), .Z(n26585) );
  IV U34205 ( .A(n26584), .Z(n34165) );
  XNOR U34206 ( .A(n26582), .B(n34167), .Z(n26584) );
  XNOR U34207 ( .A(q[2]), .B(DB[1087]), .Z(n34167) );
  XNOR U34208 ( .A(q[1]), .B(DB[1086]), .Z(n26582) );
  XOR U34209 ( .A(n34168), .B(n26547), .Z(n26510) );
  XOR U34210 ( .A(n34169), .B(n26535), .Z(n26547) );
  XNOR U34211 ( .A(q[6]), .B(DB[1098]), .Z(n26535) );
  IV U34212 ( .A(n26534), .Z(n34169) );
  XNOR U34213 ( .A(n26532), .B(n34170), .Z(n26534) );
  XNOR U34214 ( .A(q[5]), .B(DB[1097]), .Z(n34170) );
  XNOR U34215 ( .A(q[4]), .B(DB[1096]), .Z(n26532) );
  IV U34216 ( .A(n26546), .Z(n34168) );
  XOR U34217 ( .A(n34171), .B(n34172), .Z(n26546) );
  XNOR U34218 ( .A(n26542), .B(n26544), .Z(n34172) );
  XNOR U34219 ( .A(q[0]), .B(DB[1092]), .Z(n26544) );
  XNOR U34220 ( .A(q[3]), .B(DB[1095]), .Z(n26542) );
  IV U34221 ( .A(n26541), .Z(n34171) );
  XNOR U34222 ( .A(n26539), .B(n34173), .Z(n26541) );
  XNOR U34223 ( .A(q[2]), .B(DB[1094]), .Z(n34173) );
  XNOR U34224 ( .A(q[1]), .B(DB[1093]), .Z(n26539) );
  XOR U34225 ( .A(n34174), .B(n26504), .Z(n26467) );
  XOR U34226 ( .A(n34175), .B(n26492), .Z(n26504) );
  XNOR U34227 ( .A(q[6]), .B(DB[1105]), .Z(n26492) );
  IV U34228 ( .A(n26491), .Z(n34175) );
  XNOR U34229 ( .A(n26489), .B(n34176), .Z(n26491) );
  XNOR U34230 ( .A(q[5]), .B(DB[1104]), .Z(n34176) );
  XNOR U34231 ( .A(q[4]), .B(DB[1103]), .Z(n26489) );
  IV U34232 ( .A(n26503), .Z(n34174) );
  XOR U34233 ( .A(n34177), .B(n34178), .Z(n26503) );
  XNOR U34234 ( .A(n26499), .B(n26501), .Z(n34178) );
  XNOR U34235 ( .A(q[0]), .B(DB[1099]), .Z(n26501) );
  XNOR U34236 ( .A(q[3]), .B(DB[1102]), .Z(n26499) );
  IV U34237 ( .A(n26498), .Z(n34177) );
  XNOR U34238 ( .A(n26496), .B(n34179), .Z(n26498) );
  XNOR U34239 ( .A(q[2]), .B(DB[1101]), .Z(n34179) );
  XNOR U34240 ( .A(q[1]), .B(DB[1100]), .Z(n26496) );
  XOR U34241 ( .A(n34180), .B(n26461), .Z(n26424) );
  XOR U34242 ( .A(n34181), .B(n26449), .Z(n26461) );
  XNOR U34243 ( .A(q[6]), .B(DB[1112]), .Z(n26449) );
  IV U34244 ( .A(n26448), .Z(n34181) );
  XNOR U34245 ( .A(n26446), .B(n34182), .Z(n26448) );
  XNOR U34246 ( .A(q[5]), .B(DB[1111]), .Z(n34182) );
  XNOR U34247 ( .A(q[4]), .B(DB[1110]), .Z(n26446) );
  IV U34248 ( .A(n26460), .Z(n34180) );
  XOR U34249 ( .A(n34183), .B(n34184), .Z(n26460) );
  XNOR U34250 ( .A(n26456), .B(n26458), .Z(n34184) );
  XNOR U34251 ( .A(q[0]), .B(DB[1106]), .Z(n26458) );
  XNOR U34252 ( .A(q[3]), .B(DB[1109]), .Z(n26456) );
  IV U34253 ( .A(n26455), .Z(n34183) );
  XNOR U34254 ( .A(n26453), .B(n34185), .Z(n26455) );
  XNOR U34255 ( .A(q[2]), .B(DB[1108]), .Z(n34185) );
  XNOR U34256 ( .A(q[1]), .B(DB[1107]), .Z(n26453) );
  XOR U34257 ( .A(n34186), .B(n26418), .Z(n26381) );
  XOR U34258 ( .A(n34187), .B(n26406), .Z(n26418) );
  XNOR U34259 ( .A(q[6]), .B(DB[1119]), .Z(n26406) );
  IV U34260 ( .A(n26405), .Z(n34187) );
  XNOR U34261 ( .A(n26403), .B(n34188), .Z(n26405) );
  XNOR U34262 ( .A(q[5]), .B(DB[1118]), .Z(n34188) );
  XNOR U34263 ( .A(q[4]), .B(DB[1117]), .Z(n26403) );
  IV U34264 ( .A(n26417), .Z(n34186) );
  XOR U34265 ( .A(n34189), .B(n34190), .Z(n26417) );
  XNOR U34266 ( .A(n26413), .B(n26415), .Z(n34190) );
  XNOR U34267 ( .A(q[0]), .B(DB[1113]), .Z(n26415) );
  XNOR U34268 ( .A(q[3]), .B(DB[1116]), .Z(n26413) );
  IV U34269 ( .A(n26412), .Z(n34189) );
  XNOR U34270 ( .A(n26410), .B(n34191), .Z(n26412) );
  XNOR U34271 ( .A(q[2]), .B(DB[1115]), .Z(n34191) );
  XNOR U34272 ( .A(q[1]), .B(DB[1114]), .Z(n26410) );
  XOR U34273 ( .A(n34192), .B(n26375), .Z(n26338) );
  XOR U34274 ( .A(n34193), .B(n26363), .Z(n26375) );
  XNOR U34275 ( .A(q[6]), .B(DB[1126]), .Z(n26363) );
  IV U34276 ( .A(n26362), .Z(n34193) );
  XNOR U34277 ( .A(n26360), .B(n34194), .Z(n26362) );
  XNOR U34278 ( .A(q[5]), .B(DB[1125]), .Z(n34194) );
  XNOR U34279 ( .A(q[4]), .B(DB[1124]), .Z(n26360) );
  IV U34280 ( .A(n26374), .Z(n34192) );
  XOR U34281 ( .A(n34195), .B(n34196), .Z(n26374) );
  XNOR U34282 ( .A(n26370), .B(n26372), .Z(n34196) );
  XNOR U34283 ( .A(q[0]), .B(DB[1120]), .Z(n26372) );
  XNOR U34284 ( .A(q[3]), .B(DB[1123]), .Z(n26370) );
  IV U34285 ( .A(n26369), .Z(n34195) );
  XNOR U34286 ( .A(n26367), .B(n34197), .Z(n26369) );
  XNOR U34287 ( .A(q[2]), .B(DB[1122]), .Z(n34197) );
  XNOR U34288 ( .A(q[1]), .B(DB[1121]), .Z(n26367) );
  XOR U34289 ( .A(n34198), .B(n26332), .Z(n26295) );
  XOR U34290 ( .A(n34199), .B(n26320), .Z(n26332) );
  XNOR U34291 ( .A(q[6]), .B(DB[1133]), .Z(n26320) );
  IV U34292 ( .A(n26319), .Z(n34199) );
  XNOR U34293 ( .A(n26317), .B(n34200), .Z(n26319) );
  XNOR U34294 ( .A(q[5]), .B(DB[1132]), .Z(n34200) );
  XNOR U34295 ( .A(q[4]), .B(DB[1131]), .Z(n26317) );
  IV U34296 ( .A(n26331), .Z(n34198) );
  XOR U34297 ( .A(n34201), .B(n34202), .Z(n26331) );
  XNOR U34298 ( .A(n26327), .B(n26329), .Z(n34202) );
  XNOR U34299 ( .A(q[0]), .B(DB[1127]), .Z(n26329) );
  XNOR U34300 ( .A(q[3]), .B(DB[1130]), .Z(n26327) );
  IV U34301 ( .A(n26326), .Z(n34201) );
  XNOR U34302 ( .A(n26324), .B(n34203), .Z(n26326) );
  XNOR U34303 ( .A(q[2]), .B(DB[1129]), .Z(n34203) );
  XNOR U34304 ( .A(q[1]), .B(DB[1128]), .Z(n26324) );
  XOR U34305 ( .A(n34204), .B(n26289), .Z(n26252) );
  XOR U34306 ( .A(n34205), .B(n26277), .Z(n26289) );
  XNOR U34307 ( .A(q[6]), .B(DB[1140]), .Z(n26277) );
  IV U34308 ( .A(n26276), .Z(n34205) );
  XNOR U34309 ( .A(n26274), .B(n34206), .Z(n26276) );
  XNOR U34310 ( .A(q[5]), .B(DB[1139]), .Z(n34206) );
  XNOR U34311 ( .A(q[4]), .B(DB[1138]), .Z(n26274) );
  IV U34312 ( .A(n26288), .Z(n34204) );
  XOR U34313 ( .A(n34207), .B(n34208), .Z(n26288) );
  XNOR U34314 ( .A(n26284), .B(n26286), .Z(n34208) );
  XNOR U34315 ( .A(q[0]), .B(DB[1134]), .Z(n26286) );
  XNOR U34316 ( .A(q[3]), .B(DB[1137]), .Z(n26284) );
  IV U34317 ( .A(n26283), .Z(n34207) );
  XNOR U34318 ( .A(n26281), .B(n34209), .Z(n26283) );
  XNOR U34319 ( .A(q[2]), .B(DB[1136]), .Z(n34209) );
  XNOR U34320 ( .A(q[1]), .B(DB[1135]), .Z(n26281) );
  XOR U34321 ( .A(n34210), .B(n26246), .Z(n26209) );
  XOR U34322 ( .A(n34211), .B(n26234), .Z(n26246) );
  XNOR U34323 ( .A(q[6]), .B(DB[1147]), .Z(n26234) );
  IV U34324 ( .A(n26233), .Z(n34211) );
  XNOR U34325 ( .A(n26231), .B(n34212), .Z(n26233) );
  XNOR U34326 ( .A(q[5]), .B(DB[1146]), .Z(n34212) );
  XNOR U34327 ( .A(q[4]), .B(DB[1145]), .Z(n26231) );
  IV U34328 ( .A(n26245), .Z(n34210) );
  XOR U34329 ( .A(n34213), .B(n34214), .Z(n26245) );
  XNOR U34330 ( .A(n26241), .B(n26243), .Z(n34214) );
  XNOR U34331 ( .A(q[0]), .B(DB[1141]), .Z(n26243) );
  XNOR U34332 ( .A(q[3]), .B(DB[1144]), .Z(n26241) );
  IV U34333 ( .A(n26240), .Z(n34213) );
  XNOR U34334 ( .A(n26238), .B(n34215), .Z(n26240) );
  XNOR U34335 ( .A(q[2]), .B(DB[1143]), .Z(n34215) );
  XNOR U34336 ( .A(q[1]), .B(DB[1142]), .Z(n26238) );
  XOR U34337 ( .A(n34216), .B(n26203), .Z(n26166) );
  XOR U34338 ( .A(n34217), .B(n26191), .Z(n26203) );
  XNOR U34339 ( .A(q[6]), .B(DB[1154]), .Z(n26191) );
  IV U34340 ( .A(n26190), .Z(n34217) );
  XNOR U34341 ( .A(n26188), .B(n34218), .Z(n26190) );
  XNOR U34342 ( .A(q[5]), .B(DB[1153]), .Z(n34218) );
  XNOR U34343 ( .A(q[4]), .B(DB[1152]), .Z(n26188) );
  IV U34344 ( .A(n26202), .Z(n34216) );
  XOR U34345 ( .A(n34219), .B(n34220), .Z(n26202) );
  XNOR U34346 ( .A(n26198), .B(n26200), .Z(n34220) );
  XNOR U34347 ( .A(q[0]), .B(DB[1148]), .Z(n26200) );
  XNOR U34348 ( .A(q[3]), .B(DB[1151]), .Z(n26198) );
  IV U34349 ( .A(n26197), .Z(n34219) );
  XNOR U34350 ( .A(n26195), .B(n34221), .Z(n26197) );
  XNOR U34351 ( .A(q[2]), .B(DB[1150]), .Z(n34221) );
  XNOR U34352 ( .A(q[1]), .B(DB[1149]), .Z(n26195) );
  XOR U34353 ( .A(n34222), .B(n26160), .Z(n26123) );
  XOR U34354 ( .A(n34223), .B(n26148), .Z(n26160) );
  XNOR U34355 ( .A(q[6]), .B(DB[1161]), .Z(n26148) );
  IV U34356 ( .A(n26147), .Z(n34223) );
  XNOR U34357 ( .A(n26145), .B(n34224), .Z(n26147) );
  XNOR U34358 ( .A(q[5]), .B(DB[1160]), .Z(n34224) );
  XNOR U34359 ( .A(q[4]), .B(DB[1159]), .Z(n26145) );
  IV U34360 ( .A(n26159), .Z(n34222) );
  XOR U34361 ( .A(n34225), .B(n34226), .Z(n26159) );
  XNOR U34362 ( .A(n26155), .B(n26157), .Z(n34226) );
  XNOR U34363 ( .A(q[0]), .B(DB[1155]), .Z(n26157) );
  XNOR U34364 ( .A(q[3]), .B(DB[1158]), .Z(n26155) );
  IV U34365 ( .A(n26154), .Z(n34225) );
  XNOR U34366 ( .A(n26152), .B(n34227), .Z(n26154) );
  XNOR U34367 ( .A(q[2]), .B(DB[1157]), .Z(n34227) );
  XNOR U34368 ( .A(q[1]), .B(DB[1156]), .Z(n26152) );
  XOR U34369 ( .A(n34228), .B(n26117), .Z(n26080) );
  XOR U34370 ( .A(n34229), .B(n26105), .Z(n26117) );
  XNOR U34371 ( .A(q[6]), .B(DB[1168]), .Z(n26105) );
  IV U34372 ( .A(n26104), .Z(n34229) );
  XNOR U34373 ( .A(n26102), .B(n34230), .Z(n26104) );
  XNOR U34374 ( .A(q[5]), .B(DB[1167]), .Z(n34230) );
  XNOR U34375 ( .A(q[4]), .B(DB[1166]), .Z(n26102) );
  IV U34376 ( .A(n26116), .Z(n34228) );
  XOR U34377 ( .A(n34231), .B(n34232), .Z(n26116) );
  XNOR U34378 ( .A(n26112), .B(n26114), .Z(n34232) );
  XNOR U34379 ( .A(q[0]), .B(DB[1162]), .Z(n26114) );
  XNOR U34380 ( .A(q[3]), .B(DB[1165]), .Z(n26112) );
  IV U34381 ( .A(n26111), .Z(n34231) );
  XNOR U34382 ( .A(n26109), .B(n34233), .Z(n26111) );
  XNOR U34383 ( .A(q[2]), .B(DB[1164]), .Z(n34233) );
  XNOR U34384 ( .A(q[1]), .B(DB[1163]), .Z(n26109) );
  XOR U34385 ( .A(n34234), .B(n26074), .Z(n26037) );
  XOR U34386 ( .A(n34235), .B(n26062), .Z(n26074) );
  XNOR U34387 ( .A(q[6]), .B(DB[1175]), .Z(n26062) );
  IV U34388 ( .A(n26061), .Z(n34235) );
  XNOR U34389 ( .A(n26059), .B(n34236), .Z(n26061) );
  XNOR U34390 ( .A(q[5]), .B(DB[1174]), .Z(n34236) );
  XNOR U34391 ( .A(q[4]), .B(DB[1173]), .Z(n26059) );
  IV U34392 ( .A(n26073), .Z(n34234) );
  XOR U34393 ( .A(n34237), .B(n34238), .Z(n26073) );
  XNOR U34394 ( .A(n26069), .B(n26071), .Z(n34238) );
  XNOR U34395 ( .A(q[0]), .B(DB[1169]), .Z(n26071) );
  XNOR U34396 ( .A(q[3]), .B(DB[1172]), .Z(n26069) );
  IV U34397 ( .A(n26068), .Z(n34237) );
  XNOR U34398 ( .A(n26066), .B(n34239), .Z(n26068) );
  XNOR U34399 ( .A(q[2]), .B(DB[1171]), .Z(n34239) );
  XNOR U34400 ( .A(q[1]), .B(DB[1170]), .Z(n26066) );
  XOR U34401 ( .A(n34240), .B(n26031), .Z(n25994) );
  XOR U34402 ( .A(n34241), .B(n26019), .Z(n26031) );
  XNOR U34403 ( .A(q[6]), .B(DB[1182]), .Z(n26019) );
  IV U34404 ( .A(n26018), .Z(n34241) );
  XNOR U34405 ( .A(n26016), .B(n34242), .Z(n26018) );
  XNOR U34406 ( .A(q[5]), .B(DB[1181]), .Z(n34242) );
  XNOR U34407 ( .A(q[4]), .B(DB[1180]), .Z(n26016) );
  IV U34408 ( .A(n26030), .Z(n34240) );
  XOR U34409 ( .A(n34243), .B(n34244), .Z(n26030) );
  XNOR U34410 ( .A(n26026), .B(n26028), .Z(n34244) );
  XNOR U34411 ( .A(q[0]), .B(DB[1176]), .Z(n26028) );
  XNOR U34412 ( .A(q[3]), .B(DB[1179]), .Z(n26026) );
  IV U34413 ( .A(n26025), .Z(n34243) );
  XNOR U34414 ( .A(n26023), .B(n34245), .Z(n26025) );
  XNOR U34415 ( .A(q[2]), .B(DB[1178]), .Z(n34245) );
  XNOR U34416 ( .A(q[1]), .B(DB[1177]), .Z(n26023) );
  XOR U34417 ( .A(n34246), .B(n25988), .Z(n25951) );
  XOR U34418 ( .A(n34247), .B(n25976), .Z(n25988) );
  XNOR U34419 ( .A(q[6]), .B(DB[1189]), .Z(n25976) );
  IV U34420 ( .A(n25975), .Z(n34247) );
  XNOR U34421 ( .A(n25973), .B(n34248), .Z(n25975) );
  XNOR U34422 ( .A(q[5]), .B(DB[1188]), .Z(n34248) );
  XNOR U34423 ( .A(q[4]), .B(DB[1187]), .Z(n25973) );
  IV U34424 ( .A(n25987), .Z(n34246) );
  XOR U34425 ( .A(n34249), .B(n34250), .Z(n25987) );
  XNOR U34426 ( .A(n25983), .B(n25985), .Z(n34250) );
  XNOR U34427 ( .A(q[0]), .B(DB[1183]), .Z(n25985) );
  XNOR U34428 ( .A(q[3]), .B(DB[1186]), .Z(n25983) );
  IV U34429 ( .A(n25982), .Z(n34249) );
  XNOR U34430 ( .A(n25980), .B(n34251), .Z(n25982) );
  XNOR U34431 ( .A(q[2]), .B(DB[1185]), .Z(n34251) );
  XNOR U34432 ( .A(q[1]), .B(DB[1184]), .Z(n25980) );
  XOR U34433 ( .A(n34252), .B(n25945), .Z(n25908) );
  XOR U34434 ( .A(n34253), .B(n25933), .Z(n25945) );
  XNOR U34435 ( .A(q[6]), .B(DB[1196]), .Z(n25933) );
  IV U34436 ( .A(n25932), .Z(n34253) );
  XNOR U34437 ( .A(n25930), .B(n34254), .Z(n25932) );
  XNOR U34438 ( .A(q[5]), .B(DB[1195]), .Z(n34254) );
  XNOR U34439 ( .A(q[4]), .B(DB[1194]), .Z(n25930) );
  IV U34440 ( .A(n25944), .Z(n34252) );
  XOR U34441 ( .A(n34255), .B(n34256), .Z(n25944) );
  XNOR U34442 ( .A(n25940), .B(n25942), .Z(n34256) );
  XNOR U34443 ( .A(q[0]), .B(DB[1190]), .Z(n25942) );
  XNOR U34444 ( .A(q[3]), .B(DB[1193]), .Z(n25940) );
  IV U34445 ( .A(n25939), .Z(n34255) );
  XNOR U34446 ( .A(n25937), .B(n34257), .Z(n25939) );
  XNOR U34447 ( .A(q[2]), .B(DB[1192]), .Z(n34257) );
  XNOR U34448 ( .A(q[1]), .B(DB[1191]), .Z(n25937) );
  XOR U34449 ( .A(n34258), .B(n25902), .Z(n25865) );
  XOR U34450 ( .A(n34259), .B(n25890), .Z(n25902) );
  XNOR U34451 ( .A(q[6]), .B(DB[1203]), .Z(n25890) );
  IV U34452 ( .A(n25889), .Z(n34259) );
  XNOR U34453 ( .A(n25887), .B(n34260), .Z(n25889) );
  XNOR U34454 ( .A(q[5]), .B(DB[1202]), .Z(n34260) );
  XNOR U34455 ( .A(q[4]), .B(DB[1201]), .Z(n25887) );
  IV U34456 ( .A(n25901), .Z(n34258) );
  XOR U34457 ( .A(n34261), .B(n34262), .Z(n25901) );
  XNOR U34458 ( .A(n25897), .B(n25899), .Z(n34262) );
  XNOR U34459 ( .A(q[0]), .B(DB[1197]), .Z(n25899) );
  XNOR U34460 ( .A(q[3]), .B(DB[1200]), .Z(n25897) );
  IV U34461 ( .A(n25896), .Z(n34261) );
  XNOR U34462 ( .A(n25894), .B(n34263), .Z(n25896) );
  XNOR U34463 ( .A(q[2]), .B(DB[1199]), .Z(n34263) );
  XNOR U34464 ( .A(q[1]), .B(DB[1198]), .Z(n25894) );
  XOR U34465 ( .A(n34264), .B(n25859), .Z(n25822) );
  XOR U34466 ( .A(n34265), .B(n25847), .Z(n25859) );
  XNOR U34467 ( .A(q[6]), .B(DB[1210]), .Z(n25847) );
  IV U34468 ( .A(n25846), .Z(n34265) );
  XNOR U34469 ( .A(n25844), .B(n34266), .Z(n25846) );
  XNOR U34470 ( .A(q[5]), .B(DB[1209]), .Z(n34266) );
  XNOR U34471 ( .A(q[4]), .B(DB[1208]), .Z(n25844) );
  IV U34472 ( .A(n25858), .Z(n34264) );
  XOR U34473 ( .A(n34267), .B(n34268), .Z(n25858) );
  XNOR U34474 ( .A(n25854), .B(n25856), .Z(n34268) );
  XNOR U34475 ( .A(q[0]), .B(DB[1204]), .Z(n25856) );
  XNOR U34476 ( .A(q[3]), .B(DB[1207]), .Z(n25854) );
  IV U34477 ( .A(n25853), .Z(n34267) );
  XNOR U34478 ( .A(n25851), .B(n34269), .Z(n25853) );
  XNOR U34479 ( .A(q[2]), .B(DB[1206]), .Z(n34269) );
  XNOR U34480 ( .A(q[1]), .B(DB[1205]), .Z(n25851) );
  XOR U34481 ( .A(n34270), .B(n25816), .Z(n25779) );
  XOR U34482 ( .A(n34271), .B(n25804), .Z(n25816) );
  XNOR U34483 ( .A(q[6]), .B(DB[1217]), .Z(n25804) );
  IV U34484 ( .A(n25803), .Z(n34271) );
  XNOR U34485 ( .A(n25801), .B(n34272), .Z(n25803) );
  XNOR U34486 ( .A(q[5]), .B(DB[1216]), .Z(n34272) );
  XNOR U34487 ( .A(q[4]), .B(DB[1215]), .Z(n25801) );
  IV U34488 ( .A(n25815), .Z(n34270) );
  XOR U34489 ( .A(n34273), .B(n34274), .Z(n25815) );
  XNOR U34490 ( .A(n25811), .B(n25813), .Z(n34274) );
  XNOR U34491 ( .A(q[0]), .B(DB[1211]), .Z(n25813) );
  XNOR U34492 ( .A(q[3]), .B(DB[1214]), .Z(n25811) );
  IV U34493 ( .A(n25810), .Z(n34273) );
  XNOR U34494 ( .A(n25808), .B(n34275), .Z(n25810) );
  XNOR U34495 ( .A(q[2]), .B(DB[1213]), .Z(n34275) );
  XNOR U34496 ( .A(q[1]), .B(DB[1212]), .Z(n25808) );
  XOR U34497 ( .A(n34276), .B(n25773), .Z(n25736) );
  XOR U34498 ( .A(n34277), .B(n25761), .Z(n25773) );
  XNOR U34499 ( .A(q[6]), .B(DB[1224]), .Z(n25761) );
  IV U34500 ( .A(n25760), .Z(n34277) );
  XNOR U34501 ( .A(n25758), .B(n34278), .Z(n25760) );
  XNOR U34502 ( .A(q[5]), .B(DB[1223]), .Z(n34278) );
  XNOR U34503 ( .A(q[4]), .B(DB[1222]), .Z(n25758) );
  IV U34504 ( .A(n25772), .Z(n34276) );
  XOR U34505 ( .A(n34279), .B(n34280), .Z(n25772) );
  XNOR U34506 ( .A(n25768), .B(n25770), .Z(n34280) );
  XNOR U34507 ( .A(q[0]), .B(DB[1218]), .Z(n25770) );
  XNOR U34508 ( .A(q[3]), .B(DB[1221]), .Z(n25768) );
  IV U34509 ( .A(n25767), .Z(n34279) );
  XNOR U34510 ( .A(n25765), .B(n34281), .Z(n25767) );
  XNOR U34511 ( .A(q[2]), .B(DB[1220]), .Z(n34281) );
  XNOR U34512 ( .A(q[1]), .B(DB[1219]), .Z(n25765) );
  XOR U34513 ( .A(n34282), .B(n25730), .Z(n25693) );
  XOR U34514 ( .A(n34283), .B(n25718), .Z(n25730) );
  XNOR U34515 ( .A(q[6]), .B(DB[1231]), .Z(n25718) );
  IV U34516 ( .A(n25717), .Z(n34283) );
  XNOR U34517 ( .A(n25715), .B(n34284), .Z(n25717) );
  XNOR U34518 ( .A(q[5]), .B(DB[1230]), .Z(n34284) );
  XNOR U34519 ( .A(q[4]), .B(DB[1229]), .Z(n25715) );
  IV U34520 ( .A(n25729), .Z(n34282) );
  XOR U34521 ( .A(n34285), .B(n34286), .Z(n25729) );
  XNOR U34522 ( .A(n25725), .B(n25727), .Z(n34286) );
  XNOR U34523 ( .A(q[0]), .B(DB[1225]), .Z(n25727) );
  XNOR U34524 ( .A(q[3]), .B(DB[1228]), .Z(n25725) );
  IV U34525 ( .A(n25724), .Z(n34285) );
  XNOR U34526 ( .A(n25722), .B(n34287), .Z(n25724) );
  XNOR U34527 ( .A(q[2]), .B(DB[1227]), .Z(n34287) );
  XNOR U34528 ( .A(q[1]), .B(DB[1226]), .Z(n25722) );
  XOR U34529 ( .A(n34288), .B(n25687), .Z(n25650) );
  XOR U34530 ( .A(n34289), .B(n25675), .Z(n25687) );
  XNOR U34531 ( .A(q[6]), .B(DB[1238]), .Z(n25675) );
  IV U34532 ( .A(n25674), .Z(n34289) );
  XNOR U34533 ( .A(n25672), .B(n34290), .Z(n25674) );
  XNOR U34534 ( .A(q[5]), .B(DB[1237]), .Z(n34290) );
  XNOR U34535 ( .A(q[4]), .B(DB[1236]), .Z(n25672) );
  IV U34536 ( .A(n25686), .Z(n34288) );
  XOR U34537 ( .A(n34291), .B(n34292), .Z(n25686) );
  XNOR U34538 ( .A(n25682), .B(n25684), .Z(n34292) );
  XNOR U34539 ( .A(q[0]), .B(DB[1232]), .Z(n25684) );
  XNOR U34540 ( .A(q[3]), .B(DB[1235]), .Z(n25682) );
  IV U34541 ( .A(n25681), .Z(n34291) );
  XNOR U34542 ( .A(n25679), .B(n34293), .Z(n25681) );
  XNOR U34543 ( .A(q[2]), .B(DB[1234]), .Z(n34293) );
  XNOR U34544 ( .A(q[1]), .B(DB[1233]), .Z(n25679) );
  XOR U34545 ( .A(n34294), .B(n25644), .Z(n25607) );
  XOR U34546 ( .A(n34295), .B(n25632), .Z(n25644) );
  XNOR U34547 ( .A(q[6]), .B(DB[1245]), .Z(n25632) );
  IV U34548 ( .A(n25631), .Z(n34295) );
  XNOR U34549 ( .A(n25629), .B(n34296), .Z(n25631) );
  XNOR U34550 ( .A(q[5]), .B(DB[1244]), .Z(n34296) );
  XNOR U34551 ( .A(q[4]), .B(DB[1243]), .Z(n25629) );
  IV U34552 ( .A(n25643), .Z(n34294) );
  XOR U34553 ( .A(n34297), .B(n34298), .Z(n25643) );
  XNOR U34554 ( .A(n25639), .B(n25641), .Z(n34298) );
  XNOR U34555 ( .A(q[0]), .B(DB[1239]), .Z(n25641) );
  XNOR U34556 ( .A(q[3]), .B(DB[1242]), .Z(n25639) );
  IV U34557 ( .A(n25638), .Z(n34297) );
  XNOR U34558 ( .A(n25636), .B(n34299), .Z(n25638) );
  XNOR U34559 ( .A(q[2]), .B(DB[1241]), .Z(n34299) );
  XNOR U34560 ( .A(q[1]), .B(DB[1240]), .Z(n25636) );
  XOR U34561 ( .A(n34300), .B(n25601), .Z(n25564) );
  XOR U34562 ( .A(n34301), .B(n25589), .Z(n25601) );
  XNOR U34563 ( .A(q[6]), .B(DB[1252]), .Z(n25589) );
  IV U34564 ( .A(n25588), .Z(n34301) );
  XNOR U34565 ( .A(n25586), .B(n34302), .Z(n25588) );
  XNOR U34566 ( .A(q[5]), .B(DB[1251]), .Z(n34302) );
  XNOR U34567 ( .A(q[4]), .B(DB[1250]), .Z(n25586) );
  IV U34568 ( .A(n25600), .Z(n34300) );
  XOR U34569 ( .A(n34303), .B(n34304), .Z(n25600) );
  XNOR U34570 ( .A(n25596), .B(n25598), .Z(n34304) );
  XNOR U34571 ( .A(q[0]), .B(DB[1246]), .Z(n25598) );
  XNOR U34572 ( .A(q[3]), .B(DB[1249]), .Z(n25596) );
  IV U34573 ( .A(n25595), .Z(n34303) );
  XNOR U34574 ( .A(n25593), .B(n34305), .Z(n25595) );
  XNOR U34575 ( .A(q[2]), .B(DB[1248]), .Z(n34305) );
  XNOR U34576 ( .A(q[1]), .B(DB[1247]), .Z(n25593) );
  XOR U34577 ( .A(n34306), .B(n25558), .Z(n25521) );
  XOR U34578 ( .A(n34307), .B(n25546), .Z(n25558) );
  XNOR U34579 ( .A(q[6]), .B(DB[1259]), .Z(n25546) );
  IV U34580 ( .A(n25545), .Z(n34307) );
  XNOR U34581 ( .A(n25543), .B(n34308), .Z(n25545) );
  XNOR U34582 ( .A(q[5]), .B(DB[1258]), .Z(n34308) );
  XNOR U34583 ( .A(q[4]), .B(DB[1257]), .Z(n25543) );
  IV U34584 ( .A(n25557), .Z(n34306) );
  XOR U34585 ( .A(n34309), .B(n34310), .Z(n25557) );
  XNOR U34586 ( .A(n25553), .B(n25555), .Z(n34310) );
  XNOR U34587 ( .A(q[0]), .B(DB[1253]), .Z(n25555) );
  XNOR U34588 ( .A(q[3]), .B(DB[1256]), .Z(n25553) );
  IV U34589 ( .A(n25552), .Z(n34309) );
  XNOR U34590 ( .A(n25550), .B(n34311), .Z(n25552) );
  XNOR U34591 ( .A(q[2]), .B(DB[1255]), .Z(n34311) );
  XNOR U34592 ( .A(q[1]), .B(DB[1254]), .Z(n25550) );
  XOR U34593 ( .A(n34312), .B(n25515), .Z(n25478) );
  XOR U34594 ( .A(n34313), .B(n25503), .Z(n25515) );
  XNOR U34595 ( .A(q[6]), .B(DB[1266]), .Z(n25503) );
  IV U34596 ( .A(n25502), .Z(n34313) );
  XNOR U34597 ( .A(n25500), .B(n34314), .Z(n25502) );
  XNOR U34598 ( .A(q[5]), .B(DB[1265]), .Z(n34314) );
  XNOR U34599 ( .A(q[4]), .B(DB[1264]), .Z(n25500) );
  IV U34600 ( .A(n25514), .Z(n34312) );
  XOR U34601 ( .A(n34315), .B(n34316), .Z(n25514) );
  XNOR U34602 ( .A(n25510), .B(n25512), .Z(n34316) );
  XNOR U34603 ( .A(q[0]), .B(DB[1260]), .Z(n25512) );
  XNOR U34604 ( .A(q[3]), .B(DB[1263]), .Z(n25510) );
  IV U34605 ( .A(n25509), .Z(n34315) );
  XNOR U34606 ( .A(n25507), .B(n34317), .Z(n25509) );
  XNOR U34607 ( .A(q[2]), .B(DB[1262]), .Z(n34317) );
  XNOR U34608 ( .A(q[1]), .B(DB[1261]), .Z(n25507) );
  XOR U34609 ( .A(n34318), .B(n25472), .Z(n25435) );
  XOR U34610 ( .A(n34319), .B(n25460), .Z(n25472) );
  XNOR U34611 ( .A(q[6]), .B(DB[1273]), .Z(n25460) );
  IV U34612 ( .A(n25459), .Z(n34319) );
  XNOR U34613 ( .A(n25457), .B(n34320), .Z(n25459) );
  XNOR U34614 ( .A(q[5]), .B(DB[1272]), .Z(n34320) );
  XNOR U34615 ( .A(q[4]), .B(DB[1271]), .Z(n25457) );
  IV U34616 ( .A(n25471), .Z(n34318) );
  XOR U34617 ( .A(n34321), .B(n34322), .Z(n25471) );
  XNOR U34618 ( .A(n25467), .B(n25469), .Z(n34322) );
  XNOR U34619 ( .A(q[0]), .B(DB[1267]), .Z(n25469) );
  XNOR U34620 ( .A(q[3]), .B(DB[1270]), .Z(n25467) );
  IV U34621 ( .A(n25466), .Z(n34321) );
  XNOR U34622 ( .A(n25464), .B(n34323), .Z(n25466) );
  XNOR U34623 ( .A(q[2]), .B(DB[1269]), .Z(n34323) );
  XNOR U34624 ( .A(q[1]), .B(DB[1268]), .Z(n25464) );
  XOR U34625 ( .A(n34324), .B(n25429), .Z(n25392) );
  XOR U34626 ( .A(n34325), .B(n25417), .Z(n25429) );
  XNOR U34627 ( .A(q[6]), .B(DB[1280]), .Z(n25417) );
  IV U34628 ( .A(n25416), .Z(n34325) );
  XNOR U34629 ( .A(n25414), .B(n34326), .Z(n25416) );
  XNOR U34630 ( .A(q[5]), .B(DB[1279]), .Z(n34326) );
  XNOR U34631 ( .A(q[4]), .B(DB[1278]), .Z(n25414) );
  IV U34632 ( .A(n25428), .Z(n34324) );
  XOR U34633 ( .A(n34327), .B(n34328), .Z(n25428) );
  XNOR U34634 ( .A(n25424), .B(n25426), .Z(n34328) );
  XNOR U34635 ( .A(q[0]), .B(DB[1274]), .Z(n25426) );
  XNOR U34636 ( .A(q[3]), .B(DB[1277]), .Z(n25424) );
  IV U34637 ( .A(n25423), .Z(n34327) );
  XNOR U34638 ( .A(n25421), .B(n34329), .Z(n25423) );
  XNOR U34639 ( .A(q[2]), .B(DB[1276]), .Z(n34329) );
  XNOR U34640 ( .A(q[1]), .B(DB[1275]), .Z(n25421) );
  XOR U34641 ( .A(n34330), .B(n25386), .Z(n25349) );
  XOR U34642 ( .A(n34331), .B(n25374), .Z(n25386) );
  XNOR U34643 ( .A(q[6]), .B(DB[1287]), .Z(n25374) );
  IV U34644 ( .A(n25373), .Z(n34331) );
  XNOR U34645 ( .A(n25371), .B(n34332), .Z(n25373) );
  XNOR U34646 ( .A(q[5]), .B(DB[1286]), .Z(n34332) );
  XNOR U34647 ( .A(q[4]), .B(DB[1285]), .Z(n25371) );
  IV U34648 ( .A(n25385), .Z(n34330) );
  XOR U34649 ( .A(n34333), .B(n34334), .Z(n25385) );
  XNOR U34650 ( .A(n25381), .B(n25383), .Z(n34334) );
  XNOR U34651 ( .A(q[0]), .B(DB[1281]), .Z(n25383) );
  XNOR U34652 ( .A(q[3]), .B(DB[1284]), .Z(n25381) );
  IV U34653 ( .A(n25380), .Z(n34333) );
  XNOR U34654 ( .A(n25378), .B(n34335), .Z(n25380) );
  XNOR U34655 ( .A(q[2]), .B(DB[1283]), .Z(n34335) );
  XNOR U34656 ( .A(q[1]), .B(DB[1282]), .Z(n25378) );
  XOR U34657 ( .A(n34336), .B(n25343), .Z(n25306) );
  XOR U34658 ( .A(n34337), .B(n25331), .Z(n25343) );
  XNOR U34659 ( .A(q[6]), .B(DB[1294]), .Z(n25331) );
  IV U34660 ( .A(n25330), .Z(n34337) );
  XNOR U34661 ( .A(n25328), .B(n34338), .Z(n25330) );
  XNOR U34662 ( .A(q[5]), .B(DB[1293]), .Z(n34338) );
  XNOR U34663 ( .A(q[4]), .B(DB[1292]), .Z(n25328) );
  IV U34664 ( .A(n25342), .Z(n34336) );
  XOR U34665 ( .A(n34339), .B(n34340), .Z(n25342) );
  XNOR U34666 ( .A(n25338), .B(n25340), .Z(n34340) );
  XNOR U34667 ( .A(q[0]), .B(DB[1288]), .Z(n25340) );
  XNOR U34668 ( .A(q[3]), .B(DB[1291]), .Z(n25338) );
  IV U34669 ( .A(n25337), .Z(n34339) );
  XNOR U34670 ( .A(n25335), .B(n34341), .Z(n25337) );
  XNOR U34671 ( .A(q[2]), .B(DB[1290]), .Z(n34341) );
  XNOR U34672 ( .A(q[1]), .B(DB[1289]), .Z(n25335) );
  XOR U34673 ( .A(n34342), .B(n25300), .Z(n25263) );
  XOR U34674 ( .A(n34343), .B(n25288), .Z(n25300) );
  XNOR U34675 ( .A(q[6]), .B(DB[1301]), .Z(n25288) );
  IV U34676 ( .A(n25287), .Z(n34343) );
  XNOR U34677 ( .A(n25285), .B(n34344), .Z(n25287) );
  XNOR U34678 ( .A(q[5]), .B(DB[1300]), .Z(n34344) );
  XNOR U34679 ( .A(q[4]), .B(DB[1299]), .Z(n25285) );
  IV U34680 ( .A(n25299), .Z(n34342) );
  XOR U34681 ( .A(n34345), .B(n34346), .Z(n25299) );
  XNOR U34682 ( .A(n25295), .B(n25297), .Z(n34346) );
  XNOR U34683 ( .A(q[0]), .B(DB[1295]), .Z(n25297) );
  XNOR U34684 ( .A(q[3]), .B(DB[1298]), .Z(n25295) );
  IV U34685 ( .A(n25294), .Z(n34345) );
  XNOR U34686 ( .A(n25292), .B(n34347), .Z(n25294) );
  XNOR U34687 ( .A(q[2]), .B(DB[1297]), .Z(n34347) );
  XNOR U34688 ( .A(q[1]), .B(DB[1296]), .Z(n25292) );
  XOR U34689 ( .A(n34348), .B(n25257), .Z(n25220) );
  XOR U34690 ( .A(n34349), .B(n25245), .Z(n25257) );
  XNOR U34691 ( .A(q[6]), .B(DB[1308]), .Z(n25245) );
  IV U34692 ( .A(n25244), .Z(n34349) );
  XNOR U34693 ( .A(n25242), .B(n34350), .Z(n25244) );
  XNOR U34694 ( .A(q[5]), .B(DB[1307]), .Z(n34350) );
  XNOR U34695 ( .A(q[4]), .B(DB[1306]), .Z(n25242) );
  IV U34696 ( .A(n25256), .Z(n34348) );
  XOR U34697 ( .A(n34351), .B(n34352), .Z(n25256) );
  XNOR U34698 ( .A(n25252), .B(n25254), .Z(n34352) );
  XNOR U34699 ( .A(q[0]), .B(DB[1302]), .Z(n25254) );
  XNOR U34700 ( .A(q[3]), .B(DB[1305]), .Z(n25252) );
  IV U34701 ( .A(n25251), .Z(n34351) );
  XNOR U34702 ( .A(n25249), .B(n34353), .Z(n25251) );
  XNOR U34703 ( .A(q[2]), .B(DB[1304]), .Z(n34353) );
  XNOR U34704 ( .A(q[1]), .B(DB[1303]), .Z(n25249) );
  XOR U34705 ( .A(n34354), .B(n25214), .Z(n25177) );
  XOR U34706 ( .A(n34355), .B(n25202), .Z(n25214) );
  XNOR U34707 ( .A(q[6]), .B(DB[1315]), .Z(n25202) );
  IV U34708 ( .A(n25201), .Z(n34355) );
  XNOR U34709 ( .A(n25199), .B(n34356), .Z(n25201) );
  XNOR U34710 ( .A(q[5]), .B(DB[1314]), .Z(n34356) );
  XNOR U34711 ( .A(q[4]), .B(DB[1313]), .Z(n25199) );
  IV U34712 ( .A(n25213), .Z(n34354) );
  XOR U34713 ( .A(n34357), .B(n34358), .Z(n25213) );
  XNOR U34714 ( .A(n25209), .B(n25211), .Z(n34358) );
  XNOR U34715 ( .A(q[0]), .B(DB[1309]), .Z(n25211) );
  XNOR U34716 ( .A(q[3]), .B(DB[1312]), .Z(n25209) );
  IV U34717 ( .A(n25208), .Z(n34357) );
  XNOR U34718 ( .A(n25206), .B(n34359), .Z(n25208) );
  XNOR U34719 ( .A(q[2]), .B(DB[1311]), .Z(n34359) );
  XNOR U34720 ( .A(q[1]), .B(DB[1310]), .Z(n25206) );
  XOR U34721 ( .A(n34360), .B(n25171), .Z(n25134) );
  XOR U34722 ( .A(n34361), .B(n25159), .Z(n25171) );
  XNOR U34723 ( .A(q[6]), .B(DB[1322]), .Z(n25159) );
  IV U34724 ( .A(n25158), .Z(n34361) );
  XNOR U34725 ( .A(n25156), .B(n34362), .Z(n25158) );
  XNOR U34726 ( .A(q[5]), .B(DB[1321]), .Z(n34362) );
  XNOR U34727 ( .A(q[4]), .B(DB[1320]), .Z(n25156) );
  IV U34728 ( .A(n25170), .Z(n34360) );
  XOR U34729 ( .A(n34363), .B(n34364), .Z(n25170) );
  XNOR U34730 ( .A(n25166), .B(n25168), .Z(n34364) );
  XNOR U34731 ( .A(q[0]), .B(DB[1316]), .Z(n25168) );
  XNOR U34732 ( .A(q[3]), .B(DB[1319]), .Z(n25166) );
  IV U34733 ( .A(n25165), .Z(n34363) );
  XNOR U34734 ( .A(n25163), .B(n34365), .Z(n25165) );
  XNOR U34735 ( .A(q[2]), .B(DB[1318]), .Z(n34365) );
  XNOR U34736 ( .A(q[1]), .B(DB[1317]), .Z(n25163) );
  XOR U34737 ( .A(n34366), .B(n25128), .Z(n25091) );
  XOR U34738 ( .A(n34367), .B(n25116), .Z(n25128) );
  XNOR U34739 ( .A(q[6]), .B(DB[1329]), .Z(n25116) );
  IV U34740 ( .A(n25115), .Z(n34367) );
  XNOR U34741 ( .A(n25113), .B(n34368), .Z(n25115) );
  XNOR U34742 ( .A(q[5]), .B(DB[1328]), .Z(n34368) );
  XNOR U34743 ( .A(q[4]), .B(DB[1327]), .Z(n25113) );
  IV U34744 ( .A(n25127), .Z(n34366) );
  XOR U34745 ( .A(n34369), .B(n34370), .Z(n25127) );
  XNOR U34746 ( .A(n25123), .B(n25125), .Z(n34370) );
  XNOR U34747 ( .A(q[0]), .B(DB[1323]), .Z(n25125) );
  XNOR U34748 ( .A(q[3]), .B(DB[1326]), .Z(n25123) );
  IV U34749 ( .A(n25122), .Z(n34369) );
  XNOR U34750 ( .A(n25120), .B(n34371), .Z(n25122) );
  XNOR U34751 ( .A(q[2]), .B(DB[1325]), .Z(n34371) );
  XNOR U34752 ( .A(q[1]), .B(DB[1324]), .Z(n25120) );
  XOR U34753 ( .A(n34372), .B(n25085), .Z(n25048) );
  XOR U34754 ( .A(n34373), .B(n25073), .Z(n25085) );
  XNOR U34755 ( .A(q[6]), .B(DB[1336]), .Z(n25073) );
  IV U34756 ( .A(n25072), .Z(n34373) );
  XNOR U34757 ( .A(n25070), .B(n34374), .Z(n25072) );
  XNOR U34758 ( .A(q[5]), .B(DB[1335]), .Z(n34374) );
  XNOR U34759 ( .A(q[4]), .B(DB[1334]), .Z(n25070) );
  IV U34760 ( .A(n25084), .Z(n34372) );
  XOR U34761 ( .A(n34375), .B(n34376), .Z(n25084) );
  XNOR U34762 ( .A(n25080), .B(n25082), .Z(n34376) );
  XNOR U34763 ( .A(q[0]), .B(DB[1330]), .Z(n25082) );
  XNOR U34764 ( .A(q[3]), .B(DB[1333]), .Z(n25080) );
  IV U34765 ( .A(n25079), .Z(n34375) );
  XNOR U34766 ( .A(n25077), .B(n34377), .Z(n25079) );
  XNOR U34767 ( .A(q[2]), .B(DB[1332]), .Z(n34377) );
  XNOR U34768 ( .A(q[1]), .B(DB[1331]), .Z(n25077) );
  XOR U34769 ( .A(n34378), .B(n25042), .Z(n25005) );
  XOR U34770 ( .A(n34379), .B(n25030), .Z(n25042) );
  XNOR U34771 ( .A(q[6]), .B(DB[1343]), .Z(n25030) );
  IV U34772 ( .A(n25029), .Z(n34379) );
  XNOR U34773 ( .A(n25027), .B(n34380), .Z(n25029) );
  XNOR U34774 ( .A(q[5]), .B(DB[1342]), .Z(n34380) );
  XNOR U34775 ( .A(q[4]), .B(DB[1341]), .Z(n25027) );
  IV U34776 ( .A(n25041), .Z(n34378) );
  XOR U34777 ( .A(n34381), .B(n34382), .Z(n25041) );
  XNOR U34778 ( .A(n25037), .B(n25039), .Z(n34382) );
  XNOR U34779 ( .A(q[0]), .B(DB[1337]), .Z(n25039) );
  XNOR U34780 ( .A(q[3]), .B(DB[1340]), .Z(n25037) );
  IV U34781 ( .A(n25036), .Z(n34381) );
  XNOR U34782 ( .A(n25034), .B(n34383), .Z(n25036) );
  XNOR U34783 ( .A(q[2]), .B(DB[1339]), .Z(n34383) );
  XNOR U34784 ( .A(q[1]), .B(DB[1338]), .Z(n25034) );
  XOR U34785 ( .A(n34384), .B(n24999), .Z(n24962) );
  XOR U34786 ( .A(n34385), .B(n24987), .Z(n24999) );
  XNOR U34787 ( .A(q[6]), .B(DB[1350]), .Z(n24987) );
  IV U34788 ( .A(n24986), .Z(n34385) );
  XNOR U34789 ( .A(n24984), .B(n34386), .Z(n24986) );
  XNOR U34790 ( .A(q[5]), .B(DB[1349]), .Z(n34386) );
  XNOR U34791 ( .A(q[4]), .B(DB[1348]), .Z(n24984) );
  IV U34792 ( .A(n24998), .Z(n34384) );
  XOR U34793 ( .A(n34387), .B(n34388), .Z(n24998) );
  XNOR U34794 ( .A(n24994), .B(n24996), .Z(n34388) );
  XNOR U34795 ( .A(q[0]), .B(DB[1344]), .Z(n24996) );
  XNOR U34796 ( .A(q[3]), .B(DB[1347]), .Z(n24994) );
  IV U34797 ( .A(n24993), .Z(n34387) );
  XNOR U34798 ( .A(n24991), .B(n34389), .Z(n24993) );
  XNOR U34799 ( .A(q[2]), .B(DB[1346]), .Z(n34389) );
  XNOR U34800 ( .A(q[1]), .B(DB[1345]), .Z(n24991) );
  XOR U34801 ( .A(n34390), .B(n24956), .Z(n24919) );
  XOR U34802 ( .A(n34391), .B(n24944), .Z(n24956) );
  XNOR U34803 ( .A(q[6]), .B(DB[1357]), .Z(n24944) );
  IV U34804 ( .A(n24943), .Z(n34391) );
  XNOR U34805 ( .A(n24941), .B(n34392), .Z(n24943) );
  XNOR U34806 ( .A(q[5]), .B(DB[1356]), .Z(n34392) );
  XNOR U34807 ( .A(q[4]), .B(DB[1355]), .Z(n24941) );
  IV U34808 ( .A(n24955), .Z(n34390) );
  XOR U34809 ( .A(n34393), .B(n34394), .Z(n24955) );
  XNOR U34810 ( .A(n24951), .B(n24953), .Z(n34394) );
  XNOR U34811 ( .A(q[0]), .B(DB[1351]), .Z(n24953) );
  XNOR U34812 ( .A(q[3]), .B(DB[1354]), .Z(n24951) );
  IV U34813 ( .A(n24950), .Z(n34393) );
  XNOR U34814 ( .A(n24948), .B(n34395), .Z(n24950) );
  XNOR U34815 ( .A(q[2]), .B(DB[1353]), .Z(n34395) );
  XNOR U34816 ( .A(q[1]), .B(DB[1352]), .Z(n24948) );
  XOR U34817 ( .A(n34396), .B(n24913), .Z(n24876) );
  XOR U34818 ( .A(n34397), .B(n24901), .Z(n24913) );
  XNOR U34819 ( .A(q[6]), .B(DB[1364]), .Z(n24901) );
  IV U34820 ( .A(n24900), .Z(n34397) );
  XNOR U34821 ( .A(n24898), .B(n34398), .Z(n24900) );
  XNOR U34822 ( .A(q[5]), .B(DB[1363]), .Z(n34398) );
  XNOR U34823 ( .A(q[4]), .B(DB[1362]), .Z(n24898) );
  IV U34824 ( .A(n24912), .Z(n34396) );
  XOR U34825 ( .A(n34399), .B(n34400), .Z(n24912) );
  XNOR U34826 ( .A(n24908), .B(n24910), .Z(n34400) );
  XNOR U34827 ( .A(q[0]), .B(DB[1358]), .Z(n24910) );
  XNOR U34828 ( .A(q[3]), .B(DB[1361]), .Z(n24908) );
  IV U34829 ( .A(n24907), .Z(n34399) );
  XNOR U34830 ( .A(n24905), .B(n34401), .Z(n24907) );
  XNOR U34831 ( .A(q[2]), .B(DB[1360]), .Z(n34401) );
  XNOR U34832 ( .A(q[1]), .B(DB[1359]), .Z(n24905) );
  XOR U34833 ( .A(n34402), .B(n24870), .Z(n24833) );
  XOR U34834 ( .A(n34403), .B(n24858), .Z(n24870) );
  XNOR U34835 ( .A(q[6]), .B(DB[1371]), .Z(n24858) );
  IV U34836 ( .A(n24857), .Z(n34403) );
  XNOR U34837 ( .A(n24855), .B(n34404), .Z(n24857) );
  XNOR U34838 ( .A(q[5]), .B(DB[1370]), .Z(n34404) );
  XNOR U34839 ( .A(q[4]), .B(DB[1369]), .Z(n24855) );
  IV U34840 ( .A(n24869), .Z(n34402) );
  XOR U34841 ( .A(n34405), .B(n34406), .Z(n24869) );
  XNOR U34842 ( .A(n24865), .B(n24867), .Z(n34406) );
  XNOR U34843 ( .A(q[0]), .B(DB[1365]), .Z(n24867) );
  XNOR U34844 ( .A(q[3]), .B(DB[1368]), .Z(n24865) );
  IV U34845 ( .A(n24864), .Z(n34405) );
  XNOR U34846 ( .A(n24862), .B(n34407), .Z(n24864) );
  XNOR U34847 ( .A(q[2]), .B(DB[1367]), .Z(n34407) );
  XNOR U34848 ( .A(q[1]), .B(DB[1366]), .Z(n24862) );
  XOR U34849 ( .A(n34408), .B(n24827), .Z(n24790) );
  XOR U34850 ( .A(n34409), .B(n24815), .Z(n24827) );
  XNOR U34851 ( .A(q[6]), .B(DB[1378]), .Z(n24815) );
  IV U34852 ( .A(n24814), .Z(n34409) );
  XNOR U34853 ( .A(n24812), .B(n34410), .Z(n24814) );
  XNOR U34854 ( .A(q[5]), .B(DB[1377]), .Z(n34410) );
  XNOR U34855 ( .A(q[4]), .B(DB[1376]), .Z(n24812) );
  IV U34856 ( .A(n24826), .Z(n34408) );
  XOR U34857 ( .A(n34411), .B(n34412), .Z(n24826) );
  XNOR U34858 ( .A(n24822), .B(n24824), .Z(n34412) );
  XNOR U34859 ( .A(q[0]), .B(DB[1372]), .Z(n24824) );
  XNOR U34860 ( .A(q[3]), .B(DB[1375]), .Z(n24822) );
  IV U34861 ( .A(n24821), .Z(n34411) );
  XNOR U34862 ( .A(n24819), .B(n34413), .Z(n24821) );
  XNOR U34863 ( .A(q[2]), .B(DB[1374]), .Z(n34413) );
  XNOR U34864 ( .A(q[1]), .B(DB[1373]), .Z(n24819) );
  XOR U34865 ( .A(n34414), .B(n24784), .Z(n24747) );
  XOR U34866 ( .A(n34415), .B(n24772), .Z(n24784) );
  XNOR U34867 ( .A(q[6]), .B(DB[1385]), .Z(n24772) );
  IV U34868 ( .A(n24771), .Z(n34415) );
  XNOR U34869 ( .A(n24769), .B(n34416), .Z(n24771) );
  XNOR U34870 ( .A(q[5]), .B(DB[1384]), .Z(n34416) );
  XNOR U34871 ( .A(q[4]), .B(DB[1383]), .Z(n24769) );
  IV U34872 ( .A(n24783), .Z(n34414) );
  XOR U34873 ( .A(n34417), .B(n34418), .Z(n24783) );
  XNOR U34874 ( .A(n24779), .B(n24781), .Z(n34418) );
  XNOR U34875 ( .A(q[0]), .B(DB[1379]), .Z(n24781) );
  XNOR U34876 ( .A(q[3]), .B(DB[1382]), .Z(n24779) );
  IV U34877 ( .A(n24778), .Z(n34417) );
  XNOR U34878 ( .A(n24776), .B(n34419), .Z(n24778) );
  XNOR U34879 ( .A(q[2]), .B(DB[1381]), .Z(n34419) );
  XNOR U34880 ( .A(q[1]), .B(DB[1380]), .Z(n24776) );
  XOR U34881 ( .A(n34420), .B(n24741), .Z(n24704) );
  XOR U34882 ( .A(n34421), .B(n24729), .Z(n24741) );
  XNOR U34883 ( .A(q[6]), .B(DB[1392]), .Z(n24729) );
  IV U34884 ( .A(n24728), .Z(n34421) );
  XNOR U34885 ( .A(n24726), .B(n34422), .Z(n24728) );
  XNOR U34886 ( .A(q[5]), .B(DB[1391]), .Z(n34422) );
  XNOR U34887 ( .A(q[4]), .B(DB[1390]), .Z(n24726) );
  IV U34888 ( .A(n24740), .Z(n34420) );
  XOR U34889 ( .A(n34423), .B(n34424), .Z(n24740) );
  XNOR U34890 ( .A(n24736), .B(n24738), .Z(n34424) );
  XNOR U34891 ( .A(q[0]), .B(DB[1386]), .Z(n24738) );
  XNOR U34892 ( .A(q[3]), .B(DB[1389]), .Z(n24736) );
  IV U34893 ( .A(n24735), .Z(n34423) );
  XNOR U34894 ( .A(n24733), .B(n34425), .Z(n24735) );
  XNOR U34895 ( .A(q[2]), .B(DB[1388]), .Z(n34425) );
  XNOR U34896 ( .A(q[1]), .B(DB[1387]), .Z(n24733) );
  XOR U34897 ( .A(n34426), .B(n24698), .Z(n24661) );
  XOR U34898 ( .A(n34427), .B(n24686), .Z(n24698) );
  XNOR U34899 ( .A(q[6]), .B(DB[1399]), .Z(n24686) );
  IV U34900 ( .A(n24685), .Z(n34427) );
  XNOR U34901 ( .A(n24683), .B(n34428), .Z(n24685) );
  XNOR U34902 ( .A(q[5]), .B(DB[1398]), .Z(n34428) );
  XNOR U34903 ( .A(q[4]), .B(DB[1397]), .Z(n24683) );
  IV U34904 ( .A(n24697), .Z(n34426) );
  XOR U34905 ( .A(n34429), .B(n34430), .Z(n24697) );
  XNOR U34906 ( .A(n24693), .B(n24695), .Z(n34430) );
  XNOR U34907 ( .A(q[0]), .B(DB[1393]), .Z(n24695) );
  XNOR U34908 ( .A(q[3]), .B(DB[1396]), .Z(n24693) );
  IV U34909 ( .A(n24692), .Z(n34429) );
  XNOR U34910 ( .A(n24690), .B(n34431), .Z(n24692) );
  XNOR U34911 ( .A(q[2]), .B(DB[1395]), .Z(n34431) );
  XNOR U34912 ( .A(q[1]), .B(DB[1394]), .Z(n24690) );
  XOR U34913 ( .A(n34432), .B(n24655), .Z(n24618) );
  XOR U34914 ( .A(n34433), .B(n24643), .Z(n24655) );
  XNOR U34915 ( .A(q[6]), .B(DB[1406]), .Z(n24643) );
  IV U34916 ( .A(n24642), .Z(n34433) );
  XNOR U34917 ( .A(n24640), .B(n34434), .Z(n24642) );
  XNOR U34918 ( .A(q[5]), .B(DB[1405]), .Z(n34434) );
  XNOR U34919 ( .A(q[4]), .B(DB[1404]), .Z(n24640) );
  IV U34920 ( .A(n24654), .Z(n34432) );
  XOR U34921 ( .A(n34435), .B(n34436), .Z(n24654) );
  XNOR U34922 ( .A(n24650), .B(n24652), .Z(n34436) );
  XNOR U34923 ( .A(q[0]), .B(DB[1400]), .Z(n24652) );
  XNOR U34924 ( .A(q[3]), .B(DB[1403]), .Z(n24650) );
  IV U34925 ( .A(n24649), .Z(n34435) );
  XNOR U34926 ( .A(n24647), .B(n34437), .Z(n24649) );
  XNOR U34927 ( .A(q[2]), .B(DB[1402]), .Z(n34437) );
  XNOR U34928 ( .A(q[1]), .B(DB[1401]), .Z(n24647) );
  XOR U34929 ( .A(n34438), .B(n24612), .Z(n24575) );
  XOR U34930 ( .A(n34439), .B(n24600), .Z(n24612) );
  XNOR U34931 ( .A(q[6]), .B(DB[1413]), .Z(n24600) );
  IV U34932 ( .A(n24599), .Z(n34439) );
  XNOR U34933 ( .A(n24597), .B(n34440), .Z(n24599) );
  XNOR U34934 ( .A(q[5]), .B(DB[1412]), .Z(n34440) );
  XNOR U34935 ( .A(q[4]), .B(DB[1411]), .Z(n24597) );
  IV U34936 ( .A(n24611), .Z(n34438) );
  XOR U34937 ( .A(n34441), .B(n34442), .Z(n24611) );
  XNOR U34938 ( .A(n24607), .B(n24609), .Z(n34442) );
  XNOR U34939 ( .A(q[0]), .B(DB[1407]), .Z(n24609) );
  XNOR U34940 ( .A(q[3]), .B(DB[1410]), .Z(n24607) );
  IV U34941 ( .A(n24606), .Z(n34441) );
  XNOR U34942 ( .A(n24604), .B(n34443), .Z(n24606) );
  XNOR U34943 ( .A(q[2]), .B(DB[1409]), .Z(n34443) );
  XNOR U34944 ( .A(q[1]), .B(DB[1408]), .Z(n24604) );
  XOR U34945 ( .A(n34444), .B(n24569), .Z(n24532) );
  XOR U34946 ( .A(n34445), .B(n24557), .Z(n24569) );
  XNOR U34947 ( .A(q[6]), .B(DB[1420]), .Z(n24557) );
  IV U34948 ( .A(n24556), .Z(n34445) );
  XNOR U34949 ( .A(n24554), .B(n34446), .Z(n24556) );
  XNOR U34950 ( .A(q[5]), .B(DB[1419]), .Z(n34446) );
  XNOR U34951 ( .A(q[4]), .B(DB[1418]), .Z(n24554) );
  IV U34952 ( .A(n24568), .Z(n34444) );
  XOR U34953 ( .A(n34447), .B(n34448), .Z(n24568) );
  XNOR U34954 ( .A(n24564), .B(n24566), .Z(n34448) );
  XNOR U34955 ( .A(q[0]), .B(DB[1414]), .Z(n24566) );
  XNOR U34956 ( .A(q[3]), .B(DB[1417]), .Z(n24564) );
  IV U34957 ( .A(n24563), .Z(n34447) );
  XNOR U34958 ( .A(n24561), .B(n34449), .Z(n24563) );
  XNOR U34959 ( .A(q[2]), .B(DB[1416]), .Z(n34449) );
  XNOR U34960 ( .A(q[1]), .B(DB[1415]), .Z(n24561) );
  XOR U34961 ( .A(n34450), .B(n24526), .Z(n24489) );
  XOR U34962 ( .A(n34451), .B(n24514), .Z(n24526) );
  XNOR U34963 ( .A(q[6]), .B(DB[1427]), .Z(n24514) );
  IV U34964 ( .A(n24513), .Z(n34451) );
  XNOR U34965 ( .A(n24511), .B(n34452), .Z(n24513) );
  XNOR U34966 ( .A(q[5]), .B(DB[1426]), .Z(n34452) );
  XNOR U34967 ( .A(q[4]), .B(DB[1425]), .Z(n24511) );
  IV U34968 ( .A(n24525), .Z(n34450) );
  XOR U34969 ( .A(n34453), .B(n34454), .Z(n24525) );
  XNOR U34970 ( .A(n24521), .B(n24523), .Z(n34454) );
  XNOR U34971 ( .A(q[0]), .B(DB[1421]), .Z(n24523) );
  XNOR U34972 ( .A(q[3]), .B(DB[1424]), .Z(n24521) );
  IV U34973 ( .A(n24520), .Z(n34453) );
  XNOR U34974 ( .A(n24518), .B(n34455), .Z(n24520) );
  XNOR U34975 ( .A(q[2]), .B(DB[1423]), .Z(n34455) );
  XNOR U34976 ( .A(q[1]), .B(DB[1422]), .Z(n24518) );
  XOR U34977 ( .A(n34456), .B(n24483), .Z(n24446) );
  XOR U34978 ( .A(n34457), .B(n24471), .Z(n24483) );
  XNOR U34979 ( .A(q[6]), .B(DB[1434]), .Z(n24471) );
  IV U34980 ( .A(n24470), .Z(n34457) );
  XNOR U34981 ( .A(n24468), .B(n34458), .Z(n24470) );
  XNOR U34982 ( .A(q[5]), .B(DB[1433]), .Z(n34458) );
  XNOR U34983 ( .A(q[4]), .B(DB[1432]), .Z(n24468) );
  IV U34984 ( .A(n24482), .Z(n34456) );
  XOR U34985 ( .A(n34459), .B(n34460), .Z(n24482) );
  XNOR U34986 ( .A(n24478), .B(n24480), .Z(n34460) );
  XNOR U34987 ( .A(q[0]), .B(DB[1428]), .Z(n24480) );
  XNOR U34988 ( .A(q[3]), .B(DB[1431]), .Z(n24478) );
  IV U34989 ( .A(n24477), .Z(n34459) );
  XNOR U34990 ( .A(n24475), .B(n34461), .Z(n24477) );
  XNOR U34991 ( .A(q[2]), .B(DB[1430]), .Z(n34461) );
  XNOR U34992 ( .A(q[1]), .B(DB[1429]), .Z(n24475) );
  XOR U34993 ( .A(n34462), .B(n24440), .Z(n24403) );
  XOR U34994 ( .A(n34463), .B(n24428), .Z(n24440) );
  XNOR U34995 ( .A(q[6]), .B(DB[1441]), .Z(n24428) );
  IV U34996 ( .A(n24427), .Z(n34463) );
  XNOR U34997 ( .A(n24425), .B(n34464), .Z(n24427) );
  XNOR U34998 ( .A(q[5]), .B(DB[1440]), .Z(n34464) );
  XNOR U34999 ( .A(q[4]), .B(DB[1439]), .Z(n24425) );
  IV U35000 ( .A(n24439), .Z(n34462) );
  XOR U35001 ( .A(n34465), .B(n34466), .Z(n24439) );
  XNOR U35002 ( .A(n24435), .B(n24437), .Z(n34466) );
  XNOR U35003 ( .A(q[0]), .B(DB[1435]), .Z(n24437) );
  XNOR U35004 ( .A(q[3]), .B(DB[1438]), .Z(n24435) );
  IV U35005 ( .A(n24434), .Z(n34465) );
  XNOR U35006 ( .A(n24432), .B(n34467), .Z(n24434) );
  XNOR U35007 ( .A(q[2]), .B(DB[1437]), .Z(n34467) );
  XNOR U35008 ( .A(q[1]), .B(DB[1436]), .Z(n24432) );
  XOR U35009 ( .A(n34468), .B(n24397), .Z(n24360) );
  XOR U35010 ( .A(n34469), .B(n24385), .Z(n24397) );
  XNOR U35011 ( .A(q[6]), .B(DB[1448]), .Z(n24385) );
  IV U35012 ( .A(n24384), .Z(n34469) );
  XNOR U35013 ( .A(n24382), .B(n34470), .Z(n24384) );
  XNOR U35014 ( .A(q[5]), .B(DB[1447]), .Z(n34470) );
  XNOR U35015 ( .A(q[4]), .B(DB[1446]), .Z(n24382) );
  IV U35016 ( .A(n24396), .Z(n34468) );
  XOR U35017 ( .A(n34471), .B(n34472), .Z(n24396) );
  XNOR U35018 ( .A(n24392), .B(n24394), .Z(n34472) );
  XNOR U35019 ( .A(q[0]), .B(DB[1442]), .Z(n24394) );
  XNOR U35020 ( .A(q[3]), .B(DB[1445]), .Z(n24392) );
  IV U35021 ( .A(n24391), .Z(n34471) );
  XNOR U35022 ( .A(n24389), .B(n34473), .Z(n24391) );
  XNOR U35023 ( .A(q[2]), .B(DB[1444]), .Z(n34473) );
  XNOR U35024 ( .A(q[1]), .B(DB[1443]), .Z(n24389) );
  XOR U35025 ( .A(n34474), .B(n24354), .Z(n24317) );
  XOR U35026 ( .A(n34475), .B(n24342), .Z(n24354) );
  XNOR U35027 ( .A(q[6]), .B(DB[1455]), .Z(n24342) );
  IV U35028 ( .A(n24341), .Z(n34475) );
  XNOR U35029 ( .A(n24339), .B(n34476), .Z(n24341) );
  XNOR U35030 ( .A(q[5]), .B(DB[1454]), .Z(n34476) );
  XNOR U35031 ( .A(q[4]), .B(DB[1453]), .Z(n24339) );
  IV U35032 ( .A(n24353), .Z(n34474) );
  XOR U35033 ( .A(n34477), .B(n34478), .Z(n24353) );
  XNOR U35034 ( .A(n24349), .B(n24351), .Z(n34478) );
  XNOR U35035 ( .A(q[0]), .B(DB[1449]), .Z(n24351) );
  XNOR U35036 ( .A(q[3]), .B(DB[1452]), .Z(n24349) );
  IV U35037 ( .A(n24348), .Z(n34477) );
  XNOR U35038 ( .A(n24346), .B(n34479), .Z(n24348) );
  XNOR U35039 ( .A(q[2]), .B(DB[1451]), .Z(n34479) );
  XNOR U35040 ( .A(q[1]), .B(DB[1450]), .Z(n24346) );
  XOR U35041 ( .A(n34480), .B(n24311), .Z(n24274) );
  XOR U35042 ( .A(n34481), .B(n24299), .Z(n24311) );
  XNOR U35043 ( .A(q[6]), .B(DB[1462]), .Z(n24299) );
  IV U35044 ( .A(n24298), .Z(n34481) );
  XNOR U35045 ( .A(n24296), .B(n34482), .Z(n24298) );
  XNOR U35046 ( .A(q[5]), .B(DB[1461]), .Z(n34482) );
  XNOR U35047 ( .A(q[4]), .B(DB[1460]), .Z(n24296) );
  IV U35048 ( .A(n24310), .Z(n34480) );
  XOR U35049 ( .A(n34483), .B(n34484), .Z(n24310) );
  XNOR U35050 ( .A(n24306), .B(n24308), .Z(n34484) );
  XNOR U35051 ( .A(q[0]), .B(DB[1456]), .Z(n24308) );
  XNOR U35052 ( .A(q[3]), .B(DB[1459]), .Z(n24306) );
  IV U35053 ( .A(n24305), .Z(n34483) );
  XNOR U35054 ( .A(n24303), .B(n34485), .Z(n24305) );
  XNOR U35055 ( .A(q[2]), .B(DB[1458]), .Z(n34485) );
  XNOR U35056 ( .A(q[1]), .B(DB[1457]), .Z(n24303) );
  XOR U35057 ( .A(n34486), .B(n24268), .Z(n24231) );
  XOR U35058 ( .A(n34487), .B(n24256), .Z(n24268) );
  XNOR U35059 ( .A(q[6]), .B(DB[1469]), .Z(n24256) );
  IV U35060 ( .A(n24255), .Z(n34487) );
  XNOR U35061 ( .A(n24253), .B(n34488), .Z(n24255) );
  XNOR U35062 ( .A(q[5]), .B(DB[1468]), .Z(n34488) );
  XNOR U35063 ( .A(q[4]), .B(DB[1467]), .Z(n24253) );
  IV U35064 ( .A(n24267), .Z(n34486) );
  XOR U35065 ( .A(n34489), .B(n34490), .Z(n24267) );
  XNOR U35066 ( .A(n24263), .B(n24265), .Z(n34490) );
  XNOR U35067 ( .A(q[0]), .B(DB[1463]), .Z(n24265) );
  XNOR U35068 ( .A(q[3]), .B(DB[1466]), .Z(n24263) );
  IV U35069 ( .A(n24262), .Z(n34489) );
  XNOR U35070 ( .A(n24260), .B(n34491), .Z(n24262) );
  XNOR U35071 ( .A(q[2]), .B(DB[1465]), .Z(n34491) );
  XNOR U35072 ( .A(q[1]), .B(DB[1464]), .Z(n24260) );
  XOR U35073 ( .A(n34492), .B(n24225), .Z(n24188) );
  XOR U35074 ( .A(n34493), .B(n24213), .Z(n24225) );
  XNOR U35075 ( .A(q[6]), .B(DB[1476]), .Z(n24213) );
  IV U35076 ( .A(n24212), .Z(n34493) );
  XNOR U35077 ( .A(n24210), .B(n34494), .Z(n24212) );
  XNOR U35078 ( .A(q[5]), .B(DB[1475]), .Z(n34494) );
  XNOR U35079 ( .A(q[4]), .B(DB[1474]), .Z(n24210) );
  IV U35080 ( .A(n24224), .Z(n34492) );
  XOR U35081 ( .A(n34495), .B(n34496), .Z(n24224) );
  XNOR U35082 ( .A(n24220), .B(n24222), .Z(n34496) );
  XNOR U35083 ( .A(q[0]), .B(DB[1470]), .Z(n24222) );
  XNOR U35084 ( .A(q[3]), .B(DB[1473]), .Z(n24220) );
  IV U35085 ( .A(n24219), .Z(n34495) );
  XNOR U35086 ( .A(n24217), .B(n34497), .Z(n24219) );
  XNOR U35087 ( .A(q[2]), .B(DB[1472]), .Z(n34497) );
  XNOR U35088 ( .A(q[1]), .B(DB[1471]), .Z(n24217) );
  XOR U35089 ( .A(n34498), .B(n24182), .Z(n24145) );
  XOR U35090 ( .A(n34499), .B(n24170), .Z(n24182) );
  XNOR U35091 ( .A(q[6]), .B(DB[1483]), .Z(n24170) );
  IV U35092 ( .A(n24169), .Z(n34499) );
  XNOR U35093 ( .A(n24167), .B(n34500), .Z(n24169) );
  XNOR U35094 ( .A(q[5]), .B(DB[1482]), .Z(n34500) );
  XNOR U35095 ( .A(q[4]), .B(DB[1481]), .Z(n24167) );
  IV U35096 ( .A(n24181), .Z(n34498) );
  XOR U35097 ( .A(n34501), .B(n34502), .Z(n24181) );
  XNOR U35098 ( .A(n24177), .B(n24179), .Z(n34502) );
  XNOR U35099 ( .A(q[0]), .B(DB[1477]), .Z(n24179) );
  XNOR U35100 ( .A(q[3]), .B(DB[1480]), .Z(n24177) );
  IV U35101 ( .A(n24176), .Z(n34501) );
  XNOR U35102 ( .A(n24174), .B(n34503), .Z(n24176) );
  XNOR U35103 ( .A(q[2]), .B(DB[1479]), .Z(n34503) );
  XNOR U35104 ( .A(q[1]), .B(DB[1478]), .Z(n24174) );
  XOR U35105 ( .A(n34504), .B(n24139), .Z(n24102) );
  XOR U35106 ( .A(n34505), .B(n24127), .Z(n24139) );
  XNOR U35107 ( .A(q[6]), .B(DB[1490]), .Z(n24127) );
  IV U35108 ( .A(n24126), .Z(n34505) );
  XNOR U35109 ( .A(n24124), .B(n34506), .Z(n24126) );
  XNOR U35110 ( .A(q[5]), .B(DB[1489]), .Z(n34506) );
  XNOR U35111 ( .A(q[4]), .B(DB[1488]), .Z(n24124) );
  IV U35112 ( .A(n24138), .Z(n34504) );
  XOR U35113 ( .A(n34507), .B(n34508), .Z(n24138) );
  XNOR U35114 ( .A(n24134), .B(n24136), .Z(n34508) );
  XNOR U35115 ( .A(q[0]), .B(DB[1484]), .Z(n24136) );
  XNOR U35116 ( .A(q[3]), .B(DB[1487]), .Z(n24134) );
  IV U35117 ( .A(n24133), .Z(n34507) );
  XNOR U35118 ( .A(n24131), .B(n34509), .Z(n24133) );
  XNOR U35119 ( .A(q[2]), .B(DB[1486]), .Z(n34509) );
  XNOR U35120 ( .A(q[1]), .B(DB[1485]), .Z(n24131) );
  XOR U35121 ( .A(n34510), .B(n24096), .Z(n24059) );
  XOR U35122 ( .A(n34511), .B(n24084), .Z(n24096) );
  XNOR U35123 ( .A(q[6]), .B(DB[1497]), .Z(n24084) );
  IV U35124 ( .A(n24083), .Z(n34511) );
  XNOR U35125 ( .A(n24081), .B(n34512), .Z(n24083) );
  XNOR U35126 ( .A(q[5]), .B(DB[1496]), .Z(n34512) );
  XNOR U35127 ( .A(q[4]), .B(DB[1495]), .Z(n24081) );
  IV U35128 ( .A(n24095), .Z(n34510) );
  XOR U35129 ( .A(n34513), .B(n34514), .Z(n24095) );
  XNOR U35130 ( .A(n24091), .B(n24093), .Z(n34514) );
  XNOR U35131 ( .A(q[0]), .B(DB[1491]), .Z(n24093) );
  XNOR U35132 ( .A(q[3]), .B(DB[1494]), .Z(n24091) );
  IV U35133 ( .A(n24090), .Z(n34513) );
  XNOR U35134 ( .A(n24088), .B(n34515), .Z(n24090) );
  XNOR U35135 ( .A(q[2]), .B(DB[1493]), .Z(n34515) );
  XNOR U35136 ( .A(q[1]), .B(DB[1492]), .Z(n24088) );
  XOR U35137 ( .A(n34516), .B(n24053), .Z(n24016) );
  XOR U35138 ( .A(n34517), .B(n24041), .Z(n24053) );
  XNOR U35139 ( .A(q[6]), .B(DB[1504]), .Z(n24041) );
  IV U35140 ( .A(n24040), .Z(n34517) );
  XNOR U35141 ( .A(n24038), .B(n34518), .Z(n24040) );
  XNOR U35142 ( .A(q[5]), .B(DB[1503]), .Z(n34518) );
  XNOR U35143 ( .A(q[4]), .B(DB[1502]), .Z(n24038) );
  IV U35144 ( .A(n24052), .Z(n34516) );
  XOR U35145 ( .A(n34519), .B(n34520), .Z(n24052) );
  XNOR U35146 ( .A(n24048), .B(n24050), .Z(n34520) );
  XNOR U35147 ( .A(q[0]), .B(DB[1498]), .Z(n24050) );
  XNOR U35148 ( .A(q[3]), .B(DB[1501]), .Z(n24048) );
  IV U35149 ( .A(n24047), .Z(n34519) );
  XNOR U35150 ( .A(n24045), .B(n34521), .Z(n24047) );
  XNOR U35151 ( .A(q[2]), .B(DB[1500]), .Z(n34521) );
  XNOR U35152 ( .A(q[1]), .B(DB[1499]), .Z(n24045) );
  XOR U35153 ( .A(n34522), .B(n24010), .Z(n23973) );
  XOR U35154 ( .A(n34523), .B(n23998), .Z(n24010) );
  XNOR U35155 ( .A(q[6]), .B(DB[1511]), .Z(n23998) );
  IV U35156 ( .A(n23997), .Z(n34523) );
  XNOR U35157 ( .A(n23995), .B(n34524), .Z(n23997) );
  XNOR U35158 ( .A(q[5]), .B(DB[1510]), .Z(n34524) );
  XNOR U35159 ( .A(q[4]), .B(DB[1509]), .Z(n23995) );
  IV U35160 ( .A(n24009), .Z(n34522) );
  XOR U35161 ( .A(n34525), .B(n34526), .Z(n24009) );
  XNOR U35162 ( .A(n24005), .B(n24007), .Z(n34526) );
  XNOR U35163 ( .A(q[0]), .B(DB[1505]), .Z(n24007) );
  XNOR U35164 ( .A(q[3]), .B(DB[1508]), .Z(n24005) );
  IV U35165 ( .A(n24004), .Z(n34525) );
  XNOR U35166 ( .A(n24002), .B(n34527), .Z(n24004) );
  XNOR U35167 ( .A(q[2]), .B(DB[1507]), .Z(n34527) );
  XNOR U35168 ( .A(q[1]), .B(DB[1506]), .Z(n24002) );
  XOR U35169 ( .A(n34528), .B(n23967), .Z(n23930) );
  XOR U35170 ( .A(n34529), .B(n23955), .Z(n23967) );
  XNOR U35171 ( .A(q[6]), .B(DB[1518]), .Z(n23955) );
  IV U35172 ( .A(n23954), .Z(n34529) );
  XNOR U35173 ( .A(n23952), .B(n34530), .Z(n23954) );
  XNOR U35174 ( .A(q[5]), .B(DB[1517]), .Z(n34530) );
  XNOR U35175 ( .A(q[4]), .B(DB[1516]), .Z(n23952) );
  IV U35176 ( .A(n23966), .Z(n34528) );
  XOR U35177 ( .A(n34531), .B(n34532), .Z(n23966) );
  XNOR U35178 ( .A(n23962), .B(n23964), .Z(n34532) );
  XNOR U35179 ( .A(q[0]), .B(DB[1512]), .Z(n23964) );
  XNOR U35180 ( .A(q[3]), .B(DB[1515]), .Z(n23962) );
  IV U35181 ( .A(n23961), .Z(n34531) );
  XNOR U35182 ( .A(n23959), .B(n34533), .Z(n23961) );
  XNOR U35183 ( .A(q[2]), .B(DB[1514]), .Z(n34533) );
  XNOR U35184 ( .A(q[1]), .B(DB[1513]), .Z(n23959) );
  XOR U35185 ( .A(n34534), .B(n23924), .Z(n23887) );
  XOR U35186 ( .A(n34535), .B(n23912), .Z(n23924) );
  XNOR U35187 ( .A(q[6]), .B(DB[1525]), .Z(n23912) );
  IV U35188 ( .A(n23911), .Z(n34535) );
  XNOR U35189 ( .A(n23909), .B(n34536), .Z(n23911) );
  XNOR U35190 ( .A(q[5]), .B(DB[1524]), .Z(n34536) );
  XNOR U35191 ( .A(q[4]), .B(DB[1523]), .Z(n23909) );
  IV U35192 ( .A(n23923), .Z(n34534) );
  XOR U35193 ( .A(n34537), .B(n34538), .Z(n23923) );
  XNOR U35194 ( .A(n23919), .B(n23921), .Z(n34538) );
  XNOR U35195 ( .A(q[0]), .B(DB[1519]), .Z(n23921) );
  XNOR U35196 ( .A(q[3]), .B(DB[1522]), .Z(n23919) );
  IV U35197 ( .A(n23918), .Z(n34537) );
  XNOR U35198 ( .A(n23916), .B(n34539), .Z(n23918) );
  XNOR U35199 ( .A(q[2]), .B(DB[1521]), .Z(n34539) );
  XNOR U35200 ( .A(q[1]), .B(DB[1520]), .Z(n23916) );
  XOR U35201 ( .A(n34540), .B(n23881), .Z(n23844) );
  XOR U35202 ( .A(n34541), .B(n23869), .Z(n23881) );
  XNOR U35203 ( .A(q[6]), .B(DB[1532]), .Z(n23869) );
  IV U35204 ( .A(n23868), .Z(n34541) );
  XNOR U35205 ( .A(n23866), .B(n34542), .Z(n23868) );
  XNOR U35206 ( .A(q[5]), .B(DB[1531]), .Z(n34542) );
  XNOR U35207 ( .A(q[4]), .B(DB[1530]), .Z(n23866) );
  IV U35208 ( .A(n23880), .Z(n34540) );
  XOR U35209 ( .A(n34543), .B(n34544), .Z(n23880) );
  XNOR U35210 ( .A(n23876), .B(n23878), .Z(n34544) );
  XNOR U35211 ( .A(q[0]), .B(DB[1526]), .Z(n23878) );
  XNOR U35212 ( .A(q[3]), .B(DB[1529]), .Z(n23876) );
  IV U35213 ( .A(n23875), .Z(n34543) );
  XNOR U35214 ( .A(n23873), .B(n34545), .Z(n23875) );
  XNOR U35215 ( .A(q[2]), .B(DB[1528]), .Z(n34545) );
  XNOR U35216 ( .A(q[1]), .B(DB[1527]), .Z(n23873) );
  XOR U35217 ( .A(n34546), .B(n23838), .Z(n23801) );
  XOR U35218 ( .A(n34547), .B(n23826), .Z(n23838) );
  XNOR U35219 ( .A(q[6]), .B(DB[1539]), .Z(n23826) );
  IV U35220 ( .A(n23825), .Z(n34547) );
  XNOR U35221 ( .A(n23823), .B(n34548), .Z(n23825) );
  XNOR U35222 ( .A(q[5]), .B(DB[1538]), .Z(n34548) );
  XNOR U35223 ( .A(q[4]), .B(DB[1537]), .Z(n23823) );
  IV U35224 ( .A(n23837), .Z(n34546) );
  XOR U35225 ( .A(n34549), .B(n34550), .Z(n23837) );
  XNOR U35226 ( .A(n23833), .B(n23835), .Z(n34550) );
  XNOR U35227 ( .A(q[0]), .B(DB[1533]), .Z(n23835) );
  XNOR U35228 ( .A(q[3]), .B(DB[1536]), .Z(n23833) );
  IV U35229 ( .A(n23832), .Z(n34549) );
  XNOR U35230 ( .A(n23830), .B(n34551), .Z(n23832) );
  XNOR U35231 ( .A(q[2]), .B(DB[1535]), .Z(n34551) );
  XNOR U35232 ( .A(q[1]), .B(DB[1534]), .Z(n23830) );
  XOR U35233 ( .A(n34552), .B(n23795), .Z(n23758) );
  XOR U35234 ( .A(n34553), .B(n23783), .Z(n23795) );
  XNOR U35235 ( .A(q[6]), .B(DB[1546]), .Z(n23783) );
  IV U35236 ( .A(n23782), .Z(n34553) );
  XNOR U35237 ( .A(n23780), .B(n34554), .Z(n23782) );
  XNOR U35238 ( .A(q[5]), .B(DB[1545]), .Z(n34554) );
  XNOR U35239 ( .A(q[4]), .B(DB[1544]), .Z(n23780) );
  IV U35240 ( .A(n23794), .Z(n34552) );
  XOR U35241 ( .A(n34555), .B(n34556), .Z(n23794) );
  XNOR U35242 ( .A(n23790), .B(n23792), .Z(n34556) );
  XNOR U35243 ( .A(q[0]), .B(DB[1540]), .Z(n23792) );
  XNOR U35244 ( .A(q[3]), .B(DB[1543]), .Z(n23790) );
  IV U35245 ( .A(n23789), .Z(n34555) );
  XNOR U35246 ( .A(n23787), .B(n34557), .Z(n23789) );
  XNOR U35247 ( .A(q[2]), .B(DB[1542]), .Z(n34557) );
  XNOR U35248 ( .A(q[1]), .B(DB[1541]), .Z(n23787) );
  XOR U35249 ( .A(n34558), .B(n23752), .Z(n23715) );
  XOR U35250 ( .A(n34559), .B(n23740), .Z(n23752) );
  XNOR U35251 ( .A(q[6]), .B(DB[1553]), .Z(n23740) );
  IV U35252 ( .A(n23739), .Z(n34559) );
  XNOR U35253 ( .A(n23737), .B(n34560), .Z(n23739) );
  XNOR U35254 ( .A(q[5]), .B(DB[1552]), .Z(n34560) );
  XNOR U35255 ( .A(q[4]), .B(DB[1551]), .Z(n23737) );
  IV U35256 ( .A(n23751), .Z(n34558) );
  XOR U35257 ( .A(n34561), .B(n34562), .Z(n23751) );
  XNOR U35258 ( .A(n23747), .B(n23749), .Z(n34562) );
  XNOR U35259 ( .A(q[0]), .B(DB[1547]), .Z(n23749) );
  XNOR U35260 ( .A(q[3]), .B(DB[1550]), .Z(n23747) );
  IV U35261 ( .A(n23746), .Z(n34561) );
  XNOR U35262 ( .A(n23744), .B(n34563), .Z(n23746) );
  XNOR U35263 ( .A(q[2]), .B(DB[1549]), .Z(n34563) );
  XNOR U35264 ( .A(q[1]), .B(DB[1548]), .Z(n23744) );
  XOR U35265 ( .A(n34564), .B(n23709), .Z(n23672) );
  XOR U35266 ( .A(n34565), .B(n23697), .Z(n23709) );
  XNOR U35267 ( .A(q[6]), .B(DB[1560]), .Z(n23697) );
  IV U35268 ( .A(n23696), .Z(n34565) );
  XNOR U35269 ( .A(n23694), .B(n34566), .Z(n23696) );
  XNOR U35270 ( .A(q[5]), .B(DB[1559]), .Z(n34566) );
  XNOR U35271 ( .A(q[4]), .B(DB[1558]), .Z(n23694) );
  IV U35272 ( .A(n23708), .Z(n34564) );
  XOR U35273 ( .A(n34567), .B(n34568), .Z(n23708) );
  XNOR U35274 ( .A(n23704), .B(n23706), .Z(n34568) );
  XNOR U35275 ( .A(q[0]), .B(DB[1554]), .Z(n23706) );
  XNOR U35276 ( .A(q[3]), .B(DB[1557]), .Z(n23704) );
  IV U35277 ( .A(n23703), .Z(n34567) );
  XNOR U35278 ( .A(n23701), .B(n34569), .Z(n23703) );
  XNOR U35279 ( .A(q[2]), .B(DB[1556]), .Z(n34569) );
  XNOR U35280 ( .A(q[1]), .B(DB[1555]), .Z(n23701) );
  XOR U35281 ( .A(n34570), .B(n23666), .Z(n23629) );
  XOR U35282 ( .A(n34571), .B(n23654), .Z(n23666) );
  XNOR U35283 ( .A(q[6]), .B(DB[1567]), .Z(n23654) );
  IV U35284 ( .A(n23653), .Z(n34571) );
  XNOR U35285 ( .A(n23651), .B(n34572), .Z(n23653) );
  XNOR U35286 ( .A(q[5]), .B(DB[1566]), .Z(n34572) );
  XNOR U35287 ( .A(q[4]), .B(DB[1565]), .Z(n23651) );
  IV U35288 ( .A(n23665), .Z(n34570) );
  XOR U35289 ( .A(n34573), .B(n34574), .Z(n23665) );
  XNOR U35290 ( .A(n23661), .B(n23663), .Z(n34574) );
  XNOR U35291 ( .A(q[0]), .B(DB[1561]), .Z(n23663) );
  XNOR U35292 ( .A(q[3]), .B(DB[1564]), .Z(n23661) );
  IV U35293 ( .A(n23660), .Z(n34573) );
  XNOR U35294 ( .A(n23658), .B(n34575), .Z(n23660) );
  XNOR U35295 ( .A(q[2]), .B(DB[1563]), .Z(n34575) );
  XNOR U35296 ( .A(q[1]), .B(DB[1562]), .Z(n23658) );
  XOR U35297 ( .A(n34576), .B(n23623), .Z(n23586) );
  XOR U35298 ( .A(n34577), .B(n23611), .Z(n23623) );
  XNOR U35299 ( .A(q[6]), .B(DB[1574]), .Z(n23611) );
  IV U35300 ( .A(n23610), .Z(n34577) );
  XNOR U35301 ( .A(n23608), .B(n34578), .Z(n23610) );
  XNOR U35302 ( .A(q[5]), .B(DB[1573]), .Z(n34578) );
  XNOR U35303 ( .A(q[4]), .B(DB[1572]), .Z(n23608) );
  IV U35304 ( .A(n23622), .Z(n34576) );
  XOR U35305 ( .A(n34579), .B(n34580), .Z(n23622) );
  XNOR U35306 ( .A(n23618), .B(n23620), .Z(n34580) );
  XNOR U35307 ( .A(q[0]), .B(DB[1568]), .Z(n23620) );
  XNOR U35308 ( .A(q[3]), .B(DB[1571]), .Z(n23618) );
  IV U35309 ( .A(n23617), .Z(n34579) );
  XNOR U35310 ( .A(n23615), .B(n34581), .Z(n23617) );
  XNOR U35311 ( .A(q[2]), .B(DB[1570]), .Z(n34581) );
  XNOR U35312 ( .A(q[1]), .B(DB[1569]), .Z(n23615) );
  XOR U35313 ( .A(n34582), .B(n23580), .Z(n23543) );
  XOR U35314 ( .A(n34583), .B(n23568), .Z(n23580) );
  XNOR U35315 ( .A(q[6]), .B(DB[1581]), .Z(n23568) );
  IV U35316 ( .A(n23567), .Z(n34583) );
  XNOR U35317 ( .A(n23565), .B(n34584), .Z(n23567) );
  XNOR U35318 ( .A(q[5]), .B(DB[1580]), .Z(n34584) );
  XNOR U35319 ( .A(q[4]), .B(DB[1579]), .Z(n23565) );
  IV U35320 ( .A(n23579), .Z(n34582) );
  XOR U35321 ( .A(n34585), .B(n34586), .Z(n23579) );
  XNOR U35322 ( .A(n23575), .B(n23577), .Z(n34586) );
  XNOR U35323 ( .A(q[0]), .B(DB[1575]), .Z(n23577) );
  XNOR U35324 ( .A(q[3]), .B(DB[1578]), .Z(n23575) );
  IV U35325 ( .A(n23574), .Z(n34585) );
  XNOR U35326 ( .A(n23572), .B(n34587), .Z(n23574) );
  XNOR U35327 ( .A(q[2]), .B(DB[1577]), .Z(n34587) );
  XNOR U35328 ( .A(q[1]), .B(DB[1576]), .Z(n23572) );
  XOR U35329 ( .A(n34588), .B(n23537), .Z(n23500) );
  XOR U35330 ( .A(n34589), .B(n23525), .Z(n23537) );
  XNOR U35331 ( .A(q[6]), .B(DB[1588]), .Z(n23525) );
  IV U35332 ( .A(n23524), .Z(n34589) );
  XNOR U35333 ( .A(n23522), .B(n34590), .Z(n23524) );
  XNOR U35334 ( .A(q[5]), .B(DB[1587]), .Z(n34590) );
  XNOR U35335 ( .A(q[4]), .B(DB[1586]), .Z(n23522) );
  IV U35336 ( .A(n23536), .Z(n34588) );
  XOR U35337 ( .A(n34591), .B(n34592), .Z(n23536) );
  XNOR U35338 ( .A(n23532), .B(n23534), .Z(n34592) );
  XNOR U35339 ( .A(q[0]), .B(DB[1582]), .Z(n23534) );
  XNOR U35340 ( .A(q[3]), .B(DB[1585]), .Z(n23532) );
  IV U35341 ( .A(n23531), .Z(n34591) );
  XNOR U35342 ( .A(n23529), .B(n34593), .Z(n23531) );
  XNOR U35343 ( .A(q[2]), .B(DB[1584]), .Z(n34593) );
  XNOR U35344 ( .A(q[1]), .B(DB[1583]), .Z(n23529) );
  XOR U35345 ( .A(n34594), .B(n23494), .Z(n23457) );
  XOR U35346 ( .A(n34595), .B(n23482), .Z(n23494) );
  XNOR U35347 ( .A(q[6]), .B(DB[1595]), .Z(n23482) );
  IV U35348 ( .A(n23481), .Z(n34595) );
  XNOR U35349 ( .A(n23479), .B(n34596), .Z(n23481) );
  XNOR U35350 ( .A(q[5]), .B(DB[1594]), .Z(n34596) );
  XNOR U35351 ( .A(q[4]), .B(DB[1593]), .Z(n23479) );
  IV U35352 ( .A(n23493), .Z(n34594) );
  XOR U35353 ( .A(n34597), .B(n34598), .Z(n23493) );
  XNOR U35354 ( .A(n23489), .B(n23491), .Z(n34598) );
  XNOR U35355 ( .A(q[0]), .B(DB[1589]), .Z(n23491) );
  XNOR U35356 ( .A(q[3]), .B(DB[1592]), .Z(n23489) );
  IV U35357 ( .A(n23488), .Z(n34597) );
  XNOR U35358 ( .A(n23486), .B(n34599), .Z(n23488) );
  XNOR U35359 ( .A(q[2]), .B(DB[1591]), .Z(n34599) );
  XNOR U35360 ( .A(q[1]), .B(DB[1590]), .Z(n23486) );
  XOR U35361 ( .A(n34600), .B(n23451), .Z(n23414) );
  XOR U35362 ( .A(n34601), .B(n23439), .Z(n23451) );
  XNOR U35363 ( .A(q[6]), .B(DB[1602]), .Z(n23439) );
  IV U35364 ( .A(n23438), .Z(n34601) );
  XNOR U35365 ( .A(n23436), .B(n34602), .Z(n23438) );
  XNOR U35366 ( .A(q[5]), .B(DB[1601]), .Z(n34602) );
  XNOR U35367 ( .A(q[4]), .B(DB[1600]), .Z(n23436) );
  IV U35368 ( .A(n23450), .Z(n34600) );
  XOR U35369 ( .A(n34603), .B(n34604), .Z(n23450) );
  XNOR U35370 ( .A(n23446), .B(n23448), .Z(n34604) );
  XNOR U35371 ( .A(q[0]), .B(DB[1596]), .Z(n23448) );
  XNOR U35372 ( .A(q[3]), .B(DB[1599]), .Z(n23446) );
  IV U35373 ( .A(n23445), .Z(n34603) );
  XNOR U35374 ( .A(n23443), .B(n34605), .Z(n23445) );
  XNOR U35375 ( .A(q[2]), .B(DB[1598]), .Z(n34605) );
  XNOR U35376 ( .A(q[1]), .B(DB[1597]), .Z(n23443) );
  XOR U35377 ( .A(n34606), .B(n23408), .Z(n23371) );
  XOR U35378 ( .A(n34607), .B(n23396), .Z(n23408) );
  XNOR U35379 ( .A(q[6]), .B(DB[1609]), .Z(n23396) );
  IV U35380 ( .A(n23395), .Z(n34607) );
  XNOR U35381 ( .A(n23393), .B(n34608), .Z(n23395) );
  XNOR U35382 ( .A(q[5]), .B(DB[1608]), .Z(n34608) );
  XNOR U35383 ( .A(q[4]), .B(DB[1607]), .Z(n23393) );
  IV U35384 ( .A(n23407), .Z(n34606) );
  XOR U35385 ( .A(n34609), .B(n34610), .Z(n23407) );
  XNOR U35386 ( .A(n23403), .B(n23405), .Z(n34610) );
  XNOR U35387 ( .A(q[0]), .B(DB[1603]), .Z(n23405) );
  XNOR U35388 ( .A(q[3]), .B(DB[1606]), .Z(n23403) );
  IV U35389 ( .A(n23402), .Z(n34609) );
  XNOR U35390 ( .A(n23400), .B(n34611), .Z(n23402) );
  XNOR U35391 ( .A(q[2]), .B(DB[1605]), .Z(n34611) );
  XNOR U35392 ( .A(q[1]), .B(DB[1604]), .Z(n23400) );
  XOR U35393 ( .A(n34612), .B(n23365), .Z(n23328) );
  XOR U35394 ( .A(n34613), .B(n23353), .Z(n23365) );
  XNOR U35395 ( .A(q[6]), .B(DB[1616]), .Z(n23353) );
  IV U35396 ( .A(n23352), .Z(n34613) );
  XNOR U35397 ( .A(n23350), .B(n34614), .Z(n23352) );
  XNOR U35398 ( .A(q[5]), .B(DB[1615]), .Z(n34614) );
  XNOR U35399 ( .A(q[4]), .B(DB[1614]), .Z(n23350) );
  IV U35400 ( .A(n23364), .Z(n34612) );
  XOR U35401 ( .A(n34615), .B(n34616), .Z(n23364) );
  XNOR U35402 ( .A(n23360), .B(n23362), .Z(n34616) );
  XNOR U35403 ( .A(q[0]), .B(DB[1610]), .Z(n23362) );
  XNOR U35404 ( .A(q[3]), .B(DB[1613]), .Z(n23360) );
  IV U35405 ( .A(n23359), .Z(n34615) );
  XNOR U35406 ( .A(n23357), .B(n34617), .Z(n23359) );
  XNOR U35407 ( .A(q[2]), .B(DB[1612]), .Z(n34617) );
  XNOR U35408 ( .A(q[1]), .B(DB[1611]), .Z(n23357) );
  XOR U35409 ( .A(n34618), .B(n23322), .Z(n23285) );
  XOR U35410 ( .A(n34619), .B(n23310), .Z(n23322) );
  XNOR U35411 ( .A(q[6]), .B(DB[1623]), .Z(n23310) );
  IV U35412 ( .A(n23309), .Z(n34619) );
  XNOR U35413 ( .A(n23307), .B(n34620), .Z(n23309) );
  XNOR U35414 ( .A(q[5]), .B(DB[1622]), .Z(n34620) );
  XNOR U35415 ( .A(q[4]), .B(DB[1621]), .Z(n23307) );
  IV U35416 ( .A(n23321), .Z(n34618) );
  XOR U35417 ( .A(n34621), .B(n34622), .Z(n23321) );
  XNOR U35418 ( .A(n23317), .B(n23319), .Z(n34622) );
  XNOR U35419 ( .A(q[0]), .B(DB[1617]), .Z(n23319) );
  XNOR U35420 ( .A(q[3]), .B(DB[1620]), .Z(n23317) );
  IV U35421 ( .A(n23316), .Z(n34621) );
  XNOR U35422 ( .A(n23314), .B(n34623), .Z(n23316) );
  XNOR U35423 ( .A(q[2]), .B(DB[1619]), .Z(n34623) );
  XNOR U35424 ( .A(q[1]), .B(DB[1618]), .Z(n23314) );
  XOR U35425 ( .A(n34624), .B(n23279), .Z(n23242) );
  XOR U35426 ( .A(n34625), .B(n23267), .Z(n23279) );
  XNOR U35427 ( .A(q[6]), .B(DB[1630]), .Z(n23267) );
  IV U35428 ( .A(n23266), .Z(n34625) );
  XNOR U35429 ( .A(n23264), .B(n34626), .Z(n23266) );
  XNOR U35430 ( .A(q[5]), .B(DB[1629]), .Z(n34626) );
  XNOR U35431 ( .A(q[4]), .B(DB[1628]), .Z(n23264) );
  IV U35432 ( .A(n23278), .Z(n34624) );
  XOR U35433 ( .A(n34627), .B(n34628), .Z(n23278) );
  XNOR U35434 ( .A(n23274), .B(n23276), .Z(n34628) );
  XNOR U35435 ( .A(q[0]), .B(DB[1624]), .Z(n23276) );
  XNOR U35436 ( .A(q[3]), .B(DB[1627]), .Z(n23274) );
  IV U35437 ( .A(n23273), .Z(n34627) );
  XNOR U35438 ( .A(n23271), .B(n34629), .Z(n23273) );
  XNOR U35439 ( .A(q[2]), .B(DB[1626]), .Z(n34629) );
  XNOR U35440 ( .A(q[1]), .B(DB[1625]), .Z(n23271) );
  XOR U35441 ( .A(n34630), .B(n23236), .Z(n23199) );
  XOR U35442 ( .A(n34631), .B(n23224), .Z(n23236) );
  XNOR U35443 ( .A(q[6]), .B(DB[1637]), .Z(n23224) );
  IV U35444 ( .A(n23223), .Z(n34631) );
  XNOR U35445 ( .A(n23221), .B(n34632), .Z(n23223) );
  XNOR U35446 ( .A(q[5]), .B(DB[1636]), .Z(n34632) );
  XNOR U35447 ( .A(q[4]), .B(DB[1635]), .Z(n23221) );
  IV U35448 ( .A(n23235), .Z(n34630) );
  XOR U35449 ( .A(n34633), .B(n34634), .Z(n23235) );
  XNOR U35450 ( .A(n23231), .B(n23233), .Z(n34634) );
  XNOR U35451 ( .A(q[0]), .B(DB[1631]), .Z(n23233) );
  XNOR U35452 ( .A(q[3]), .B(DB[1634]), .Z(n23231) );
  IV U35453 ( .A(n23230), .Z(n34633) );
  XNOR U35454 ( .A(n23228), .B(n34635), .Z(n23230) );
  XNOR U35455 ( .A(q[2]), .B(DB[1633]), .Z(n34635) );
  XNOR U35456 ( .A(q[1]), .B(DB[1632]), .Z(n23228) );
  XOR U35457 ( .A(n34636), .B(n23193), .Z(n23156) );
  XOR U35458 ( .A(n34637), .B(n23181), .Z(n23193) );
  XNOR U35459 ( .A(q[6]), .B(DB[1644]), .Z(n23181) );
  IV U35460 ( .A(n23180), .Z(n34637) );
  XNOR U35461 ( .A(n23178), .B(n34638), .Z(n23180) );
  XNOR U35462 ( .A(q[5]), .B(DB[1643]), .Z(n34638) );
  XNOR U35463 ( .A(q[4]), .B(DB[1642]), .Z(n23178) );
  IV U35464 ( .A(n23192), .Z(n34636) );
  XOR U35465 ( .A(n34639), .B(n34640), .Z(n23192) );
  XNOR U35466 ( .A(n23188), .B(n23190), .Z(n34640) );
  XNOR U35467 ( .A(q[0]), .B(DB[1638]), .Z(n23190) );
  XNOR U35468 ( .A(q[3]), .B(DB[1641]), .Z(n23188) );
  IV U35469 ( .A(n23187), .Z(n34639) );
  XNOR U35470 ( .A(n23185), .B(n34641), .Z(n23187) );
  XNOR U35471 ( .A(q[2]), .B(DB[1640]), .Z(n34641) );
  XNOR U35472 ( .A(q[1]), .B(DB[1639]), .Z(n23185) );
  XOR U35473 ( .A(n34642), .B(n23150), .Z(n23113) );
  XOR U35474 ( .A(n34643), .B(n23138), .Z(n23150) );
  XNOR U35475 ( .A(q[6]), .B(DB[1651]), .Z(n23138) );
  IV U35476 ( .A(n23137), .Z(n34643) );
  XNOR U35477 ( .A(n23135), .B(n34644), .Z(n23137) );
  XNOR U35478 ( .A(q[5]), .B(DB[1650]), .Z(n34644) );
  XNOR U35479 ( .A(q[4]), .B(DB[1649]), .Z(n23135) );
  IV U35480 ( .A(n23149), .Z(n34642) );
  XOR U35481 ( .A(n34645), .B(n34646), .Z(n23149) );
  XNOR U35482 ( .A(n23145), .B(n23147), .Z(n34646) );
  XNOR U35483 ( .A(q[0]), .B(DB[1645]), .Z(n23147) );
  XNOR U35484 ( .A(q[3]), .B(DB[1648]), .Z(n23145) );
  IV U35485 ( .A(n23144), .Z(n34645) );
  XNOR U35486 ( .A(n23142), .B(n34647), .Z(n23144) );
  XNOR U35487 ( .A(q[2]), .B(DB[1647]), .Z(n34647) );
  XNOR U35488 ( .A(q[1]), .B(DB[1646]), .Z(n23142) );
  XOR U35489 ( .A(n34648), .B(n23107), .Z(n23070) );
  XOR U35490 ( .A(n34649), .B(n23095), .Z(n23107) );
  XNOR U35491 ( .A(q[6]), .B(DB[1658]), .Z(n23095) );
  IV U35492 ( .A(n23094), .Z(n34649) );
  XNOR U35493 ( .A(n23092), .B(n34650), .Z(n23094) );
  XNOR U35494 ( .A(q[5]), .B(DB[1657]), .Z(n34650) );
  XNOR U35495 ( .A(q[4]), .B(DB[1656]), .Z(n23092) );
  IV U35496 ( .A(n23106), .Z(n34648) );
  XOR U35497 ( .A(n34651), .B(n34652), .Z(n23106) );
  XNOR U35498 ( .A(n23102), .B(n23104), .Z(n34652) );
  XNOR U35499 ( .A(q[0]), .B(DB[1652]), .Z(n23104) );
  XNOR U35500 ( .A(q[3]), .B(DB[1655]), .Z(n23102) );
  IV U35501 ( .A(n23101), .Z(n34651) );
  XNOR U35502 ( .A(n23099), .B(n34653), .Z(n23101) );
  XNOR U35503 ( .A(q[2]), .B(DB[1654]), .Z(n34653) );
  XNOR U35504 ( .A(q[1]), .B(DB[1653]), .Z(n23099) );
  XOR U35505 ( .A(n34654), .B(n23064), .Z(n23027) );
  XOR U35506 ( .A(n34655), .B(n23052), .Z(n23064) );
  XNOR U35507 ( .A(q[6]), .B(DB[1665]), .Z(n23052) );
  IV U35508 ( .A(n23051), .Z(n34655) );
  XNOR U35509 ( .A(n23049), .B(n34656), .Z(n23051) );
  XNOR U35510 ( .A(q[5]), .B(DB[1664]), .Z(n34656) );
  XNOR U35511 ( .A(q[4]), .B(DB[1663]), .Z(n23049) );
  IV U35512 ( .A(n23063), .Z(n34654) );
  XOR U35513 ( .A(n34657), .B(n34658), .Z(n23063) );
  XNOR U35514 ( .A(n23059), .B(n23061), .Z(n34658) );
  XNOR U35515 ( .A(q[0]), .B(DB[1659]), .Z(n23061) );
  XNOR U35516 ( .A(q[3]), .B(DB[1662]), .Z(n23059) );
  IV U35517 ( .A(n23058), .Z(n34657) );
  XNOR U35518 ( .A(n23056), .B(n34659), .Z(n23058) );
  XNOR U35519 ( .A(q[2]), .B(DB[1661]), .Z(n34659) );
  XNOR U35520 ( .A(q[1]), .B(DB[1660]), .Z(n23056) );
  XOR U35521 ( .A(n34660), .B(n23021), .Z(n22984) );
  XOR U35522 ( .A(n34661), .B(n23009), .Z(n23021) );
  XNOR U35523 ( .A(q[6]), .B(DB[1672]), .Z(n23009) );
  IV U35524 ( .A(n23008), .Z(n34661) );
  XNOR U35525 ( .A(n23006), .B(n34662), .Z(n23008) );
  XNOR U35526 ( .A(q[5]), .B(DB[1671]), .Z(n34662) );
  XNOR U35527 ( .A(q[4]), .B(DB[1670]), .Z(n23006) );
  IV U35528 ( .A(n23020), .Z(n34660) );
  XOR U35529 ( .A(n34663), .B(n34664), .Z(n23020) );
  XNOR U35530 ( .A(n23016), .B(n23018), .Z(n34664) );
  XNOR U35531 ( .A(q[0]), .B(DB[1666]), .Z(n23018) );
  XNOR U35532 ( .A(q[3]), .B(DB[1669]), .Z(n23016) );
  IV U35533 ( .A(n23015), .Z(n34663) );
  XNOR U35534 ( .A(n23013), .B(n34665), .Z(n23015) );
  XNOR U35535 ( .A(q[2]), .B(DB[1668]), .Z(n34665) );
  XNOR U35536 ( .A(q[1]), .B(DB[1667]), .Z(n23013) );
  XOR U35537 ( .A(n34666), .B(n22978), .Z(n22941) );
  XOR U35538 ( .A(n34667), .B(n22966), .Z(n22978) );
  XNOR U35539 ( .A(q[6]), .B(DB[1679]), .Z(n22966) );
  IV U35540 ( .A(n22965), .Z(n34667) );
  XNOR U35541 ( .A(n22963), .B(n34668), .Z(n22965) );
  XNOR U35542 ( .A(q[5]), .B(DB[1678]), .Z(n34668) );
  XNOR U35543 ( .A(q[4]), .B(DB[1677]), .Z(n22963) );
  IV U35544 ( .A(n22977), .Z(n34666) );
  XOR U35545 ( .A(n34669), .B(n34670), .Z(n22977) );
  XNOR U35546 ( .A(n22973), .B(n22975), .Z(n34670) );
  XNOR U35547 ( .A(q[0]), .B(DB[1673]), .Z(n22975) );
  XNOR U35548 ( .A(q[3]), .B(DB[1676]), .Z(n22973) );
  IV U35549 ( .A(n22972), .Z(n34669) );
  XNOR U35550 ( .A(n22970), .B(n34671), .Z(n22972) );
  XNOR U35551 ( .A(q[2]), .B(DB[1675]), .Z(n34671) );
  XNOR U35552 ( .A(q[1]), .B(DB[1674]), .Z(n22970) );
  XOR U35553 ( .A(n34672), .B(n22935), .Z(n22898) );
  XOR U35554 ( .A(n34673), .B(n22923), .Z(n22935) );
  XNOR U35555 ( .A(q[6]), .B(DB[1686]), .Z(n22923) );
  IV U35556 ( .A(n22922), .Z(n34673) );
  XNOR U35557 ( .A(n22920), .B(n34674), .Z(n22922) );
  XNOR U35558 ( .A(q[5]), .B(DB[1685]), .Z(n34674) );
  XNOR U35559 ( .A(q[4]), .B(DB[1684]), .Z(n22920) );
  IV U35560 ( .A(n22934), .Z(n34672) );
  XOR U35561 ( .A(n34675), .B(n34676), .Z(n22934) );
  XNOR U35562 ( .A(n22930), .B(n22932), .Z(n34676) );
  XNOR U35563 ( .A(q[0]), .B(DB[1680]), .Z(n22932) );
  XNOR U35564 ( .A(q[3]), .B(DB[1683]), .Z(n22930) );
  IV U35565 ( .A(n22929), .Z(n34675) );
  XNOR U35566 ( .A(n22927), .B(n34677), .Z(n22929) );
  XNOR U35567 ( .A(q[2]), .B(DB[1682]), .Z(n34677) );
  XNOR U35568 ( .A(q[1]), .B(DB[1681]), .Z(n22927) );
  XOR U35569 ( .A(n34678), .B(n22892), .Z(n22855) );
  XOR U35570 ( .A(n34679), .B(n22880), .Z(n22892) );
  XNOR U35571 ( .A(q[6]), .B(DB[1693]), .Z(n22880) );
  IV U35572 ( .A(n22879), .Z(n34679) );
  XNOR U35573 ( .A(n22877), .B(n34680), .Z(n22879) );
  XNOR U35574 ( .A(q[5]), .B(DB[1692]), .Z(n34680) );
  XNOR U35575 ( .A(q[4]), .B(DB[1691]), .Z(n22877) );
  IV U35576 ( .A(n22891), .Z(n34678) );
  XOR U35577 ( .A(n34681), .B(n34682), .Z(n22891) );
  XNOR U35578 ( .A(n22887), .B(n22889), .Z(n34682) );
  XNOR U35579 ( .A(q[0]), .B(DB[1687]), .Z(n22889) );
  XNOR U35580 ( .A(q[3]), .B(DB[1690]), .Z(n22887) );
  IV U35581 ( .A(n22886), .Z(n34681) );
  XNOR U35582 ( .A(n22884), .B(n34683), .Z(n22886) );
  XNOR U35583 ( .A(q[2]), .B(DB[1689]), .Z(n34683) );
  XNOR U35584 ( .A(q[1]), .B(DB[1688]), .Z(n22884) );
  XOR U35585 ( .A(n34684), .B(n22849), .Z(n22812) );
  XOR U35586 ( .A(n34685), .B(n22837), .Z(n22849) );
  XNOR U35587 ( .A(q[6]), .B(DB[1700]), .Z(n22837) );
  IV U35588 ( .A(n22836), .Z(n34685) );
  XNOR U35589 ( .A(n22834), .B(n34686), .Z(n22836) );
  XNOR U35590 ( .A(q[5]), .B(DB[1699]), .Z(n34686) );
  XNOR U35591 ( .A(q[4]), .B(DB[1698]), .Z(n22834) );
  IV U35592 ( .A(n22848), .Z(n34684) );
  XOR U35593 ( .A(n34687), .B(n34688), .Z(n22848) );
  XNOR U35594 ( .A(n22844), .B(n22846), .Z(n34688) );
  XNOR U35595 ( .A(q[0]), .B(DB[1694]), .Z(n22846) );
  XNOR U35596 ( .A(q[3]), .B(DB[1697]), .Z(n22844) );
  IV U35597 ( .A(n22843), .Z(n34687) );
  XNOR U35598 ( .A(n22841), .B(n34689), .Z(n22843) );
  XNOR U35599 ( .A(q[2]), .B(DB[1696]), .Z(n34689) );
  XNOR U35600 ( .A(q[1]), .B(DB[1695]), .Z(n22841) );
  XOR U35601 ( .A(n34690), .B(n22806), .Z(n22769) );
  XOR U35602 ( .A(n34691), .B(n22794), .Z(n22806) );
  XNOR U35603 ( .A(q[6]), .B(DB[1707]), .Z(n22794) );
  IV U35604 ( .A(n22793), .Z(n34691) );
  XNOR U35605 ( .A(n22791), .B(n34692), .Z(n22793) );
  XNOR U35606 ( .A(q[5]), .B(DB[1706]), .Z(n34692) );
  XNOR U35607 ( .A(q[4]), .B(DB[1705]), .Z(n22791) );
  IV U35608 ( .A(n22805), .Z(n34690) );
  XOR U35609 ( .A(n34693), .B(n34694), .Z(n22805) );
  XNOR U35610 ( .A(n22801), .B(n22803), .Z(n34694) );
  XNOR U35611 ( .A(q[0]), .B(DB[1701]), .Z(n22803) );
  XNOR U35612 ( .A(q[3]), .B(DB[1704]), .Z(n22801) );
  IV U35613 ( .A(n22800), .Z(n34693) );
  XNOR U35614 ( .A(n22798), .B(n34695), .Z(n22800) );
  XNOR U35615 ( .A(q[2]), .B(DB[1703]), .Z(n34695) );
  XNOR U35616 ( .A(q[1]), .B(DB[1702]), .Z(n22798) );
  XOR U35617 ( .A(n34696), .B(n22763), .Z(n22726) );
  XOR U35618 ( .A(n34697), .B(n22751), .Z(n22763) );
  XNOR U35619 ( .A(q[6]), .B(DB[1714]), .Z(n22751) );
  IV U35620 ( .A(n22750), .Z(n34697) );
  XNOR U35621 ( .A(n22748), .B(n34698), .Z(n22750) );
  XNOR U35622 ( .A(q[5]), .B(DB[1713]), .Z(n34698) );
  XNOR U35623 ( .A(q[4]), .B(DB[1712]), .Z(n22748) );
  IV U35624 ( .A(n22762), .Z(n34696) );
  XOR U35625 ( .A(n34699), .B(n34700), .Z(n22762) );
  XNOR U35626 ( .A(n22758), .B(n22760), .Z(n34700) );
  XNOR U35627 ( .A(q[0]), .B(DB[1708]), .Z(n22760) );
  XNOR U35628 ( .A(q[3]), .B(DB[1711]), .Z(n22758) );
  IV U35629 ( .A(n22757), .Z(n34699) );
  XNOR U35630 ( .A(n22755), .B(n34701), .Z(n22757) );
  XNOR U35631 ( .A(q[2]), .B(DB[1710]), .Z(n34701) );
  XNOR U35632 ( .A(q[1]), .B(DB[1709]), .Z(n22755) );
  XOR U35633 ( .A(n34702), .B(n22720), .Z(n22683) );
  XOR U35634 ( .A(n34703), .B(n22708), .Z(n22720) );
  XNOR U35635 ( .A(q[6]), .B(DB[1721]), .Z(n22708) );
  IV U35636 ( .A(n22707), .Z(n34703) );
  XNOR U35637 ( .A(n22705), .B(n34704), .Z(n22707) );
  XNOR U35638 ( .A(q[5]), .B(DB[1720]), .Z(n34704) );
  XNOR U35639 ( .A(q[4]), .B(DB[1719]), .Z(n22705) );
  IV U35640 ( .A(n22719), .Z(n34702) );
  XOR U35641 ( .A(n34705), .B(n34706), .Z(n22719) );
  XNOR U35642 ( .A(n22715), .B(n22717), .Z(n34706) );
  XNOR U35643 ( .A(q[0]), .B(DB[1715]), .Z(n22717) );
  XNOR U35644 ( .A(q[3]), .B(DB[1718]), .Z(n22715) );
  IV U35645 ( .A(n22714), .Z(n34705) );
  XNOR U35646 ( .A(n22712), .B(n34707), .Z(n22714) );
  XNOR U35647 ( .A(q[2]), .B(DB[1717]), .Z(n34707) );
  XNOR U35648 ( .A(q[1]), .B(DB[1716]), .Z(n22712) );
  XOR U35649 ( .A(n34708), .B(n22677), .Z(n22640) );
  XOR U35650 ( .A(n34709), .B(n22665), .Z(n22677) );
  XNOR U35651 ( .A(q[6]), .B(DB[1728]), .Z(n22665) );
  IV U35652 ( .A(n22664), .Z(n34709) );
  XNOR U35653 ( .A(n22662), .B(n34710), .Z(n22664) );
  XNOR U35654 ( .A(q[5]), .B(DB[1727]), .Z(n34710) );
  XNOR U35655 ( .A(q[4]), .B(DB[1726]), .Z(n22662) );
  IV U35656 ( .A(n22676), .Z(n34708) );
  XOR U35657 ( .A(n34711), .B(n34712), .Z(n22676) );
  XNOR U35658 ( .A(n22672), .B(n22674), .Z(n34712) );
  XNOR U35659 ( .A(q[0]), .B(DB[1722]), .Z(n22674) );
  XNOR U35660 ( .A(q[3]), .B(DB[1725]), .Z(n22672) );
  IV U35661 ( .A(n22671), .Z(n34711) );
  XNOR U35662 ( .A(n22669), .B(n34713), .Z(n22671) );
  XNOR U35663 ( .A(q[2]), .B(DB[1724]), .Z(n34713) );
  XNOR U35664 ( .A(q[1]), .B(DB[1723]), .Z(n22669) );
  XOR U35665 ( .A(n34714), .B(n22634), .Z(n22597) );
  XOR U35666 ( .A(n34715), .B(n22622), .Z(n22634) );
  XNOR U35667 ( .A(q[6]), .B(DB[1735]), .Z(n22622) );
  IV U35668 ( .A(n22621), .Z(n34715) );
  XNOR U35669 ( .A(n22619), .B(n34716), .Z(n22621) );
  XNOR U35670 ( .A(q[5]), .B(DB[1734]), .Z(n34716) );
  XNOR U35671 ( .A(q[4]), .B(DB[1733]), .Z(n22619) );
  IV U35672 ( .A(n22633), .Z(n34714) );
  XOR U35673 ( .A(n34717), .B(n34718), .Z(n22633) );
  XNOR U35674 ( .A(n22629), .B(n22631), .Z(n34718) );
  XNOR U35675 ( .A(q[0]), .B(DB[1729]), .Z(n22631) );
  XNOR U35676 ( .A(q[3]), .B(DB[1732]), .Z(n22629) );
  IV U35677 ( .A(n22628), .Z(n34717) );
  XNOR U35678 ( .A(n22626), .B(n34719), .Z(n22628) );
  XNOR U35679 ( .A(q[2]), .B(DB[1731]), .Z(n34719) );
  XNOR U35680 ( .A(q[1]), .B(DB[1730]), .Z(n22626) );
  XOR U35681 ( .A(n34720), .B(n22591), .Z(n22554) );
  XOR U35682 ( .A(n34721), .B(n22579), .Z(n22591) );
  XNOR U35683 ( .A(q[6]), .B(DB[1742]), .Z(n22579) );
  IV U35684 ( .A(n22578), .Z(n34721) );
  XNOR U35685 ( .A(n22576), .B(n34722), .Z(n22578) );
  XNOR U35686 ( .A(q[5]), .B(DB[1741]), .Z(n34722) );
  XNOR U35687 ( .A(q[4]), .B(DB[1740]), .Z(n22576) );
  IV U35688 ( .A(n22590), .Z(n34720) );
  XOR U35689 ( .A(n34723), .B(n34724), .Z(n22590) );
  XNOR U35690 ( .A(n22586), .B(n22588), .Z(n34724) );
  XNOR U35691 ( .A(q[0]), .B(DB[1736]), .Z(n22588) );
  XNOR U35692 ( .A(q[3]), .B(DB[1739]), .Z(n22586) );
  IV U35693 ( .A(n22585), .Z(n34723) );
  XNOR U35694 ( .A(n22583), .B(n34725), .Z(n22585) );
  XNOR U35695 ( .A(q[2]), .B(DB[1738]), .Z(n34725) );
  XNOR U35696 ( .A(q[1]), .B(DB[1737]), .Z(n22583) );
  XOR U35697 ( .A(n34726), .B(n22548), .Z(n22511) );
  XOR U35698 ( .A(n34727), .B(n22536), .Z(n22548) );
  XNOR U35699 ( .A(q[6]), .B(DB[1749]), .Z(n22536) );
  IV U35700 ( .A(n22535), .Z(n34727) );
  XNOR U35701 ( .A(n22533), .B(n34728), .Z(n22535) );
  XNOR U35702 ( .A(q[5]), .B(DB[1748]), .Z(n34728) );
  XNOR U35703 ( .A(q[4]), .B(DB[1747]), .Z(n22533) );
  IV U35704 ( .A(n22547), .Z(n34726) );
  XOR U35705 ( .A(n34729), .B(n34730), .Z(n22547) );
  XNOR U35706 ( .A(n22543), .B(n22545), .Z(n34730) );
  XNOR U35707 ( .A(q[0]), .B(DB[1743]), .Z(n22545) );
  XNOR U35708 ( .A(q[3]), .B(DB[1746]), .Z(n22543) );
  IV U35709 ( .A(n22542), .Z(n34729) );
  XNOR U35710 ( .A(n22540), .B(n34731), .Z(n22542) );
  XNOR U35711 ( .A(q[2]), .B(DB[1745]), .Z(n34731) );
  XNOR U35712 ( .A(q[1]), .B(DB[1744]), .Z(n22540) );
  XOR U35713 ( .A(n34732), .B(n22505), .Z(n22468) );
  XOR U35714 ( .A(n34733), .B(n22493), .Z(n22505) );
  XNOR U35715 ( .A(q[6]), .B(DB[1756]), .Z(n22493) );
  IV U35716 ( .A(n22492), .Z(n34733) );
  XNOR U35717 ( .A(n22490), .B(n34734), .Z(n22492) );
  XNOR U35718 ( .A(q[5]), .B(DB[1755]), .Z(n34734) );
  XNOR U35719 ( .A(q[4]), .B(DB[1754]), .Z(n22490) );
  IV U35720 ( .A(n22504), .Z(n34732) );
  XOR U35721 ( .A(n34735), .B(n34736), .Z(n22504) );
  XNOR U35722 ( .A(n22500), .B(n22502), .Z(n34736) );
  XNOR U35723 ( .A(q[0]), .B(DB[1750]), .Z(n22502) );
  XNOR U35724 ( .A(q[3]), .B(DB[1753]), .Z(n22500) );
  IV U35725 ( .A(n22499), .Z(n34735) );
  XNOR U35726 ( .A(n22497), .B(n34737), .Z(n22499) );
  XNOR U35727 ( .A(q[2]), .B(DB[1752]), .Z(n34737) );
  XNOR U35728 ( .A(q[1]), .B(DB[1751]), .Z(n22497) );
  XOR U35729 ( .A(n34738), .B(n22462), .Z(n22425) );
  XOR U35730 ( .A(n34739), .B(n22450), .Z(n22462) );
  XNOR U35731 ( .A(q[6]), .B(DB[1763]), .Z(n22450) );
  IV U35732 ( .A(n22449), .Z(n34739) );
  XNOR U35733 ( .A(n22447), .B(n34740), .Z(n22449) );
  XNOR U35734 ( .A(q[5]), .B(DB[1762]), .Z(n34740) );
  XNOR U35735 ( .A(q[4]), .B(DB[1761]), .Z(n22447) );
  IV U35736 ( .A(n22461), .Z(n34738) );
  XOR U35737 ( .A(n34741), .B(n34742), .Z(n22461) );
  XNOR U35738 ( .A(n22457), .B(n22459), .Z(n34742) );
  XNOR U35739 ( .A(q[0]), .B(DB[1757]), .Z(n22459) );
  XNOR U35740 ( .A(q[3]), .B(DB[1760]), .Z(n22457) );
  IV U35741 ( .A(n22456), .Z(n34741) );
  XNOR U35742 ( .A(n22454), .B(n34743), .Z(n22456) );
  XNOR U35743 ( .A(q[2]), .B(DB[1759]), .Z(n34743) );
  XNOR U35744 ( .A(q[1]), .B(DB[1758]), .Z(n22454) );
  XOR U35745 ( .A(n34744), .B(n22419), .Z(n22382) );
  XOR U35746 ( .A(n34745), .B(n22407), .Z(n22419) );
  XNOR U35747 ( .A(q[6]), .B(DB[1770]), .Z(n22407) );
  IV U35748 ( .A(n22406), .Z(n34745) );
  XNOR U35749 ( .A(n22404), .B(n34746), .Z(n22406) );
  XNOR U35750 ( .A(q[5]), .B(DB[1769]), .Z(n34746) );
  XNOR U35751 ( .A(q[4]), .B(DB[1768]), .Z(n22404) );
  IV U35752 ( .A(n22418), .Z(n34744) );
  XOR U35753 ( .A(n34747), .B(n34748), .Z(n22418) );
  XNOR U35754 ( .A(n22414), .B(n22416), .Z(n34748) );
  XNOR U35755 ( .A(q[0]), .B(DB[1764]), .Z(n22416) );
  XNOR U35756 ( .A(q[3]), .B(DB[1767]), .Z(n22414) );
  IV U35757 ( .A(n22413), .Z(n34747) );
  XNOR U35758 ( .A(n22411), .B(n34749), .Z(n22413) );
  XNOR U35759 ( .A(q[2]), .B(DB[1766]), .Z(n34749) );
  XNOR U35760 ( .A(q[1]), .B(DB[1765]), .Z(n22411) );
  XOR U35761 ( .A(n34750), .B(n22376), .Z(n22339) );
  XOR U35762 ( .A(n34751), .B(n22364), .Z(n22376) );
  XNOR U35763 ( .A(q[6]), .B(DB[1777]), .Z(n22364) );
  IV U35764 ( .A(n22363), .Z(n34751) );
  XNOR U35765 ( .A(n22361), .B(n34752), .Z(n22363) );
  XNOR U35766 ( .A(q[5]), .B(DB[1776]), .Z(n34752) );
  XNOR U35767 ( .A(q[4]), .B(DB[1775]), .Z(n22361) );
  IV U35768 ( .A(n22375), .Z(n34750) );
  XOR U35769 ( .A(n34753), .B(n34754), .Z(n22375) );
  XNOR U35770 ( .A(n22371), .B(n22373), .Z(n34754) );
  XNOR U35771 ( .A(q[0]), .B(DB[1771]), .Z(n22373) );
  XNOR U35772 ( .A(q[3]), .B(DB[1774]), .Z(n22371) );
  IV U35773 ( .A(n22370), .Z(n34753) );
  XNOR U35774 ( .A(n22368), .B(n34755), .Z(n22370) );
  XNOR U35775 ( .A(q[2]), .B(DB[1773]), .Z(n34755) );
  XNOR U35776 ( .A(q[1]), .B(DB[1772]), .Z(n22368) );
  XOR U35777 ( .A(n34756), .B(n22333), .Z(n22296) );
  XOR U35778 ( .A(n34757), .B(n22321), .Z(n22333) );
  XNOR U35779 ( .A(q[6]), .B(DB[1784]), .Z(n22321) );
  IV U35780 ( .A(n22320), .Z(n34757) );
  XNOR U35781 ( .A(n22318), .B(n34758), .Z(n22320) );
  XNOR U35782 ( .A(q[5]), .B(DB[1783]), .Z(n34758) );
  XNOR U35783 ( .A(q[4]), .B(DB[1782]), .Z(n22318) );
  IV U35784 ( .A(n22332), .Z(n34756) );
  XOR U35785 ( .A(n34759), .B(n34760), .Z(n22332) );
  XNOR U35786 ( .A(n22328), .B(n22330), .Z(n34760) );
  XNOR U35787 ( .A(q[0]), .B(DB[1778]), .Z(n22330) );
  XNOR U35788 ( .A(q[3]), .B(DB[1781]), .Z(n22328) );
  IV U35789 ( .A(n22327), .Z(n34759) );
  XNOR U35790 ( .A(n22325), .B(n34761), .Z(n22327) );
  XNOR U35791 ( .A(q[2]), .B(DB[1780]), .Z(n34761) );
  XNOR U35792 ( .A(q[1]), .B(DB[1779]), .Z(n22325) );
  XOR U35793 ( .A(n34762), .B(n22290), .Z(n22253) );
  XOR U35794 ( .A(n34763), .B(n22278), .Z(n22290) );
  XNOR U35795 ( .A(q[6]), .B(DB[1791]), .Z(n22278) );
  IV U35796 ( .A(n22277), .Z(n34763) );
  XNOR U35797 ( .A(n22275), .B(n34764), .Z(n22277) );
  XNOR U35798 ( .A(q[5]), .B(DB[1790]), .Z(n34764) );
  XNOR U35799 ( .A(q[4]), .B(DB[1789]), .Z(n22275) );
  IV U35800 ( .A(n22289), .Z(n34762) );
  XOR U35801 ( .A(n34765), .B(n34766), .Z(n22289) );
  XNOR U35802 ( .A(n22285), .B(n22287), .Z(n34766) );
  XNOR U35803 ( .A(q[0]), .B(DB[1785]), .Z(n22287) );
  XNOR U35804 ( .A(q[3]), .B(DB[1788]), .Z(n22285) );
  IV U35805 ( .A(n22284), .Z(n34765) );
  XNOR U35806 ( .A(n22282), .B(n34767), .Z(n22284) );
  XNOR U35807 ( .A(q[2]), .B(DB[1787]), .Z(n34767) );
  XNOR U35808 ( .A(q[1]), .B(DB[1786]), .Z(n22282) );
  XOR U35809 ( .A(n34768), .B(n22247), .Z(n22210) );
  XOR U35810 ( .A(n34769), .B(n22235), .Z(n22247) );
  XNOR U35811 ( .A(q[6]), .B(DB[1798]), .Z(n22235) );
  IV U35812 ( .A(n22234), .Z(n34769) );
  XNOR U35813 ( .A(n22232), .B(n34770), .Z(n22234) );
  XNOR U35814 ( .A(q[5]), .B(DB[1797]), .Z(n34770) );
  XNOR U35815 ( .A(q[4]), .B(DB[1796]), .Z(n22232) );
  IV U35816 ( .A(n22246), .Z(n34768) );
  XOR U35817 ( .A(n34771), .B(n34772), .Z(n22246) );
  XNOR U35818 ( .A(n22242), .B(n22244), .Z(n34772) );
  XNOR U35819 ( .A(q[0]), .B(DB[1792]), .Z(n22244) );
  XNOR U35820 ( .A(q[3]), .B(DB[1795]), .Z(n22242) );
  IV U35821 ( .A(n22241), .Z(n34771) );
  XNOR U35822 ( .A(n22239), .B(n34773), .Z(n22241) );
  XNOR U35823 ( .A(q[2]), .B(DB[1794]), .Z(n34773) );
  XNOR U35824 ( .A(q[1]), .B(DB[1793]), .Z(n22239) );
  XOR U35825 ( .A(n34774), .B(n22204), .Z(n22167) );
  XOR U35826 ( .A(n34775), .B(n22192), .Z(n22204) );
  XNOR U35827 ( .A(q[6]), .B(DB[1805]), .Z(n22192) );
  IV U35828 ( .A(n22191), .Z(n34775) );
  XNOR U35829 ( .A(n22189), .B(n34776), .Z(n22191) );
  XNOR U35830 ( .A(q[5]), .B(DB[1804]), .Z(n34776) );
  XNOR U35831 ( .A(q[4]), .B(DB[1803]), .Z(n22189) );
  IV U35832 ( .A(n22203), .Z(n34774) );
  XOR U35833 ( .A(n34777), .B(n34778), .Z(n22203) );
  XNOR U35834 ( .A(n22199), .B(n22201), .Z(n34778) );
  XNOR U35835 ( .A(q[0]), .B(DB[1799]), .Z(n22201) );
  XNOR U35836 ( .A(q[3]), .B(DB[1802]), .Z(n22199) );
  IV U35837 ( .A(n22198), .Z(n34777) );
  XNOR U35838 ( .A(n22196), .B(n34779), .Z(n22198) );
  XNOR U35839 ( .A(q[2]), .B(DB[1801]), .Z(n34779) );
  XNOR U35840 ( .A(q[1]), .B(DB[1800]), .Z(n22196) );
  XOR U35841 ( .A(n34780), .B(n22161), .Z(n22124) );
  XOR U35842 ( .A(n34781), .B(n22149), .Z(n22161) );
  XNOR U35843 ( .A(q[6]), .B(DB[1812]), .Z(n22149) );
  IV U35844 ( .A(n22148), .Z(n34781) );
  XNOR U35845 ( .A(n22146), .B(n34782), .Z(n22148) );
  XNOR U35846 ( .A(q[5]), .B(DB[1811]), .Z(n34782) );
  XNOR U35847 ( .A(q[4]), .B(DB[1810]), .Z(n22146) );
  IV U35848 ( .A(n22160), .Z(n34780) );
  XOR U35849 ( .A(n34783), .B(n34784), .Z(n22160) );
  XNOR U35850 ( .A(n22156), .B(n22158), .Z(n34784) );
  XNOR U35851 ( .A(q[0]), .B(DB[1806]), .Z(n22158) );
  XNOR U35852 ( .A(q[3]), .B(DB[1809]), .Z(n22156) );
  IV U35853 ( .A(n22155), .Z(n34783) );
  XNOR U35854 ( .A(n22153), .B(n34785), .Z(n22155) );
  XNOR U35855 ( .A(q[2]), .B(DB[1808]), .Z(n34785) );
  XNOR U35856 ( .A(q[1]), .B(DB[1807]), .Z(n22153) );
  XOR U35857 ( .A(n34786), .B(n22118), .Z(n22081) );
  XOR U35858 ( .A(n34787), .B(n22106), .Z(n22118) );
  XNOR U35859 ( .A(q[6]), .B(DB[1819]), .Z(n22106) );
  IV U35860 ( .A(n22105), .Z(n34787) );
  XNOR U35861 ( .A(n22103), .B(n34788), .Z(n22105) );
  XNOR U35862 ( .A(q[5]), .B(DB[1818]), .Z(n34788) );
  XNOR U35863 ( .A(q[4]), .B(DB[1817]), .Z(n22103) );
  IV U35864 ( .A(n22117), .Z(n34786) );
  XOR U35865 ( .A(n34789), .B(n34790), .Z(n22117) );
  XNOR U35866 ( .A(n22113), .B(n22115), .Z(n34790) );
  XNOR U35867 ( .A(q[0]), .B(DB[1813]), .Z(n22115) );
  XNOR U35868 ( .A(q[3]), .B(DB[1816]), .Z(n22113) );
  IV U35869 ( .A(n22112), .Z(n34789) );
  XNOR U35870 ( .A(n22110), .B(n34791), .Z(n22112) );
  XNOR U35871 ( .A(q[2]), .B(DB[1815]), .Z(n34791) );
  XNOR U35872 ( .A(q[1]), .B(DB[1814]), .Z(n22110) );
  XOR U35873 ( .A(n34792), .B(n22075), .Z(n22038) );
  XOR U35874 ( .A(n34793), .B(n22063), .Z(n22075) );
  XNOR U35875 ( .A(q[6]), .B(DB[1826]), .Z(n22063) );
  IV U35876 ( .A(n22062), .Z(n34793) );
  XNOR U35877 ( .A(n22060), .B(n34794), .Z(n22062) );
  XNOR U35878 ( .A(q[5]), .B(DB[1825]), .Z(n34794) );
  XNOR U35879 ( .A(q[4]), .B(DB[1824]), .Z(n22060) );
  IV U35880 ( .A(n22074), .Z(n34792) );
  XOR U35881 ( .A(n34795), .B(n34796), .Z(n22074) );
  XNOR U35882 ( .A(n22070), .B(n22072), .Z(n34796) );
  XNOR U35883 ( .A(q[0]), .B(DB[1820]), .Z(n22072) );
  XNOR U35884 ( .A(q[3]), .B(DB[1823]), .Z(n22070) );
  IV U35885 ( .A(n22069), .Z(n34795) );
  XNOR U35886 ( .A(n22067), .B(n34797), .Z(n22069) );
  XNOR U35887 ( .A(q[2]), .B(DB[1822]), .Z(n34797) );
  XNOR U35888 ( .A(q[1]), .B(DB[1821]), .Z(n22067) );
  XOR U35889 ( .A(n34798), .B(n22032), .Z(n21995) );
  XOR U35890 ( .A(n34799), .B(n22020), .Z(n22032) );
  XNOR U35891 ( .A(q[6]), .B(DB[1833]), .Z(n22020) );
  IV U35892 ( .A(n22019), .Z(n34799) );
  XNOR U35893 ( .A(n22017), .B(n34800), .Z(n22019) );
  XNOR U35894 ( .A(q[5]), .B(DB[1832]), .Z(n34800) );
  XNOR U35895 ( .A(q[4]), .B(DB[1831]), .Z(n22017) );
  IV U35896 ( .A(n22031), .Z(n34798) );
  XOR U35897 ( .A(n34801), .B(n34802), .Z(n22031) );
  XNOR U35898 ( .A(n22027), .B(n22029), .Z(n34802) );
  XNOR U35899 ( .A(q[0]), .B(DB[1827]), .Z(n22029) );
  XNOR U35900 ( .A(q[3]), .B(DB[1830]), .Z(n22027) );
  IV U35901 ( .A(n22026), .Z(n34801) );
  XNOR U35902 ( .A(n22024), .B(n34803), .Z(n22026) );
  XNOR U35903 ( .A(q[2]), .B(DB[1829]), .Z(n34803) );
  XNOR U35904 ( .A(q[1]), .B(DB[1828]), .Z(n22024) );
  XOR U35905 ( .A(n34804), .B(n21989), .Z(n21952) );
  XOR U35906 ( .A(n34805), .B(n21977), .Z(n21989) );
  XNOR U35907 ( .A(q[6]), .B(DB[1840]), .Z(n21977) );
  IV U35908 ( .A(n21976), .Z(n34805) );
  XNOR U35909 ( .A(n21974), .B(n34806), .Z(n21976) );
  XNOR U35910 ( .A(q[5]), .B(DB[1839]), .Z(n34806) );
  XNOR U35911 ( .A(q[4]), .B(DB[1838]), .Z(n21974) );
  IV U35912 ( .A(n21988), .Z(n34804) );
  XOR U35913 ( .A(n34807), .B(n34808), .Z(n21988) );
  XNOR U35914 ( .A(n21984), .B(n21986), .Z(n34808) );
  XNOR U35915 ( .A(q[0]), .B(DB[1834]), .Z(n21986) );
  XNOR U35916 ( .A(q[3]), .B(DB[1837]), .Z(n21984) );
  IV U35917 ( .A(n21983), .Z(n34807) );
  XNOR U35918 ( .A(n21981), .B(n34809), .Z(n21983) );
  XNOR U35919 ( .A(q[2]), .B(DB[1836]), .Z(n34809) );
  XNOR U35920 ( .A(q[1]), .B(DB[1835]), .Z(n21981) );
  XOR U35921 ( .A(n34810), .B(n21946), .Z(n21909) );
  XOR U35922 ( .A(n34811), .B(n21934), .Z(n21946) );
  XNOR U35923 ( .A(q[6]), .B(DB[1847]), .Z(n21934) );
  IV U35924 ( .A(n21933), .Z(n34811) );
  XNOR U35925 ( .A(n21931), .B(n34812), .Z(n21933) );
  XNOR U35926 ( .A(q[5]), .B(DB[1846]), .Z(n34812) );
  XNOR U35927 ( .A(q[4]), .B(DB[1845]), .Z(n21931) );
  IV U35928 ( .A(n21945), .Z(n34810) );
  XOR U35929 ( .A(n34813), .B(n34814), .Z(n21945) );
  XNOR U35930 ( .A(n21941), .B(n21943), .Z(n34814) );
  XNOR U35931 ( .A(q[0]), .B(DB[1841]), .Z(n21943) );
  XNOR U35932 ( .A(q[3]), .B(DB[1844]), .Z(n21941) );
  IV U35933 ( .A(n21940), .Z(n34813) );
  XNOR U35934 ( .A(n21938), .B(n34815), .Z(n21940) );
  XNOR U35935 ( .A(q[2]), .B(DB[1843]), .Z(n34815) );
  XNOR U35936 ( .A(q[1]), .B(DB[1842]), .Z(n21938) );
  XOR U35937 ( .A(n34816), .B(n21903), .Z(n21866) );
  XOR U35938 ( .A(n34817), .B(n21891), .Z(n21903) );
  XNOR U35939 ( .A(q[6]), .B(DB[1854]), .Z(n21891) );
  IV U35940 ( .A(n21890), .Z(n34817) );
  XNOR U35941 ( .A(n21888), .B(n34818), .Z(n21890) );
  XNOR U35942 ( .A(q[5]), .B(DB[1853]), .Z(n34818) );
  XNOR U35943 ( .A(q[4]), .B(DB[1852]), .Z(n21888) );
  IV U35944 ( .A(n21902), .Z(n34816) );
  XOR U35945 ( .A(n34819), .B(n34820), .Z(n21902) );
  XNOR U35946 ( .A(n21898), .B(n21900), .Z(n34820) );
  XNOR U35947 ( .A(q[0]), .B(DB[1848]), .Z(n21900) );
  XNOR U35948 ( .A(q[3]), .B(DB[1851]), .Z(n21898) );
  IV U35949 ( .A(n21897), .Z(n34819) );
  XNOR U35950 ( .A(n21895), .B(n34821), .Z(n21897) );
  XNOR U35951 ( .A(q[2]), .B(DB[1850]), .Z(n34821) );
  XNOR U35952 ( .A(q[1]), .B(DB[1849]), .Z(n21895) );
  XOR U35953 ( .A(n34822), .B(n21860), .Z(n21823) );
  XOR U35954 ( .A(n34823), .B(n21848), .Z(n21860) );
  XNOR U35955 ( .A(q[6]), .B(DB[1861]), .Z(n21848) );
  IV U35956 ( .A(n21847), .Z(n34823) );
  XNOR U35957 ( .A(n21845), .B(n34824), .Z(n21847) );
  XNOR U35958 ( .A(q[5]), .B(DB[1860]), .Z(n34824) );
  XNOR U35959 ( .A(q[4]), .B(DB[1859]), .Z(n21845) );
  IV U35960 ( .A(n21859), .Z(n34822) );
  XOR U35961 ( .A(n34825), .B(n34826), .Z(n21859) );
  XNOR U35962 ( .A(n21855), .B(n21857), .Z(n34826) );
  XNOR U35963 ( .A(q[0]), .B(DB[1855]), .Z(n21857) );
  XNOR U35964 ( .A(q[3]), .B(DB[1858]), .Z(n21855) );
  IV U35965 ( .A(n21854), .Z(n34825) );
  XNOR U35966 ( .A(n21852), .B(n34827), .Z(n21854) );
  XNOR U35967 ( .A(q[2]), .B(DB[1857]), .Z(n34827) );
  XNOR U35968 ( .A(q[1]), .B(DB[1856]), .Z(n21852) );
  XOR U35969 ( .A(n34828), .B(n21817), .Z(n21780) );
  XOR U35970 ( .A(n34829), .B(n21805), .Z(n21817) );
  XNOR U35971 ( .A(q[6]), .B(DB[1868]), .Z(n21805) );
  IV U35972 ( .A(n21804), .Z(n34829) );
  XNOR U35973 ( .A(n21802), .B(n34830), .Z(n21804) );
  XNOR U35974 ( .A(q[5]), .B(DB[1867]), .Z(n34830) );
  XNOR U35975 ( .A(q[4]), .B(DB[1866]), .Z(n21802) );
  IV U35976 ( .A(n21816), .Z(n34828) );
  XOR U35977 ( .A(n34831), .B(n34832), .Z(n21816) );
  XNOR U35978 ( .A(n21812), .B(n21814), .Z(n34832) );
  XNOR U35979 ( .A(q[0]), .B(DB[1862]), .Z(n21814) );
  XNOR U35980 ( .A(q[3]), .B(DB[1865]), .Z(n21812) );
  IV U35981 ( .A(n21811), .Z(n34831) );
  XNOR U35982 ( .A(n21809), .B(n34833), .Z(n21811) );
  XNOR U35983 ( .A(q[2]), .B(DB[1864]), .Z(n34833) );
  XNOR U35984 ( .A(q[1]), .B(DB[1863]), .Z(n21809) );
  XOR U35985 ( .A(n34834), .B(n21774), .Z(n21737) );
  XOR U35986 ( .A(n34835), .B(n21762), .Z(n21774) );
  XNOR U35987 ( .A(q[6]), .B(DB[1875]), .Z(n21762) );
  IV U35988 ( .A(n21761), .Z(n34835) );
  XNOR U35989 ( .A(n21759), .B(n34836), .Z(n21761) );
  XNOR U35990 ( .A(q[5]), .B(DB[1874]), .Z(n34836) );
  XNOR U35991 ( .A(q[4]), .B(DB[1873]), .Z(n21759) );
  IV U35992 ( .A(n21773), .Z(n34834) );
  XOR U35993 ( .A(n34837), .B(n34838), .Z(n21773) );
  XNOR U35994 ( .A(n21769), .B(n21771), .Z(n34838) );
  XNOR U35995 ( .A(q[0]), .B(DB[1869]), .Z(n21771) );
  XNOR U35996 ( .A(q[3]), .B(DB[1872]), .Z(n21769) );
  IV U35997 ( .A(n21768), .Z(n34837) );
  XNOR U35998 ( .A(n21766), .B(n34839), .Z(n21768) );
  XNOR U35999 ( .A(q[2]), .B(DB[1871]), .Z(n34839) );
  XNOR U36000 ( .A(q[1]), .B(DB[1870]), .Z(n21766) );
  XOR U36001 ( .A(n34840), .B(n21731), .Z(n21694) );
  XOR U36002 ( .A(n34841), .B(n21719), .Z(n21731) );
  XNOR U36003 ( .A(q[6]), .B(DB[1882]), .Z(n21719) );
  IV U36004 ( .A(n21718), .Z(n34841) );
  XNOR U36005 ( .A(n21716), .B(n34842), .Z(n21718) );
  XNOR U36006 ( .A(q[5]), .B(DB[1881]), .Z(n34842) );
  XNOR U36007 ( .A(q[4]), .B(DB[1880]), .Z(n21716) );
  IV U36008 ( .A(n21730), .Z(n34840) );
  XOR U36009 ( .A(n34843), .B(n34844), .Z(n21730) );
  XNOR U36010 ( .A(n21726), .B(n21728), .Z(n34844) );
  XNOR U36011 ( .A(q[0]), .B(DB[1876]), .Z(n21728) );
  XNOR U36012 ( .A(q[3]), .B(DB[1879]), .Z(n21726) );
  IV U36013 ( .A(n21725), .Z(n34843) );
  XNOR U36014 ( .A(n21723), .B(n34845), .Z(n21725) );
  XNOR U36015 ( .A(q[2]), .B(DB[1878]), .Z(n34845) );
  XNOR U36016 ( .A(q[1]), .B(DB[1877]), .Z(n21723) );
  XOR U36017 ( .A(n34846), .B(n21688), .Z(n21651) );
  XOR U36018 ( .A(n34847), .B(n21676), .Z(n21688) );
  XNOR U36019 ( .A(q[6]), .B(DB[1889]), .Z(n21676) );
  IV U36020 ( .A(n21675), .Z(n34847) );
  XNOR U36021 ( .A(n21673), .B(n34848), .Z(n21675) );
  XNOR U36022 ( .A(q[5]), .B(DB[1888]), .Z(n34848) );
  XNOR U36023 ( .A(q[4]), .B(DB[1887]), .Z(n21673) );
  IV U36024 ( .A(n21687), .Z(n34846) );
  XOR U36025 ( .A(n34849), .B(n34850), .Z(n21687) );
  XNOR U36026 ( .A(n21683), .B(n21685), .Z(n34850) );
  XNOR U36027 ( .A(q[0]), .B(DB[1883]), .Z(n21685) );
  XNOR U36028 ( .A(q[3]), .B(DB[1886]), .Z(n21683) );
  IV U36029 ( .A(n21682), .Z(n34849) );
  XNOR U36030 ( .A(n21680), .B(n34851), .Z(n21682) );
  XNOR U36031 ( .A(q[2]), .B(DB[1885]), .Z(n34851) );
  XNOR U36032 ( .A(q[1]), .B(DB[1884]), .Z(n21680) );
  XOR U36033 ( .A(n34852), .B(n21645), .Z(n21608) );
  XOR U36034 ( .A(n34853), .B(n21633), .Z(n21645) );
  XNOR U36035 ( .A(q[6]), .B(DB[1896]), .Z(n21633) );
  IV U36036 ( .A(n21632), .Z(n34853) );
  XNOR U36037 ( .A(n21630), .B(n34854), .Z(n21632) );
  XNOR U36038 ( .A(q[5]), .B(DB[1895]), .Z(n34854) );
  XNOR U36039 ( .A(q[4]), .B(DB[1894]), .Z(n21630) );
  IV U36040 ( .A(n21644), .Z(n34852) );
  XOR U36041 ( .A(n34855), .B(n34856), .Z(n21644) );
  XNOR U36042 ( .A(n21640), .B(n21642), .Z(n34856) );
  XNOR U36043 ( .A(q[0]), .B(DB[1890]), .Z(n21642) );
  XNOR U36044 ( .A(q[3]), .B(DB[1893]), .Z(n21640) );
  IV U36045 ( .A(n21639), .Z(n34855) );
  XNOR U36046 ( .A(n21637), .B(n34857), .Z(n21639) );
  XNOR U36047 ( .A(q[2]), .B(DB[1892]), .Z(n34857) );
  XNOR U36048 ( .A(q[1]), .B(DB[1891]), .Z(n21637) );
  XOR U36049 ( .A(n34858), .B(n21602), .Z(n21565) );
  XOR U36050 ( .A(n34859), .B(n21590), .Z(n21602) );
  XNOR U36051 ( .A(q[6]), .B(DB[1903]), .Z(n21590) );
  IV U36052 ( .A(n21589), .Z(n34859) );
  XNOR U36053 ( .A(n21587), .B(n34860), .Z(n21589) );
  XNOR U36054 ( .A(q[5]), .B(DB[1902]), .Z(n34860) );
  XNOR U36055 ( .A(q[4]), .B(DB[1901]), .Z(n21587) );
  IV U36056 ( .A(n21601), .Z(n34858) );
  XOR U36057 ( .A(n34861), .B(n34862), .Z(n21601) );
  XNOR U36058 ( .A(n21597), .B(n21599), .Z(n34862) );
  XNOR U36059 ( .A(q[0]), .B(DB[1897]), .Z(n21599) );
  XNOR U36060 ( .A(q[3]), .B(DB[1900]), .Z(n21597) );
  IV U36061 ( .A(n21596), .Z(n34861) );
  XNOR U36062 ( .A(n21594), .B(n34863), .Z(n21596) );
  XNOR U36063 ( .A(q[2]), .B(DB[1899]), .Z(n34863) );
  XNOR U36064 ( .A(q[1]), .B(DB[1898]), .Z(n21594) );
  XOR U36065 ( .A(n34864), .B(n21559), .Z(n21522) );
  XOR U36066 ( .A(n34865), .B(n21547), .Z(n21559) );
  XNOR U36067 ( .A(q[6]), .B(DB[1910]), .Z(n21547) );
  IV U36068 ( .A(n21546), .Z(n34865) );
  XNOR U36069 ( .A(n21544), .B(n34866), .Z(n21546) );
  XNOR U36070 ( .A(q[5]), .B(DB[1909]), .Z(n34866) );
  XNOR U36071 ( .A(q[4]), .B(DB[1908]), .Z(n21544) );
  IV U36072 ( .A(n21558), .Z(n34864) );
  XOR U36073 ( .A(n34867), .B(n34868), .Z(n21558) );
  XNOR U36074 ( .A(n21554), .B(n21556), .Z(n34868) );
  XNOR U36075 ( .A(q[0]), .B(DB[1904]), .Z(n21556) );
  XNOR U36076 ( .A(q[3]), .B(DB[1907]), .Z(n21554) );
  IV U36077 ( .A(n21553), .Z(n34867) );
  XNOR U36078 ( .A(n21551), .B(n34869), .Z(n21553) );
  XNOR U36079 ( .A(q[2]), .B(DB[1906]), .Z(n34869) );
  XNOR U36080 ( .A(q[1]), .B(DB[1905]), .Z(n21551) );
  XOR U36081 ( .A(n34870), .B(n21516), .Z(n21479) );
  XOR U36082 ( .A(n34871), .B(n21504), .Z(n21516) );
  XNOR U36083 ( .A(q[6]), .B(DB[1917]), .Z(n21504) );
  IV U36084 ( .A(n21503), .Z(n34871) );
  XNOR U36085 ( .A(n21501), .B(n34872), .Z(n21503) );
  XNOR U36086 ( .A(q[5]), .B(DB[1916]), .Z(n34872) );
  XNOR U36087 ( .A(q[4]), .B(DB[1915]), .Z(n21501) );
  IV U36088 ( .A(n21515), .Z(n34870) );
  XOR U36089 ( .A(n34873), .B(n34874), .Z(n21515) );
  XNOR U36090 ( .A(n21511), .B(n21513), .Z(n34874) );
  XNOR U36091 ( .A(q[0]), .B(DB[1911]), .Z(n21513) );
  XNOR U36092 ( .A(q[3]), .B(DB[1914]), .Z(n21511) );
  IV U36093 ( .A(n21510), .Z(n34873) );
  XNOR U36094 ( .A(n21508), .B(n34875), .Z(n21510) );
  XNOR U36095 ( .A(q[2]), .B(DB[1913]), .Z(n34875) );
  XNOR U36096 ( .A(q[1]), .B(DB[1912]), .Z(n21508) );
  XOR U36097 ( .A(n34876), .B(n21473), .Z(n21436) );
  XOR U36098 ( .A(n34877), .B(n21461), .Z(n21473) );
  XNOR U36099 ( .A(q[6]), .B(DB[1924]), .Z(n21461) );
  IV U36100 ( .A(n21460), .Z(n34877) );
  XNOR U36101 ( .A(n21458), .B(n34878), .Z(n21460) );
  XNOR U36102 ( .A(q[5]), .B(DB[1923]), .Z(n34878) );
  XNOR U36103 ( .A(q[4]), .B(DB[1922]), .Z(n21458) );
  IV U36104 ( .A(n21472), .Z(n34876) );
  XOR U36105 ( .A(n34879), .B(n34880), .Z(n21472) );
  XNOR U36106 ( .A(n21468), .B(n21470), .Z(n34880) );
  XNOR U36107 ( .A(q[0]), .B(DB[1918]), .Z(n21470) );
  XNOR U36108 ( .A(q[3]), .B(DB[1921]), .Z(n21468) );
  IV U36109 ( .A(n21467), .Z(n34879) );
  XNOR U36110 ( .A(n21465), .B(n34881), .Z(n21467) );
  XNOR U36111 ( .A(q[2]), .B(DB[1920]), .Z(n34881) );
  XNOR U36112 ( .A(q[1]), .B(DB[1919]), .Z(n21465) );
  XOR U36113 ( .A(n34882), .B(n21430), .Z(n21393) );
  XOR U36114 ( .A(n34883), .B(n21418), .Z(n21430) );
  XNOR U36115 ( .A(q[6]), .B(DB[1931]), .Z(n21418) );
  IV U36116 ( .A(n21417), .Z(n34883) );
  XNOR U36117 ( .A(n21415), .B(n34884), .Z(n21417) );
  XNOR U36118 ( .A(q[5]), .B(DB[1930]), .Z(n34884) );
  XNOR U36119 ( .A(q[4]), .B(DB[1929]), .Z(n21415) );
  IV U36120 ( .A(n21429), .Z(n34882) );
  XOR U36121 ( .A(n34885), .B(n34886), .Z(n21429) );
  XNOR U36122 ( .A(n21425), .B(n21427), .Z(n34886) );
  XNOR U36123 ( .A(q[0]), .B(DB[1925]), .Z(n21427) );
  XNOR U36124 ( .A(q[3]), .B(DB[1928]), .Z(n21425) );
  IV U36125 ( .A(n21424), .Z(n34885) );
  XNOR U36126 ( .A(n21422), .B(n34887), .Z(n21424) );
  XNOR U36127 ( .A(q[2]), .B(DB[1927]), .Z(n34887) );
  XNOR U36128 ( .A(q[1]), .B(DB[1926]), .Z(n21422) );
  XOR U36129 ( .A(n34888), .B(n21387), .Z(n21350) );
  XOR U36130 ( .A(n34889), .B(n21375), .Z(n21387) );
  XNOR U36131 ( .A(q[6]), .B(DB[1938]), .Z(n21375) );
  IV U36132 ( .A(n21374), .Z(n34889) );
  XNOR U36133 ( .A(n21372), .B(n34890), .Z(n21374) );
  XNOR U36134 ( .A(q[5]), .B(DB[1937]), .Z(n34890) );
  XNOR U36135 ( .A(q[4]), .B(DB[1936]), .Z(n21372) );
  IV U36136 ( .A(n21386), .Z(n34888) );
  XOR U36137 ( .A(n34891), .B(n34892), .Z(n21386) );
  XNOR U36138 ( .A(n21382), .B(n21384), .Z(n34892) );
  XNOR U36139 ( .A(q[0]), .B(DB[1932]), .Z(n21384) );
  XNOR U36140 ( .A(q[3]), .B(DB[1935]), .Z(n21382) );
  IV U36141 ( .A(n21381), .Z(n34891) );
  XNOR U36142 ( .A(n21379), .B(n34893), .Z(n21381) );
  XNOR U36143 ( .A(q[2]), .B(DB[1934]), .Z(n34893) );
  XNOR U36144 ( .A(q[1]), .B(DB[1933]), .Z(n21379) );
  XOR U36145 ( .A(n34894), .B(n21344), .Z(n21307) );
  XOR U36146 ( .A(n34895), .B(n21332), .Z(n21344) );
  XNOR U36147 ( .A(q[6]), .B(DB[1945]), .Z(n21332) );
  IV U36148 ( .A(n21331), .Z(n34895) );
  XNOR U36149 ( .A(n21329), .B(n34896), .Z(n21331) );
  XNOR U36150 ( .A(q[5]), .B(DB[1944]), .Z(n34896) );
  XNOR U36151 ( .A(q[4]), .B(DB[1943]), .Z(n21329) );
  IV U36152 ( .A(n21343), .Z(n34894) );
  XOR U36153 ( .A(n34897), .B(n34898), .Z(n21343) );
  XNOR U36154 ( .A(n21339), .B(n21341), .Z(n34898) );
  XNOR U36155 ( .A(q[0]), .B(DB[1939]), .Z(n21341) );
  XNOR U36156 ( .A(q[3]), .B(DB[1942]), .Z(n21339) );
  IV U36157 ( .A(n21338), .Z(n34897) );
  XNOR U36158 ( .A(n21336), .B(n34899), .Z(n21338) );
  XNOR U36159 ( .A(q[2]), .B(DB[1941]), .Z(n34899) );
  XNOR U36160 ( .A(q[1]), .B(DB[1940]), .Z(n21336) );
  XOR U36161 ( .A(n34900), .B(n21301), .Z(n21264) );
  XOR U36162 ( .A(n34901), .B(n21289), .Z(n21301) );
  XNOR U36163 ( .A(q[6]), .B(DB[1952]), .Z(n21289) );
  IV U36164 ( .A(n21288), .Z(n34901) );
  XNOR U36165 ( .A(n21286), .B(n34902), .Z(n21288) );
  XNOR U36166 ( .A(q[5]), .B(DB[1951]), .Z(n34902) );
  XNOR U36167 ( .A(q[4]), .B(DB[1950]), .Z(n21286) );
  IV U36168 ( .A(n21300), .Z(n34900) );
  XOR U36169 ( .A(n34903), .B(n34904), .Z(n21300) );
  XNOR U36170 ( .A(n21296), .B(n21298), .Z(n34904) );
  XNOR U36171 ( .A(q[0]), .B(DB[1946]), .Z(n21298) );
  XNOR U36172 ( .A(q[3]), .B(DB[1949]), .Z(n21296) );
  IV U36173 ( .A(n21295), .Z(n34903) );
  XNOR U36174 ( .A(n21293), .B(n34905), .Z(n21295) );
  XNOR U36175 ( .A(q[2]), .B(DB[1948]), .Z(n34905) );
  XNOR U36176 ( .A(q[1]), .B(DB[1947]), .Z(n21293) );
  XOR U36177 ( .A(n34906), .B(n21258), .Z(n21221) );
  XOR U36178 ( .A(n34907), .B(n21246), .Z(n21258) );
  XNOR U36179 ( .A(q[6]), .B(DB[1959]), .Z(n21246) );
  IV U36180 ( .A(n21245), .Z(n34907) );
  XNOR U36181 ( .A(n21243), .B(n34908), .Z(n21245) );
  XNOR U36182 ( .A(q[5]), .B(DB[1958]), .Z(n34908) );
  XNOR U36183 ( .A(q[4]), .B(DB[1957]), .Z(n21243) );
  IV U36184 ( .A(n21257), .Z(n34906) );
  XOR U36185 ( .A(n34909), .B(n34910), .Z(n21257) );
  XNOR U36186 ( .A(n21253), .B(n21255), .Z(n34910) );
  XNOR U36187 ( .A(q[0]), .B(DB[1953]), .Z(n21255) );
  XNOR U36188 ( .A(q[3]), .B(DB[1956]), .Z(n21253) );
  IV U36189 ( .A(n21252), .Z(n34909) );
  XNOR U36190 ( .A(n21250), .B(n34911), .Z(n21252) );
  XNOR U36191 ( .A(q[2]), .B(DB[1955]), .Z(n34911) );
  XNOR U36192 ( .A(q[1]), .B(DB[1954]), .Z(n21250) );
  XOR U36193 ( .A(n34912), .B(n21215), .Z(n21178) );
  XOR U36194 ( .A(n34913), .B(n21203), .Z(n21215) );
  XNOR U36195 ( .A(q[6]), .B(DB[1966]), .Z(n21203) );
  IV U36196 ( .A(n21202), .Z(n34913) );
  XNOR U36197 ( .A(n21200), .B(n34914), .Z(n21202) );
  XNOR U36198 ( .A(q[5]), .B(DB[1965]), .Z(n34914) );
  XNOR U36199 ( .A(q[4]), .B(DB[1964]), .Z(n21200) );
  IV U36200 ( .A(n21214), .Z(n34912) );
  XOR U36201 ( .A(n34915), .B(n34916), .Z(n21214) );
  XNOR U36202 ( .A(n21210), .B(n21212), .Z(n34916) );
  XNOR U36203 ( .A(q[0]), .B(DB[1960]), .Z(n21212) );
  XNOR U36204 ( .A(q[3]), .B(DB[1963]), .Z(n21210) );
  IV U36205 ( .A(n21209), .Z(n34915) );
  XNOR U36206 ( .A(n21207), .B(n34917), .Z(n21209) );
  XNOR U36207 ( .A(q[2]), .B(DB[1962]), .Z(n34917) );
  XNOR U36208 ( .A(q[1]), .B(DB[1961]), .Z(n21207) );
  XOR U36209 ( .A(n34918), .B(n21172), .Z(n21135) );
  XOR U36210 ( .A(n34919), .B(n21160), .Z(n21172) );
  XNOR U36211 ( .A(q[6]), .B(DB[1973]), .Z(n21160) );
  IV U36212 ( .A(n21159), .Z(n34919) );
  XNOR U36213 ( .A(n21157), .B(n34920), .Z(n21159) );
  XNOR U36214 ( .A(q[5]), .B(DB[1972]), .Z(n34920) );
  XNOR U36215 ( .A(q[4]), .B(DB[1971]), .Z(n21157) );
  IV U36216 ( .A(n21171), .Z(n34918) );
  XOR U36217 ( .A(n34921), .B(n34922), .Z(n21171) );
  XNOR U36218 ( .A(n21167), .B(n21169), .Z(n34922) );
  XNOR U36219 ( .A(q[0]), .B(DB[1967]), .Z(n21169) );
  XNOR U36220 ( .A(q[3]), .B(DB[1970]), .Z(n21167) );
  IV U36221 ( .A(n21166), .Z(n34921) );
  XNOR U36222 ( .A(n21164), .B(n34923), .Z(n21166) );
  XNOR U36223 ( .A(q[2]), .B(DB[1969]), .Z(n34923) );
  XNOR U36224 ( .A(q[1]), .B(DB[1968]), .Z(n21164) );
  XOR U36225 ( .A(n34924), .B(n21129), .Z(n21092) );
  XOR U36226 ( .A(n34925), .B(n21117), .Z(n21129) );
  XNOR U36227 ( .A(q[6]), .B(DB[1980]), .Z(n21117) );
  IV U36228 ( .A(n21116), .Z(n34925) );
  XNOR U36229 ( .A(n21114), .B(n34926), .Z(n21116) );
  XNOR U36230 ( .A(q[5]), .B(DB[1979]), .Z(n34926) );
  XNOR U36231 ( .A(q[4]), .B(DB[1978]), .Z(n21114) );
  IV U36232 ( .A(n21128), .Z(n34924) );
  XOR U36233 ( .A(n34927), .B(n34928), .Z(n21128) );
  XNOR U36234 ( .A(n21124), .B(n21126), .Z(n34928) );
  XNOR U36235 ( .A(q[0]), .B(DB[1974]), .Z(n21126) );
  XNOR U36236 ( .A(q[3]), .B(DB[1977]), .Z(n21124) );
  IV U36237 ( .A(n21123), .Z(n34927) );
  XNOR U36238 ( .A(n21121), .B(n34929), .Z(n21123) );
  XNOR U36239 ( .A(q[2]), .B(DB[1976]), .Z(n34929) );
  XNOR U36240 ( .A(q[1]), .B(DB[1975]), .Z(n21121) );
  XOR U36241 ( .A(n34930), .B(n21086), .Z(n21049) );
  XOR U36242 ( .A(n34931), .B(n21074), .Z(n21086) );
  XNOR U36243 ( .A(q[6]), .B(DB[1987]), .Z(n21074) );
  IV U36244 ( .A(n21073), .Z(n34931) );
  XNOR U36245 ( .A(n21071), .B(n34932), .Z(n21073) );
  XNOR U36246 ( .A(q[5]), .B(DB[1986]), .Z(n34932) );
  XNOR U36247 ( .A(q[4]), .B(DB[1985]), .Z(n21071) );
  IV U36248 ( .A(n21085), .Z(n34930) );
  XOR U36249 ( .A(n34933), .B(n34934), .Z(n21085) );
  XNOR U36250 ( .A(n21081), .B(n21083), .Z(n34934) );
  XNOR U36251 ( .A(q[0]), .B(DB[1981]), .Z(n21083) );
  XNOR U36252 ( .A(q[3]), .B(DB[1984]), .Z(n21081) );
  IV U36253 ( .A(n21080), .Z(n34933) );
  XNOR U36254 ( .A(n21078), .B(n34935), .Z(n21080) );
  XNOR U36255 ( .A(q[2]), .B(DB[1983]), .Z(n34935) );
  XNOR U36256 ( .A(q[1]), .B(DB[1982]), .Z(n21078) );
  XOR U36257 ( .A(n34936), .B(n21043), .Z(n21006) );
  XOR U36258 ( .A(n34937), .B(n21031), .Z(n21043) );
  XNOR U36259 ( .A(q[6]), .B(DB[1994]), .Z(n21031) );
  IV U36260 ( .A(n21030), .Z(n34937) );
  XNOR U36261 ( .A(n21028), .B(n34938), .Z(n21030) );
  XNOR U36262 ( .A(q[5]), .B(DB[1993]), .Z(n34938) );
  XNOR U36263 ( .A(q[4]), .B(DB[1992]), .Z(n21028) );
  IV U36264 ( .A(n21042), .Z(n34936) );
  XOR U36265 ( .A(n34939), .B(n34940), .Z(n21042) );
  XNOR U36266 ( .A(n21038), .B(n21040), .Z(n34940) );
  XNOR U36267 ( .A(q[0]), .B(DB[1988]), .Z(n21040) );
  XNOR U36268 ( .A(q[3]), .B(DB[1991]), .Z(n21038) );
  IV U36269 ( .A(n21037), .Z(n34939) );
  XNOR U36270 ( .A(n21035), .B(n34941), .Z(n21037) );
  XNOR U36271 ( .A(q[2]), .B(DB[1990]), .Z(n34941) );
  XNOR U36272 ( .A(q[1]), .B(DB[1989]), .Z(n21035) );
  XOR U36273 ( .A(n34942), .B(n21000), .Z(n20963) );
  XOR U36274 ( .A(n34943), .B(n20988), .Z(n21000) );
  XNOR U36275 ( .A(q[6]), .B(DB[2001]), .Z(n20988) );
  IV U36276 ( .A(n20987), .Z(n34943) );
  XNOR U36277 ( .A(n20985), .B(n34944), .Z(n20987) );
  XNOR U36278 ( .A(q[5]), .B(DB[2000]), .Z(n34944) );
  XNOR U36279 ( .A(q[4]), .B(DB[1999]), .Z(n20985) );
  IV U36280 ( .A(n20999), .Z(n34942) );
  XOR U36281 ( .A(n34945), .B(n34946), .Z(n20999) );
  XNOR U36282 ( .A(n20995), .B(n20997), .Z(n34946) );
  XNOR U36283 ( .A(q[0]), .B(DB[1995]), .Z(n20997) );
  XNOR U36284 ( .A(q[3]), .B(DB[1998]), .Z(n20995) );
  IV U36285 ( .A(n20994), .Z(n34945) );
  XNOR U36286 ( .A(n20992), .B(n34947), .Z(n20994) );
  XNOR U36287 ( .A(q[2]), .B(DB[1997]), .Z(n34947) );
  XNOR U36288 ( .A(q[1]), .B(DB[1996]), .Z(n20992) );
  XOR U36289 ( .A(n34948), .B(n20957), .Z(n20920) );
  XOR U36290 ( .A(n34949), .B(n20945), .Z(n20957) );
  XNOR U36291 ( .A(q[6]), .B(DB[2008]), .Z(n20945) );
  IV U36292 ( .A(n20944), .Z(n34949) );
  XNOR U36293 ( .A(n20942), .B(n34950), .Z(n20944) );
  XNOR U36294 ( .A(q[5]), .B(DB[2007]), .Z(n34950) );
  XNOR U36295 ( .A(q[4]), .B(DB[2006]), .Z(n20942) );
  IV U36296 ( .A(n20956), .Z(n34948) );
  XOR U36297 ( .A(n34951), .B(n34952), .Z(n20956) );
  XNOR U36298 ( .A(n20952), .B(n20954), .Z(n34952) );
  XNOR U36299 ( .A(q[0]), .B(DB[2002]), .Z(n20954) );
  XNOR U36300 ( .A(q[3]), .B(DB[2005]), .Z(n20952) );
  IV U36301 ( .A(n20951), .Z(n34951) );
  XNOR U36302 ( .A(n20949), .B(n34953), .Z(n20951) );
  XNOR U36303 ( .A(q[2]), .B(DB[2004]), .Z(n34953) );
  XNOR U36304 ( .A(q[1]), .B(DB[2003]), .Z(n20949) );
  XOR U36305 ( .A(n34954), .B(n20914), .Z(n20877) );
  XOR U36306 ( .A(n34955), .B(n20902), .Z(n20914) );
  XNOR U36307 ( .A(q[6]), .B(DB[2015]), .Z(n20902) );
  IV U36308 ( .A(n20901), .Z(n34955) );
  XNOR U36309 ( .A(n20899), .B(n34956), .Z(n20901) );
  XNOR U36310 ( .A(q[5]), .B(DB[2014]), .Z(n34956) );
  XNOR U36311 ( .A(q[4]), .B(DB[2013]), .Z(n20899) );
  IV U36312 ( .A(n20913), .Z(n34954) );
  XOR U36313 ( .A(n34957), .B(n34958), .Z(n20913) );
  XNOR U36314 ( .A(n20909), .B(n20911), .Z(n34958) );
  XNOR U36315 ( .A(q[0]), .B(DB[2009]), .Z(n20911) );
  XNOR U36316 ( .A(q[3]), .B(DB[2012]), .Z(n20909) );
  IV U36317 ( .A(n20908), .Z(n34957) );
  XNOR U36318 ( .A(n20906), .B(n34959), .Z(n20908) );
  XNOR U36319 ( .A(q[2]), .B(DB[2011]), .Z(n34959) );
  XNOR U36320 ( .A(q[1]), .B(DB[2010]), .Z(n20906) );
  XOR U36321 ( .A(n34960), .B(n20871), .Z(n20834) );
  XOR U36322 ( .A(n34961), .B(n20859), .Z(n20871) );
  XNOR U36323 ( .A(q[6]), .B(DB[2022]), .Z(n20859) );
  IV U36324 ( .A(n20858), .Z(n34961) );
  XNOR U36325 ( .A(n20856), .B(n34962), .Z(n20858) );
  XNOR U36326 ( .A(q[5]), .B(DB[2021]), .Z(n34962) );
  XNOR U36327 ( .A(q[4]), .B(DB[2020]), .Z(n20856) );
  IV U36328 ( .A(n20870), .Z(n34960) );
  XOR U36329 ( .A(n34963), .B(n34964), .Z(n20870) );
  XNOR U36330 ( .A(n20866), .B(n20868), .Z(n34964) );
  XNOR U36331 ( .A(q[0]), .B(DB[2016]), .Z(n20868) );
  XNOR U36332 ( .A(q[3]), .B(DB[2019]), .Z(n20866) );
  IV U36333 ( .A(n20865), .Z(n34963) );
  XNOR U36334 ( .A(n20863), .B(n34965), .Z(n20865) );
  XNOR U36335 ( .A(q[2]), .B(DB[2018]), .Z(n34965) );
  XNOR U36336 ( .A(q[1]), .B(DB[2017]), .Z(n20863) );
  XOR U36337 ( .A(n34966), .B(n20828), .Z(n20791) );
  XOR U36338 ( .A(n34967), .B(n20816), .Z(n20828) );
  XNOR U36339 ( .A(q[6]), .B(DB[2029]), .Z(n20816) );
  IV U36340 ( .A(n20815), .Z(n34967) );
  XNOR U36341 ( .A(n20813), .B(n34968), .Z(n20815) );
  XNOR U36342 ( .A(q[5]), .B(DB[2028]), .Z(n34968) );
  XNOR U36343 ( .A(q[4]), .B(DB[2027]), .Z(n20813) );
  IV U36344 ( .A(n20827), .Z(n34966) );
  XOR U36345 ( .A(n34969), .B(n34970), .Z(n20827) );
  XNOR U36346 ( .A(n20823), .B(n20825), .Z(n34970) );
  XNOR U36347 ( .A(q[0]), .B(DB[2023]), .Z(n20825) );
  XNOR U36348 ( .A(q[3]), .B(DB[2026]), .Z(n20823) );
  IV U36349 ( .A(n20822), .Z(n34969) );
  XNOR U36350 ( .A(n20820), .B(n34971), .Z(n20822) );
  XNOR U36351 ( .A(q[2]), .B(DB[2025]), .Z(n34971) );
  XNOR U36352 ( .A(q[1]), .B(DB[2024]), .Z(n20820) );
  XOR U36353 ( .A(n34972), .B(n20785), .Z(n20748) );
  XOR U36354 ( .A(n34973), .B(n20773), .Z(n20785) );
  XNOR U36355 ( .A(q[6]), .B(DB[2036]), .Z(n20773) );
  IV U36356 ( .A(n20772), .Z(n34973) );
  XNOR U36357 ( .A(n20770), .B(n34974), .Z(n20772) );
  XNOR U36358 ( .A(q[5]), .B(DB[2035]), .Z(n34974) );
  XNOR U36359 ( .A(q[4]), .B(DB[2034]), .Z(n20770) );
  IV U36360 ( .A(n20784), .Z(n34972) );
  XOR U36361 ( .A(n34975), .B(n34976), .Z(n20784) );
  XNOR U36362 ( .A(n20780), .B(n20782), .Z(n34976) );
  XNOR U36363 ( .A(q[0]), .B(DB[2030]), .Z(n20782) );
  XNOR U36364 ( .A(q[3]), .B(DB[2033]), .Z(n20780) );
  IV U36365 ( .A(n20779), .Z(n34975) );
  XNOR U36366 ( .A(n20777), .B(n34977), .Z(n20779) );
  XNOR U36367 ( .A(q[2]), .B(DB[2032]), .Z(n34977) );
  XNOR U36368 ( .A(q[1]), .B(DB[2031]), .Z(n20777) );
  XOR U36369 ( .A(n34978), .B(n20742), .Z(n20705) );
  XOR U36370 ( .A(n34979), .B(n20730), .Z(n20742) );
  XNOR U36371 ( .A(q[6]), .B(DB[2043]), .Z(n20730) );
  IV U36372 ( .A(n20729), .Z(n34979) );
  XNOR U36373 ( .A(n20727), .B(n34980), .Z(n20729) );
  XNOR U36374 ( .A(q[5]), .B(DB[2042]), .Z(n34980) );
  XNOR U36375 ( .A(q[4]), .B(DB[2041]), .Z(n20727) );
  IV U36376 ( .A(n20741), .Z(n34978) );
  XOR U36377 ( .A(n34981), .B(n34982), .Z(n20741) );
  XNOR U36378 ( .A(n20737), .B(n20739), .Z(n34982) );
  XNOR U36379 ( .A(q[0]), .B(DB[2037]), .Z(n20739) );
  XNOR U36380 ( .A(q[3]), .B(DB[2040]), .Z(n20737) );
  IV U36381 ( .A(n20736), .Z(n34981) );
  XNOR U36382 ( .A(n20734), .B(n34983), .Z(n20736) );
  XNOR U36383 ( .A(q[2]), .B(DB[2039]), .Z(n34983) );
  XNOR U36384 ( .A(q[1]), .B(DB[2038]), .Z(n20734) );
  XOR U36385 ( .A(n34984), .B(n20699), .Z(n20662) );
  XOR U36386 ( .A(n34985), .B(n20687), .Z(n20699) );
  XNOR U36387 ( .A(q[6]), .B(DB[2050]), .Z(n20687) );
  IV U36388 ( .A(n20686), .Z(n34985) );
  XNOR U36389 ( .A(n20684), .B(n34986), .Z(n20686) );
  XNOR U36390 ( .A(q[5]), .B(DB[2049]), .Z(n34986) );
  XNOR U36391 ( .A(q[4]), .B(DB[2048]), .Z(n20684) );
  IV U36392 ( .A(n20698), .Z(n34984) );
  XOR U36393 ( .A(n34987), .B(n34988), .Z(n20698) );
  XNOR U36394 ( .A(n20694), .B(n20696), .Z(n34988) );
  XNOR U36395 ( .A(q[0]), .B(DB[2044]), .Z(n20696) );
  XNOR U36396 ( .A(q[3]), .B(DB[2047]), .Z(n20694) );
  IV U36397 ( .A(n20693), .Z(n34987) );
  XNOR U36398 ( .A(n20691), .B(n34989), .Z(n20693) );
  XNOR U36399 ( .A(q[2]), .B(DB[2046]), .Z(n34989) );
  XNOR U36400 ( .A(q[1]), .B(DB[2045]), .Z(n20691) );
  XOR U36401 ( .A(n34990), .B(n20656), .Z(n20619) );
  XOR U36402 ( .A(n34991), .B(n20644), .Z(n20656) );
  XNOR U36403 ( .A(q[6]), .B(DB[2057]), .Z(n20644) );
  IV U36404 ( .A(n20643), .Z(n34991) );
  XNOR U36405 ( .A(n20641), .B(n34992), .Z(n20643) );
  XNOR U36406 ( .A(q[5]), .B(DB[2056]), .Z(n34992) );
  XNOR U36407 ( .A(q[4]), .B(DB[2055]), .Z(n20641) );
  IV U36408 ( .A(n20655), .Z(n34990) );
  XOR U36409 ( .A(n34993), .B(n34994), .Z(n20655) );
  XNOR U36410 ( .A(n20651), .B(n20653), .Z(n34994) );
  XNOR U36411 ( .A(q[0]), .B(DB[2051]), .Z(n20653) );
  XNOR U36412 ( .A(q[3]), .B(DB[2054]), .Z(n20651) );
  IV U36413 ( .A(n20650), .Z(n34993) );
  XNOR U36414 ( .A(n20648), .B(n34995), .Z(n20650) );
  XNOR U36415 ( .A(q[2]), .B(DB[2053]), .Z(n34995) );
  XNOR U36416 ( .A(q[1]), .B(DB[2052]), .Z(n20648) );
  XOR U36417 ( .A(n34996), .B(n20613), .Z(n20576) );
  XOR U36418 ( .A(n34997), .B(n20601), .Z(n20613) );
  XNOR U36419 ( .A(q[6]), .B(DB[2064]), .Z(n20601) );
  IV U36420 ( .A(n20600), .Z(n34997) );
  XNOR U36421 ( .A(n20598), .B(n34998), .Z(n20600) );
  XNOR U36422 ( .A(q[5]), .B(DB[2063]), .Z(n34998) );
  XNOR U36423 ( .A(q[4]), .B(DB[2062]), .Z(n20598) );
  IV U36424 ( .A(n20612), .Z(n34996) );
  XOR U36425 ( .A(n34999), .B(n35000), .Z(n20612) );
  XNOR U36426 ( .A(n20608), .B(n20610), .Z(n35000) );
  XNOR U36427 ( .A(q[0]), .B(DB[2058]), .Z(n20610) );
  XNOR U36428 ( .A(q[3]), .B(DB[2061]), .Z(n20608) );
  IV U36429 ( .A(n20607), .Z(n34999) );
  XNOR U36430 ( .A(n20605), .B(n35001), .Z(n20607) );
  XNOR U36431 ( .A(q[2]), .B(DB[2060]), .Z(n35001) );
  XNOR U36432 ( .A(q[1]), .B(DB[2059]), .Z(n20605) );
  XOR U36433 ( .A(n35002), .B(n20570), .Z(n20533) );
  XOR U36434 ( .A(n35003), .B(n20558), .Z(n20570) );
  XNOR U36435 ( .A(q[6]), .B(DB[2071]), .Z(n20558) );
  IV U36436 ( .A(n20557), .Z(n35003) );
  XNOR U36437 ( .A(n20555), .B(n35004), .Z(n20557) );
  XNOR U36438 ( .A(q[5]), .B(DB[2070]), .Z(n35004) );
  XNOR U36439 ( .A(q[4]), .B(DB[2069]), .Z(n20555) );
  IV U36440 ( .A(n20569), .Z(n35002) );
  XOR U36441 ( .A(n35005), .B(n35006), .Z(n20569) );
  XNOR U36442 ( .A(n20565), .B(n20567), .Z(n35006) );
  XNOR U36443 ( .A(q[0]), .B(DB[2065]), .Z(n20567) );
  XNOR U36444 ( .A(q[3]), .B(DB[2068]), .Z(n20565) );
  IV U36445 ( .A(n20564), .Z(n35005) );
  XNOR U36446 ( .A(n20562), .B(n35007), .Z(n20564) );
  XNOR U36447 ( .A(q[2]), .B(DB[2067]), .Z(n35007) );
  XNOR U36448 ( .A(q[1]), .B(DB[2066]), .Z(n20562) );
  XOR U36449 ( .A(n35008), .B(n20527), .Z(n20490) );
  XOR U36450 ( .A(n35009), .B(n20515), .Z(n20527) );
  XNOR U36451 ( .A(q[6]), .B(DB[2078]), .Z(n20515) );
  IV U36452 ( .A(n20514), .Z(n35009) );
  XNOR U36453 ( .A(n20512), .B(n35010), .Z(n20514) );
  XNOR U36454 ( .A(q[5]), .B(DB[2077]), .Z(n35010) );
  XNOR U36455 ( .A(q[4]), .B(DB[2076]), .Z(n20512) );
  IV U36456 ( .A(n20526), .Z(n35008) );
  XOR U36457 ( .A(n35011), .B(n35012), .Z(n20526) );
  XNOR U36458 ( .A(n20522), .B(n20524), .Z(n35012) );
  XNOR U36459 ( .A(q[0]), .B(DB[2072]), .Z(n20524) );
  XNOR U36460 ( .A(q[3]), .B(DB[2075]), .Z(n20522) );
  IV U36461 ( .A(n20521), .Z(n35011) );
  XNOR U36462 ( .A(n20519), .B(n35013), .Z(n20521) );
  XNOR U36463 ( .A(q[2]), .B(DB[2074]), .Z(n35013) );
  XNOR U36464 ( .A(q[1]), .B(DB[2073]), .Z(n20519) );
  XOR U36465 ( .A(n35014), .B(n20484), .Z(n20447) );
  XOR U36466 ( .A(n35015), .B(n20472), .Z(n20484) );
  XNOR U36467 ( .A(q[6]), .B(DB[2085]), .Z(n20472) );
  IV U36468 ( .A(n20471), .Z(n35015) );
  XNOR U36469 ( .A(n20469), .B(n35016), .Z(n20471) );
  XNOR U36470 ( .A(q[5]), .B(DB[2084]), .Z(n35016) );
  XNOR U36471 ( .A(q[4]), .B(DB[2083]), .Z(n20469) );
  IV U36472 ( .A(n20483), .Z(n35014) );
  XOR U36473 ( .A(n35017), .B(n35018), .Z(n20483) );
  XNOR U36474 ( .A(n20479), .B(n20481), .Z(n35018) );
  XNOR U36475 ( .A(q[0]), .B(DB[2079]), .Z(n20481) );
  XNOR U36476 ( .A(q[3]), .B(DB[2082]), .Z(n20479) );
  IV U36477 ( .A(n20478), .Z(n35017) );
  XNOR U36478 ( .A(n20476), .B(n35019), .Z(n20478) );
  XNOR U36479 ( .A(q[2]), .B(DB[2081]), .Z(n35019) );
  XNOR U36480 ( .A(q[1]), .B(DB[2080]), .Z(n20476) );
  XOR U36481 ( .A(n35020), .B(n20441), .Z(n20404) );
  XOR U36482 ( .A(n35021), .B(n20429), .Z(n20441) );
  XNOR U36483 ( .A(q[6]), .B(DB[2092]), .Z(n20429) );
  IV U36484 ( .A(n20428), .Z(n35021) );
  XNOR U36485 ( .A(n20426), .B(n35022), .Z(n20428) );
  XNOR U36486 ( .A(q[5]), .B(DB[2091]), .Z(n35022) );
  XNOR U36487 ( .A(q[4]), .B(DB[2090]), .Z(n20426) );
  IV U36488 ( .A(n20440), .Z(n35020) );
  XOR U36489 ( .A(n35023), .B(n35024), .Z(n20440) );
  XNOR U36490 ( .A(n20436), .B(n20438), .Z(n35024) );
  XNOR U36491 ( .A(q[0]), .B(DB[2086]), .Z(n20438) );
  XNOR U36492 ( .A(q[3]), .B(DB[2089]), .Z(n20436) );
  IV U36493 ( .A(n20435), .Z(n35023) );
  XNOR U36494 ( .A(n20433), .B(n35025), .Z(n20435) );
  XNOR U36495 ( .A(q[2]), .B(DB[2088]), .Z(n35025) );
  XNOR U36496 ( .A(q[1]), .B(DB[2087]), .Z(n20433) );
  XOR U36497 ( .A(n35026), .B(n20398), .Z(n20361) );
  XOR U36498 ( .A(n35027), .B(n20386), .Z(n20398) );
  XNOR U36499 ( .A(q[6]), .B(DB[2099]), .Z(n20386) );
  IV U36500 ( .A(n20385), .Z(n35027) );
  XNOR U36501 ( .A(n20383), .B(n35028), .Z(n20385) );
  XNOR U36502 ( .A(q[5]), .B(DB[2098]), .Z(n35028) );
  XNOR U36503 ( .A(q[4]), .B(DB[2097]), .Z(n20383) );
  IV U36504 ( .A(n20397), .Z(n35026) );
  XOR U36505 ( .A(n35029), .B(n35030), .Z(n20397) );
  XNOR U36506 ( .A(n20393), .B(n20395), .Z(n35030) );
  XNOR U36507 ( .A(q[0]), .B(DB[2093]), .Z(n20395) );
  XNOR U36508 ( .A(q[3]), .B(DB[2096]), .Z(n20393) );
  IV U36509 ( .A(n20392), .Z(n35029) );
  XNOR U36510 ( .A(n20390), .B(n35031), .Z(n20392) );
  XNOR U36511 ( .A(q[2]), .B(DB[2095]), .Z(n35031) );
  XNOR U36512 ( .A(q[1]), .B(DB[2094]), .Z(n20390) );
  XOR U36513 ( .A(n35032), .B(n20355), .Z(n20318) );
  XOR U36514 ( .A(n35033), .B(n20343), .Z(n20355) );
  XNOR U36515 ( .A(q[6]), .B(DB[2106]), .Z(n20343) );
  IV U36516 ( .A(n20342), .Z(n35033) );
  XNOR U36517 ( .A(n20340), .B(n35034), .Z(n20342) );
  XNOR U36518 ( .A(q[5]), .B(DB[2105]), .Z(n35034) );
  XNOR U36519 ( .A(q[4]), .B(DB[2104]), .Z(n20340) );
  IV U36520 ( .A(n20354), .Z(n35032) );
  XOR U36521 ( .A(n35035), .B(n35036), .Z(n20354) );
  XNOR U36522 ( .A(n20350), .B(n20352), .Z(n35036) );
  XNOR U36523 ( .A(q[0]), .B(DB[2100]), .Z(n20352) );
  XNOR U36524 ( .A(q[3]), .B(DB[2103]), .Z(n20350) );
  IV U36525 ( .A(n20349), .Z(n35035) );
  XNOR U36526 ( .A(n20347), .B(n35037), .Z(n20349) );
  XNOR U36527 ( .A(q[2]), .B(DB[2102]), .Z(n35037) );
  XNOR U36528 ( .A(q[1]), .B(DB[2101]), .Z(n20347) );
  XOR U36529 ( .A(n35038), .B(n20312), .Z(n20275) );
  XOR U36530 ( .A(n35039), .B(n20300), .Z(n20312) );
  XNOR U36531 ( .A(q[6]), .B(DB[2113]), .Z(n20300) );
  IV U36532 ( .A(n20299), .Z(n35039) );
  XNOR U36533 ( .A(n20297), .B(n35040), .Z(n20299) );
  XNOR U36534 ( .A(q[5]), .B(DB[2112]), .Z(n35040) );
  XNOR U36535 ( .A(q[4]), .B(DB[2111]), .Z(n20297) );
  IV U36536 ( .A(n20311), .Z(n35038) );
  XOR U36537 ( .A(n35041), .B(n35042), .Z(n20311) );
  XNOR U36538 ( .A(n20307), .B(n20309), .Z(n35042) );
  XNOR U36539 ( .A(q[0]), .B(DB[2107]), .Z(n20309) );
  XNOR U36540 ( .A(q[3]), .B(DB[2110]), .Z(n20307) );
  IV U36541 ( .A(n20306), .Z(n35041) );
  XNOR U36542 ( .A(n20304), .B(n35043), .Z(n20306) );
  XNOR U36543 ( .A(q[2]), .B(DB[2109]), .Z(n35043) );
  XNOR U36544 ( .A(q[1]), .B(DB[2108]), .Z(n20304) );
  XOR U36545 ( .A(n35044), .B(n20269), .Z(n20232) );
  XOR U36546 ( .A(n35045), .B(n20257), .Z(n20269) );
  XNOR U36547 ( .A(q[6]), .B(DB[2120]), .Z(n20257) );
  IV U36548 ( .A(n20256), .Z(n35045) );
  XNOR U36549 ( .A(n20254), .B(n35046), .Z(n20256) );
  XNOR U36550 ( .A(q[5]), .B(DB[2119]), .Z(n35046) );
  XNOR U36551 ( .A(q[4]), .B(DB[2118]), .Z(n20254) );
  IV U36552 ( .A(n20268), .Z(n35044) );
  XOR U36553 ( .A(n35047), .B(n35048), .Z(n20268) );
  XNOR U36554 ( .A(n20264), .B(n20266), .Z(n35048) );
  XNOR U36555 ( .A(q[0]), .B(DB[2114]), .Z(n20266) );
  XNOR U36556 ( .A(q[3]), .B(DB[2117]), .Z(n20264) );
  IV U36557 ( .A(n20263), .Z(n35047) );
  XNOR U36558 ( .A(n20261), .B(n35049), .Z(n20263) );
  XNOR U36559 ( .A(q[2]), .B(DB[2116]), .Z(n35049) );
  XNOR U36560 ( .A(q[1]), .B(DB[2115]), .Z(n20261) );
  XOR U36561 ( .A(n35050), .B(n20226), .Z(n20189) );
  XOR U36562 ( .A(n35051), .B(n20214), .Z(n20226) );
  XNOR U36563 ( .A(q[6]), .B(DB[2127]), .Z(n20214) );
  IV U36564 ( .A(n20213), .Z(n35051) );
  XNOR U36565 ( .A(n20211), .B(n35052), .Z(n20213) );
  XNOR U36566 ( .A(q[5]), .B(DB[2126]), .Z(n35052) );
  XNOR U36567 ( .A(q[4]), .B(DB[2125]), .Z(n20211) );
  IV U36568 ( .A(n20225), .Z(n35050) );
  XOR U36569 ( .A(n35053), .B(n35054), .Z(n20225) );
  XNOR U36570 ( .A(n20221), .B(n20223), .Z(n35054) );
  XNOR U36571 ( .A(q[0]), .B(DB[2121]), .Z(n20223) );
  XNOR U36572 ( .A(q[3]), .B(DB[2124]), .Z(n20221) );
  IV U36573 ( .A(n20220), .Z(n35053) );
  XNOR U36574 ( .A(n20218), .B(n35055), .Z(n20220) );
  XNOR U36575 ( .A(q[2]), .B(DB[2123]), .Z(n35055) );
  XNOR U36576 ( .A(q[1]), .B(DB[2122]), .Z(n20218) );
  XOR U36577 ( .A(n35056), .B(n20183), .Z(n20146) );
  XOR U36578 ( .A(n35057), .B(n20171), .Z(n20183) );
  XNOR U36579 ( .A(q[6]), .B(DB[2134]), .Z(n20171) );
  IV U36580 ( .A(n20170), .Z(n35057) );
  XNOR U36581 ( .A(n20168), .B(n35058), .Z(n20170) );
  XNOR U36582 ( .A(q[5]), .B(DB[2133]), .Z(n35058) );
  XNOR U36583 ( .A(q[4]), .B(DB[2132]), .Z(n20168) );
  IV U36584 ( .A(n20182), .Z(n35056) );
  XOR U36585 ( .A(n35059), .B(n35060), .Z(n20182) );
  XNOR U36586 ( .A(n20178), .B(n20180), .Z(n35060) );
  XNOR U36587 ( .A(q[0]), .B(DB[2128]), .Z(n20180) );
  XNOR U36588 ( .A(q[3]), .B(DB[2131]), .Z(n20178) );
  IV U36589 ( .A(n20177), .Z(n35059) );
  XNOR U36590 ( .A(n20175), .B(n35061), .Z(n20177) );
  XNOR U36591 ( .A(q[2]), .B(DB[2130]), .Z(n35061) );
  XNOR U36592 ( .A(q[1]), .B(DB[2129]), .Z(n20175) );
  XOR U36593 ( .A(n35062), .B(n20140), .Z(n20103) );
  XOR U36594 ( .A(n35063), .B(n20128), .Z(n20140) );
  XNOR U36595 ( .A(q[6]), .B(DB[2141]), .Z(n20128) );
  IV U36596 ( .A(n20127), .Z(n35063) );
  XNOR U36597 ( .A(n20125), .B(n35064), .Z(n20127) );
  XNOR U36598 ( .A(q[5]), .B(DB[2140]), .Z(n35064) );
  XNOR U36599 ( .A(q[4]), .B(DB[2139]), .Z(n20125) );
  IV U36600 ( .A(n20139), .Z(n35062) );
  XOR U36601 ( .A(n35065), .B(n35066), .Z(n20139) );
  XNOR U36602 ( .A(n20135), .B(n20137), .Z(n35066) );
  XNOR U36603 ( .A(q[0]), .B(DB[2135]), .Z(n20137) );
  XNOR U36604 ( .A(q[3]), .B(DB[2138]), .Z(n20135) );
  IV U36605 ( .A(n20134), .Z(n35065) );
  XNOR U36606 ( .A(n20132), .B(n35067), .Z(n20134) );
  XNOR U36607 ( .A(q[2]), .B(DB[2137]), .Z(n35067) );
  XNOR U36608 ( .A(q[1]), .B(DB[2136]), .Z(n20132) );
  XOR U36609 ( .A(n35068), .B(n20097), .Z(n20060) );
  XOR U36610 ( .A(n35069), .B(n20085), .Z(n20097) );
  XNOR U36611 ( .A(q[6]), .B(DB[2148]), .Z(n20085) );
  IV U36612 ( .A(n20084), .Z(n35069) );
  XNOR U36613 ( .A(n20082), .B(n35070), .Z(n20084) );
  XNOR U36614 ( .A(q[5]), .B(DB[2147]), .Z(n35070) );
  XNOR U36615 ( .A(q[4]), .B(DB[2146]), .Z(n20082) );
  IV U36616 ( .A(n20096), .Z(n35068) );
  XOR U36617 ( .A(n35071), .B(n35072), .Z(n20096) );
  XNOR U36618 ( .A(n20092), .B(n20094), .Z(n35072) );
  XNOR U36619 ( .A(q[0]), .B(DB[2142]), .Z(n20094) );
  XNOR U36620 ( .A(q[3]), .B(DB[2145]), .Z(n20092) );
  IV U36621 ( .A(n20091), .Z(n35071) );
  XNOR U36622 ( .A(n20089), .B(n35073), .Z(n20091) );
  XNOR U36623 ( .A(q[2]), .B(DB[2144]), .Z(n35073) );
  XNOR U36624 ( .A(q[1]), .B(DB[2143]), .Z(n20089) );
  XOR U36625 ( .A(n35074), .B(n20054), .Z(n20017) );
  XOR U36626 ( .A(n35075), .B(n20042), .Z(n20054) );
  XNOR U36627 ( .A(q[6]), .B(DB[2155]), .Z(n20042) );
  IV U36628 ( .A(n20041), .Z(n35075) );
  XNOR U36629 ( .A(n20039), .B(n35076), .Z(n20041) );
  XNOR U36630 ( .A(q[5]), .B(DB[2154]), .Z(n35076) );
  XNOR U36631 ( .A(q[4]), .B(DB[2153]), .Z(n20039) );
  IV U36632 ( .A(n20053), .Z(n35074) );
  XOR U36633 ( .A(n35077), .B(n35078), .Z(n20053) );
  XNOR U36634 ( .A(n20049), .B(n20051), .Z(n35078) );
  XNOR U36635 ( .A(q[0]), .B(DB[2149]), .Z(n20051) );
  XNOR U36636 ( .A(q[3]), .B(DB[2152]), .Z(n20049) );
  IV U36637 ( .A(n20048), .Z(n35077) );
  XNOR U36638 ( .A(n20046), .B(n35079), .Z(n20048) );
  XNOR U36639 ( .A(q[2]), .B(DB[2151]), .Z(n35079) );
  XNOR U36640 ( .A(q[1]), .B(DB[2150]), .Z(n20046) );
  XOR U36641 ( .A(n35080), .B(n20011), .Z(n19974) );
  XOR U36642 ( .A(n35081), .B(n19999), .Z(n20011) );
  XNOR U36643 ( .A(q[6]), .B(DB[2162]), .Z(n19999) );
  IV U36644 ( .A(n19998), .Z(n35081) );
  XNOR U36645 ( .A(n19996), .B(n35082), .Z(n19998) );
  XNOR U36646 ( .A(q[5]), .B(DB[2161]), .Z(n35082) );
  XNOR U36647 ( .A(q[4]), .B(DB[2160]), .Z(n19996) );
  IV U36648 ( .A(n20010), .Z(n35080) );
  XOR U36649 ( .A(n35083), .B(n35084), .Z(n20010) );
  XNOR U36650 ( .A(n20006), .B(n20008), .Z(n35084) );
  XNOR U36651 ( .A(q[0]), .B(DB[2156]), .Z(n20008) );
  XNOR U36652 ( .A(q[3]), .B(DB[2159]), .Z(n20006) );
  IV U36653 ( .A(n20005), .Z(n35083) );
  XNOR U36654 ( .A(n20003), .B(n35085), .Z(n20005) );
  XNOR U36655 ( .A(q[2]), .B(DB[2158]), .Z(n35085) );
  XNOR U36656 ( .A(q[1]), .B(DB[2157]), .Z(n20003) );
  XOR U36657 ( .A(n35086), .B(n19968), .Z(n19931) );
  XOR U36658 ( .A(n35087), .B(n19956), .Z(n19968) );
  XNOR U36659 ( .A(q[6]), .B(DB[2169]), .Z(n19956) );
  IV U36660 ( .A(n19955), .Z(n35087) );
  XNOR U36661 ( .A(n19953), .B(n35088), .Z(n19955) );
  XNOR U36662 ( .A(q[5]), .B(DB[2168]), .Z(n35088) );
  XNOR U36663 ( .A(q[4]), .B(DB[2167]), .Z(n19953) );
  IV U36664 ( .A(n19967), .Z(n35086) );
  XOR U36665 ( .A(n35089), .B(n35090), .Z(n19967) );
  XNOR U36666 ( .A(n19963), .B(n19965), .Z(n35090) );
  XNOR U36667 ( .A(q[0]), .B(DB[2163]), .Z(n19965) );
  XNOR U36668 ( .A(q[3]), .B(DB[2166]), .Z(n19963) );
  IV U36669 ( .A(n19962), .Z(n35089) );
  XNOR U36670 ( .A(n19960), .B(n35091), .Z(n19962) );
  XNOR U36671 ( .A(q[2]), .B(DB[2165]), .Z(n35091) );
  XNOR U36672 ( .A(q[1]), .B(DB[2164]), .Z(n19960) );
  XOR U36673 ( .A(n35092), .B(n19925), .Z(n19888) );
  XOR U36674 ( .A(n35093), .B(n19913), .Z(n19925) );
  XNOR U36675 ( .A(q[6]), .B(DB[2176]), .Z(n19913) );
  IV U36676 ( .A(n19912), .Z(n35093) );
  XNOR U36677 ( .A(n19910), .B(n35094), .Z(n19912) );
  XNOR U36678 ( .A(q[5]), .B(DB[2175]), .Z(n35094) );
  XNOR U36679 ( .A(q[4]), .B(DB[2174]), .Z(n19910) );
  IV U36680 ( .A(n19924), .Z(n35092) );
  XOR U36681 ( .A(n35095), .B(n35096), .Z(n19924) );
  XNOR U36682 ( .A(n19920), .B(n19922), .Z(n35096) );
  XNOR U36683 ( .A(q[0]), .B(DB[2170]), .Z(n19922) );
  XNOR U36684 ( .A(q[3]), .B(DB[2173]), .Z(n19920) );
  IV U36685 ( .A(n19919), .Z(n35095) );
  XNOR U36686 ( .A(n19917), .B(n35097), .Z(n19919) );
  XNOR U36687 ( .A(q[2]), .B(DB[2172]), .Z(n35097) );
  XNOR U36688 ( .A(q[1]), .B(DB[2171]), .Z(n19917) );
  XOR U36689 ( .A(n35098), .B(n19882), .Z(n19845) );
  XOR U36690 ( .A(n35099), .B(n19870), .Z(n19882) );
  XNOR U36691 ( .A(q[6]), .B(DB[2183]), .Z(n19870) );
  IV U36692 ( .A(n19869), .Z(n35099) );
  XNOR U36693 ( .A(n19867), .B(n35100), .Z(n19869) );
  XNOR U36694 ( .A(q[5]), .B(DB[2182]), .Z(n35100) );
  XNOR U36695 ( .A(q[4]), .B(DB[2181]), .Z(n19867) );
  IV U36696 ( .A(n19881), .Z(n35098) );
  XOR U36697 ( .A(n35101), .B(n35102), .Z(n19881) );
  XNOR U36698 ( .A(n19877), .B(n19879), .Z(n35102) );
  XNOR U36699 ( .A(q[0]), .B(DB[2177]), .Z(n19879) );
  XNOR U36700 ( .A(q[3]), .B(DB[2180]), .Z(n19877) );
  IV U36701 ( .A(n19876), .Z(n35101) );
  XNOR U36702 ( .A(n19874), .B(n35103), .Z(n19876) );
  XNOR U36703 ( .A(q[2]), .B(DB[2179]), .Z(n35103) );
  XNOR U36704 ( .A(q[1]), .B(DB[2178]), .Z(n19874) );
  XOR U36705 ( .A(n35104), .B(n19839), .Z(n19802) );
  XOR U36706 ( .A(n35105), .B(n19827), .Z(n19839) );
  XNOR U36707 ( .A(q[6]), .B(DB[2190]), .Z(n19827) );
  IV U36708 ( .A(n19826), .Z(n35105) );
  XNOR U36709 ( .A(n19824), .B(n35106), .Z(n19826) );
  XNOR U36710 ( .A(q[5]), .B(DB[2189]), .Z(n35106) );
  XNOR U36711 ( .A(q[4]), .B(DB[2188]), .Z(n19824) );
  IV U36712 ( .A(n19838), .Z(n35104) );
  XOR U36713 ( .A(n35107), .B(n35108), .Z(n19838) );
  XNOR U36714 ( .A(n19834), .B(n19836), .Z(n35108) );
  XNOR U36715 ( .A(q[0]), .B(DB[2184]), .Z(n19836) );
  XNOR U36716 ( .A(q[3]), .B(DB[2187]), .Z(n19834) );
  IV U36717 ( .A(n19833), .Z(n35107) );
  XNOR U36718 ( .A(n19831), .B(n35109), .Z(n19833) );
  XNOR U36719 ( .A(q[2]), .B(DB[2186]), .Z(n35109) );
  XNOR U36720 ( .A(q[1]), .B(DB[2185]), .Z(n19831) );
  XOR U36721 ( .A(n35110), .B(n19796), .Z(n19759) );
  XOR U36722 ( .A(n35111), .B(n19784), .Z(n19796) );
  XNOR U36723 ( .A(q[6]), .B(DB[2197]), .Z(n19784) );
  IV U36724 ( .A(n19783), .Z(n35111) );
  XNOR U36725 ( .A(n19781), .B(n35112), .Z(n19783) );
  XNOR U36726 ( .A(q[5]), .B(DB[2196]), .Z(n35112) );
  XNOR U36727 ( .A(q[4]), .B(DB[2195]), .Z(n19781) );
  IV U36728 ( .A(n19795), .Z(n35110) );
  XOR U36729 ( .A(n35113), .B(n35114), .Z(n19795) );
  XNOR U36730 ( .A(n19791), .B(n19793), .Z(n35114) );
  XNOR U36731 ( .A(q[0]), .B(DB[2191]), .Z(n19793) );
  XNOR U36732 ( .A(q[3]), .B(DB[2194]), .Z(n19791) );
  IV U36733 ( .A(n19790), .Z(n35113) );
  XNOR U36734 ( .A(n19788), .B(n35115), .Z(n19790) );
  XNOR U36735 ( .A(q[2]), .B(DB[2193]), .Z(n35115) );
  XNOR U36736 ( .A(q[1]), .B(DB[2192]), .Z(n19788) );
  XOR U36737 ( .A(n35116), .B(n19753), .Z(n19716) );
  XOR U36738 ( .A(n35117), .B(n19741), .Z(n19753) );
  XNOR U36739 ( .A(q[6]), .B(DB[2204]), .Z(n19741) );
  IV U36740 ( .A(n19740), .Z(n35117) );
  XNOR U36741 ( .A(n19738), .B(n35118), .Z(n19740) );
  XNOR U36742 ( .A(q[5]), .B(DB[2203]), .Z(n35118) );
  XNOR U36743 ( .A(q[4]), .B(DB[2202]), .Z(n19738) );
  IV U36744 ( .A(n19752), .Z(n35116) );
  XOR U36745 ( .A(n35119), .B(n35120), .Z(n19752) );
  XNOR U36746 ( .A(n19748), .B(n19750), .Z(n35120) );
  XNOR U36747 ( .A(q[0]), .B(DB[2198]), .Z(n19750) );
  XNOR U36748 ( .A(q[3]), .B(DB[2201]), .Z(n19748) );
  IV U36749 ( .A(n19747), .Z(n35119) );
  XNOR U36750 ( .A(n19745), .B(n35121), .Z(n19747) );
  XNOR U36751 ( .A(q[2]), .B(DB[2200]), .Z(n35121) );
  XNOR U36752 ( .A(q[1]), .B(DB[2199]), .Z(n19745) );
  XOR U36753 ( .A(n35122), .B(n19710), .Z(n19673) );
  XOR U36754 ( .A(n35123), .B(n19698), .Z(n19710) );
  XNOR U36755 ( .A(q[6]), .B(DB[2211]), .Z(n19698) );
  IV U36756 ( .A(n19697), .Z(n35123) );
  XNOR U36757 ( .A(n19695), .B(n35124), .Z(n19697) );
  XNOR U36758 ( .A(q[5]), .B(DB[2210]), .Z(n35124) );
  XNOR U36759 ( .A(q[4]), .B(DB[2209]), .Z(n19695) );
  IV U36760 ( .A(n19709), .Z(n35122) );
  XOR U36761 ( .A(n35125), .B(n35126), .Z(n19709) );
  XNOR U36762 ( .A(n19705), .B(n19707), .Z(n35126) );
  XNOR U36763 ( .A(q[0]), .B(DB[2205]), .Z(n19707) );
  XNOR U36764 ( .A(q[3]), .B(DB[2208]), .Z(n19705) );
  IV U36765 ( .A(n19704), .Z(n35125) );
  XNOR U36766 ( .A(n19702), .B(n35127), .Z(n19704) );
  XNOR U36767 ( .A(q[2]), .B(DB[2207]), .Z(n35127) );
  XNOR U36768 ( .A(q[1]), .B(DB[2206]), .Z(n19702) );
  XOR U36769 ( .A(n35128), .B(n19667), .Z(n19630) );
  XOR U36770 ( .A(n35129), .B(n19655), .Z(n19667) );
  XNOR U36771 ( .A(q[6]), .B(DB[2218]), .Z(n19655) );
  IV U36772 ( .A(n19654), .Z(n35129) );
  XNOR U36773 ( .A(n19652), .B(n35130), .Z(n19654) );
  XNOR U36774 ( .A(q[5]), .B(DB[2217]), .Z(n35130) );
  XNOR U36775 ( .A(q[4]), .B(DB[2216]), .Z(n19652) );
  IV U36776 ( .A(n19666), .Z(n35128) );
  XOR U36777 ( .A(n35131), .B(n35132), .Z(n19666) );
  XNOR U36778 ( .A(n19662), .B(n19664), .Z(n35132) );
  XNOR U36779 ( .A(q[0]), .B(DB[2212]), .Z(n19664) );
  XNOR U36780 ( .A(q[3]), .B(DB[2215]), .Z(n19662) );
  IV U36781 ( .A(n19661), .Z(n35131) );
  XNOR U36782 ( .A(n19659), .B(n35133), .Z(n19661) );
  XNOR U36783 ( .A(q[2]), .B(DB[2214]), .Z(n35133) );
  XNOR U36784 ( .A(q[1]), .B(DB[2213]), .Z(n19659) );
  XOR U36785 ( .A(n35134), .B(n19624), .Z(n19587) );
  XOR U36786 ( .A(n35135), .B(n19612), .Z(n19624) );
  XNOR U36787 ( .A(q[6]), .B(DB[2225]), .Z(n19612) );
  IV U36788 ( .A(n19611), .Z(n35135) );
  XNOR U36789 ( .A(n19609), .B(n35136), .Z(n19611) );
  XNOR U36790 ( .A(q[5]), .B(DB[2224]), .Z(n35136) );
  XNOR U36791 ( .A(q[4]), .B(DB[2223]), .Z(n19609) );
  IV U36792 ( .A(n19623), .Z(n35134) );
  XOR U36793 ( .A(n35137), .B(n35138), .Z(n19623) );
  XNOR U36794 ( .A(n19619), .B(n19621), .Z(n35138) );
  XNOR U36795 ( .A(q[0]), .B(DB[2219]), .Z(n19621) );
  XNOR U36796 ( .A(q[3]), .B(DB[2222]), .Z(n19619) );
  IV U36797 ( .A(n19618), .Z(n35137) );
  XNOR U36798 ( .A(n19616), .B(n35139), .Z(n19618) );
  XNOR U36799 ( .A(q[2]), .B(DB[2221]), .Z(n35139) );
  XNOR U36800 ( .A(q[1]), .B(DB[2220]), .Z(n19616) );
  XOR U36801 ( .A(n35140), .B(n19581), .Z(n19544) );
  XOR U36802 ( .A(n35141), .B(n19569), .Z(n19581) );
  XNOR U36803 ( .A(q[6]), .B(DB[2232]), .Z(n19569) );
  IV U36804 ( .A(n19568), .Z(n35141) );
  XNOR U36805 ( .A(n19566), .B(n35142), .Z(n19568) );
  XNOR U36806 ( .A(q[5]), .B(DB[2231]), .Z(n35142) );
  XNOR U36807 ( .A(q[4]), .B(DB[2230]), .Z(n19566) );
  IV U36808 ( .A(n19580), .Z(n35140) );
  XOR U36809 ( .A(n35143), .B(n35144), .Z(n19580) );
  XNOR U36810 ( .A(n19576), .B(n19578), .Z(n35144) );
  XNOR U36811 ( .A(q[0]), .B(DB[2226]), .Z(n19578) );
  XNOR U36812 ( .A(q[3]), .B(DB[2229]), .Z(n19576) );
  IV U36813 ( .A(n19575), .Z(n35143) );
  XNOR U36814 ( .A(n19573), .B(n35145), .Z(n19575) );
  XNOR U36815 ( .A(q[2]), .B(DB[2228]), .Z(n35145) );
  XNOR U36816 ( .A(q[1]), .B(DB[2227]), .Z(n19573) );
  XOR U36817 ( .A(n35146), .B(n19538), .Z(n19501) );
  XOR U36818 ( .A(n35147), .B(n19526), .Z(n19538) );
  XNOR U36819 ( .A(q[6]), .B(DB[2239]), .Z(n19526) );
  IV U36820 ( .A(n19525), .Z(n35147) );
  XNOR U36821 ( .A(n19523), .B(n35148), .Z(n19525) );
  XNOR U36822 ( .A(q[5]), .B(DB[2238]), .Z(n35148) );
  XNOR U36823 ( .A(q[4]), .B(DB[2237]), .Z(n19523) );
  IV U36824 ( .A(n19537), .Z(n35146) );
  XOR U36825 ( .A(n35149), .B(n35150), .Z(n19537) );
  XNOR U36826 ( .A(n19533), .B(n19535), .Z(n35150) );
  XNOR U36827 ( .A(q[0]), .B(DB[2233]), .Z(n19535) );
  XNOR U36828 ( .A(q[3]), .B(DB[2236]), .Z(n19533) );
  IV U36829 ( .A(n19532), .Z(n35149) );
  XNOR U36830 ( .A(n19530), .B(n35151), .Z(n19532) );
  XNOR U36831 ( .A(q[2]), .B(DB[2235]), .Z(n35151) );
  XNOR U36832 ( .A(q[1]), .B(DB[2234]), .Z(n19530) );
  XOR U36833 ( .A(n35152), .B(n19495), .Z(n19458) );
  XOR U36834 ( .A(n35153), .B(n19483), .Z(n19495) );
  XNOR U36835 ( .A(q[6]), .B(DB[2246]), .Z(n19483) );
  IV U36836 ( .A(n19482), .Z(n35153) );
  XNOR U36837 ( .A(n19480), .B(n35154), .Z(n19482) );
  XNOR U36838 ( .A(q[5]), .B(DB[2245]), .Z(n35154) );
  XNOR U36839 ( .A(q[4]), .B(DB[2244]), .Z(n19480) );
  IV U36840 ( .A(n19494), .Z(n35152) );
  XOR U36841 ( .A(n35155), .B(n35156), .Z(n19494) );
  XNOR U36842 ( .A(n19490), .B(n19492), .Z(n35156) );
  XNOR U36843 ( .A(q[0]), .B(DB[2240]), .Z(n19492) );
  XNOR U36844 ( .A(q[3]), .B(DB[2243]), .Z(n19490) );
  IV U36845 ( .A(n19489), .Z(n35155) );
  XNOR U36846 ( .A(n19487), .B(n35157), .Z(n19489) );
  XNOR U36847 ( .A(q[2]), .B(DB[2242]), .Z(n35157) );
  XNOR U36848 ( .A(q[1]), .B(DB[2241]), .Z(n19487) );
  XOR U36849 ( .A(n35158), .B(n19452), .Z(n19415) );
  XOR U36850 ( .A(n35159), .B(n19440), .Z(n19452) );
  XNOR U36851 ( .A(q[6]), .B(DB[2253]), .Z(n19440) );
  IV U36852 ( .A(n19439), .Z(n35159) );
  XNOR U36853 ( .A(n19437), .B(n35160), .Z(n19439) );
  XNOR U36854 ( .A(q[5]), .B(DB[2252]), .Z(n35160) );
  XNOR U36855 ( .A(q[4]), .B(DB[2251]), .Z(n19437) );
  IV U36856 ( .A(n19451), .Z(n35158) );
  XOR U36857 ( .A(n35161), .B(n35162), .Z(n19451) );
  XNOR U36858 ( .A(n19447), .B(n19449), .Z(n35162) );
  XNOR U36859 ( .A(q[0]), .B(DB[2247]), .Z(n19449) );
  XNOR U36860 ( .A(q[3]), .B(DB[2250]), .Z(n19447) );
  IV U36861 ( .A(n19446), .Z(n35161) );
  XNOR U36862 ( .A(n19444), .B(n35163), .Z(n19446) );
  XNOR U36863 ( .A(q[2]), .B(DB[2249]), .Z(n35163) );
  XNOR U36864 ( .A(q[1]), .B(DB[2248]), .Z(n19444) );
  XOR U36865 ( .A(n35164), .B(n19409), .Z(n19372) );
  XOR U36866 ( .A(n35165), .B(n19397), .Z(n19409) );
  XNOR U36867 ( .A(q[6]), .B(DB[2260]), .Z(n19397) );
  IV U36868 ( .A(n19396), .Z(n35165) );
  XNOR U36869 ( .A(n19394), .B(n35166), .Z(n19396) );
  XNOR U36870 ( .A(q[5]), .B(DB[2259]), .Z(n35166) );
  XNOR U36871 ( .A(q[4]), .B(DB[2258]), .Z(n19394) );
  IV U36872 ( .A(n19408), .Z(n35164) );
  XOR U36873 ( .A(n35167), .B(n35168), .Z(n19408) );
  XNOR U36874 ( .A(n19404), .B(n19406), .Z(n35168) );
  XNOR U36875 ( .A(q[0]), .B(DB[2254]), .Z(n19406) );
  XNOR U36876 ( .A(q[3]), .B(DB[2257]), .Z(n19404) );
  IV U36877 ( .A(n19403), .Z(n35167) );
  XNOR U36878 ( .A(n19401), .B(n35169), .Z(n19403) );
  XNOR U36879 ( .A(q[2]), .B(DB[2256]), .Z(n35169) );
  XNOR U36880 ( .A(q[1]), .B(DB[2255]), .Z(n19401) );
  XOR U36881 ( .A(n35170), .B(n19366), .Z(n19329) );
  XOR U36882 ( .A(n35171), .B(n19354), .Z(n19366) );
  XNOR U36883 ( .A(q[6]), .B(DB[2267]), .Z(n19354) );
  IV U36884 ( .A(n19353), .Z(n35171) );
  XNOR U36885 ( .A(n19351), .B(n35172), .Z(n19353) );
  XNOR U36886 ( .A(q[5]), .B(DB[2266]), .Z(n35172) );
  XNOR U36887 ( .A(q[4]), .B(DB[2265]), .Z(n19351) );
  IV U36888 ( .A(n19365), .Z(n35170) );
  XOR U36889 ( .A(n35173), .B(n35174), .Z(n19365) );
  XNOR U36890 ( .A(n19361), .B(n19363), .Z(n35174) );
  XNOR U36891 ( .A(q[0]), .B(DB[2261]), .Z(n19363) );
  XNOR U36892 ( .A(q[3]), .B(DB[2264]), .Z(n19361) );
  IV U36893 ( .A(n19360), .Z(n35173) );
  XNOR U36894 ( .A(n19358), .B(n35175), .Z(n19360) );
  XNOR U36895 ( .A(q[2]), .B(DB[2263]), .Z(n35175) );
  XNOR U36896 ( .A(q[1]), .B(DB[2262]), .Z(n19358) );
  XOR U36897 ( .A(n35176), .B(n19323), .Z(n19286) );
  XOR U36898 ( .A(n35177), .B(n19311), .Z(n19323) );
  XNOR U36899 ( .A(q[6]), .B(DB[2274]), .Z(n19311) );
  IV U36900 ( .A(n19310), .Z(n35177) );
  XNOR U36901 ( .A(n19308), .B(n35178), .Z(n19310) );
  XNOR U36902 ( .A(q[5]), .B(DB[2273]), .Z(n35178) );
  XNOR U36903 ( .A(q[4]), .B(DB[2272]), .Z(n19308) );
  IV U36904 ( .A(n19322), .Z(n35176) );
  XOR U36905 ( .A(n35179), .B(n35180), .Z(n19322) );
  XNOR U36906 ( .A(n19318), .B(n19320), .Z(n35180) );
  XNOR U36907 ( .A(q[0]), .B(DB[2268]), .Z(n19320) );
  XNOR U36908 ( .A(q[3]), .B(DB[2271]), .Z(n19318) );
  IV U36909 ( .A(n19317), .Z(n35179) );
  XNOR U36910 ( .A(n19315), .B(n35181), .Z(n19317) );
  XNOR U36911 ( .A(q[2]), .B(DB[2270]), .Z(n35181) );
  XNOR U36912 ( .A(q[1]), .B(DB[2269]), .Z(n19315) );
  XOR U36913 ( .A(n35182), .B(n19280), .Z(n19243) );
  XOR U36914 ( .A(n35183), .B(n19268), .Z(n19280) );
  XNOR U36915 ( .A(q[6]), .B(DB[2281]), .Z(n19268) );
  IV U36916 ( .A(n19267), .Z(n35183) );
  XNOR U36917 ( .A(n19265), .B(n35184), .Z(n19267) );
  XNOR U36918 ( .A(q[5]), .B(DB[2280]), .Z(n35184) );
  XNOR U36919 ( .A(q[4]), .B(DB[2279]), .Z(n19265) );
  IV U36920 ( .A(n19279), .Z(n35182) );
  XOR U36921 ( .A(n35185), .B(n35186), .Z(n19279) );
  XNOR U36922 ( .A(n19275), .B(n19277), .Z(n35186) );
  XNOR U36923 ( .A(q[0]), .B(DB[2275]), .Z(n19277) );
  XNOR U36924 ( .A(q[3]), .B(DB[2278]), .Z(n19275) );
  IV U36925 ( .A(n19274), .Z(n35185) );
  XNOR U36926 ( .A(n19272), .B(n35187), .Z(n19274) );
  XNOR U36927 ( .A(q[2]), .B(DB[2277]), .Z(n35187) );
  XNOR U36928 ( .A(q[1]), .B(DB[2276]), .Z(n19272) );
  XOR U36929 ( .A(n35188), .B(n19237), .Z(n19200) );
  XOR U36930 ( .A(n35189), .B(n19225), .Z(n19237) );
  XNOR U36931 ( .A(q[6]), .B(DB[2288]), .Z(n19225) );
  IV U36932 ( .A(n19224), .Z(n35189) );
  XNOR U36933 ( .A(n19222), .B(n35190), .Z(n19224) );
  XNOR U36934 ( .A(q[5]), .B(DB[2287]), .Z(n35190) );
  XNOR U36935 ( .A(q[4]), .B(DB[2286]), .Z(n19222) );
  IV U36936 ( .A(n19236), .Z(n35188) );
  XOR U36937 ( .A(n35191), .B(n35192), .Z(n19236) );
  XNOR U36938 ( .A(n19232), .B(n19234), .Z(n35192) );
  XNOR U36939 ( .A(q[0]), .B(DB[2282]), .Z(n19234) );
  XNOR U36940 ( .A(q[3]), .B(DB[2285]), .Z(n19232) );
  IV U36941 ( .A(n19231), .Z(n35191) );
  XNOR U36942 ( .A(n19229), .B(n35193), .Z(n19231) );
  XNOR U36943 ( .A(q[2]), .B(DB[2284]), .Z(n35193) );
  XNOR U36944 ( .A(q[1]), .B(DB[2283]), .Z(n19229) );
  XOR U36945 ( .A(n35194), .B(n19194), .Z(n19157) );
  XOR U36946 ( .A(n35195), .B(n19182), .Z(n19194) );
  XNOR U36947 ( .A(q[6]), .B(DB[2295]), .Z(n19182) );
  IV U36948 ( .A(n19181), .Z(n35195) );
  XNOR U36949 ( .A(n19179), .B(n35196), .Z(n19181) );
  XNOR U36950 ( .A(q[5]), .B(DB[2294]), .Z(n35196) );
  XNOR U36951 ( .A(q[4]), .B(DB[2293]), .Z(n19179) );
  IV U36952 ( .A(n19193), .Z(n35194) );
  XOR U36953 ( .A(n35197), .B(n35198), .Z(n19193) );
  XNOR U36954 ( .A(n19189), .B(n19191), .Z(n35198) );
  XNOR U36955 ( .A(q[0]), .B(DB[2289]), .Z(n19191) );
  XNOR U36956 ( .A(q[3]), .B(DB[2292]), .Z(n19189) );
  IV U36957 ( .A(n19188), .Z(n35197) );
  XNOR U36958 ( .A(n19186), .B(n35199), .Z(n19188) );
  XNOR U36959 ( .A(q[2]), .B(DB[2291]), .Z(n35199) );
  XNOR U36960 ( .A(q[1]), .B(DB[2290]), .Z(n19186) );
  XOR U36961 ( .A(n35200), .B(n19151), .Z(n19114) );
  XOR U36962 ( .A(n35201), .B(n19139), .Z(n19151) );
  XNOR U36963 ( .A(q[6]), .B(DB[2302]), .Z(n19139) );
  IV U36964 ( .A(n19138), .Z(n35201) );
  XNOR U36965 ( .A(n19136), .B(n35202), .Z(n19138) );
  XNOR U36966 ( .A(q[5]), .B(DB[2301]), .Z(n35202) );
  XNOR U36967 ( .A(q[4]), .B(DB[2300]), .Z(n19136) );
  IV U36968 ( .A(n19150), .Z(n35200) );
  XOR U36969 ( .A(n35203), .B(n35204), .Z(n19150) );
  XNOR U36970 ( .A(n19146), .B(n19148), .Z(n35204) );
  XNOR U36971 ( .A(q[0]), .B(DB[2296]), .Z(n19148) );
  XNOR U36972 ( .A(q[3]), .B(DB[2299]), .Z(n19146) );
  IV U36973 ( .A(n19145), .Z(n35203) );
  XNOR U36974 ( .A(n19143), .B(n35205), .Z(n19145) );
  XNOR U36975 ( .A(q[2]), .B(DB[2298]), .Z(n35205) );
  XNOR U36976 ( .A(q[1]), .B(DB[2297]), .Z(n19143) );
  XOR U36977 ( .A(n35206), .B(n19108), .Z(n19071) );
  XOR U36978 ( .A(n35207), .B(n19096), .Z(n19108) );
  XNOR U36979 ( .A(q[6]), .B(DB[2309]), .Z(n19096) );
  IV U36980 ( .A(n19095), .Z(n35207) );
  XNOR U36981 ( .A(n19093), .B(n35208), .Z(n19095) );
  XNOR U36982 ( .A(q[5]), .B(DB[2308]), .Z(n35208) );
  XNOR U36983 ( .A(q[4]), .B(DB[2307]), .Z(n19093) );
  IV U36984 ( .A(n19107), .Z(n35206) );
  XOR U36985 ( .A(n35209), .B(n35210), .Z(n19107) );
  XNOR U36986 ( .A(n19103), .B(n19105), .Z(n35210) );
  XNOR U36987 ( .A(q[0]), .B(DB[2303]), .Z(n19105) );
  XNOR U36988 ( .A(q[3]), .B(DB[2306]), .Z(n19103) );
  IV U36989 ( .A(n19102), .Z(n35209) );
  XNOR U36990 ( .A(n19100), .B(n35211), .Z(n19102) );
  XNOR U36991 ( .A(q[2]), .B(DB[2305]), .Z(n35211) );
  XNOR U36992 ( .A(q[1]), .B(DB[2304]), .Z(n19100) );
  XOR U36993 ( .A(n35212), .B(n19065), .Z(n19028) );
  XOR U36994 ( .A(n35213), .B(n19053), .Z(n19065) );
  XNOR U36995 ( .A(q[6]), .B(DB[2316]), .Z(n19053) );
  IV U36996 ( .A(n19052), .Z(n35213) );
  XNOR U36997 ( .A(n19050), .B(n35214), .Z(n19052) );
  XNOR U36998 ( .A(q[5]), .B(DB[2315]), .Z(n35214) );
  XNOR U36999 ( .A(q[4]), .B(DB[2314]), .Z(n19050) );
  IV U37000 ( .A(n19064), .Z(n35212) );
  XOR U37001 ( .A(n35215), .B(n35216), .Z(n19064) );
  XNOR U37002 ( .A(n19060), .B(n19062), .Z(n35216) );
  XNOR U37003 ( .A(q[0]), .B(DB[2310]), .Z(n19062) );
  XNOR U37004 ( .A(q[3]), .B(DB[2313]), .Z(n19060) );
  IV U37005 ( .A(n19059), .Z(n35215) );
  XNOR U37006 ( .A(n19057), .B(n35217), .Z(n19059) );
  XNOR U37007 ( .A(q[2]), .B(DB[2312]), .Z(n35217) );
  XNOR U37008 ( .A(q[1]), .B(DB[2311]), .Z(n19057) );
  XOR U37009 ( .A(n35218), .B(n19022), .Z(n18985) );
  XOR U37010 ( .A(n35219), .B(n19010), .Z(n19022) );
  XNOR U37011 ( .A(q[6]), .B(DB[2323]), .Z(n19010) );
  IV U37012 ( .A(n19009), .Z(n35219) );
  XNOR U37013 ( .A(n19007), .B(n35220), .Z(n19009) );
  XNOR U37014 ( .A(q[5]), .B(DB[2322]), .Z(n35220) );
  XNOR U37015 ( .A(q[4]), .B(DB[2321]), .Z(n19007) );
  IV U37016 ( .A(n19021), .Z(n35218) );
  XOR U37017 ( .A(n35221), .B(n35222), .Z(n19021) );
  XNOR U37018 ( .A(n19017), .B(n19019), .Z(n35222) );
  XNOR U37019 ( .A(q[0]), .B(DB[2317]), .Z(n19019) );
  XNOR U37020 ( .A(q[3]), .B(DB[2320]), .Z(n19017) );
  IV U37021 ( .A(n19016), .Z(n35221) );
  XNOR U37022 ( .A(n19014), .B(n35223), .Z(n19016) );
  XNOR U37023 ( .A(q[2]), .B(DB[2319]), .Z(n35223) );
  XNOR U37024 ( .A(q[1]), .B(DB[2318]), .Z(n19014) );
  XOR U37025 ( .A(n35224), .B(n18979), .Z(n18942) );
  XOR U37026 ( .A(n35225), .B(n18967), .Z(n18979) );
  XNOR U37027 ( .A(q[6]), .B(DB[2330]), .Z(n18967) );
  IV U37028 ( .A(n18966), .Z(n35225) );
  XNOR U37029 ( .A(n18964), .B(n35226), .Z(n18966) );
  XNOR U37030 ( .A(q[5]), .B(DB[2329]), .Z(n35226) );
  XNOR U37031 ( .A(q[4]), .B(DB[2328]), .Z(n18964) );
  IV U37032 ( .A(n18978), .Z(n35224) );
  XOR U37033 ( .A(n35227), .B(n35228), .Z(n18978) );
  XNOR U37034 ( .A(n18974), .B(n18976), .Z(n35228) );
  XNOR U37035 ( .A(q[0]), .B(DB[2324]), .Z(n18976) );
  XNOR U37036 ( .A(q[3]), .B(DB[2327]), .Z(n18974) );
  IV U37037 ( .A(n18973), .Z(n35227) );
  XNOR U37038 ( .A(n18971), .B(n35229), .Z(n18973) );
  XNOR U37039 ( .A(q[2]), .B(DB[2326]), .Z(n35229) );
  XNOR U37040 ( .A(q[1]), .B(DB[2325]), .Z(n18971) );
  XOR U37041 ( .A(n35230), .B(n18936), .Z(n18899) );
  XOR U37042 ( .A(n35231), .B(n18924), .Z(n18936) );
  XNOR U37043 ( .A(q[6]), .B(DB[2337]), .Z(n18924) );
  IV U37044 ( .A(n18923), .Z(n35231) );
  XNOR U37045 ( .A(n18921), .B(n35232), .Z(n18923) );
  XNOR U37046 ( .A(q[5]), .B(DB[2336]), .Z(n35232) );
  XNOR U37047 ( .A(q[4]), .B(DB[2335]), .Z(n18921) );
  IV U37048 ( .A(n18935), .Z(n35230) );
  XOR U37049 ( .A(n35233), .B(n35234), .Z(n18935) );
  XNOR U37050 ( .A(n18931), .B(n18933), .Z(n35234) );
  XNOR U37051 ( .A(q[0]), .B(DB[2331]), .Z(n18933) );
  XNOR U37052 ( .A(q[3]), .B(DB[2334]), .Z(n18931) );
  IV U37053 ( .A(n18930), .Z(n35233) );
  XNOR U37054 ( .A(n18928), .B(n35235), .Z(n18930) );
  XNOR U37055 ( .A(q[2]), .B(DB[2333]), .Z(n35235) );
  XNOR U37056 ( .A(q[1]), .B(DB[2332]), .Z(n18928) );
  XOR U37057 ( .A(n35236), .B(n18893), .Z(n18856) );
  XOR U37058 ( .A(n35237), .B(n18881), .Z(n18893) );
  XNOR U37059 ( .A(q[6]), .B(DB[2344]), .Z(n18881) );
  IV U37060 ( .A(n18880), .Z(n35237) );
  XNOR U37061 ( .A(n18878), .B(n35238), .Z(n18880) );
  XNOR U37062 ( .A(q[5]), .B(DB[2343]), .Z(n35238) );
  XNOR U37063 ( .A(q[4]), .B(DB[2342]), .Z(n18878) );
  IV U37064 ( .A(n18892), .Z(n35236) );
  XOR U37065 ( .A(n35239), .B(n35240), .Z(n18892) );
  XNOR U37066 ( .A(n18888), .B(n18890), .Z(n35240) );
  XNOR U37067 ( .A(q[0]), .B(DB[2338]), .Z(n18890) );
  XNOR U37068 ( .A(q[3]), .B(DB[2341]), .Z(n18888) );
  IV U37069 ( .A(n18887), .Z(n35239) );
  XNOR U37070 ( .A(n18885), .B(n35241), .Z(n18887) );
  XNOR U37071 ( .A(q[2]), .B(DB[2340]), .Z(n35241) );
  XNOR U37072 ( .A(q[1]), .B(DB[2339]), .Z(n18885) );
  XOR U37073 ( .A(n35242), .B(n18850), .Z(n18813) );
  XOR U37074 ( .A(n35243), .B(n18838), .Z(n18850) );
  XNOR U37075 ( .A(q[6]), .B(DB[2351]), .Z(n18838) );
  IV U37076 ( .A(n18837), .Z(n35243) );
  XNOR U37077 ( .A(n18835), .B(n35244), .Z(n18837) );
  XNOR U37078 ( .A(q[5]), .B(DB[2350]), .Z(n35244) );
  XNOR U37079 ( .A(q[4]), .B(DB[2349]), .Z(n18835) );
  IV U37080 ( .A(n18849), .Z(n35242) );
  XOR U37081 ( .A(n35245), .B(n35246), .Z(n18849) );
  XNOR U37082 ( .A(n18845), .B(n18847), .Z(n35246) );
  XNOR U37083 ( .A(q[0]), .B(DB[2345]), .Z(n18847) );
  XNOR U37084 ( .A(q[3]), .B(DB[2348]), .Z(n18845) );
  IV U37085 ( .A(n18844), .Z(n35245) );
  XNOR U37086 ( .A(n18842), .B(n35247), .Z(n18844) );
  XNOR U37087 ( .A(q[2]), .B(DB[2347]), .Z(n35247) );
  XNOR U37088 ( .A(q[1]), .B(DB[2346]), .Z(n18842) );
  XOR U37089 ( .A(n35248), .B(n18807), .Z(n18770) );
  XOR U37090 ( .A(n35249), .B(n18795), .Z(n18807) );
  XNOR U37091 ( .A(q[6]), .B(DB[2358]), .Z(n18795) );
  IV U37092 ( .A(n18794), .Z(n35249) );
  XNOR U37093 ( .A(n18792), .B(n35250), .Z(n18794) );
  XNOR U37094 ( .A(q[5]), .B(DB[2357]), .Z(n35250) );
  XNOR U37095 ( .A(q[4]), .B(DB[2356]), .Z(n18792) );
  IV U37096 ( .A(n18806), .Z(n35248) );
  XOR U37097 ( .A(n35251), .B(n35252), .Z(n18806) );
  XNOR U37098 ( .A(n18802), .B(n18804), .Z(n35252) );
  XNOR U37099 ( .A(q[0]), .B(DB[2352]), .Z(n18804) );
  XNOR U37100 ( .A(q[3]), .B(DB[2355]), .Z(n18802) );
  IV U37101 ( .A(n18801), .Z(n35251) );
  XNOR U37102 ( .A(n18799), .B(n35253), .Z(n18801) );
  XNOR U37103 ( .A(q[2]), .B(DB[2354]), .Z(n35253) );
  XNOR U37104 ( .A(q[1]), .B(DB[2353]), .Z(n18799) );
  XOR U37105 ( .A(n35254), .B(n18764), .Z(n18727) );
  XOR U37106 ( .A(n35255), .B(n18752), .Z(n18764) );
  XNOR U37107 ( .A(q[6]), .B(DB[2365]), .Z(n18752) );
  IV U37108 ( .A(n18751), .Z(n35255) );
  XNOR U37109 ( .A(n18749), .B(n35256), .Z(n18751) );
  XNOR U37110 ( .A(q[5]), .B(DB[2364]), .Z(n35256) );
  XNOR U37111 ( .A(q[4]), .B(DB[2363]), .Z(n18749) );
  IV U37112 ( .A(n18763), .Z(n35254) );
  XOR U37113 ( .A(n35257), .B(n35258), .Z(n18763) );
  XNOR U37114 ( .A(n18759), .B(n18761), .Z(n35258) );
  XNOR U37115 ( .A(q[0]), .B(DB[2359]), .Z(n18761) );
  XNOR U37116 ( .A(q[3]), .B(DB[2362]), .Z(n18759) );
  IV U37117 ( .A(n18758), .Z(n35257) );
  XNOR U37118 ( .A(n18756), .B(n35259), .Z(n18758) );
  XNOR U37119 ( .A(q[2]), .B(DB[2361]), .Z(n35259) );
  XNOR U37120 ( .A(q[1]), .B(DB[2360]), .Z(n18756) );
  XOR U37121 ( .A(n35260), .B(n18721), .Z(n18684) );
  XOR U37122 ( .A(n35261), .B(n18709), .Z(n18721) );
  XNOR U37123 ( .A(q[6]), .B(DB[2372]), .Z(n18709) );
  IV U37124 ( .A(n18708), .Z(n35261) );
  XNOR U37125 ( .A(n18706), .B(n35262), .Z(n18708) );
  XNOR U37126 ( .A(q[5]), .B(DB[2371]), .Z(n35262) );
  XNOR U37127 ( .A(q[4]), .B(DB[2370]), .Z(n18706) );
  IV U37128 ( .A(n18720), .Z(n35260) );
  XOR U37129 ( .A(n35263), .B(n35264), .Z(n18720) );
  XNOR U37130 ( .A(n18716), .B(n18718), .Z(n35264) );
  XNOR U37131 ( .A(q[0]), .B(DB[2366]), .Z(n18718) );
  XNOR U37132 ( .A(q[3]), .B(DB[2369]), .Z(n18716) );
  IV U37133 ( .A(n18715), .Z(n35263) );
  XNOR U37134 ( .A(n18713), .B(n35265), .Z(n18715) );
  XNOR U37135 ( .A(q[2]), .B(DB[2368]), .Z(n35265) );
  XNOR U37136 ( .A(q[1]), .B(DB[2367]), .Z(n18713) );
  XOR U37137 ( .A(n35266), .B(n18678), .Z(n18641) );
  XOR U37138 ( .A(n35267), .B(n18666), .Z(n18678) );
  XNOR U37139 ( .A(q[6]), .B(DB[2379]), .Z(n18666) );
  IV U37140 ( .A(n18665), .Z(n35267) );
  XNOR U37141 ( .A(n18663), .B(n35268), .Z(n18665) );
  XNOR U37142 ( .A(q[5]), .B(DB[2378]), .Z(n35268) );
  XNOR U37143 ( .A(q[4]), .B(DB[2377]), .Z(n18663) );
  IV U37144 ( .A(n18677), .Z(n35266) );
  XOR U37145 ( .A(n35269), .B(n35270), .Z(n18677) );
  XNOR U37146 ( .A(n18673), .B(n18675), .Z(n35270) );
  XNOR U37147 ( .A(q[0]), .B(DB[2373]), .Z(n18675) );
  XNOR U37148 ( .A(q[3]), .B(DB[2376]), .Z(n18673) );
  IV U37149 ( .A(n18672), .Z(n35269) );
  XNOR U37150 ( .A(n18670), .B(n35271), .Z(n18672) );
  XNOR U37151 ( .A(q[2]), .B(DB[2375]), .Z(n35271) );
  XNOR U37152 ( .A(q[1]), .B(DB[2374]), .Z(n18670) );
  XOR U37153 ( .A(n35272), .B(n18635), .Z(n18598) );
  XOR U37154 ( .A(n35273), .B(n18623), .Z(n18635) );
  XNOR U37155 ( .A(q[6]), .B(DB[2386]), .Z(n18623) );
  IV U37156 ( .A(n18622), .Z(n35273) );
  XNOR U37157 ( .A(n18620), .B(n35274), .Z(n18622) );
  XNOR U37158 ( .A(q[5]), .B(DB[2385]), .Z(n35274) );
  XNOR U37159 ( .A(q[4]), .B(DB[2384]), .Z(n18620) );
  IV U37160 ( .A(n18634), .Z(n35272) );
  XOR U37161 ( .A(n35275), .B(n35276), .Z(n18634) );
  XNOR U37162 ( .A(n18630), .B(n18632), .Z(n35276) );
  XNOR U37163 ( .A(q[0]), .B(DB[2380]), .Z(n18632) );
  XNOR U37164 ( .A(q[3]), .B(DB[2383]), .Z(n18630) );
  IV U37165 ( .A(n18629), .Z(n35275) );
  XNOR U37166 ( .A(n18627), .B(n35277), .Z(n18629) );
  XNOR U37167 ( .A(q[2]), .B(DB[2382]), .Z(n35277) );
  XNOR U37168 ( .A(q[1]), .B(DB[2381]), .Z(n18627) );
  XOR U37169 ( .A(n35278), .B(n18592), .Z(n18555) );
  XOR U37170 ( .A(n35279), .B(n18580), .Z(n18592) );
  XNOR U37171 ( .A(q[6]), .B(DB[2393]), .Z(n18580) );
  IV U37172 ( .A(n18579), .Z(n35279) );
  XNOR U37173 ( .A(n18577), .B(n35280), .Z(n18579) );
  XNOR U37174 ( .A(q[5]), .B(DB[2392]), .Z(n35280) );
  XNOR U37175 ( .A(q[4]), .B(DB[2391]), .Z(n18577) );
  IV U37176 ( .A(n18591), .Z(n35278) );
  XOR U37177 ( .A(n35281), .B(n35282), .Z(n18591) );
  XNOR U37178 ( .A(n18587), .B(n18589), .Z(n35282) );
  XNOR U37179 ( .A(q[0]), .B(DB[2387]), .Z(n18589) );
  XNOR U37180 ( .A(q[3]), .B(DB[2390]), .Z(n18587) );
  IV U37181 ( .A(n18586), .Z(n35281) );
  XNOR U37182 ( .A(n18584), .B(n35283), .Z(n18586) );
  XNOR U37183 ( .A(q[2]), .B(DB[2389]), .Z(n35283) );
  XNOR U37184 ( .A(q[1]), .B(DB[2388]), .Z(n18584) );
  XOR U37185 ( .A(n35284), .B(n18549), .Z(n18512) );
  XOR U37186 ( .A(n35285), .B(n18537), .Z(n18549) );
  XNOR U37187 ( .A(q[6]), .B(DB[2400]), .Z(n18537) );
  IV U37188 ( .A(n18536), .Z(n35285) );
  XNOR U37189 ( .A(n18534), .B(n35286), .Z(n18536) );
  XNOR U37190 ( .A(q[5]), .B(DB[2399]), .Z(n35286) );
  XNOR U37191 ( .A(q[4]), .B(DB[2398]), .Z(n18534) );
  IV U37192 ( .A(n18548), .Z(n35284) );
  XOR U37193 ( .A(n35287), .B(n35288), .Z(n18548) );
  XNOR U37194 ( .A(n18544), .B(n18546), .Z(n35288) );
  XNOR U37195 ( .A(q[0]), .B(DB[2394]), .Z(n18546) );
  XNOR U37196 ( .A(q[3]), .B(DB[2397]), .Z(n18544) );
  IV U37197 ( .A(n18543), .Z(n35287) );
  XNOR U37198 ( .A(n18541), .B(n35289), .Z(n18543) );
  XNOR U37199 ( .A(q[2]), .B(DB[2396]), .Z(n35289) );
  XNOR U37200 ( .A(q[1]), .B(DB[2395]), .Z(n18541) );
  XOR U37201 ( .A(n35290), .B(n18506), .Z(n18469) );
  XOR U37202 ( .A(n35291), .B(n18494), .Z(n18506) );
  XNOR U37203 ( .A(q[6]), .B(DB[2407]), .Z(n18494) );
  IV U37204 ( .A(n18493), .Z(n35291) );
  XNOR U37205 ( .A(n18491), .B(n35292), .Z(n18493) );
  XNOR U37206 ( .A(q[5]), .B(DB[2406]), .Z(n35292) );
  XNOR U37207 ( .A(q[4]), .B(DB[2405]), .Z(n18491) );
  IV U37208 ( .A(n18505), .Z(n35290) );
  XOR U37209 ( .A(n35293), .B(n35294), .Z(n18505) );
  XNOR U37210 ( .A(n18501), .B(n18503), .Z(n35294) );
  XNOR U37211 ( .A(q[0]), .B(DB[2401]), .Z(n18503) );
  XNOR U37212 ( .A(q[3]), .B(DB[2404]), .Z(n18501) );
  IV U37213 ( .A(n18500), .Z(n35293) );
  XNOR U37214 ( .A(n18498), .B(n35295), .Z(n18500) );
  XNOR U37215 ( .A(q[2]), .B(DB[2403]), .Z(n35295) );
  XNOR U37216 ( .A(q[1]), .B(DB[2402]), .Z(n18498) );
  XOR U37217 ( .A(n35296), .B(n18463), .Z(n18426) );
  XOR U37218 ( .A(n35297), .B(n18451), .Z(n18463) );
  XNOR U37219 ( .A(q[6]), .B(DB[2414]), .Z(n18451) );
  IV U37220 ( .A(n18450), .Z(n35297) );
  XNOR U37221 ( .A(n18448), .B(n35298), .Z(n18450) );
  XNOR U37222 ( .A(q[5]), .B(DB[2413]), .Z(n35298) );
  XNOR U37223 ( .A(q[4]), .B(DB[2412]), .Z(n18448) );
  IV U37224 ( .A(n18462), .Z(n35296) );
  XOR U37225 ( .A(n35299), .B(n35300), .Z(n18462) );
  XNOR U37226 ( .A(n18458), .B(n18460), .Z(n35300) );
  XNOR U37227 ( .A(q[0]), .B(DB[2408]), .Z(n18460) );
  XNOR U37228 ( .A(q[3]), .B(DB[2411]), .Z(n18458) );
  IV U37229 ( .A(n18457), .Z(n35299) );
  XNOR U37230 ( .A(n18455), .B(n35301), .Z(n18457) );
  XNOR U37231 ( .A(q[2]), .B(DB[2410]), .Z(n35301) );
  XNOR U37232 ( .A(q[1]), .B(DB[2409]), .Z(n18455) );
  XOR U37233 ( .A(n35302), .B(n18420), .Z(n18383) );
  XOR U37234 ( .A(n35303), .B(n18408), .Z(n18420) );
  XNOR U37235 ( .A(q[6]), .B(DB[2421]), .Z(n18408) );
  IV U37236 ( .A(n18407), .Z(n35303) );
  XNOR U37237 ( .A(n18405), .B(n35304), .Z(n18407) );
  XNOR U37238 ( .A(q[5]), .B(DB[2420]), .Z(n35304) );
  XNOR U37239 ( .A(q[4]), .B(DB[2419]), .Z(n18405) );
  IV U37240 ( .A(n18419), .Z(n35302) );
  XOR U37241 ( .A(n35305), .B(n35306), .Z(n18419) );
  XNOR U37242 ( .A(n18415), .B(n18417), .Z(n35306) );
  XNOR U37243 ( .A(q[0]), .B(DB[2415]), .Z(n18417) );
  XNOR U37244 ( .A(q[3]), .B(DB[2418]), .Z(n18415) );
  IV U37245 ( .A(n18414), .Z(n35305) );
  XNOR U37246 ( .A(n18412), .B(n35307), .Z(n18414) );
  XNOR U37247 ( .A(q[2]), .B(DB[2417]), .Z(n35307) );
  XNOR U37248 ( .A(q[1]), .B(DB[2416]), .Z(n18412) );
  XOR U37249 ( .A(n35308), .B(n18377), .Z(n18340) );
  XOR U37250 ( .A(n35309), .B(n18365), .Z(n18377) );
  XNOR U37251 ( .A(q[6]), .B(DB[2428]), .Z(n18365) );
  IV U37252 ( .A(n18364), .Z(n35309) );
  XNOR U37253 ( .A(n18362), .B(n35310), .Z(n18364) );
  XNOR U37254 ( .A(q[5]), .B(DB[2427]), .Z(n35310) );
  XNOR U37255 ( .A(q[4]), .B(DB[2426]), .Z(n18362) );
  IV U37256 ( .A(n18376), .Z(n35308) );
  XOR U37257 ( .A(n35311), .B(n35312), .Z(n18376) );
  XNOR U37258 ( .A(n18372), .B(n18374), .Z(n35312) );
  XNOR U37259 ( .A(q[0]), .B(DB[2422]), .Z(n18374) );
  XNOR U37260 ( .A(q[3]), .B(DB[2425]), .Z(n18372) );
  IV U37261 ( .A(n18371), .Z(n35311) );
  XNOR U37262 ( .A(n18369), .B(n35313), .Z(n18371) );
  XNOR U37263 ( .A(q[2]), .B(DB[2424]), .Z(n35313) );
  XNOR U37264 ( .A(q[1]), .B(DB[2423]), .Z(n18369) );
  XOR U37265 ( .A(n35314), .B(n18334), .Z(n18297) );
  XOR U37266 ( .A(n35315), .B(n18322), .Z(n18334) );
  XNOR U37267 ( .A(q[6]), .B(DB[2435]), .Z(n18322) );
  IV U37268 ( .A(n18321), .Z(n35315) );
  XNOR U37269 ( .A(n18319), .B(n35316), .Z(n18321) );
  XNOR U37270 ( .A(q[5]), .B(DB[2434]), .Z(n35316) );
  XNOR U37271 ( .A(q[4]), .B(DB[2433]), .Z(n18319) );
  IV U37272 ( .A(n18333), .Z(n35314) );
  XOR U37273 ( .A(n35317), .B(n35318), .Z(n18333) );
  XNOR U37274 ( .A(n18329), .B(n18331), .Z(n35318) );
  XNOR U37275 ( .A(q[0]), .B(DB[2429]), .Z(n18331) );
  XNOR U37276 ( .A(q[3]), .B(DB[2432]), .Z(n18329) );
  IV U37277 ( .A(n18328), .Z(n35317) );
  XNOR U37278 ( .A(n18326), .B(n35319), .Z(n18328) );
  XNOR U37279 ( .A(q[2]), .B(DB[2431]), .Z(n35319) );
  XNOR U37280 ( .A(q[1]), .B(DB[2430]), .Z(n18326) );
  XOR U37281 ( .A(n35320), .B(n18291), .Z(n18254) );
  XOR U37282 ( .A(n35321), .B(n18279), .Z(n18291) );
  XNOR U37283 ( .A(q[6]), .B(DB[2442]), .Z(n18279) );
  IV U37284 ( .A(n18278), .Z(n35321) );
  XNOR U37285 ( .A(n18276), .B(n35322), .Z(n18278) );
  XNOR U37286 ( .A(q[5]), .B(DB[2441]), .Z(n35322) );
  XNOR U37287 ( .A(q[4]), .B(DB[2440]), .Z(n18276) );
  IV U37288 ( .A(n18290), .Z(n35320) );
  XOR U37289 ( .A(n35323), .B(n35324), .Z(n18290) );
  XNOR U37290 ( .A(n18286), .B(n18288), .Z(n35324) );
  XNOR U37291 ( .A(q[0]), .B(DB[2436]), .Z(n18288) );
  XNOR U37292 ( .A(q[3]), .B(DB[2439]), .Z(n18286) );
  IV U37293 ( .A(n18285), .Z(n35323) );
  XNOR U37294 ( .A(n18283), .B(n35325), .Z(n18285) );
  XNOR U37295 ( .A(q[2]), .B(DB[2438]), .Z(n35325) );
  XNOR U37296 ( .A(q[1]), .B(DB[2437]), .Z(n18283) );
  XOR U37297 ( .A(n35326), .B(n18248), .Z(n18211) );
  XOR U37298 ( .A(n35327), .B(n18236), .Z(n18248) );
  XNOR U37299 ( .A(q[6]), .B(DB[2449]), .Z(n18236) );
  IV U37300 ( .A(n18235), .Z(n35327) );
  XNOR U37301 ( .A(n18233), .B(n35328), .Z(n18235) );
  XNOR U37302 ( .A(q[5]), .B(DB[2448]), .Z(n35328) );
  XNOR U37303 ( .A(q[4]), .B(DB[2447]), .Z(n18233) );
  IV U37304 ( .A(n18247), .Z(n35326) );
  XOR U37305 ( .A(n35329), .B(n35330), .Z(n18247) );
  XNOR U37306 ( .A(n18243), .B(n18245), .Z(n35330) );
  XNOR U37307 ( .A(q[0]), .B(DB[2443]), .Z(n18245) );
  XNOR U37308 ( .A(q[3]), .B(DB[2446]), .Z(n18243) );
  IV U37309 ( .A(n18242), .Z(n35329) );
  XNOR U37310 ( .A(n18240), .B(n35331), .Z(n18242) );
  XNOR U37311 ( .A(q[2]), .B(DB[2445]), .Z(n35331) );
  XNOR U37312 ( .A(q[1]), .B(DB[2444]), .Z(n18240) );
  XOR U37313 ( .A(n35332), .B(n18205), .Z(n18168) );
  XOR U37314 ( .A(n35333), .B(n18193), .Z(n18205) );
  XNOR U37315 ( .A(q[6]), .B(DB[2456]), .Z(n18193) );
  IV U37316 ( .A(n18192), .Z(n35333) );
  XNOR U37317 ( .A(n18190), .B(n35334), .Z(n18192) );
  XNOR U37318 ( .A(q[5]), .B(DB[2455]), .Z(n35334) );
  XNOR U37319 ( .A(q[4]), .B(DB[2454]), .Z(n18190) );
  IV U37320 ( .A(n18204), .Z(n35332) );
  XOR U37321 ( .A(n35335), .B(n35336), .Z(n18204) );
  XNOR U37322 ( .A(n18200), .B(n18202), .Z(n35336) );
  XNOR U37323 ( .A(q[0]), .B(DB[2450]), .Z(n18202) );
  XNOR U37324 ( .A(q[3]), .B(DB[2453]), .Z(n18200) );
  IV U37325 ( .A(n18199), .Z(n35335) );
  XNOR U37326 ( .A(n18197), .B(n35337), .Z(n18199) );
  XNOR U37327 ( .A(q[2]), .B(DB[2452]), .Z(n35337) );
  XNOR U37328 ( .A(q[1]), .B(DB[2451]), .Z(n18197) );
  XOR U37329 ( .A(n35338), .B(n18162), .Z(n18125) );
  XOR U37330 ( .A(n35339), .B(n18150), .Z(n18162) );
  XNOR U37331 ( .A(q[6]), .B(DB[2463]), .Z(n18150) );
  IV U37332 ( .A(n18149), .Z(n35339) );
  XNOR U37333 ( .A(n18147), .B(n35340), .Z(n18149) );
  XNOR U37334 ( .A(q[5]), .B(DB[2462]), .Z(n35340) );
  XNOR U37335 ( .A(q[4]), .B(DB[2461]), .Z(n18147) );
  IV U37336 ( .A(n18161), .Z(n35338) );
  XOR U37337 ( .A(n35341), .B(n35342), .Z(n18161) );
  XNOR U37338 ( .A(n18157), .B(n18159), .Z(n35342) );
  XNOR U37339 ( .A(q[0]), .B(DB[2457]), .Z(n18159) );
  XNOR U37340 ( .A(q[3]), .B(DB[2460]), .Z(n18157) );
  IV U37341 ( .A(n18156), .Z(n35341) );
  XNOR U37342 ( .A(n18154), .B(n35343), .Z(n18156) );
  XNOR U37343 ( .A(q[2]), .B(DB[2459]), .Z(n35343) );
  XNOR U37344 ( .A(q[1]), .B(DB[2458]), .Z(n18154) );
  XOR U37345 ( .A(n35344), .B(n18119), .Z(n18082) );
  XOR U37346 ( .A(n35345), .B(n18107), .Z(n18119) );
  XNOR U37347 ( .A(q[6]), .B(DB[2470]), .Z(n18107) );
  IV U37348 ( .A(n18106), .Z(n35345) );
  XNOR U37349 ( .A(n18104), .B(n35346), .Z(n18106) );
  XNOR U37350 ( .A(q[5]), .B(DB[2469]), .Z(n35346) );
  XNOR U37351 ( .A(q[4]), .B(DB[2468]), .Z(n18104) );
  IV U37352 ( .A(n18118), .Z(n35344) );
  XOR U37353 ( .A(n35347), .B(n35348), .Z(n18118) );
  XNOR U37354 ( .A(n18114), .B(n18116), .Z(n35348) );
  XNOR U37355 ( .A(q[0]), .B(DB[2464]), .Z(n18116) );
  XNOR U37356 ( .A(q[3]), .B(DB[2467]), .Z(n18114) );
  IV U37357 ( .A(n18113), .Z(n35347) );
  XNOR U37358 ( .A(n18111), .B(n35349), .Z(n18113) );
  XNOR U37359 ( .A(q[2]), .B(DB[2466]), .Z(n35349) );
  XNOR U37360 ( .A(q[1]), .B(DB[2465]), .Z(n18111) );
  XOR U37361 ( .A(n35350), .B(n18076), .Z(n18039) );
  XOR U37362 ( .A(n35351), .B(n18064), .Z(n18076) );
  XNOR U37363 ( .A(q[6]), .B(DB[2477]), .Z(n18064) );
  IV U37364 ( .A(n18063), .Z(n35351) );
  XNOR U37365 ( .A(n18061), .B(n35352), .Z(n18063) );
  XNOR U37366 ( .A(q[5]), .B(DB[2476]), .Z(n35352) );
  XNOR U37367 ( .A(q[4]), .B(DB[2475]), .Z(n18061) );
  IV U37368 ( .A(n18075), .Z(n35350) );
  XOR U37369 ( .A(n35353), .B(n35354), .Z(n18075) );
  XNOR U37370 ( .A(n18071), .B(n18073), .Z(n35354) );
  XNOR U37371 ( .A(q[0]), .B(DB[2471]), .Z(n18073) );
  XNOR U37372 ( .A(q[3]), .B(DB[2474]), .Z(n18071) );
  IV U37373 ( .A(n18070), .Z(n35353) );
  XNOR U37374 ( .A(n18068), .B(n35355), .Z(n18070) );
  XNOR U37375 ( .A(q[2]), .B(DB[2473]), .Z(n35355) );
  XNOR U37376 ( .A(q[1]), .B(DB[2472]), .Z(n18068) );
  XOR U37377 ( .A(n35356), .B(n18033), .Z(n17996) );
  XOR U37378 ( .A(n35357), .B(n18021), .Z(n18033) );
  XNOR U37379 ( .A(q[6]), .B(DB[2484]), .Z(n18021) );
  IV U37380 ( .A(n18020), .Z(n35357) );
  XNOR U37381 ( .A(n18018), .B(n35358), .Z(n18020) );
  XNOR U37382 ( .A(q[5]), .B(DB[2483]), .Z(n35358) );
  XNOR U37383 ( .A(q[4]), .B(DB[2482]), .Z(n18018) );
  IV U37384 ( .A(n18032), .Z(n35356) );
  XOR U37385 ( .A(n35359), .B(n35360), .Z(n18032) );
  XNOR U37386 ( .A(n18028), .B(n18030), .Z(n35360) );
  XNOR U37387 ( .A(q[0]), .B(DB[2478]), .Z(n18030) );
  XNOR U37388 ( .A(q[3]), .B(DB[2481]), .Z(n18028) );
  IV U37389 ( .A(n18027), .Z(n35359) );
  XNOR U37390 ( .A(n18025), .B(n35361), .Z(n18027) );
  XNOR U37391 ( .A(q[2]), .B(DB[2480]), .Z(n35361) );
  XNOR U37392 ( .A(q[1]), .B(DB[2479]), .Z(n18025) );
  XOR U37393 ( .A(n35362), .B(n17990), .Z(n17953) );
  XOR U37394 ( .A(n35363), .B(n17978), .Z(n17990) );
  XNOR U37395 ( .A(q[6]), .B(DB[2491]), .Z(n17978) );
  IV U37396 ( .A(n17977), .Z(n35363) );
  XNOR U37397 ( .A(n17975), .B(n35364), .Z(n17977) );
  XNOR U37398 ( .A(q[5]), .B(DB[2490]), .Z(n35364) );
  XNOR U37399 ( .A(q[4]), .B(DB[2489]), .Z(n17975) );
  IV U37400 ( .A(n17989), .Z(n35362) );
  XOR U37401 ( .A(n35365), .B(n35366), .Z(n17989) );
  XNOR U37402 ( .A(n17985), .B(n17987), .Z(n35366) );
  XNOR U37403 ( .A(q[0]), .B(DB[2485]), .Z(n17987) );
  XNOR U37404 ( .A(q[3]), .B(DB[2488]), .Z(n17985) );
  IV U37405 ( .A(n17984), .Z(n35365) );
  XNOR U37406 ( .A(n17982), .B(n35367), .Z(n17984) );
  XNOR U37407 ( .A(q[2]), .B(DB[2487]), .Z(n35367) );
  XNOR U37408 ( .A(q[1]), .B(DB[2486]), .Z(n17982) );
  XOR U37409 ( .A(n35368), .B(n17947), .Z(n17910) );
  XOR U37410 ( .A(n35369), .B(n17935), .Z(n17947) );
  XNOR U37411 ( .A(q[6]), .B(DB[2498]), .Z(n17935) );
  IV U37412 ( .A(n17934), .Z(n35369) );
  XNOR U37413 ( .A(n17932), .B(n35370), .Z(n17934) );
  XNOR U37414 ( .A(q[5]), .B(DB[2497]), .Z(n35370) );
  XNOR U37415 ( .A(q[4]), .B(DB[2496]), .Z(n17932) );
  IV U37416 ( .A(n17946), .Z(n35368) );
  XOR U37417 ( .A(n35371), .B(n35372), .Z(n17946) );
  XNOR U37418 ( .A(n17942), .B(n17944), .Z(n35372) );
  XNOR U37419 ( .A(q[0]), .B(DB[2492]), .Z(n17944) );
  XNOR U37420 ( .A(q[3]), .B(DB[2495]), .Z(n17942) );
  IV U37421 ( .A(n17941), .Z(n35371) );
  XNOR U37422 ( .A(n17939), .B(n35373), .Z(n17941) );
  XNOR U37423 ( .A(q[2]), .B(DB[2494]), .Z(n35373) );
  XNOR U37424 ( .A(q[1]), .B(DB[2493]), .Z(n17939) );
  XOR U37425 ( .A(n35374), .B(n17904), .Z(n17867) );
  XOR U37426 ( .A(n35375), .B(n17892), .Z(n17904) );
  XNOR U37427 ( .A(q[6]), .B(DB[2505]), .Z(n17892) );
  IV U37428 ( .A(n17891), .Z(n35375) );
  XNOR U37429 ( .A(n17889), .B(n35376), .Z(n17891) );
  XNOR U37430 ( .A(q[5]), .B(DB[2504]), .Z(n35376) );
  XNOR U37431 ( .A(q[4]), .B(DB[2503]), .Z(n17889) );
  IV U37432 ( .A(n17903), .Z(n35374) );
  XOR U37433 ( .A(n35377), .B(n35378), .Z(n17903) );
  XNOR U37434 ( .A(n17899), .B(n17901), .Z(n35378) );
  XNOR U37435 ( .A(q[0]), .B(DB[2499]), .Z(n17901) );
  XNOR U37436 ( .A(q[3]), .B(DB[2502]), .Z(n17899) );
  IV U37437 ( .A(n17898), .Z(n35377) );
  XNOR U37438 ( .A(n17896), .B(n35379), .Z(n17898) );
  XNOR U37439 ( .A(q[2]), .B(DB[2501]), .Z(n35379) );
  XNOR U37440 ( .A(q[1]), .B(DB[2500]), .Z(n17896) );
  XOR U37441 ( .A(n35380), .B(n17861), .Z(n17824) );
  XOR U37442 ( .A(n35381), .B(n17849), .Z(n17861) );
  XNOR U37443 ( .A(q[6]), .B(DB[2512]), .Z(n17849) );
  IV U37444 ( .A(n17848), .Z(n35381) );
  XNOR U37445 ( .A(n17846), .B(n35382), .Z(n17848) );
  XNOR U37446 ( .A(q[5]), .B(DB[2511]), .Z(n35382) );
  XNOR U37447 ( .A(q[4]), .B(DB[2510]), .Z(n17846) );
  IV U37448 ( .A(n17860), .Z(n35380) );
  XOR U37449 ( .A(n35383), .B(n35384), .Z(n17860) );
  XNOR U37450 ( .A(n17856), .B(n17858), .Z(n35384) );
  XNOR U37451 ( .A(q[0]), .B(DB[2506]), .Z(n17858) );
  XNOR U37452 ( .A(q[3]), .B(DB[2509]), .Z(n17856) );
  IV U37453 ( .A(n17855), .Z(n35383) );
  XNOR U37454 ( .A(n17853), .B(n35385), .Z(n17855) );
  XNOR U37455 ( .A(q[2]), .B(DB[2508]), .Z(n35385) );
  XNOR U37456 ( .A(q[1]), .B(DB[2507]), .Z(n17853) );
  XOR U37457 ( .A(n35386), .B(n17818), .Z(n17781) );
  XOR U37458 ( .A(n35387), .B(n17806), .Z(n17818) );
  XNOR U37459 ( .A(q[6]), .B(DB[2519]), .Z(n17806) );
  IV U37460 ( .A(n17805), .Z(n35387) );
  XNOR U37461 ( .A(n17803), .B(n35388), .Z(n17805) );
  XNOR U37462 ( .A(q[5]), .B(DB[2518]), .Z(n35388) );
  XNOR U37463 ( .A(q[4]), .B(DB[2517]), .Z(n17803) );
  IV U37464 ( .A(n17817), .Z(n35386) );
  XOR U37465 ( .A(n35389), .B(n35390), .Z(n17817) );
  XNOR U37466 ( .A(n17813), .B(n17815), .Z(n35390) );
  XNOR U37467 ( .A(q[0]), .B(DB[2513]), .Z(n17815) );
  XNOR U37468 ( .A(q[3]), .B(DB[2516]), .Z(n17813) );
  IV U37469 ( .A(n17812), .Z(n35389) );
  XNOR U37470 ( .A(n17810), .B(n35391), .Z(n17812) );
  XNOR U37471 ( .A(q[2]), .B(DB[2515]), .Z(n35391) );
  XNOR U37472 ( .A(q[1]), .B(DB[2514]), .Z(n17810) );
  XOR U37473 ( .A(n35392), .B(n17775), .Z(n17738) );
  XOR U37474 ( .A(n35393), .B(n17763), .Z(n17775) );
  XNOR U37475 ( .A(q[6]), .B(DB[2526]), .Z(n17763) );
  IV U37476 ( .A(n17762), .Z(n35393) );
  XNOR U37477 ( .A(n17760), .B(n35394), .Z(n17762) );
  XNOR U37478 ( .A(q[5]), .B(DB[2525]), .Z(n35394) );
  XNOR U37479 ( .A(q[4]), .B(DB[2524]), .Z(n17760) );
  IV U37480 ( .A(n17774), .Z(n35392) );
  XOR U37481 ( .A(n35395), .B(n35396), .Z(n17774) );
  XNOR U37482 ( .A(n17770), .B(n17772), .Z(n35396) );
  XNOR U37483 ( .A(q[0]), .B(DB[2520]), .Z(n17772) );
  XNOR U37484 ( .A(q[3]), .B(DB[2523]), .Z(n17770) );
  IV U37485 ( .A(n17769), .Z(n35395) );
  XNOR U37486 ( .A(n17767), .B(n35397), .Z(n17769) );
  XNOR U37487 ( .A(q[2]), .B(DB[2522]), .Z(n35397) );
  XNOR U37488 ( .A(q[1]), .B(DB[2521]), .Z(n17767) );
  XOR U37489 ( .A(n35398), .B(n17732), .Z(n17695) );
  XOR U37490 ( .A(n35399), .B(n17720), .Z(n17732) );
  XNOR U37491 ( .A(q[6]), .B(DB[2533]), .Z(n17720) );
  IV U37492 ( .A(n17719), .Z(n35399) );
  XNOR U37493 ( .A(n17717), .B(n35400), .Z(n17719) );
  XNOR U37494 ( .A(q[5]), .B(DB[2532]), .Z(n35400) );
  XNOR U37495 ( .A(q[4]), .B(DB[2531]), .Z(n17717) );
  IV U37496 ( .A(n17731), .Z(n35398) );
  XOR U37497 ( .A(n35401), .B(n35402), .Z(n17731) );
  XNOR U37498 ( .A(n17727), .B(n17729), .Z(n35402) );
  XNOR U37499 ( .A(q[0]), .B(DB[2527]), .Z(n17729) );
  XNOR U37500 ( .A(q[3]), .B(DB[2530]), .Z(n17727) );
  IV U37501 ( .A(n17726), .Z(n35401) );
  XNOR U37502 ( .A(n17724), .B(n35403), .Z(n17726) );
  XNOR U37503 ( .A(q[2]), .B(DB[2529]), .Z(n35403) );
  XNOR U37504 ( .A(q[1]), .B(DB[2528]), .Z(n17724) );
  XOR U37505 ( .A(n35404), .B(n17689), .Z(n17652) );
  XOR U37506 ( .A(n35405), .B(n17677), .Z(n17689) );
  XNOR U37507 ( .A(q[6]), .B(DB[2540]), .Z(n17677) );
  IV U37508 ( .A(n17676), .Z(n35405) );
  XNOR U37509 ( .A(n17674), .B(n35406), .Z(n17676) );
  XNOR U37510 ( .A(q[5]), .B(DB[2539]), .Z(n35406) );
  XNOR U37511 ( .A(q[4]), .B(DB[2538]), .Z(n17674) );
  IV U37512 ( .A(n17688), .Z(n35404) );
  XOR U37513 ( .A(n35407), .B(n35408), .Z(n17688) );
  XNOR U37514 ( .A(n17684), .B(n17686), .Z(n35408) );
  XNOR U37515 ( .A(q[0]), .B(DB[2534]), .Z(n17686) );
  XNOR U37516 ( .A(q[3]), .B(DB[2537]), .Z(n17684) );
  IV U37517 ( .A(n17683), .Z(n35407) );
  XNOR U37518 ( .A(n17681), .B(n35409), .Z(n17683) );
  XNOR U37519 ( .A(q[2]), .B(DB[2536]), .Z(n35409) );
  XNOR U37520 ( .A(q[1]), .B(DB[2535]), .Z(n17681) );
  XOR U37521 ( .A(n35410), .B(n17646), .Z(n17609) );
  XOR U37522 ( .A(n35411), .B(n17634), .Z(n17646) );
  XNOR U37523 ( .A(q[6]), .B(DB[2547]), .Z(n17634) );
  IV U37524 ( .A(n17633), .Z(n35411) );
  XNOR U37525 ( .A(n17631), .B(n35412), .Z(n17633) );
  XNOR U37526 ( .A(q[5]), .B(DB[2546]), .Z(n35412) );
  XNOR U37527 ( .A(q[4]), .B(DB[2545]), .Z(n17631) );
  IV U37528 ( .A(n17645), .Z(n35410) );
  XOR U37529 ( .A(n35413), .B(n35414), .Z(n17645) );
  XNOR U37530 ( .A(n17641), .B(n17643), .Z(n35414) );
  XNOR U37531 ( .A(q[0]), .B(DB[2541]), .Z(n17643) );
  XNOR U37532 ( .A(q[3]), .B(DB[2544]), .Z(n17641) );
  IV U37533 ( .A(n17640), .Z(n35413) );
  XNOR U37534 ( .A(n17638), .B(n35415), .Z(n17640) );
  XNOR U37535 ( .A(q[2]), .B(DB[2543]), .Z(n35415) );
  XNOR U37536 ( .A(q[1]), .B(DB[2542]), .Z(n17638) );
  XOR U37537 ( .A(n35416), .B(n17603), .Z(n17566) );
  XOR U37538 ( .A(n35417), .B(n17591), .Z(n17603) );
  XNOR U37539 ( .A(q[6]), .B(DB[2554]), .Z(n17591) );
  IV U37540 ( .A(n17590), .Z(n35417) );
  XNOR U37541 ( .A(n17588), .B(n35418), .Z(n17590) );
  XNOR U37542 ( .A(q[5]), .B(DB[2553]), .Z(n35418) );
  XNOR U37543 ( .A(q[4]), .B(DB[2552]), .Z(n17588) );
  IV U37544 ( .A(n17602), .Z(n35416) );
  XOR U37545 ( .A(n35419), .B(n35420), .Z(n17602) );
  XNOR U37546 ( .A(n17598), .B(n17600), .Z(n35420) );
  XNOR U37547 ( .A(q[0]), .B(DB[2548]), .Z(n17600) );
  XNOR U37548 ( .A(q[3]), .B(DB[2551]), .Z(n17598) );
  IV U37549 ( .A(n17597), .Z(n35419) );
  XNOR U37550 ( .A(n17595), .B(n35421), .Z(n17597) );
  XNOR U37551 ( .A(q[2]), .B(DB[2550]), .Z(n35421) );
  XNOR U37552 ( .A(q[1]), .B(DB[2549]), .Z(n17595) );
  XOR U37553 ( .A(n35422), .B(n17560), .Z(n17523) );
  XOR U37554 ( .A(n35423), .B(n17548), .Z(n17560) );
  XNOR U37555 ( .A(q[6]), .B(DB[2561]), .Z(n17548) );
  IV U37556 ( .A(n17547), .Z(n35423) );
  XNOR U37557 ( .A(n17545), .B(n35424), .Z(n17547) );
  XNOR U37558 ( .A(q[5]), .B(DB[2560]), .Z(n35424) );
  XNOR U37559 ( .A(q[4]), .B(DB[2559]), .Z(n17545) );
  IV U37560 ( .A(n17559), .Z(n35422) );
  XOR U37561 ( .A(n35425), .B(n35426), .Z(n17559) );
  XNOR U37562 ( .A(n17555), .B(n17557), .Z(n35426) );
  XNOR U37563 ( .A(q[0]), .B(DB[2555]), .Z(n17557) );
  XNOR U37564 ( .A(q[3]), .B(DB[2558]), .Z(n17555) );
  IV U37565 ( .A(n17554), .Z(n35425) );
  XNOR U37566 ( .A(n17552), .B(n35427), .Z(n17554) );
  XNOR U37567 ( .A(q[2]), .B(DB[2557]), .Z(n35427) );
  XNOR U37568 ( .A(q[1]), .B(DB[2556]), .Z(n17552) );
  XOR U37569 ( .A(n35428), .B(n17517), .Z(n17480) );
  XOR U37570 ( .A(n35429), .B(n17505), .Z(n17517) );
  XNOR U37571 ( .A(q[6]), .B(DB[2568]), .Z(n17505) );
  IV U37572 ( .A(n17504), .Z(n35429) );
  XNOR U37573 ( .A(n17502), .B(n35430), .Z(n17504) );
  XNOR U37574 ( .A(q[5]), .B(DB[2567]), .Z(n35430) );
  XNOR U37575 ( .A(q[4]), .B(DB[2566]), .Z(n17502) );
  IV U37576 ( .A(n17516), .Z(n35428) );
  XOR U37577 ( .A(n35431), .B(n35432), .Z(n17516) );
  XNOR U37578 ( .A(n17512), .B(n17514), .Z(n35432) );
  XNOR U37579 ( .A(q[0]), .B(DB[2562]), .Z(n17514) );
  XNOR U37580 ( .A(q[3]), .B(DB[2565]), .Z(n17512) );
  IV U37581 ( .A(n17511), .Z(n35431) );
  XNOR U37582 ( .A(n17509), .B(n35433), .Z(n17511) );
  XNOR U37583 ( .A(q[2]), .B(DB[2564]), .Z(n35433) );
  XNOR U37584 ( .A(q[1]), .B(DB[2563]), .Z(n17509) );
  XOR U37585 ( .A(n35434), .B(n17474), .Z(n17437) );
  XOR U37586 ( .A(n35435), .B(n17462), .Z(n17474) );
  XNOR U37587 ( .A(q[6]), .B(DB[2575]), .Z(n17462) );
  IV U37588 ( .A(n17461), .Z(n35435) );
  XNOR U37589 ( .A(n17459), .B(n35436), .Z(n17461) );
  XNOR U37590 ( .A(q[5]), .B(DB[2574]), .Z(n35436) );
  XNOR U37591 ( .A(q[4]), .B(DB[2573]), .Z(n17459) );
  IV U37592 ( .A(n17473), .Z(n35434) );
  XOR U37593 ( .A(n35437), .B(n35438), .Z(n17473) );
  XNOR U37594 ( .A(n17469), .B(n17471), .Z(n35438) );
  XNOR U37595 ( .A(q[0]), .B(DB[2569]), .Z(n17471) );
  XNOR U37596 ( .A(q[3]), .B(DB[2572]), .Z(n17469) );
  IV U37597 ( .A(n17468), .Z(n35437) );
  XNOR U37598 ( .A(n17466), .B(n35439), .Z(n17468) );
  XNOR U37599 ( .A(q[2]), .B(DB[2571]), .Z(n35439) );
  XNOR U37600 ( .A(q[1]), .B(DB[2570]), .Z(n17466) );
  XOR U37601 ( .A(n35440), .B(n17431), .Z(n17394) );
  XOR U37602 ( .A(n35441), .B(n17419), .Z(n17431) );
  XNOR U37603 ( .A(q[6]), .B(DB[2582]), .Z(n17419) );
  IV U37604 ( .A(n17418), .Z(n35441) );
  XNOR U37605 ( .A(n17416), .B(n35442), .Z(n17418) );
  XNOR U37606 ( .A(q[5]), .B(DB[2581]), .Z(n35442) );
  XNOR U37607 ( .A(q[4]), .B(DB[2580]), .Z(n17416) );
  IV U37608 ( .A(n17430), .Z(n35440) );
  XOR U37609 ( .A(n35443), .B(n35444), .Z(n17430) );
  XNOR U37610 ( .A(n17426), .B(n17428), .Z(n35444) );
  XNOR U37611 ( .A(q[0]), .B(DB[2576]), .Z(n17428) );
  XNOR U37612 ( .A(q[3]), .B(DB[2579]), .Z(n17426) );
  IV U37613 ( .A(n17425), .Z(n35443) );
  XNOR U37614 ( .A(n17423), .B(n35445), .Z(n17425) );
  XNOR U37615 ( .A(q[2]), .B(DB[2578]), .Z(n35445) );
  XNOR U37616 ( .A(q[1]), .B(DB[2577]), .Z(n17423) );
  XOR U37617 ( .A(n35446), .B(n17388), .Z(n17351) );
  XOR U37618 ( .A(n35447), .B(n17376), .Z(n17388) );
  XNOR U37619 ( .A(q[6]), .B(DB[2589]), .Z(n17376) );
  IV U37620 ( .A(n17375), .Z(n35447) );
  XNOR U37621 ( .A(n17373), .B(n35448), .Z(n17375) );
  XNOR U37622 ( .A(q[5]), .B(DB[2588]), .Z(n35448) );
  XNOR U37623 ( .A(q[4]), .B(DB[2587]), .Z(n17373) );
  IV U37624 ( .A(n17387), .Z(n35446) );
  XOR U37625 ( .A(n35449), .B(n35450), .Z(n17387) );
  XNOR U37626 ( .A(n17383), .B(n17385), .Z(n35450) );
  XNOR U37627 ( .A(q[0]), .B(DB[2583]), .Z(n17385) );
  XNOR U37628 ( .A(q[3]), .B(DB[2586]), .Z(n17383) );
  IV U37629 ( .A(n17382), .Z(n35449) );
  XNOR U37630 ( .A(n17380), .B(n35451), .Z(n17382) );
  XNOR U37631 ( .A(q[2]), .B(DB[2585]), .Z(n35451) );
  XNOR U37632 ( .A(q[1]), .B(DB[2584]), .Z(n17380) );
  XOR U37633 ( .A(n35452), .B(n17345), .Z(n17308) );
  XOR U37634 ( .A(n35453), .B(n17333), .Z(n17345) );
  XNOR U37635 ( .A(q[6]), .B(DB[2596]), .Z(n17333) );
  IV U37636 ( .A(n17332), .Z(n35453) );
  XNOR U37637 ( .A(n17330), .B(n35454), .Z(n17332) );
  XNOR U37638 ( .A(q[5]), .B(DB[2595]), .Z(n35454) );
  XNOR U37639 ( .A(q[4]), .B(DB[2594]), .Z(n17330) );
  IV U37640 ( .A(n17344), .Z(n35452) );
  XOR U37641 ( .A(n35455), .B(n35456), .Z(n17344) );
  XNOR U37642 ( .A(n17340), .B(n17342), .Z(n35456) );
  XNOR U37643 ( .A(q[0]), .B(DB[2590]), .Z(n17342) );
  XNOR U37644 ( .A(q[3]), .B(DB[2593]), .Z(n17340) );
  IV U37645 ( .A(n17339), .Z(n35455) );
  XNOR U37646 ( .A(n17337), .B(n35457), .Z(n17339) );
  XNOR U37647 ( .A(q[2]), .B(DB[2592]), .Z(n35457) );
  XNOR U37648 ( .A(q[1]), .B(DB[2591]), .Z(n17337) );
  XOR U37649 ( .A(n35458), .B(n17302), .Z(n17265) );
  XOR U37650 ( .A(n35459), .B(n17290), .Z(n17302) );
  XNOR U37651 ( .A(q[6]), .B(DB[2603]), .Z(n17290) );
  IV U37652 ( .A(n17289), .Z(n35459) );
  XNOR U37653 ( .A(n17287), .B(n35460), .Z(n17289) );
  XNOR U37654 ( .A(q[5]), .B(DB[2602]), .Z(n35460) );
  XNOR U37655 ( .A(q[4]), .B(DB[2601]), .Z(n17287) );
  IV U37656 ( .A(n17301), .Z(n35458) );
  XOR U37657 ( .A(n35461), .B(n35462), .Z(n17301) );
  XNOR U37658 ( .A(n17297), .B(n17299), .Z(n35462) );
  XNOR U37659 ( .A(q[0]), .B(DB[2597]), .Z(n17299) );
  XNOR U37660 ( .A(q[3]), .B(DB[2600]), .Z(n17297) );
  IV U37661 ( .A(n17296), .Z(n35461) );
  XNOR U37662 ( .A(n17294), .B(n35463), .Z(n17296) );
  XNOR U37663 ( .A(q[2]), .B(DB[2599]), .Z(n35463) );
  XNOR U37664 ( .A(q[1]), .B(DB[2598]), .Z(n17294) );
  XOR U37665 ( .A(n35464), .B(n17259), .Z(n17222) );
  XOR U37666 ( .A(n35465), .B(n17247), .Z(n17259) );
  XNOR U37667 ( .A(q[6]), .B(DB[2610]), .Z(n17247) );
  IV U37668 ( .A(n17246), .Z(n35465) );
  XNOR U37669 ( .A(n17244), .B(n35466), .Z(n17246) );
  XNOR U37670 ( .A(q[5]), .B(DB[2609]), .Z(n35466) );
  XNOR U37671 ( .A(q[4]), .B(DB[2608]), .Z(n17244) );
  IV U37672 ( .A(n17258), .Z(n35464) );
  XOR U37673 ( .A(n35467), .B(n35468), .Z(n17258) );
  XNOR U37674 ( .A(n17254), .B(n17256), .Z(n35468) );
  XNOR U37675 ( .A(q[0]), .B(DB[2604]), .Z(n17256) );
  XNOR U37676 ( .A(q[3]), .B(DB[2607]), .Z(n17254) );
  IV U37677 ( .A(n17253), .Z(n35467) );
  XNOR U37678 ( .A(n17251), .B(n35469), .Z(n17253) );
  XNOR U37679 ( .A(q[2]), .B(DB[2606]), .Z(n35469) );
  XNOR U37680 ( .A(q[1]), .B(DB[2605]), .Z(n17251) );
  XOR U37681 ( .A(n35470), .B(n17216), .Z(n17179) );
  XOR U37682 ( .A(n35471), .B(n17204), .Z(n17216) );
  XNOR U37683 ( .A(q[6]), .B(DB[2617]), .Z(n17204) );
  IV U37684 ( .A(n17203), .Z(n35471) );
  XNOR U37685 ( .A(n17201), .B(n35472), .Z(n17203) );
  XNOR U37686 ( .A(q[5]), .B(DB[2616]), .Z(n35472) );
  XNOR U37687 ( .A(q[4]), .B(DB[2615]), .Z(n17201) );
  IV U37688 ( .A(n17215), .Z(n35470) );
  XOR U37689 ( .A(n35473), .B(n35474), .Z(n17215) );
  XNOR U37690 ( .A(n17211), .B(n17213), .Z(n35474) );
  XNOR U37691 ( .A(q[0]), .B(DB[2611]), .Z(n17213) );
  XNOR U37692 ( .A(q[3]), .B(DB[2614]), .Z(n17211) );
  IV U37693 ( .A(n17210), .Z(n35473) );
  XNOR U37694 ( .A(n17208), .B(n35475), .Z(n17210) );
  XNOR U37695 ( .A(q[2]), .B(DB[2613]), .Z(n35475) );
  XNOR U37696 ( .A(q[1]), .B(DB[2612]), .Z(n17208) );
  XOR U37697 ( .A(n35476), .B(n17173), .Z(n17136) );
  XOR U37698 ( .A(n35477), .B(n17161), .Z(n17173) );
  XNOR U37699 ( .A(q[6]), .B(DB[2624]), .Z(n17161) );
  IV U37700 ( .A(n17160), .Z(n35477) );
  XNOR U37701 ( .A(n17158), .B(n35478), .Z(n17160) );
  XNOR U37702 ( .A(q[5]), .B(DB[2623]), .Z(n35478) );
  XNOR U37703 ( .A(q[4]), .B(DB[2622]), .Z(n17158) );
  IV U37704 ( .A(n17172), .Z(n35476) );
  XOR U37705 ( .A(n35479), .B(n35480), .Z(n17172) );
  XNOR U37706 ( .A(n17168), .B(n17170), .Z(n35480) );
  XNOR U37707 ( .A(q[0]), .B(DB[2618]), .Z(n17170) );
  XNOR U37708 ( .A(q[3]), .B(DB[2621]), .Z(n17168) );
  IV U37709 ( .A(n17167), .Z(n35479) );
  XNOR U37710 ( .A(n17165), .B(n35481), .Z(n17167) );
  XNOR U37711 ( .A(q[2]), .B(DB[2620]), .Z(n35481) );
  XNOR U37712 ( .A(q[1]), .B(DB[2619]), .Z(n17165) );
  XOR U37713 ( .A(n35482), .B(n17130), .Z(n17093) );
  XOR U37714 ( .A(n35483), .B(n17118), .Z(n17130) );
  XNOR U37715 ( .A(q[6]), .B(DB[2631]), .Z(n17118) );
  IV U37716 ( .A(n17117), .Z(n35483) );
  XNOR U37717 ( .A(n17115), .B(n35484), .Z(n17117) );
  XNOR U37718 ( .A(q[5]), .B(DB[2630]), .Z(n35484) );
  XNOR U37719 ( .A(q[4]), .B(DB[2629]), .Z(n17115) );
  IV U37720 ( .A(n17129), .Z(n35482) );
  XOR U37721 ( .A(n35485), .B(n35486), .Z(n17129) );
  XNOR U37722 ( .A(n17125), .B(n17127), .Z(n35486) );
  XNOR U37723 ( .A(q[0]), .B(DB[2625]), .Z(n17127) );
  XNOR U37724 ( .A(q[3]), .B(DB[2628]), .Z(n17125) );
  IV U37725 ( .A(n17124), .Z(n35485) );
  XNOR U37726 ( .A(n17122), .B(n35487), .Z(n17124) );
  XNOR U37727 ( .A(q[2]), .B(DB[2627]), .Z(n35487) );
  XNOR U37728 ( .A(q[1]), .B(DB[2626]), .Z(n17122) );
  XOR U37729 ( .A(n35488), .B(n17087), .Z(n17050) );
  XOR U37730 ( .A(n35489), .B(n17075), .Z(n17087) );
  XNOR U37731 ( .A(q[6]), .B(DB[2638]), .Z(n17075) );
  IV U37732 ( .A(n17074), .Z(n35489) );
  XNOR U37733 ( .A(n17072), .B(n35490), .Z(n17074) );
  XNOR U37734 ( .A(q[5]), .B(DB[2637]), .Z(n35490) );
  XNOR U37735 ( .A(q[4]), .B(DB[2636]), .Z(n17072) );
  IV U37736 ( .A(n17086), .Z(n35488) );
  XOR U37737 ( .A(n35491), .B(n35492), .Z(n17086) );
  XNOR U37738 ( .A(n17082), .B(n17084), .Z(n35492) );
  XNOR U37739 ( .A(q[0]), .B(DB[2632]), .Z(n17084) );
  XNOR U37740 ( .A(q[3]), .B(DB[2635]), .Z(n17082) );
  IV U37741 ( .A(n17081), .Z(n35491) );
  XNOR U37742 ( .A(n17079), .B(n35493), .Z(n17081) );
  XNOR U37743 ( .A(q[2]), .B(DB[2634]), .Z(n35493) );
  XNOR U37744 ( .A(q[1]), .B(DB[2633]), .Z(n17079) );
  XOR U37745 ( .A(n35494), .B(n17044), .Z(n17007) );
  XOR U37746 ( .A(n35495), .B(n17032), .Z(n17044) );
  XNOR U37747 ( .A(q[6]), .B(DB[2645]), .Z(n17032) );
  IV U37748 ( .A(n17031), .Z(n35495) );
  XNOR U37749 ( .A(n17029), .B(n35496), .Z(n17031) );
  XNOR U37750 ( .A(q[5]), .B(DB[2644]), .Z(n35496) );
  XNOR U37751 ( .A(q[4]), .B(DB[2643]), .Z(n17029) );
  IV U37752 ( .A(n17043), .Z(n35494) );
  XOR U37753 ( .A(n35497), .B(n35498), .Z(n17043) );
  XNOR U37754 ( .A(n17039), .B(n17041), .Z(n35498) );
  XNOR U37755 ( .A(q[0]), .B(DB[2639]), .Z(n17041) );
  XNOR U37756 ( .A(q[3]), .B(DB[2642]), .Z(n17039) );
  IV U37757 ( .A(n17038), .Z(n35497) );
  XNOR U37758 ( .A(n17036), .B(n35499), .Z(n17038) );
  XNOR U37759 ( .A(q[2]), .B(DB[2641]), .Z(n35499) );
  XNOR U37760 ( .A(q[1]), .B(DB[2640]), .Z(n17036) );
  XOR U37761 ( .A(n35500), .B(n17001), .Z(n16964) );
  XOR U37762 ( .A(n35501), .B(n16989), .Z(n17001) );
  XNOR U37763 ( .A(q[6]), .B(DB[2652]), .Z(n16989) );
  IV U37764 ( .A(n16988), .Z(n35501) );
  XNOR U37765 ( .A(n16986), .B(n35502), .Z(n16988) );
  XNOR U37766 ( .A(q[5]), .B(DB[2651]), .Z(n35502) );
  XNOR U37767 ( .A(q[4]), .B(DB[2650]), .Z(n16986) );
  IV U37768 ( .A(n17000), .Z(n35500) );
  XOR U37769 ( .A(n35503), .B(n35504), .Z(n17000) );
  XNOR U37770 ( .A(n16996), .B(n16998), .Z(n35504) );
  XNOR U37771 ( .A(q[0]), .B(DB[2646]), .Z(n16998) );
  XNOR U37772 ( .A(q[3]), .B(DB[2649]), .Z(n16996) );
  IV U37773 ( .A(n16995), .Z(n35503) );
  XNOR U37774 ( .A(n16993), .B(n35505), .Z(n16995) );
  XNOR U37775 ( .A(q[2]), .B(DB[2648]), .Z(n35505) );
  XNOR U37776 ( .A(q[1]), .B(DB[2647]), .Z(n16993) );
  XOR U37777 ( .A(n35506), .B(n16958), .Z(n16921) );
  XOR U37778 ( .A(n35507), .B(n16946), .Z(n16958) );
  XNOR U37779 ( .A(q[6]), .B(DB[2659]), .Z(n16946) );
  IV U37780 ( .A(n16945), .Z(n35507) );
  XNOR U37781 ( .A(n16943), .B(n35508), .Z(n16945) );
  XNOR U37782 ( .A(q[5]), .B(DB[2658]), .Z(n35508) );
  XNOR U37783 ( .A(q[4]), .B(DB[2657]), .Z(n16943) );
  IV U37784 ( .A(n16957), .Z(n35506) );
  XOR U37785 ( .A(n35509), .B(n35510), .Z(n16957) );
  XNOR U37786 ( .A(n16953), .B(n16955), .Z(n35510) );
  XNOR U37787 ( .A(q[0]), .B(DB[2653]), .Z(n16955) );
  XNOR U37788 ( .A(q[3]), .B(DB[2656]), .Z(n16953) );
  IV U37789 ( .A(n16952), .Z(n35509) );
  XNOR U37790 ( .A(n16950), .B(n35511), .Z(n16952) );
  XNOR U37791 ( .A(q[2]), .B(DB[2655]), .Z(n35511) );
  XNOR U37792 ( .A(q[1]), .B(DB[2654]), .Z(n16950) );
  XOR U37793 ( .A(n35512), .B(n16915), .Z(n16878) );
  XOR U37794 ( .A(n35513), .B(n16903), .Z(n16915) );
  XNOR U37795 ( .A(q[6]), .B(DB[2666]), .Z(n16903) );
  IV U37796 ( .A(n16902), .Z(n35513) );
  XNOR U37797 ( .A(n16900), .B(n35514), .Z(n16902) );
  XNOR U37798 ( .A(q[5]), .B(DB[2665]), .Z(n35514) );
  XNOR U37799 ( .A(q[4]), .B(DB[2664]), .Z(n16900) );
  IV U37800 ( .A(n16914), .Z(n35512) );
  XOR U37801 ( .A(n35515), .B(n35516), .Z(n16914) );
  XNOR U37802 ( .A(n16910), .B(n16912), .Z(n35516) );
  XNOR U37803 ( .A(q[0]), .B(DB[2660]), .Z(n16912) );
  XNOR U37804 ( .A(q[3]), .B(DB[2663]), .Z(n16910) );
  IV U37805 ( .A(n16909), .Z(n35515) );
  XNOR U37806 ( .A(n16907), .B(n35517), .Z(n16909) );
  XNOR U37807 ( .A(q[2]), .B(DB[2662]), .Z(n35517) );
  XNOR U37808 ( .A(q[1]), .B(DB[2661]), .Z(n16907) );
  XOR U37809 ( .A(n35518), .B(n16872), .Z(n16835) );
  XOR U37810 ( .A(n35519), .B(n16860), .Z(n16872) );
  XNOR U37811 ( .A(q[6]), .B(DB[2673]), .Z(n16860) );
  IV U37812 ( .A(n16859), .Z(n35519) );
  XNOR U37813 ( .A(n16857), .B(n35520), .Z(n16859) );
  XNOR U37814 ( .A(q[5]), .B(DB[2672]), .Z(n35520) );
  XNOR U37815 ( .A(q[4]), .B(DB[2671]), .Z(n16857) );
  IV U37816 ( .A(n16871), .Z(n35518) );
  XOR U37817 ( .A(n35521), .B(n35522), .Z(n16871) );
  XNOR U37818 ( .A(n16867), .B(n16869), .Z(n35522) );
  XNOR U37819 ( .A(q[0]), .B(DB[2667]), .Z(n16869) );
  XNOR U37820 ( .A(q[3]), .B(DB[2670]), .Z(n16867) );
  IV U37821 ( .A(n16866), .Z(n35521) );
  XNOR U37822 ( .A(n16864), .B(n35523), .Z(n16866) );
  XNOR U37823 ( .A(q[2]), .B(DB[2669]), .Z(n35523) );
  XNOR U37824 ( .A(q[1]), .B(DB[2668]), .Z(n16864) );
  XOR U37825 ( .A(n35524), .B(n16829), .Z(n16792) );
  XOR U37826 ( .A(n35525), .B(n16817), .Z(n16829) );
  XNOR U37827 ( .A(q[6]), .B(DB[2680]), .Z(n16817) );
  IV U37828 ( .A(n16816), .Z(n35525) );
  XNOR U37829 ( .A(n16814), .B(n35526), .Z(n16816) );
  XNOR U37830 ( .A(q[5]), .B(DB[2679]), .Z(n35526) );
  XNOR U37831 ( .A(q[4]), .B(DB[2678]), .Z(n16814) );
  IV U37832 ( .A(n16828), .Z(n35524) );
  XOR U37833 ( .A(n35527), .B(n35528), .Z(n16828) );
  XNOR U37834 ( .A(n16824), .B(n16826), .Z(n35528) );
  XNOR U37835 ( .A(q[0]), .B(DB[2674]), .Z(n16826) );
  XNOR U37836 ( .A(q[3]), .B(DB[2677]), .Z(n16824) );
  IV U37837 ( .A(n16823), .Z(n35527) );
  XNOR U37838 ( .A(n16821), .B(n35529), .Z(n16823) );
  XNOR U37839 ( .A(q[2]), .B(DB[2676]), .Z(n35529) );
  XNOR U37840 ( .A(q[1]), .B(DB[2675]), .Z(n16821) );
  XOR U37841 ( .A(n35530), .B(n16786), .Z(n16749) );
  XOR U37842 ( .A(n35531), .B(n16774), .Z(n16786) );
  XNOR U37843 ( .A(q[6]), .B(DB[2687]), .Z(n16774) );
  IV U37844 ( .A(n16773), .Z(n35531) );
  XNOR U37845 ( .A(n16771), .B(n35532), .Z(n16773) );
  XNOR U37846 ( .A(q[5]), .B(DB[2686]), .Z(n35532) );
  XNOR U37847 ( .A(q[4]), .B(DB[2685]), .Z(n16771) );
  IV U37848 ( .A(n16785), .Z(n35530) );
  XOR U37849 ( .A(n35533), .B(n35534), .Z(n16785) );
  XNOR U37850 ( .A(n16781), .B(n16783), .Z(n35534) );
  XNOR U37851 ( .A(q[0]), .B(DB[2681]), .Z(n16783) );
  XNOR U37852 ( .A(q[3]), .B(DB[2684]), .Z(n16781) );
  IV U37853 ( .A(n16780), .Z(n35533) );
  XNOR U37854 ( .A(n16778), .B(n35535), .Z(n16780) );
  XNOR U37855 ( .A(q[2]), .B(DB[2683]), .Z(n35535) );
  XNOR U37856 ( .A(q[1]), .B(DB[2682]), .Z(n16778) );
  XOR U37857 ( .A(n35536), .B(n16743), .Z(n16706) );
  XOR U37858 ( .A(n35537), .B(n16731), .Z(n16743) );
  XNOR U37859 ( .A(q[6]), .B(DB[2694]), .Z(n16731) );
  IV U37860 ( .A(n16730), .Z(n35537) );
  XNOR U37861 ( .A(n16728), .B(n35538), .Z(n16730) );
  XNOR U37862 ( .A(q[5]), .B(DB[2693]), .Z(n35538) );
  XNOR U37863 ( .A(q[4]), .B(DB[2692]), .Z(n16728) );
  IV U37864 ( .A(n16742), .Z(n35536) );
  XOR U37865 ( .A(n35539), .B(n35540), .Z(n16742) );
  XNOR U37866 ( .A(n16738), .B(n16740), .Z(n35540) );
  XNOR U37867 ( .A(q[0]), .B(DB[2688]), .Z(n16740) );
  XNOR U37868 ( .A(q[3]), .B(DB[2691]), .Z(n16738) );
  IV U37869 ( .A(n16737), .Z(n35539) );
  XNOR U37870 ( .A(n16735), .B(n35541), .Z(n16737) );
  XNOR U37871 ( .A(q[2]), .B(DB[2690]), .Z(n35541) );
  XNOR U37872 ( .A(q[1]), .B(DB[2689]), .Z(n16735) );
  XOR U37873 ( .A(n35542), .B(n16700), .Z(n16663) );
  XOR U37874 ( .A(n35543), .B(n16688), .Z(n16700) );
  XNOR U37875 ( .A(q[6]), .B(DB[2701]), .Z(n16688) );
  IV U37876 ( .A(n16687), .Z(n35543) );
  XNOR U37877 ( .A(n16685), .B(n35544), .Z(n16687) );
  XNOR U37878 ( .A(q[5]), .B(DB[2700]), .Z(n35544) );
  XNOR U37879 ( .A(q[4]), .B(DB[2699]), .Z(n16685) );
  IV U37880 ( .A(n16699), .Z(n35542) );
  XOR U37881 ( .A(n35545), .B(n35546), .Z(n16699) );
  XNOR U37882 ( .A(n16695), .B(n16697), .Z(n35546) );
  XNOR U37883 ( .A(q[0]), .B(DB[2695]), .Z(n16697) );
  XNOR U37884 ( .A(q[3]), .B(DB[2698]), .Z(n16695) );
  IV U37885 ( .A(n16694), .Z(n35545) );
  XNOR U37886 ( .A(n16692), .B(n35547), .Z(n16694) );
  XNOR U37887 ( .A(q[2]), .B(DB[2697]), .Z(n35547) );
  XNOR U37888 ( .A(q[1]), .B(DB[2696]), .Z(n16692) );
  XOR U37889 ( .A(n35548), .B(n16657), .Z(n16620) );
  XOR U37890 ( .A(n35549), .B(n16645), .Z(n16657) );
  XNOR U37891 ( .A(q[6]), .B(DB[2708]), .Z(n16645) );
  IV U37892 ( .A(n16644), .Z(n35549) );
  XNOR U37893 ( .A(n16642), .B(n35550), .Z(n16644) );
  XNOR U37894 ( .A(q[5]), .B(DB[2707]), .Z(n35550) );
  XNOR U37895 ( .A(q[4]), .B(DB[2706]), .Z(n16642) );
  IV U37896 ( .A(n16656), .Z(n35548) );
  XOR U37897 ( .A(n35551), .B(n35552), .Z(n16656) );
  XNOR U37898 ( .A(n16652), .B(n16654), .Z(n35552) );
  XNOR U37899 ( .A(q[0]), .B(DB[2702]), .Z(n16654) );
  XNOR U37900 ( .A(q[3]), .B(DB[2705]), .Z(n16652) );
  IV U37901 ( .A(n16651), .Z(n35551) );
  XNOR U37902 ( .A(n16649), .B(n35553), .Z(n16651) );
  XNOR U37903 ( .A(q[2]), .B(DB[2704]), .Z(n35553) );
  XNOR U37904 ( .A(q[1]), .B(DB[2703]), .Z(n16649) );
  XOR U37905 ( .A(n35554), .B(n16614), .Z(n16577) );
  XOR U37906 ( .A(n35555), .B(n16602), .Z(n16614) );
  XNOR U37907 ( .A(q[6]), .B(DB[2715]), .Z(n16602) );
  IV U37908 ( .A(n16601), .Z(n35555) );
  XNOR U37909 ( .A(n16599), .B(n35556), .Z(n16601) );
  XNOR U37910 ( .A(q[5]), .B(DB[2714]), .Z(n35556) );
  XNOR U37911 ( .A(q[4]), .B(DB[2713]), .Z(n16599) );
  IV U37912 ( .A(n16613), .Z(n35554) );
  XOR U37913 ( .A(n35557), .B(n35558), .Z(n16613) );
  XNOR U37914 ( .A(n16609), .B(n16611), .Z(n35558) );
  XNOR U37915 ( .A(q[0]), .B(DB[2709]), .Z(n16611) );
  XNOR U37916 ( .A(q[3]), .B(DB[2712]), .Z(n16609) );
  IV U37917 ( .A(n16608), .Z(n35557) );
  XNOR U37918 ( .A(n16606), .B(n35559), .Z(n16608) );
  XNOR U37919 ( .A(q[2]), .B(DB[2711]), .Z(n35559) );
  XNOR U37920 ( .A(q[1]), .B(DB[2710]), .Z(n16606) );
  XOR U37921 ( .A(n35560), .B(n16571), .Z(n16534) );
  XOR U37922 ( .A(n35561), .B(n16559), .Z(n16571) );
  XNOR U37923 ( .A(q[6]), .B(DB[2722]), .Z(n16559) );
  IV U37924 ( .A(n16558), .Z(n35561) );
  XNOR U37925 ( .A(n16556), .B(n35562), .Z(n16558) );
  XNOR U37926 ( .A(q[5]), .B(DB[2721]), .Z(n35562) );
  XNOR U37927 ( .A(q[4]), .B(DB[2720]), .Z(n16556) );
  IV U37928 ( .A(n16570), .Z(n35560) );
  XOR U37929 ( .A(n35563), .B(n35564), .Z(n16570) );
  XNOR U37930 ( .A(n16566), .B(n16568), .Z(n35564) );
  XNOR U37931 ( .A(q[0]), .B(DB[2716]), .Z(n16568) );
  XNOR U37932 ( .A(q[3]), .B(DB[2719]), .Z(n16566) );
  IV U37933 ( .A(n16565), .Z(n35563) );
  XNOR U37934 ( .A(n16563), .B(n35565), .Z(n16565) );
  XNOR U37935 ( .A(q[2]), .B(DB[2718]), .Z(n35565) );
  XNOR U37936 ( .A(q[1]), .B(DB[2717]), .Z(n16563) );
  XOR U37937 ( .A(n35566), .B(n16528), .Z(n16491) );
  XOR U37938 ( .A(n35567), .B(n16516), .Z(n16528) );
  XNOR U37939 ( .A(q[6]), .B(DB[2729]), .Z(n16516) );
  IV U37940 ( .A(n16515), .Z(n35567) );
  XNOR U37941 ( .A(n16513), .B(n35568), .Z(n16515) );
  XNOR U37942 ( .A(q[5]), .B(DB[2728]), .Z(n35568) );
  XNOR U37943 ( .A(q[4]), .B(DB[2727]), .Z(n16513) );
  IV U37944 ( .A(n16527), .Z(n35566) );
  XOR U37945 ( .A(n35569), .B(n35570), .Z(n16527) );
  XNOR U37946 ( .A(n16523), .B(n16525), .Z(n35570) );
  XNOR U37947 ( .A(q[0]), .B(DB[2723]), .Z(n16525) );
  XNOR U37948 ( .A(q[3]), .B(DB[2726]), .Z(n16523) );
  IV U37949 ( .A(n16522), .Z(n35569) );
  XNOR U37950 ( .A(n16520), .B(n35571), .Z(n16522) );
  XNOR U37951 ( .A(q[2]), .B(DB[2725]), .Z(n35571) );
  XNOR U37952 ( .A(q[1]), .B(DB[2724]), .Z(n16520) );
  XOR U37953 ( .A(n35572), .B(n16485), .Z(n16448) );
  XOR U37954 ( .A(n35573), .B(n16473), .Z(n16485) );
  XNOR U37955 ( .A(q[6]), .B(DB[2736]), .Z(n16473) );
  IV U37956 ( .A(n16472), .Z(n35573) );
  XNOR U37957 ( .A(n16470), .B(n35574), .Z(n16472) );
  XNOR U37958 ( .A(q[5]), .B(DB[2735]), .Z(n35574) );
  XNOR U37959 ( .A(q[4]), .B(DB[2734]), .Z(n16470) );
  IV U37960 ( .A(n16484), .Z(n35572) );
  XOR U37961 ( .A(n35575), .B(n35576), .Z(n16484) );
  XNOR U37962 ( .A(n16480), .B(n16482), .Z(n35576) );
  XNOR U37963 ( .A(q[0]), .B(DB[2730]), .Z(n16482) );
  XNOR U37964 ( .A(q[3]), .B(DB[2733]), .Z(n16480) );
  IV U37965 ( .A(n16479), .Z(n35575) );
  XNOR U37966 ( .A(n16477), .B(n35577), .Z(n16479) );
  XNOR U37967 ( .A(q[2]), .B(DB[2732]), .Z(n35577) );
  XNOR U37968 ( .A(q[1]), .B(DB[2731]), .Z(n16477) );
  XOR U37969 ( .A(n35578), .B(n16442), .Z(n16405) );
  XOR U37970 ( .A(n35579), .B(n16430), .Z(n16442) );
  XNOR U37971 ( .A(q[6]), .B(DB[2743]), .Z(n16430) );
  IV U37972 ( .A(n16429), .Z(n35579) );
  XNOR U37973 ( .A(n16427), .B(n35580), .Z(n16429) );
  XNOR U37974 ( .A(q[5]), .B(DB[2742]), .Z(n35580) );
  XNOR U37975 ( .A(q[4]), .B(DB[2741]), .Z(n16427) );
  IV U37976 ( .A(n16441), .Z(n35578) );
  XOR U37977 ( .A(n35581), .B(n35582), .Z(n16441) );
  XNOR U37978 ( .A(n16437), .B(n16439), .Z(n35582) );
  XNOR U37979 ( .A(q[0]), .B(DB[2737]), .Z(n16439) );
  XNOR U37980 ( .A(q[3]), .B(DB[2740]), .Z(n16437) );
  IV U37981 ( .A(n16436), .Z(n35581) );
  XNOR U37982 ( .A(n16434), .B(n35583), .Z(n16436) );
  XNOR U37983 ( .A(q[2]), .B(DB[2739]), .Z(n35583) );
  XNOR U37984 ( .A(q[1]), .B(DB[2738]), .Z(n16434) );
  XOR U37985 ( .A(n35584), .B(n16399), .Z(n16362) );
  XOR U37986 ( .A(n35585), .B(n16387), .Z(n16399) );
  XNOR U37987 ( .A(q[6]), .B(DB[2750]), .Z(n16387) );
  IV U37988 ( .A(n16386), .Z(n35585) );
  XNOR U37989 ( .A(n16384), .B(n35586), .Z(n16386) );
  XNOR U37990 ( .A(q[5]), .B(DB[2749]), .Z(n35586) );
  XNOR U37991 ( .A(q[4]), .B(DB[2748]), .Z(n16384) );
  IV U37992 ( .A(n16398), .Z(n35584) );
  XOR U37993 ( .A(n35587), .B(n35588), .Z(n16398) );
  XNOR U37994 ( .A(n16394), .B(n16396), .Z(n35588) );
  XNOR U37995 ( .A(q[0]), .B(DB[2744]), .Z(n16396) );
  XNOR U37996 ( .A(q[3]), .B(DB[2747]), .Z(n16394) );
  IV U37997 ( .A(n16393), .Z(n35587) );
  XNOR U37998 ( .A(n16391), .B(n35589), .Z(n16393) );
  XNOR U37999 ( .A(q[2]), .B(DB[2746]), .Z(n35589) );
  XNOR U38000 ( .A(q[1]), .B(DB[2745]), .Z(n16391) );
  XOR U38001 ( .A(n35590), .B(n16356), .Z(n16319) );
  XOR U38002 ( .A(n35591), .B(n16344), .Z(n16356) );
  XNOR U38003 ( .A(q[6]), .B(DB[2757]), .Z(n16344) );
  IV U38004 ( .A(n16343), .Z(n35591) );
  XNOR U38005 ( .A(n16341), .B(n35592), .Z(n16343) );
  XNOR U38006 ( .A(q[5]), .B(DB[2756]), .Z(n35592) );
  XNOR U38007 ( .A(q[4]), .B(DB[2755]), .Z(n16341) );
  IV U38008 ( .A(n16355), .Z(n35590) );
  XOR U38009 ( .A(n35593), .B(n35594), .Z(n16355) );
  XNOR U38010 ( .A(n16351), .B(n16353), .Z(n35594) );
  XNOR U38011 ( .A(q[0]), .B(DB[2751]), .Z(n16353) );
  XNOR U38012 ( .A(q[3]), .B(DB[2754]), .Z(n16351) );
  IV U38013 ( .A(n16350), .Z(n35593) );
  XNOR U38014 ( .A(n16348), .B(n35595), .Z(n16350) );
  XNOR U38015 ( .A(q[2]), .B(DB[2753]), .Z(n35595) );
  XNOR U38016 ( .A(q[1]), .B(DB[2752]), .Z(n16348) );
  XOR U38017 ( .A(n35596), .B(n16313), .Z(n16276) );
  XOR U38018 ( .A(n35597), .B(n16301), .Z(n16313) );
  XNOR U38019 ( .A(q[6]), .B(DB[2764]), .Z(n16301) );
  IV U38020 ( .A(n16300), .Z(n35597) );
  XNOR U38021 ( .A(n16298), .B(n35598), .Z(n16300) );
  XNOR U38022 ( .A(q[5]), .B(DB[2763]), .Z(n35598) );
  XNOR U38023 ( .A(q[4]), .B(DB[2762]), .Z(n16298) );
  IV U38024 ( .A(n16312), .Z(n35596) );
  XOR U38025 ( .A(n35599), .B(n35600), .Z(n16312) );
  XNOR U38026 ( .A(n16308), .B(n16310), .Z(n35600) );
  XNOR U38027 ( .A(q[0]), .B(DB[2758]), .Z(n16310) );
  XNOR U38028 ( .A(q[3]), .B(DB[2761]), .Z(n16308) );
  IV U38029 ( .A(n16307), .Z(n35599) );
  XNOR U38030 ( .A(n16305), .B(n35601), .Z(n16307) );
  XNOR U38031 ( .A(q[2]), .B(DB[2760]), .Z(n35601) );
  XNOR U38032 ( .A(q[1]), .B(DB[2759]), .Z(n16305) );
  XOR U38033 ( .A(n35602), .B(n16270), .Z(n16233) );
  XOR U38034 ( .A(n35603), .B(n16258), .Z(n16270) );
  XNOR U38035 ( .A(q[6]), .B(DB[2771]), .Z(n16258) );
  IV U38036 ( .A(n16257), .Z(n35603) );
  XNOR U38037 ( .A(n16255), .B(n35604), .Z(n16257) );
  XNOR U38038 ( .A(q[5]), .B(DB[2770]), .Z(n35604) );
  XNOR U38039 ( .A(q[4]), .B(DB[2769]), .Z(n16255) );
  IV U38040 ( .A(n16269), .Z(n35602) );
  XOR U38041 ( .A(n35605), .B(n35606), .Z(n16269) );
  XNOR U38042 ( .A(n16265), .B(n16267), .Z(n35606) );
  XNOR U38043 ( .A(q[0]), .B(DB[2765]), .Z(n16267) );
  XNOR U38044 ( .A(q[3]), .B(DB[2768]), .Z(n16265) );
  IV U38045 ( .A(n16264), .Z(n35605) );
  XNOR U38046 ( .A(n16262), .B(n35607), .Z(n16264) );
  XNOR U38047 ( .A(q[2]), .B(DB[2767]), .Z(n35607) );
  XNOR U38048 ( .A(q[1]), .B(DB[2766]), .Z(n16262) );
  XOR U38049 ( .A(n35608), .B(n16227), .Z(n16190) );
  XOR U38050 ( .A(n35609), .B(n16215), .Z(n16227) );
  XNOR U38051 ( .A(q[6]), .B(DB[2778]), .Z(n16215) );
  IV U38052 ( .A(n16214), .Z(n35609) );
  XNOR U38053 ( .A(n16212), .B(n35610), .Z(n16214) );
  XNOR U38054 ( .A(q[5]), .B(DB[2777]), .Z(n35610) );
  XNOR U38055 ( .A(q[4]), .B(DB[2776]), .Z(n16212) );
  IV U38056 ( .A(n16226), .Z(n35608) );
  XOR U38057 ( .A(n35611), .B(n35612), .Z(n16226) );
  XNOR U38058 ( .A(n16222), .B(n16224), .Z(n35612) );
  XNOR U38059 ( .A(q[0]), .B(DB[2772]), .Z(n16224) );
  XNOR U38060 ( .A(q[3]), .B(DB[2775]), .Z(n16222) );
  IV U38061 ( .A(n16221), .Z(n35611) );
  XNOR U38062 ( .A(n16219), .B(n35613), .Z(n16221) );
  XNOR U38063 ( .A(q[2]), .B(DB[2774]), .Z(n35613) );
  XNOR U38064 ( .A(q[1]), .B(DB[2773]), .Z(n16219) );
  XOR U38065 ( .A(n35614), .B(n16184), .Z(n16147) );
  XOR U38066 ( .A(n35615), .B(n16172), .Z(n16184) );
  XNOR U38067 ( .A(q[6]), .B(DB[2785]), .Z(n16172) );
  IV U38068 ( .A(n16171), .Z(n35615) );
  XNOR U38069 ( .A(n16169), .B(n35616), .Z(n16171) );
  XNOR U38070 ( .A(q[5]), .B(DB[2784]), .Z(n35616) );
  XNOR U38071 ( .A(q[4]), .B(DB[2783]), .Z(n16169) );
  IV U38072 ( .A(n16183), .Z(n35614) );
  XOR U38073 ( .A(n35617), .B(n35618), .Z(n16183) );
  XNOR U38074 ( .A(n16179), .B(n16181), .Z(n35618) );
  XNOR U38075 ( .A(q[0]), .B(DB[2779]), .Z(n16181) );
  XNOR U38076 ( .A(q[3]), .B(DB[2782]), .Z(n16179) );
  IV U38077 ( .A(n16178), .Z(n35617) );
  XNOR U38078 ( .A(n16176), .B(n35619), .Z(n16178) );
  XNOR U38079 ( .A(q[2]), .B(DB[2781]), .Z(n35619) );
  XNOR U38080 ( .A(q[1]), .B(DB[2780]), .Z(n16176) );
  XOR U38081 ( .A(n35620), .B(n16141), .Z(n16104) );
  XOR U38082 ( .A(n35621), .B(n16129), .Z(n16141) );
  XNOR U38083 ( .A(q[6]), .B(DB[2792]), .Z(n16129) );
  IV U38084 ( .A(n16128), .Z(n35621) );
  XNOR U38085 ( .A(n16126), .B(n35622), .Z(n16128) );
  XNOR U38086 ( .A(q[5]), .B(DB[2791]), .Z(n35622) );
  XNOR U38087 ( .A(q[4]), .B(DB[2790]), .Z(n16126) );
  IV U38088 ( .A(n16140), .Z(n35620) );
  XOR U38089 ( .A(n35623), .B(n35624), .Z(n16140) );
  XNOR U38090 ( .A(n16136), .B(n16138), .Z(n35624) );
  XNOR U38091 ( .A(q[0]), .B(DB[2786]), .Z(n16138) );
  XNOR U38092 ( .A(q[3]), .B(DB[2789]), .Z(n16136) );
  IV U38093 ( .A(n16135), .Z(n35623) );
  XNOR U38094 ( .A(n16133), .B(n35625), .Z(n16135) );
  XNOR U38095 ( .A(q[2]), .B(DB[2788]), .Z(n35625) );
  XNOR U38096 ( .A(q[1]), .B(DB[2787]), .Z(n16133) );
  XOR U38097 ( .A(n35626), .B(n16098), .Z(n16061) );
  XOR U38098 ( .A(n35627), .B(n16086), .Z(n16098) );
  XNOR U38099 ( .A(q[6]), .B(DB[2799]), .Z(n16086) );
  IV U38100 ( .A(n16085), .Z(n35627) );
  XNOR U38101 ( .A(n16083), .B(n35628), .Z(n16085) );
  XNOR U38102 ( .A(q[5]), .B(DB[2798]), .Z(n35628) );
  XNOR U38103 ( .A(q[4]), .B(DB[2797]), .Z(n16083) );
  IV U38104 ( .A(n16097), .Z(n35626) );
  XOR U38105 ( .A(n35629), .B(n35630), .Z(n16097) );
  XNOR U38106 ( .A(n16093), .B(n16095), .Z(n35630) );
  XNOR U38107 ( .A(q[0]), .B(DB[2793]), .Z(n16095) );
  XNOR U38108 ( .A(q[3]), .B(DB[2796]), .Z(n16093) );
  IV U38109 ( .A(n16092), .Z(n35629) );
  XNOR U38110 ( .A(n16090), .B(n35631), .Z(n16092) );
  XNOR U38111 ( .A(q[2]), .B(DB[2795]), .Z(n35631) );
  XNOR U38112 ( .A(q[1]), .B(DB[2794]), .Z(n16090) );
  XOR U38113 ( .A(n35632), .B(n16055), .Z(n16018) );
  XOR U38114 ( .A(n35633), .B(n16043), .Z(n16055) );
  XNOR U38115 ( .A(q[6]), .B(DB[2806]), .Z(n16043) );
  IV U38116 ( .A(n16042), .Z(n35633) );
  XNOR U38117 ( .A(n16040), .B(n35634), .Z(n16042) );
  XNOR U38118 ( .A(q[5]), .B(DB[2805]), .Z(n35634) );
  XNOR U38119 ( .A(q[4]), .B(DB[2804]), .Z(n16040) );
  IV U38120 ( .A(n16054), .Z(n35632) );
  XOR U38121 ( .A(n35635), .B(n35636), .Z(n16054) );
  XNOR U38122 ( .A(n16050), .B(n16052), .Z(n35636) );
  XNOR U38123 ( .A(q[0]), .B(DB[2800]), .Z(n16052) );
  XNOR U38124 ( .A(q[3]), .B(DB[2803]), .Z(n16050) );
  IV U38125 ( .A(n16049), .Z(n35635) );
  XNOR U38126 ( .A(n16047), .B(n35637), .Z(n16049) );
  XNOR U38127 ( .A(q[2]), .B(DB[2802]), .Z(n35637) );
  XNOR U38128 ( .A(q[1]), .B(DB[2801]), .Z(n16047) );
  XOR U38129 ( .A(n35638), .B(n16012), .Z(n15975) );
  XOR U38130 ( .A(n35639), .B(n16000), .Z(n16012) );
  XNOR U38131 ( .A(q[6]), .B(DB[2813]), .Z(n16000) );
  IV U38132 ( .A(n15999), .Z(n35639) );
  XNOR U38133 ( .A(n15997), .B(n35640), .Z(n15999) );
  XNOR U38134 ( .A(q[5]), .B(DB[2812]), .Z(n35640) );
  XNOR U38135 ( .A(q[4]), .B(DB[2811]), .Z(n15997) );
  IV U38136 ( .A(n16011), .Z(n35638) );
  XOR U38137 ( .A(n35641), .B(n35642), .Z(n16011) );
  XNOR U38138 ( .A(n16007), .B(n16009), .Z(n35642) );
  XNOR U38139 ( .A(q[0]), .B(DB[2807]), .Z(n16009) );
  XNOR U38140 ( .A(q[3]), .B(DB[2810]), .Z(n16007) );
  IV U38141 ( .A(n16006), .Z(n35641) );
  XNOR U38142 ( .A(n16004), .B(n35643), .Z(n16006) );
  XNOR U38143 ( .A(q[2]), .B(DB[2809]), .Z(n35643) );
  XNOR U38144 ( .A(q[1]), .B(DB[2808]), .Z(n16004) );
  XOR U38145 ( .A(n35644), .B(n15969), .Z(n15932) );
  XOR U38146 ( .A(n35645), .B(n15957), .Z(n15969) );
  XNOR U38147 ( .A(q[6]), .B(DB[2820]), .Z(n15957) );
  IV U38148 ( .A(n15956), .Z(n35645) );
  XNOR U38149 ( .A(n15954), .B(n35646), .Z(n15956) );
  XNOR U38150 ( .A(q[5]), .B(DB[2819]), .Z(n35646) );
  XNOR U38151 ( .A(q[4]), .B(DB[2818]), .Z(n15954) );
  IV U38152 ( .A(n15968), .Z(n35644) );
  XOR U38153 ( .A(n35647), .B(n35648), .Z(n15968) );
  XNOR U38154 ( .A(n15964), .B(n15966), .Z(n35648) );
  XNOR U38155 ( .A(q[0]), .B(DB[2814]), .Z(n15966) );
  XNOR U38156 ( .A(q[3]), .B(DB[2817]), .Z(n15964) );
  IV U38157 ( .A(n15963), .Z(n35647) );
  XNOR U38158 ( .A(n15961), .B(n35649), .Z(n15963) );
  XNOR U38159 ( .A(q[2]), .B(DB[2816]), .Z(n35649) );
  XNOR U38160 ( .A(q[1]), .B(DB[2815]), .Z(n15961) );
  XOR U38161 ( .A(n35650), .B(n15926), .Z(n15889) );
  XOR U38162 ( .A(n35651), .B(n15914), .Z(n15926) );
  XNOR U38163 ( .A(q[6]), .B(DB[2827]), .Z(n15914) );
  IV U38164 ( .A(n15913), .Z(n35651) );
  XNOR U38165 ( .A(n15911), .B(n35652), .Z(n15913) );
  XNOR U38166 ( .A(q[5]), .B(DB[2826]), .Z(n35652) );
  XNOR U38167 ( .A(q[4]), .B(DB[2825]), .Z(n15911) );
  IV U38168 ( .A(n15925), .Z(n35650) );
  XOR U38169 ( .A(n35653), .B(n35654), .Z(n15925) );
  XNOR U38170 ( .A(n15921), .B(n15923), .Z(n35654) );
  XNOR U38171 ( .A(q[0]), .B(DB[2821]), .Z(n15923) );
  XNOR U38172 ( .A(q[3]), .B(DB[2824]), .Z(n15921) );
  IV U38173 ( .A(n15920), .Z(n35653) );
  XNOR U38174 ( .A(n15918), .B(n35655), .Z(n15920) );
  XNOR U38175 ( .A(q[2]), .B(DB[2823]), .Z(n35655) );
  XNOR U38176 ( .A(q[1]), .B(DB[2822]), .Z(n15918) );
  XOR U38177 ( .A(n35656), .B(n15883), .Z(n15846) );
  XOR U38178 ( .A(n35657), .B(n15871), .Z(n15883) );
  XNOR U38179 ( .A(q[6]), .B(DB[2834]), .Z(n15871) );
  IV U38180 ( .A(n15870), .Z(n35657) );
  XNOR U38181 ( .A(n15868), .B(n35658), .Z(n15870) );
  XNOR U38182 ( .A(q[5]), .B(DB[2833]), .Z(n35658) );
  XNOR U38183 ( .A(q[4]), .B(DB[2832]), .Z(n15868) );
  IV U38184 ( .A(n15882), .Z(n35656) );
  XOR U38185 ( .A(n35659), .B(n35660), .Z(n15882) );
  XNOR U38186 ( .A(n15878), .B(n15880), .Z(n35660) );
  XNOR U38187 ( .A(q[0]), .B(DB[2828]), .Z(n15880) );
  XNOR U38188 ( .A(q[3]), .B(DB[2831]), .Z(n15878) );
  IV U38189 ( .A(n15877), .Z(n35659) );
  XNOR U38190 ( .A(n15875), .B(n35661), .Z(n15877) );
  XNOR U38191 ( .A(q[2]), .B(DB[2830]), .Z(n35661) );
  XNOR U38192 ( .A(q[1]), .B(DB[2829]), .Z(n15875) );
  XOR U38193 ( .A(n35662), .B(n15840), .Z(n15803) );
  XOR U38194 ( .A(n35663), .B(n15828), .Z(n15840) );
  XNOR U38195 ( .A(q[6]), .B(DB[2841]), .Z(n15828) );
  IV U38196 ( .A(n15827), .Z(n35663) );
  XNOR U38197 ( .A(n15825), .B(n35664), .Z(n15827) );
  XNOR U38198 ( .A(q[5]), .B(DB[2840]), .Z(n35664) );
  XNOR U38199 ( .A(q[4]), .B(DB[2839]), .Z(n15825) );
  IV U38200 ( .A(n15839), .Z(n35662) );
  XOR U38201 ( .A(n35665), .B(n35666), .Z(n15839) );
  XNOR U38202 ( .A(n15835), .B(n15837), .Z(n35666) );
  XNOR U38203 ( .A(q[0]), .B(DB[2835]), .Z(n15837) );
  XNOR U38204 ( .A(q[3]), .B(DB[2838]), .Z(n15835) );
  IV U38205 ( .A(n15834), .Z(n35665) );
  XNOR U38206 ( .A(n15832), .B(n35667), .Z(n15834) );
  XNOR U38207 ( .A(q[2]), .B(DB[2837]), .Z(n35667) );
  XNOR U38208 ( .A(q[1]), .B(DB[2836]), .Z(n15832) );
  XOR U38209 ( .A(n35668), .B(n15797), .Z(n15760) );
  XOR U38210 ( .A(n35669), .B(n15785), .Z(n15797) );
  XNOR U38211 ( .A(q[6]), .B(DB[2848]), .Z(n15785) );
  IV U38212 ( .A(n15784), .Z(n35669) );
  XNOR U38213 ( .A(n15782), .B(n35670), .Z(n15784) );
  XNOR U38214 ( .A(q[5]), .B(DB[2847]), .Z(n35670) );
  XNOR U38215 ( .A(q[4]), .B(DB[2846]), .Z(n15782) );
  IV U38216 ( .A(n15796), .Z(n35668) );
  XOR U38217 ( .A(n35671), .B(n35672), .Z(n15796) );
  XNOR U38218 ( .A(n15792), .B(n15794), .Z(n35672) );
  XNOR U38219 ( .A(q[0]), .B(DB[2842]), .Z(n15794) );
  XNOR U38220 ( .A(q[3]), .B(DB[2845]), .Z(n15792) );
  IV U38221 ( .A(n15791), .Z(n35671) );
  XNOR U38222 ( .A(n15789), .B(n35673), .Z(n15791) );
  XNOR U38223 ( .A(q[2]), .B(DB[2844]), .Z(n35673) );
  XNOR U38224 ( .A(q[1]), .B(DB[2843]), .Z(n15789) );
  XOR U38225 ( .A(n35674), .B(n15754), .Z(n15717) );
  XOR U38226 ( .A(n35675), .B(n15742), .Z(n15754) );
  XNOR U38227 ( .A(q[6]), .B(DB[2855]), .Z(n15742) );
  IV U38228 ( .A(n15741), .Z(n35675) );
  XNOR U38229 ( .A(n15739), .B(n35676), .Z(n15741) );
  XNOR U38230 ( .A(q[5]), .B(DB[2854]), .Z(n35676) );
  XNOR U38231 ( .A(q[4]), .B(DB[2853]), .Z(n15739) );
  IV U38232 ( .A(n15753), .Z(n35674) );
  XOR U38233 ( .A(n35677), .B(n35678), .Z(n15753) );
  XNOR U38234 ( .A(n15749), .B(n15751), .Z(n35678) );
  XNOR U38235 ( .A(q[0]), .B(DB[2849]), .Z(n15751) );
  XNOR U38236 ( .A(q[3]), .B(DB[2852]), .Z(n15749) );
  IV U38237 ( .A(n15748), .Z(n35677) );
  XNOR U38238 ( .A(n15746), .B(n35679), .Z(n15748) );
  XNOR U38239 ( .A(q[2]), .B(DB[2851]), .Z(n35679) );
  XNOR U38240 ( .A(q[1]), .B(DB[2850]), .Z(n15746) );
  XOR U38241 ( .A(n35680), .B(n15711), .Z(n15674) );
  XOR U38242 ( .A(n35681), .B(n15699), .Z(n15711) );
  XNOR U38243 ( .A(q[6]), .B(DB[2862]), .Z(n15699) );
  IV U38244 ( .A(n15698), .Z(n35681) );
  XNOR U38245 ( .A(n15696), .B(n35682), .Z(n15698) );
  XNOR U38246 ( .A(q[5]), .B(DB[2861]), .Z(n35682) );
  XNOR U38247 ( .A(q[4]), .B(DB[2860]), .Z(n15696) );
  IV U38248 ( .A(n15710), .Z(n35680) );
  XOR U38249 ( .A(n35683), .B(n35684), .Z(n15710) );
  XNOR U38250 ( .A(n15706), .B(n15708), .Z(n35684) );
  XNOR U38251 ( .A(q[0]), .B(DB[2856]), .Z(n15708) );
  XNOR U38252 ( .A(q[3]), .B(DB[2859]), .Z(n15706) );
  IV U38253 ( .A(n15705), .Z(n35683) );
  XNOR U38254 ( .A(n15703), .B(n35685), .Z(n15705) );
  XNOR U38255 ( .A(q[2]), .B(DB[2858]), .Z(n35685) );
  XNOR U38256 ( .A(q[1]), .B(DB[2857]), .Z(n15703) );
  XOR U38257 ( .A(n35686), .B(n15668), .Z(n15631) );
  XOR U38258 ( .A(n35687), .B(n15656), .Z(n15668) );
  XNOR U38259 ( .A(q[6]), .B(DB[2869]), .Z(n15656) );
  IV U38260 ( .A(n15655), .Z(n35687) );
  XNOR U38261 ( .A(n15653), .B(n35688), .Z(n15655) );
  XNOR U38262 ( .A(q[5]), .B(DB[2868]), .Z(n35688) );
  XNOR U38263 ( .A(q[4]), .B(DB[2867]), .Z(n15653) );
  IV U38264 ( .A(n15667), .Z(n35686) );
  XOR U38265 ( .A(n35689), .B(n35690), .Z(n15667) );
  XNOR U38266 ( .A(n15663), .B(n15665), .Z(n35690) );
  XNOR U38267 ( .A(q[0]), .B(DB[2863]), .Z(n15665) );
  XNOR U38268 ( .A(q[3]), .B(DB[2866]), .Z(n15663) );
  IV U38269 ( .A(n15662), .Z(n35689) );
  XNOR U38270 ( .A(n15660), .B(n35691), .Z(n15662) );
  XNOR U38271 ( .A(q[2]), .B(DB[2865]), .Z(n35691) );
  XNOR U38272 ( .A(q[1]), .B(DB[2864]), .Z(n15660) );
  XOR U38273 ( .A(n35692), .B(n15625), .Z(n15588) );
  XOR U38274 ( .A(n35693), .B(n15613), .Z(n15625) );
  XNOR U38275 ( .A(q[6]), .B(DB[2876]), .Z(n15613) );
  IV U38276 ( .A(n15612), .Z(n35693) );
  XNOR U38277 ( .A(n15610), .B(n35694), .Z(n15612) );
  XNOR U38278 ( .A(q[5]), .B(DB[2875]), .Z(n35694) );
  XNOR U38279 ( .A(q[4]), .B(DB[2874]), .Z(n15610) );
  IV U38280 ( .A(n15624), .Z(n35692) );
  XOR U38281 ( .A(n35695), .B(n35696), .Z(n15624) );
  XNOR U38282 ( .A(n15620), .B(n15622), .Z(n35696) );
  XNOR U38283 ( .A(q[0]), .B(DB[2870]), .Z(n15622) );
  XNOR U38284 ( .A(q[3]), .B(DB[2873]), .Z(n15620) );
  IV U38285 ( .A(n15619), .Z(n35695) );
  XNOR U38286 ( .A(n15617), .B(n35697), .Z(n15619) );
  XNOR U38287 ( .A(q[2]), .B(DB[2872]), .Z(n35697) );
  XNOR U38288 ( .A(q[1]), .B(DB[2871]), .Z(n15617) );
  XOR U38289 ( .A(n35698), .B(n15582), .Z(n15545) );
  XOR U38290 ( .A(n35699), .B(n15570), .Z(n15582) );
  XNOR U38291 ( .A(q[6]), .B(DB[2883]), .Z(n15570) );
  IV U38292 ( .A(n15569), .Z(n35699) );
  XNOR U38293 ( .A(n15567), .B(n35700), .Z(n15569) );
  XNOR U38294 ( .A(q[5]), .B(DB[2882]), .Z(n35700) );
  XNOR U38295 ( .A(q[4]), .B(DB[2881]), .Z(n15567) );
  IV U38296 ( .A(n15581), .Z(n35698) );
  XOR U38297 ( .A(n35701), .B(n35702), .Z(n15581) );
  XNOR U38298 ( .A(n15577), .B(n15579), .Z(n35702) );
  XNOR U38299 ( .A(q[0]), .B(DB[2877]), .Z(n15579) );
  XNOR U38300 ( .A(q[3]), .B(DB[2880]), .Z(n15577) );
  IV U38301 ( .A(n15576), .Z(n35701) );
  XNOR U38302 ( .A(n15574), .B(n35703), .Z(n15576) );
  XNOR U38303 ( .A(q[2]), .B(DB[2879]), .Z(n35703) );
  XNOR U38304 ( .A(q[1]), .B(DB[2878]), .Z(n15574) );
  XOR U38305 ( .A(n35704), .B(n15539), .Z(n15502) );
  XOR U38306 ( .A(n35705), .B(n15527), .Z(n15539) );
  XNOR U38307 ( .A(q[6]), .B(DB[2890]), .Z(n15527) );
  IV U38308 ( .A(n15526), .Z(n35705) );
  XNOR U38309 ( .A(n15524), .B(n35706), .Z(n15526) );
  XNOR U38310 ( .A(q[5]), .B(DB[2889]), .Z(n35706) );
  XNOR U38311 ( .A(q[4]), .B(DB[2888]), .Z(n15524) );
  IV U38312 ( .A(n15538), .Z(n35704) );
  XOR U38313 ( .A(n35707), .B(n35708), .Z(n15538) );
  XNOR U38314 ( .A(n15534), .B(n15536), .Z(n35708) );
  XNOR U38315 ( .A(q[0]), .B(DB[2884]), .Z(n15536) );
  XNOR U38316 ( .A(q[3]), .B(DB[2887]), .Z(n15534) );
  IV U38317 ( .A(n15533), .Z(n35707) );
  XNOR U38318 ( .A(n15531), .B(n35709), .Z(n15533) );
  XNOR U38319 ( .A(q[2]), .B(DB[2886]), .Z(n35709) );
  XNOR U38320 ( .A(q[1]), .B(DB[2885]), .Z(n15531) );
  XOR U38321 ( .A(n35710), .B(n15496), .Z(n15459) );
  XOR U38322 ( .A(n35711), .B(n15484), .Z(n15496) );
  XNOR U38323 ( .A(q[6]), .B(DB[2897]), .Z(n15484) );
  IV U38324 ( .A(n15483), .Z(n35711) );
  XNOR U38325 ( .A(n15481), .B(n35712), .Z(n15483) );
  XNOR U38326 ( .A(q[5]), .B(DB[2896]), .Z(n35712) );
  XNOR U38327 ( .A(q[4]), .B(DB[2895]), .Z(n15481) );
  IV U38328 ( .A(n15495), .Z(n35710) );
  XOR U38329 ( .A(n35713), .B(n35714), .Z(n15495) );
  XNOR U38330 ( .A(n15491), .B(n15493), .Z(n35714) );
  XNOR U38331 ( .A(q[0]), .B(DB[2891]), .Z(n15493) );
  XNOR U38332 ( .A(q[3]), .B(DB[2894]), .Z(n15491) );
  IV U38333 ( .A(n15490), .Z(n35713) );
  XNOR U38334 ( .A(n15488), .B(n35715), .Z(n15490) );
  XNOR U38335 ( .A(q[2]), .B(DB[2893]), .Z(n35715) );
  XNOR U38336 ( .A(q[1]), .B(DB[2892]), .Z(n15488) );
  XOR U38337 ( .A(n35716), .B(n15453), .Z(n15416) );
  XOR U38338 ( .A(n35717), .B(n15441), .Z(n15453) );
  XNOR U38339 ( .A(q[6]), .B(DB[2904]), .Z(n15441) );
  IV U38340 ( .A(n15440), .Z(n35717) );
  XNOR U38341 ( .A(n15438), .B(n35718), .Z(n15440) );
  XNOR U38342 ( .A(q[5]), .B(DB[2903]), .Z(n35718) );
  XNOR U38343 ( .A(q[4]), .B(DB[2902]), .Z(n15438) );
  IV U38344 ( .A(n15452), .Z(n35716) );
  XOR U38345 ( .A(n35719), .B(n35720), .Z(n15452) );
  XNOR U38346 ( .A(n15448), .B(n15450), .Z(n35720) );
  XNOR U38347 ( .A(q[0]), .B(DB[2898]), .Z(n15450) );
  XNOR U38348 ( .A(q[3]), .B(DB[2901]), .Z(n15448) );
  IV U38349 ( .A(n15447), .Z(n35719) );
  XNOR U38350 ( .A(n15445), .B(n35721), .Z(n15447) );
  XNOR U38351 ( .A(q[2]), .B(DB[2900]), .Z(n35721) );
  XNOR U38352 ( .A(q[1]), .B(DB[2899]), .Z(n15445) );
  XOR U38353 ( .A(n35722), .B(n15410), .Z(n15373) );
  XOR U38354 ( .A(n35723), .B(n15398), .Z(n15410) );
  XNOR U38355 ( .A(q[6]), .B(DB[2911]), .Z(n15398) );
  IV U38356 ( .A(n15397), .Z(n35723) );
  XNOR U38357 ( .A(n15395), .B(n35724), .Z(n15397) );
  XNOR U38358 ( .A(q[5]), .B(DB[2910]), .Z(n35724) );
  XNOR U38359 ( .A(q[4]), .B(DB[2909]), .Z(n15395) );
  IV U38360 ( .A(n15409), .Z(n35722) );
  XOR U38361 ( .A(n35725), .B(n35726), .Z(n15409) );
  XNOR U38362 ( .A(n15405), .B(n15407), .Z(n35726) );
  XNOR U38363 ( .A(q[0]), .B(DB[2905]), .Z(n15407) );
  XNOR U38364 ( .A(q[3]), .B(DB[2908]), .Z(n15405) );
  IV U38365 ( .A(n15404), .Z(n35725) );
  XNOR U38366 ( .A(n15402), .B(n35727), .Z(n15404) );
  XNOR U38367 ( .A(q[2]), .B(DB[2907]), .Z(n35727) );
  XNOR U38368 ( .A(q[1]), .B(DB[2906]), .Z(n15402) );
  XOR U38369 ( .A(n35728), .B(n15367), .Z(n15330) );
  XOR U38370 ( .A(n35729), .B(n15355), .Z(n15367) );
  XNOR U38371 ( .A(q[6]), .B(DB[2918]), .Z(n15355) );
  IV U38372 ( .A(n15354), .Z(n35729) );
  XNOR U38373 ( .A(n15352), .B(n35730), .Z(n15354) );
  XNOR U38374 ( .A(q[5]), .B(DB[2917]), .Z(n35730) );
  XNOR U38375 ( .A(q[4]), .B(DB[2916]), .Z(n15352) );
  IV U38376 ( .A(n15366), .Z(n35728) );
  XOR U38377 ( .A(n35731), .B(n35732), .Z(n15366) );
  XNOR U38378 ( .A(n15362), .B(n15364), .Z(n35732) );
  XNOR U38379 ( .A(q[0]), .B(DB[2912]), .Z(n15364) );
  XNOR U38380 ( .A(q[3]), .B(DB[2915]), .Z(n15362) );
  IV U38381 ( .A(n15361), .Z(n35731) );
  XNOR U38382 ( .A(n15359), .B(n35733), .Z(n15361) );
  XNOR U38383 ( .A(q[2]), .B(DB[2914]), .Z(n35733) );
  XNOR U38384 ( .A(q[1]), .B(DB[2913]), .Z(n15359) );
  XOR U38385 ( .A(n35734), .B(n15324), .Z(n15287) );
  XOR U38386 ( .A(n35735), .B(n15312), .Z(n15324) );
  XNOR U38387 ( .A(q[6]), .B(DB[2925]), .Z(n15312) );
  IV U38388 ( .A(n15311), .Z(n35735) );
  XNOR U38389 ( .A(n15309), .B(n35736), .Z(n15311) );
  XNOR U38390 ( .A(q[5]), .B(DB[2924]), .Z(n35736) );
  XNOR U38391 ( .A(q[4]), .B(DB[2923]), .Z(n15309) );
  IV U38392 ( .A(n15323), .Z(n35734) );
  XOR U38393 ( .A(n35737), .B(n35738), .Z(n15323) );
  XNOR U38394 ( .A(n15319), .B(n15321), .Z(n35738) );
  XNOR U38395 ( .A(q[0]), .B(DB[2919]), .Z(n15321) );
  XNOR U38396 ( .A(q[3]), .B(DB[2922]), .Z(n15319) );
  IV U38397 ( .A(n15318), .Z(n35737) );
  XNOR U38398 ( .A(n15316), .B(n35739), .Z(n15318) );
  XNOR U38399 ( .A(q[2]), .B(DB[2921]), .Z(n35739) );
  XNOR U38400 ( .A(q[1]), .B(DB[2920]), .Z(n15316) );
  XOR U38401 ( .A(n35740), .B(n15281), .Z(n15244) );
  XOR U38402 ( .A(n35741), .B(n15269), .Z(n15281) );
  XNOR U38403 ( .A(q[6]), .B(DB[2932]), .Z(n15269) );
  IV U38404 ( .A(n15268), .Z(n35741) );
  XNOR U38405 ( .A(n15266), .B(n35742), .Z(n15268) );
  XNOR U38406 ( .A(q[5]), .B(DB[2931]), .Z(n35742) );
  XNOR U38407 ( .A(q[4]), .B(DB[2930]), .Z(n15266) );
  IV U38408 ( .A(n15280), .Z(n35740) );
  XOR U38409 ( .A(n35743), .B(n35744), .Z(n15280) );
  XNOR U38410 ( .A(n15276), .B(n15278), .Z(n35744) );
  XNOR U38411 ( .A(q[0]), .B(DB[2926]), .Z(n15278) );
  XNOR U38412 ( .A(q[3]), .B(DB[2929]), .Z(n15276) );
  IV U38413 ( .A(n15275), .Z(n35743) );
  XNOR U38414 ( .A(n15273), .B(n35745), .Z(n15275) );
  XNOR U38415 ( .A(q[2]), .B(DB[2928]), .Z(n35745) );
  XNOR U38416 ( .A(q[1]), .B(DB[2927]), .Z(n15273) );
  XOR U38417 ( .A(n35746), .B(n15238), .Z(n15201) );
  XOR U38418 ( .A(n35747), .B(n15226), .Z(n15238) );
  XNOR U38419 ( .A(q[6]), .B(DB[2939]), .Z(n15226) );
  IV U38420 ( .A(n15225), .Z(n35747) );
  XNOR U38421 ( .A(n15223), .B(n35748), .Z(n15225) );
  XNOR U38422 ( .A(q[5]), .B(DB[2938]), .Z(n35748) );
  XNOR U38423 ( .A(q[4]), .B(DB[2937]), .Z(n15223) );
  IV U38424 ( .A(n15237), .Z(n35746) );
  XOR U38425 ( .A(n35749), .B(n35750), .Z(n15237) );
  XNOR U38426 ( .A(n15233), .B(n15235), .Z(n35750) );
  XNOR U38427 ( .A(q[0]), .B(DB[2933]), .Z(n15235) );
  XNOR U38428 ( .A(q[3]), .B(DB[2936]), .Z(n15233) );
  IV U38429 ( .A(n15232), .Z(n35749) );
  XNOR U38430 ( .A(n15230), .B(n35751), .Z(n15232) );
  XNOR U38431 ( .A(q[2]), .B(DB[2935]), .Z(n35751) );
  XNOR U38432 ( .A(q[1]), .B(DB[2934]), .Z(n15230) );
  XOR U38433 ( .A(n35752), .B(n15195), .Z(n15158) );
  XOR U38434 ( .A(n35753), .B(n15183), .Z(n15195) );
  XNOR U38435 ( .A(q[6]), .B(DB[2946]), .Z(n15183) );
  IV U38436 ( .A(n15182), .Z(n35753) );
  XNOR U38437 ( .A(n15180), .B(n35754), .Z(n15182) );
  XNOR U38438 ( .A(q[5]), .B(DB[2945]), .Z(n35754) );
  XNOR U38439 ( .A(q[4]), .B(DB[2944]), .Z(n15180) );
  IV U38440 ( .A(n15194), .Z(n35752) );
  XOR U38441 ( .A(n35755), .B(n35756), .Z(n15194) );
  XNOR U38442 ( .A(n15190), .B(n15192), .Z(n35756) );
  XNOR U38443 ( .A(q[0]), .B(DB[2940]), .Z(n15192) );
  XNOR U38444 ( .A(q[3]), .B(DB[2943]), .Z(n15190) );
  IV U38445 ( .A(n15189), .Z(n35755) );
  XNOR U38446 ( .A(n15187), .B(n35757), .Z(n15189) );
  XNOR U38447 ( .A(q[2]), .B(DB[2942]), .Z(n35757) );
  XNOR U38448 ( .A(q[1]), .B(DB[2941]), .Z(n15187) );
  XOR U38449 ( .A(n35758), .B(n15152), .Z(n15115) );
  XOR U38450 ( .A(n35759), .B(n15140), .Z(n15152) );
  XNOR U38451 ( .A(q[6]), .B(DB[2953]), .Z(n15140) );
  IV U38452 ( .A(n15139), .Z(n35759) );
  XNOR U38453 ( .A(n15137), .B(n35760), .Z(n15139) );
  XNOR U38454 ( .A(q[5]), .B(DB[2952]), .Z(n35760) );
  XNOR U38455 ( .A(q[4]), .B(DB[2951]), .Z(n15137) );
  IV U38456 ( .A(n15151), .Z(n35758) );
  XOR U38457 ( .A(n35761), .B(n35762), .Z(n15151) );
  XNOR U38458 ( .A(n15147), .B(n15149), .Z(n35762) );
  XNOR U38459 ( .A(q[0]), .B(DB[2947]), .Z(n15149) );
  XNOR U38460 ( .A(q[3]), .B(DB[2950]), .Z(n15147) );
  IV U38461 ( .A(n15146), .Z(n35761) );
  XNOR U38462 ( .A(n15144), .B(n35763), .Z(n15146) );
  XNOR U38463 ( .A(q[2]), .B(DB[2949]), .Z(n35763) );
  XNOR U38464 ( .A(q[1]), .B(DB[2948]), .Z(n15144) );
  XOR U38465 ( .A(n35764), .B(n15109), .Z(n15072) );
  XOR U38466 ( .A(n35765), .B(n15097), .Z(n15109) );
  XNOR U38467 ( .A(q[6]), .B(DB[2960]), .Z(n15097) );
  IV U38468 ( .A(n15096), .Z(n35765) );
  XNOR U38469 ( .A(n15094), .B(n35766), .Z(n15096) );
  XNOR U38470 ( .A(q[5]), .B(DB[2959]), .Z(n35766) );
  XNOR U38471 ( .A(q[4]), .B(DB[2958]), .Z(n15094) );
  IV U38472 ( .A(n15108), .Z(n35764) );
  XOR U38473 ( .A(n35767), .B(n35768), .Z(n15108) );
  XNOR U38474 ( .A(n15104), .B(n15106), .Z(n35768) );
  XNOR U38475 ( .A(q[0]), .B(DB[2954]), .Z(n15106) );
  XNOR U38476 ( .A(q[3]), .B(DB[2957]), .Z(n15104) );
  IV U38477 ( .A(n15103), .Z(n35767) );
  XNOR U38478 ( .A(n15101), .B(n35769), .Z(n15103) );
  XNOR U38479 ( .A(q[2]), .B(DB[2956]), .Z(n35769) );
  XNOR U38480 ( .A(q[1]), .B(DB[2955]), .Z(n15101) );
  XOR U38481 ( .A(n35770), .B(n15066), .Z(n15029) );
  XOR U38482 ( .A(n35771), .B(n15054), .Z(n15066) );
  XNOR U38483 ( .A(q[6]), .B(DB[2967]), .Z(n15054) );
  IV U38484 ( .A(n15053), .Z(n35771) );
  XNOR U38485 ( .A(n15051), .B(n35772), .Z(n15053) );
  XNOR U38486 ( .A(q[5]), .B(DB[2966]), .Z(n35772) );
  XNOR U38487 ( .A(q[4]), .B(DB[2965]), .Z(n15051) );
  IV U38488 ( .A(n15065), .Z(n35770) );
  XOR U38489 ( .A(n35773), .B(n35774), .Z(n15065) );
  XNOR U38490 ( .A(n15061), .B(n15063), .Z(n35774) );
  XNOR U38491 ( .A(q[0]), .B(DB[2961]), .Z(n15063) );
  XNOR U38492 ( .A(q[3]), .B(DB[2964]), .Z(n15061) );
  IV U38493 ( .A(n15060), .Z(n35773) );
  XNOR U38494 ( .A(n15058), .B(n35775), .Z(n15060) );
  XNOR U38495 ( .A(q[2]), .B(DB[2963]), .Z(n35775) );
  XNOR U38496 ( .A(q[1]), .B(DB[2962]), .Z(n15058) );
  XOR U38497 ( .A(n35776), .B(n15023), .Z(n14986) );
  XOR U38498 ( .A(n35777), .B(n15011), .Z(n15023) );
  XNOR U38499 ( .A(q[6]), .B(DB[2974]), .Z(n15011) );
  IV U38500 ( .A(n15010), .Z(n35777) );
  XNOR U38501 ( .A(n15008), .B(n35778), .Z(n15010) );
  XNOR U38502 ( .A(q[5]), .B(DB[2973]), .Z(n35778) );
  XNOR U38503 ( .A(q[4]), .B(DB[2972]), .Z(n15008) );
  IV U38504 ( .A(n15022), .Z(n35776) );
  XOR U38505 ( .A(n35779), .B(n35780), .Z(n15022) );
  XNOR U38506 ( .A(n15018), .B(n15020), .Z(n35780) );
  XNOR U38507 ( .A(q[0]), .B(DB[2968]), .Z(n15020) );
  XNOR U38508 ( .A(q[3]), .B(DB[2971]), .Z(n15018) );
  IV U38509 ( .A(n15017), .Z(n35779) );
  XNOR U38510 ( .A(n15015), .B(n35781), .Z(n15017) );
  XNOR U38511 ( .A(q[2]), .B(DB[2970]), .Z(n35781) );
  XNOR U38512 ( .A(q[1]), .B(DB[2969]), .Z(n15015) );
  XOR U38513 ( .A(n35782), .B(n14980), .Z(n14943) );
  XOR U38514 ( .A(n35783), .B(n14968), .Z(n14980) );
  XNOR U38515 ( .A(q[6]), .B(DB[2981]), .Z(n14968) );
  IV U38516 ( .A(n14967), .Z(n35783) );
  XNOR U38517 ( .A(n14965), .B(n35784), .Z(n14967) );
  XNOR U38518 ( .A(q[5]), .B(DB[2980]), .Z(n35784) );
  XNOR U38519 ( .A(q[4]), .B(DB[2979]), .Z(n14965) );
  IV U38520 ( .A(n14979), .Z(n35782) );
  XOR U38521 ( .A(n35785), .B(n35786), .Z(n14979) );
  XNOR U38522 ( .A(n14975), .B(n14977), .Z(n35786) );
  XNOR U38523 ( .A(q[0]), .B(DB[2975]), .Z(n14977) );
  XNOR U38524 ( .A(q[3]), .B(DB[2978]), .Z(n14975) );
  IV U38525 ( .A(n14974), .Z(n35785) );
  XNOR U38526 ( .A(n14972), .B(n35787), .Z(n14974) );
  XNOR U38527 ( .A(q[2]), .B(DB[2977]), .Z(n35787) );
  XNOR U38528 ( .A(q[1]), .B(DB[2976]), .Z(n14972) );
  XOR U38529 ( .A(n35788), .B(n14937), .Z(n14900) );
  XOR U38530 ( .A(n35789), .B(n14925), .Z(n14937) );
  XNOR U38531 ( .A(q[6]), .B(DB[2988]), .Z(n14925) );
  IV U38532 ( .A(n14924), .Z(n35789) );
  XNOR U38533 ( .A(n14922), .B(n35790), .Z(n14924) );
  XNOR U38534 ( .A(q[5]), .B(DB[2987]), .Z(n35790) );
  XNOR U38535 ( .A(q[4]), .B(DB[2986]), .Z(n14922) );
  IV U38536 ( .A(n14936), .Z(n35788) );
  XOR U38537 ( .A(n35791), .B(n35792), .Z(n14936) );
  XNOR U38538 ( .A(n14932), .B(n14934), .Z(n35792) );
  XNOR U38539 ( .A(q[0]), .B(DB[2982]), .Z(n14934) );
  XNOR U38540 ( .A(q[3]), .B(DB[2985]), .Z(n14932) );
  IV U38541 ( .A(n14931), .Z(n35791) );
  XNOR U38542 ( .A(n14929), .B(n35793), .Z(n14931) );
  XNOR U38543 ( .A(q[2]), .B(DB[2984]), .Z(n35793) );
  XNOR U38544 ( .A(q[1]), .B(DB[2983]), .Z(n14929) );
  XOR U38545 ( .A(n35794), .B(n14894), .Z(n14857) );
  XOR U38546 ( .A(n35795), .B(n14882), .Z(n14894) );
  XNOR U38547 ( .A(q[6]), .B(DB[2995]), .Z(n14882) );
  IV U38548 ( .A(n14881), .Z(n35795) );
  XNOR U38549 ( .A(n14879), .B(n35796), .Z(n14881) );
  XNOR U38550 ( .A(q[5]), .B(DB[2994]), .Z(n35796) );
  XNOR U38551 ( .A(q[4]), .B(DB[2993]), .Z(n14879) );
  IV U38552 ( .A(n14893), .Z(n35794) );
  XOR U38553 ( .A(n35797), .B(n35798), .Z(n14893) );
  XNOR U38554 ( .A(n14889), .B(n14891), .Z(n35798) );
  XNOR U38555 ( .A(q[0]), .B(DB[2989]), .Z(n14891) );
  XNOR U38556 ( .A(q[3]), .B(DB[2992]), .Z(n14889) );
  IV U38557 ( .A(n14888), .Z(n35797) );
  XNOR U38558 ( .A(n14886), .B(n35799), .Z(n14888) );
  XNOR U38559 ( .A(q[2]), .B(DB[2991]), .Z(n35799) );
  XNOR U38560 ( .A(q[1]), .B(DB[2990]), .Z(n14886) );
  XOR U38561 ( .A(n35800), .B(n14851), .Z(n14814) );
  XOR U38562 ( .A(n35801), .B(n14839), .Z(n14851) );
  XNOR U38563 ( .A(q[6]), .B(DB[3002]), .Z(n14839) );
  IV U38564 ( .A(n14838), .Z(n35801) );
  XNOR U38565 ( .A(n14836), .B(n35802), .Z(n14838) );
  XNOR U38566 ( .A(q[5]), .B(DB[3001]), .Z(n35802) );
  XNOR U38567 ( .A(q[4]), .B(DB[3000]), .Z(n14836) );
  IV U38568 ( .A(n14850), .Z(n35800) );
  XOR U38569 ( .A(n35803), .B(n35804), .Z(n14850) );
  XNOR U38570 ( .A(n14846), .B(n14848), .Z(n35804) );
  XNOR U38571 ( .A(q[0]), .B(DB[2996]), .Z(n14848) );
  XNOR U38572 ( .A(q[3]), .B(DB[2999]), .Z(n14846) );
  IV U38573 ( .A(n14845), .Z(n35803) );
  XNOR U38574 ( .A(n14843), .B(n35805), .Z(n14845) );
  XNOR U38575 ( .A(q[2]), .B(DB[2998]), .Z(n35805) );
  XNOR U38576 ( .A(q[1]), .B(DB[2997]), .Z(n14843) );
  XOR U38577 ( .A(n35806), .B(n14808), .Z(n14771) );
  XOR U38578 ( .A(n35807), .B(n14796), .Z(n14808) );
  XNOR U38579 ( .A(q[6]), .B(DB[3009]), .Z(n14796) );
  IV U38580 ( .A(n14795), .Z(n35807) );
  XNOR U38581 ( .A(n14793), .B(n35808), .Z(n14795) );
  XNOR U38582 ( .A(q[5]), .B(DB[3008]), .Z(n35808) );
  XNOR U38583 ( .A(q[4]), .B(DB[3007]), .Z(n14793) );
  IV U38584 ( .A(n14807), .Z(n35806) );
  XOR U38585 ( .A(n35809), .B(n35810), .Z(n14807) );
  XNOR U38586 ( .A(n14803), .B(n14805), .Z(n35810) );
  XNOR U38587 ( .A(q[0]), .B(DB[3003]), .Z(n14805) );
  XNOR U38588 ( .A(q[3]), .B(DB[3006]), .Z(n14803) );
  IV U38589 ( .A(n14802), .Z(n35809) );
  XNOR U38590 ( .A(n14800), .B(n35811), .Z(n14802) );
  XNOR U38591 ( .A(q[2]), .B(DB[3005]), .Z(n35811) );
  XNOR U38592 ( .A(q[1]), .B(DB[3004]), .Z(n14800) );
  XOR U38593 ( .A(n35812), .B(n14765), .Z(n14728) );
  XOR U38594 ( .A(n35813), .B(n14753), .Z(n14765) );
  XNOR U38595 ( .A(q[6]), .B(DB[3016]), .Z(n14753) );
  IV U38596 ( .A(n14752), .Z(n35813) );
  XNOR U38597 ( .A(n14750), .B(n35814), .Z(n14752) );
  XNOR U38598 ( .A(q[5]), .B(DB[3015]), .Z(n35814) );
  XNOR U38599 ( .A(q[4]), .B(DB[3014]), .Z(n14750) );
  IV U38600 ( .A(n14764), .Z(n35812) );
  XOR U38601 ( .A(n35815), .B(n35816), .Z(n14764) );
  XNOR U38602 ( .A(n14760), .B(n14762), .Z(n35816) );
  XNOR U38603 ( .A(q[0]), .B(DB[3010]), .Z(n14762) );
  XNOR U38604 ( .A(q[3]), .B(DB[3013]), .Z(n14760) );
  IV U38605 ( .A(n14759), .Z(n35815) );
  XNOR U38606 ( .A(n14757), .B(n35817), .Z(n14759) );
  XNOR U38607 ( .A(q[2]), .B(DB[3012]), .Z(n35817) );
  XNOR U38608 ( .A(q[1]), .B(DB[3011]), .Z(n14757) );
  XOR U38609 ( .A(n35818), .B(n14722), .Z(n14685) );
  XOR U38610 ( .A(n35819), .B(n14710), .Z(n14722) );
  XNOR U38611 ( .A(q[6]), .B(DB[3023]), .Z(n14710) );
  IV U38612 ( .A(n14709), .Z(n35819) );
  XNOR U38613 ( .A(n14707), .B(n35820), .Z(n14709) );
  XNOR U38614 ( .A(q[5]), .B(DB[3022]), .Z(n35820) );
  XNOR U38615 ( .A(q[4]), .B(DB[3021]), .Z(n14707) );
  IV U38616 ( .A(n14721), .Z(n35818) );
  XOR U38617 ( .A(n35821), .B(n35822), .Z(n14721) );
  XNOR U38618 ( .A(n14717), .B(n14719), .Z(n35822) );
  XNOR U38619 ( .A(q[0]), .B(DB[3017]), .Z(n14719) );
  XNOR U38620 ( .A(q[3]), .B(DB[3020]), .Z(n14717) );
  IV U38621 ( .A(n14716), .Z(n35821) );
  XNOR U38622 ( .A(n14714), .B(n35823), .Z(n14716) );
  XNOR U38623 ( .A(q[2]), .B(DB[3019]), .Z(n35823) );
  XNOR U38624 ( .A(q[1]), .B(DB[3018]), .Z(n14714) );
  XOR U38625 ( .A(n35824), .B(n14679), .Z(n14642) );
  XOR U38626 ( .A(n35825), .B(n14667), .Z(n14679) );
  XNOR U38627 ( .A(q[6]), .B(DB[3030]), .Z(n14667) );
  IV U38628 ( .A(n14666), .Z(n35825) );
  XNOR U38629 ( .A(n14664), .B(n35826), .Z(n14666) );
  XNOR U38630 ( .A(q[5]), .B(DB[3029]), .Z(n35826) );
  XNOR U38631 ( .A(q[4]), .B(DB[3028]), .Z(n14664) );
  IV U38632 ( .A(n14678), .Z(n35824) );
  XOR U38633 ( .A(n35827), .B(n35828), .Z(n14678) );
  XNOR U38634 ( .A(n14674), .B(n14676), .Z(n35828) );
  XNOR U38635 ( .A(q[0]), .B(DB[3024]), .Z(n14676) );
  XNOR U38636 ( .A(q[3]), .B(DB[3027]), .Z(n14674) );
  IV U38637 ( .A(n14673), .Z(n35827) );
  XNOR U38638 ( .A(n14671), .B(n35829), .Z(n14673) );
  XNOR U38639 ( .A(q[2]), .B(DB[3026]), .Z(n35829) );
  XNOR U38640 ( .A(q[1]), .B(DB[3025]), .Z(n14671) );
  XOR U38641 ( .A(n35830), .B(n14636), .Z(n14599) );
  XOR U38642 ( .A(n35831), .B(n14624), .Z(n14636) );
  XNOR U38643 ( .A(q[6]), .B(DB[3037]), .Z(n14624) );
  IV U38644 ( .A(n14623), .Z(n35831) );
  XNOR U38645 ( .A(n14621), .B(n35832), .Z(n14623) );
  XNOR U38646 ( .A(q[5]), .B(DB[3036]), .Z(n35832) );
  XNOR U38647 ( .A(q[4]), .B(DB[3035]), .Z(n14621) );
  IV U38648 ( .A(n14635), .Z(n35830) );
  XOR U38649 ( .A(n35833), .B(n35834), .Z(n14635) );
  XNOR U38650 ( .A(n14631), .B(n14633), .Z(n35834) );
  XNOR U38651 ( .A(q[0]), .B(DB[3031]), .Z(n14633) );
  XNOR U38652 ( .A(q[3]), .B(DB[3034]), .Z(n14631) );
  IV U38653 ( .A(n14630), .Z(n35833) );
  XNOR U38654 ( .A(n14628), .B(n35835), .Z(n14630) );
  XNOR U38655 ( .A(q[2]), .B(DB[3033]), .Z(n35835) );
  XNOR U38656 ( .A(q[1]), .B(DB[3032]), .Z(n14628) );
  XOR U38657 ( .A(n35836), .B(n14593), .Z(n14556) );
  XOR U38658 ( .A(n35837), .B(n14581), .Z(n14593) );
  XNOR U38659 ( .A(q[6]), .B(DB[3044]), .Z(n14581) );
  IV U38660 ( .A(n14580), .Z(n35837) );
  XNOR U38661 ( .A(n14578), .B(n35838), .Z(n14580) );
  XNOR U38662 ( .A(q[5]), .B(DB[3043]), .Z(n35838) );
  XNOR U38663 ( .A(q[4]), .B(DB[3042]), .Z(n14578) );
  IV U38664 ( .A(n14592), .Z(n35836) );
  XOR U38665 ( .A(n35839), .B(n35840), .Z(n14592) );
  XNOR U38666 ( .A(n14588), .B(n14590), .Z(n35840) );
  XNOR U38667 ( .A(q[0]), .B(DB[3038]), .Z(n14590) );
  XNOR U38668 ( .A(q[3]), .B(DB[3041]), .Z(n14588) );
  IV U38669 ( .A(n14587), .Z(n35839) );
  XNOR U38670 ( .A(n14585), .B(n35841), .Z(n14587) );
  XNOR U38671 ( .A(q[2]), .B(DB[3040]), .Z(n35841) );
  XNOR U38672 ( .A(q[1]), .B(DB[3039]), .Z(n14585) );
  XOR U38673 ( .A(n35842), .B(n14550), .Z(n14513) );
  XOR U38674 ( .A(n35843), .B(n14538), .Z(n14550) );
  XNOR U38675 ( .A(q[6]), .B(DB[3051]), .Z(n14538) );
  IV U38676 ( .A(n14537), .Z(n35843) );
  XNOR U38677 ( .A(n14535), .B(n35844), .Z(n14537) );
  XNOR U38678 ( .A(q[5]), .B(DB[3050]), .Z(n35844) );
  XNOR U38679 ( .A(q[4]), .B(DB[3049]), .Z(n14535) );
  IV U38680 ( .A(n14549), .Z(n35842) );
  XOR U38681 ( .A(n35845), .B(n35846), .Z(n14549) );
  XNOR U38682 ( .A(n14545), .B(n14547), .Z(n35846) );
  XNOR U38683 ( .A(q[0]), .B(DB[3045]), .Z(n14547) );
  XNOR U38684 ( .A(q[3]), .B(DB[3048]), .Z(n14545) );
  IV U38685 ( .A(n14544), .Z(n35845) );
  XNOR U38686 ( .A(n14542), .B(n35847), .Z(n14544) );
  XNOR U38687 ( .A(q[2]), .B(DB[3047]), .Z(n35847) );
  XNOR U38688 ( .A(q[1]), .B(DB[3046]), .Z(n14542) );
  XOR U38689 ( .A(n35848), .B(n14507), .Z(n14470) );
  XOR U38690 ( .A(n35849), .B(n14495), .Z(n14507) );
  XNOR U38691 ( .A(q[6]), .B(DB[3058]), .Z(n14495) );
  IV U38692 ( .A(n14494), .Z(n35849) );
  XNOR U38693 ( .A(n14492), .B(n35850), .Z(n14494) );
  XNOR U38694 ( .A(q[5]), .B(DB[3057]), .Z(n35850) );
  XNOR U38695 ( .A(q[4]), .B(DB[3056]), .Z(n14492) );
  IV U38696 ( .A(n14506), .Z(n35848) );
  XOR U38697 ( .A(n35851), .B(n35852), .Z(n14506) );
  XNOR U38698 ( .A(n14502), .B(n14504), .Z(n35852) );
  XNOR U38699 ( .A(q[0]), .B(DB[3052]), .Z(n14504) );
  XNOR U38700 ( .A(q[3]), .B(DB[3055]), .Z(n14502) );
  IV U38701 ( .A(n14501), .Z(n35851) );
  XNOR U38702 ( .A(n14499), .B(n35853), .Z(n14501) );
  XNOR U38703 ( .A(q[2]), .B(DB[3054]), .Z(n35853) );
  XNOR U38704 ( .A(q[1]), .B(DB[3053]), .Z(n14499) );
  XOR U38705 ( .A(n35854), .B(n14464), .Z(n14427) );
  XOR U38706 ( .A(n35855), .B(n14452), .Z(n14464) );
  XNOR U38707 ( .A(q[6]), .B(DB[3065]), .Z(n14452) );
  IV U38708 ( .A(n14451), .Z(n35855) );
  XNOR U38709 ( .A(n14449), .B(n35856), .Z(n14451) );
  XNOR U38710 ( .A(q[5]), .B(DB[3064]), .Z(n35856) );
  XNOR U38711 ( .A(q[4]), .B(DB[3063]), .Z(n14449) );
  IV U38712 ( .A(n14463), .Z(n35854) );
  XOR U38713 ( .A(n35857), .B(n35858), .Z(n14463) );
  XNOR U38714 ( .A(n14459), .B(n14461), .Z(n35858) );
  XNOR U38715 ( .A(q[0]), .B(DB[3059]), .Z(n14461) );
  XNOR U38716 ( .A(q[3]), .B(DB[3062]), .Z(n14459) );
  IV U38717 ( .A(n14458), .Z(n35857) );
  XNOR U38718 ( .A(n14456), .B(n35859), .Z(n14458) );
  XNOR U38719 ( .A(q[2]), .B(DB[3061]), .Z(n35859) );
  XNOR U38720 ( .A(q[1]), .B(DB[3060]), .Z(n14456) );
  XOR U38721 ( .A(n35860), .B(n14421), .Z(n14384) );
  XOR U38722 ( .A(n35861), .B(n14409), .Z(n14421) );
  XNOR U38723 ( .A(q[6]), .B(DB[3072]), .Z(n14409) );
  IV U38724 ( .A(n14408), .Z(n35861) );
  XNOR U38725 ( .A(n14406), .B(n35862), .Z(n14408) );
  XNOR U38726 ( .A(q[5]), .B(DB[3071]), .Z(n35862) );
  XNOR U38727 ( .A(q[4]), .B(DB[3070]), .Z(n14406) );
  IV U38728 ( .A(n14420), .Z(n35860) );
  XOR U38729 ( .A(n35863), .B(n35864), .Z(n14420) );
  XNOR U38730 ( .A(n14416), .B(n14418), .Z(n35864) );
  XNOR U38731 ( .A(q[0]), .B(DB[3066]), .Z(n14418) );
  XNOR U38732 ( .A(q[3]), .B(DB[3069]), .Z(n14416) );
  IV U38733 ( .A(n14415), .Z(n35863) );
  XNOR U38734 ( .A(n14413), .B(n35865), .Z(n14415) );
  XNOR U38735 ( .A(q[2]), .B(DB[3068]), .Z(n35865) );
  XNOR U38736 ( .A(q[1]), .B(DB[3067]), .Z(n14413) );
  XOR U38737 ( .A(n35866), .B(n14378), .Z(n14341) );
  XOR U38738 ( .A(n35867), .B(n14366), .Z(n14378) );
  XNOR U38739 ( .A(q[6]), .B(DB[3079]), .Z(n14366) );
  IV U38740 ( .A(n14365), .Z(n35867) );
  XNOR U38741 ( .A(n14363), .B(n35868), .Z(n14365) );
  XNOR U38742 ( .A(q[5]), .B(DB[3078]), .Z(n35868) );
  XNOR U38743 ( .A(q[4]), .B(DB[3077]), .Z(n14363) );
  IV U38744 ( .A(n14377), .Z(n35866) );
  XOR U38745 ( .A(n35869), .B(n35870), .Z(n14377) );
  XNOR U38746 ( .A(n14373), .B(n14375), .Z(n35870) );
  XNOR U38747 ( .A(q[0]), .B(DB[3073]), .Z(n14375) );
  XNOR U38748 ( .A(q[3]), .B(DB[3076]), .Z(n14373) );
  IV U38749 ( .A(n14372), .Z(n35869) );
  XNOR U38750 ( .A(n14370), .B(n35871), .Z(n14372) );
  XNOR U38751 ( .A(q[2]), .B(DB[3075]), .Z(n35871) );
  XNOR U38752 ( .A(q[1]), .B(DB[3074]), .Z(n14370) );
  XOR U38753 ( .A(n35872), .B(n14335), .Z(n14298) );
  XOR U38754 ( .A(n35873), .B(n14323), .Z(n14335) );
  XNOR U38755 ( .A(q[6]), .B(DB[3086]), .Z(n14323) );
  IV U38756 ( .A(n14322), .Z(n35873) );
  XNOR U38757 ( .A(n14320), .B(n35874), .Z(n14322) );
  XNOR U38758 ( .A(q[5]), .B(DB[3085]), .Z(n35874) );
  XNOR U38759 ( .A(q[4]), .B(DB[3084]), .Z(n14320) );
  IV U38760 ( .A(n14334), .Z(n35872) );
  XOR U38761 ( .A(n35875), .B(n35876), .Z(n14334) );
  XNOR U38762 ( .A(n14330), .B(n14332), .Z(n35876) );
  XNOR U38763 ( .A(q[0]), .B(DB[3080]), .Z(n14332) );
  XNOR U38764 ( .A(q[3]), .B(DB[3083]), .Z(n14330) );
  IV U38765 ( .A(n14329), .Z(n35875) );
  XNOR U38766 ( .A(n14327), .B(n35877), .Z(n14329) );
  XNOR U38767 ( .A(q[2]), .B(DB[3082]), .Z(n35877) );
  XNOR U38768 ( .A(q[1]), .B(DB[3081]), .Z(n14327) );
  XOR U38769 ( .A(n35878), .B(n14292), .Z(n14255) );
  XOR U38770 ( .A(n35879), .B(n14280), .Z(n14292) );
  XNOR U38771 ( .A(q[6]), .B(DB[3093]), .Z(n14280) );
  IV U38772 ( .A(n14279), .Z(n35879) );
  XNOR U38773 ( .A(n14277), .B(n35880), .Z(n14279) );
  XNOR U38774 ( .A(q[5]), .B(DB[3092]), .Z(n35880) );
  XNOR U38775 ( .A(q[4]), .B(DB[3091]), .Z(n14277) );
  IV U38776 ( .A(n14291), .Z(n35878) );
  XOR U38777 ( .A(n35881), .B(n35882), .Z(n14291) );
  XNOR U38778 ( .A(n14287), .B(n14289), .Z(n35882) );
  XNOR U38779 ( .A(q[0]), .B(DB[3087]), .Z(n14289) );
  XNOR U38780 ( .A(q[3]), .B(DB[3090]), .Z(n14287) );
  IV U38781 ( .A(n14286), .Z(n35881) );
  XNOR U38782 ( .A(n14284), .B(n35883), .Z(n14286) );
  XNOR U38783 ( .A(q[2]), .B(DB[3089]), .Z(n35883) );
  XNOR U38784 ( .A(q[1]), .B(DB[3088]), .Z(n14284) );
  XOR U38785 ( .A(n35884), .B(n14249), .Z(n14212) );
  XOR U38786 ( .A(n35885), .B(n14237), .Z(n14249) );
  XNOR U38787 ( .A(q[6]), .B(DB[3100]), .Z(n14237) );
  IV U38788 ( .A(n14236), .Z(n35885) );
  XNOR U38789 ( .A(n14234), .B(n35886), .Z(n14236) );
  XNOR U38790 ( .A(q[5]), .B(DB[3099]), .Z(n35886) );
  XNOR U38791 ( .A(q[4]), .B(DB[3098]), .Z(n14234) );
  IV U38792 ( .A(n14248), .Z(n35884) );
  XOR U38793 ( .A(n35887), .B(n35888), .Z(n14248) );
  XNOR U38794 ( .A(n14244), .B(n14246), .Z(n35888) );
  XNOR U38795 ( .A(q[0]), .B(DB[3094]), .Z(n14246) );
  XNOR U38796 ( .A(q[3]), .B(DB[3097]), .Z(n14244) );
  IV U38797 ( .A(n14243), .Z(n35887) );
  XNOR U38798 ( .A(n14241), .B(n35889), .Z(n14243) );
  XNOR U38799 ( .A(q[2]), .B(DB[3096]), .Z(n35889) );
  XNOR U38800 ( .A(q[1]), .B(DB[3095]), .Z(n14241) );
  XOR U38801 ( .A(n35890), .B(n14206), .Z(n14169) );
  XOR U38802 ( .A(n35891), .B(n14194), .Z(n14206) );
  XNOR U38803 ( .A(q[6]), .B(DB[3107]), .Z(n14194) );
  IV U38804 ( .A(n14193), .Z(n35891) );
  XNOR U38805 ( .A(n14191), .B(n35892), .Z(n14193) );
  XNOR U38806 ( .A(q[5]), .B(DB[3106]), .Z(n35892) );
  XNOR U38807 ( .A(q[4]), .B(DB[3105]), .Z(n14191) );
  IV U38808 ( .A(n14205), .Z(n35890) );
  XOR U38809 ( .A(n35893), .B(n35894), .Z(n14205) );
  XNOR U38810 ( .A(n14201), .B(n14203), .Z(n35894) );
  XNOR U38811 ( .A(q[0]), .B(DB[3101]), .Z(n14203) );
  XNOR U38812 ( .A(q[3]), .B(DB[3104]), .Z(n14201) );
  IV U38813 ( .A(n14200), .Z(n35893) );
  XNOR U38814 ( .A(n14198), .B(n35895), .Z(n14200) );
  XNOR U38815 ( .A(q[2]), .B(DB[3103]), .Z(n35895) );
  XNOR U38816 ( .A(q[1]), .B(DB[3102]), .Z(n14198) );
  XOR U38817 ( .A(n35896), .B(n14163), .Z(n14126) );
  XOR U38818 ( .A(n35897), .B(n14151), .Z(n14163) );
  XNOR U38819 ( .A(q[6]), .B(DB[3114]), .Z(n14151) );
  IV U38820 ( .A(n14150), .Z(n35897) );
  XNOR U38821 ( .A(n14148), .B(n35898), .Z(n14150) );
  XNOR U38822 ( .A(q[5]), .B(DB[3113]), .Z(n35898) );
  XNOR U38823 ( .A(q[4]), .B(DB[3112]), .Z(n14148) );
  IV U38824 ( .A(n14162), .Z(n35896) );
  XOR U38825 ( .A(n35899), .B(n35900), .Z(n14162) );
  XNOR U38826 ( .A(n14158), .B(n14160), .Z(n35900) );
  XNOR U38827 ( .A(q[0]), .B(DB[3108]), .Z(n14160) );
  XNOR U38828 ( .A(q[3]), .B(DB[3111]), .Z(n14158) );
  IV U38829 ( .A(n14157), .Z(n35899) );
  XNOR U38830 ( .A(n14155), .B(n35901), .Z(n14157) );
  XNOR U38831 ( .A(q[2]), .B(DB[3110]), .Z(n35901) );
  XNOR U38832 ( .A(q[1]), .B(DB[3109]), .Z(n14155) );
  XOR U38833 ( .A(n35902), .B(n14120), .Z(n14083) );
  XOR U38834 ( .A(n35903), .B(n14108), .Z(n14120) );
  XNOR U38835 ( .A(q[6]), .B(DB[3121]), .Z(n14108) );
  IV U38836 ( .A(n14107), .Z(n35903) );
  XNOR U38837 ( .A(n14105), .B(n35904), .Z(n14107) );
  XNOR U38838 ( .A(q[5]), .B(DB[3120]), .Z(n35904) );
  XNOR U38839 ( .A(q[4]), .B(DB[3119]), .Z(n14105) );
  IV U38840 ( .A(n14119), .Z(n35902) );
  XOR U38841 ( .A(n35905), .B(n35906), .Z(n14119) );
  XNOR U38842 ( .A(n14115), .B(n14117), .Z(n35906) );
  XNOR U38843 ( .A(q[0]), .B(DB[3115]), .Z(n14117) );
  XNOR U38844 ( .A(q[3]), .B(DB[3118]), .Z(n14115) );
  IV U38845 ( .A(n14114), .Z(n35905) );
  XNOR U38846 ( .A(n14112), .B(n35907), .Z(n14114) );
  XNOR U38847 ( .A(q[2]), .B(DB[3117]), .Z(n35907) );
  XNOR U38848 ( .A(q[1]), .B(DB[3116]), .Z(n14112) );
  XOR U38849 ( .A(n35908), .B(n14077), .Z(n14040) );
  XOR U38850 ( .A(n35909), .B(n14065), .Z(n14077) );
  XNOR U38851 ( .A(q[6]), .B(DB[3128]), .Z(n14065) );
  IV U38852 ( .A(n14064), .Z(n35909) );
  XNOR U38853 ( .A(n14062), .B(n35910), .Z(n14064) );
  XNOR U38854 ( .A(q[5]), .B(DB[3127]), .Z(n35910) );
  XNOR U38855 ( .A(q[4]), .B(DB[3126]), .Z(n14062) );
  IV U38856 ( .A(n14076), .Z(n35908) );
  XOR U38857 ( .A(n35911), .B(n35912), .Z(n14076) );
  XNOR U38858 ( .A(n14072), .B(n14074), .Z(n35912) );
  XNOR U38859 ( .A(q[0]), .B(DB[3122]), .Z(n14074) );
  XNOR U38860 ( .A(q[3]), .B(DB[3125]), .Z(n14072) );
  IV U38861 ( .A(n14071), .Z(n35911) );
  XNOR U38862 ( .A(n14069), .B(n35913), .Z(n14071) );
  XNOR U38863 ( .A(q[2]), .B(DB[3124]), .Z(n35913) );
  XNOR U38864 ( .A(q[1]), .B(DB[3123]), .Z(n14069) );
  XOR U38865 ( .A(n35914), .B(n14034), .Z(n13997) );
  XOR U38866 ( .A(n35915), .B(n14022), .Z(n14034) );
  XNOR U38867 ( .A(q[6]), .B(DB[3135]), .Z(n14022) );
  IV U38868 ( .A(n14021), .Z(n35915) );
  XNOR U38869 ( .A(n14019), .B(n35916), .Z(n14021) );
  XNOR U38870 ( .A(q[5]), .B(DB[3134]), .Z(n35916) );
  XNOR U38871 ( .A(q[4]), .B(DB[3133]), .Z(n14019) );
  IV U38872 ( .A(n14033), .Z(n35914) );
  XOR U38873 ( .A(n35917), .B(n35918), .Z(n14033) );
  XNOR U38874 ( .A(n14029), .B(n14031), .Z(n35918) );
  XNOR U38875 ( .A(q[0]), .B(DB[3129]), .Z(n14031) );
  XNOR U38876 ( .A(q[3]), .B(DB[3132]), .Z(n14029) );
  IV U38877 ( .A(n14028), .Z(n35917) );
  XNOR U38878 ( .A(n14026), .B(n35919), .Z(n14028) );
  XNOR U38879 ( .A(q[2]), .B(DB[3131]), .Z(n35919) );
  XNOR U38880 ( .A(q[1]), .B(DB[3130]), .Z(n14026) );
  XOR U38881 ( .A(n35920), .B(n13991), .Z(n13954) );
  XOR U38882 ( .A(n35921), .B(n13979), .Z(n13991) );
  XNOR U38883 ( .A(q[6]), .B(DB[3142]), .Z(n13979) );
  IV U38884 ( .A(n13978), .Z(n35921) );
  XNOR U38885 ( .A(n13976), .B(n35922), .Z(n13978) );
  XNOR U38886 ( .A(q[5]), .B(DB[3141]), .Z(n35922) );
  XNOR U38887 ( .A(q[4]), .B(DB[3140]), .Z(n13976) );
  IV U38888 ( .A(n13990), .Z(n35920) );
  XOR U38889 ( .A(n35923), .B(n35924), .Z(n13990) );
  XNOR U38890 ( .A(n13986), .B(n13988), .Z(n35924) );
  XNOR U38891 ( .A(q[0]), .B(DB[3136]), .Z(n13988) );
  XNOR U38892 ( .A(q[3]), .B(DB[3139]), .Z(n13986) );
  IV U38893 ( .A(n13985), .Z(n35923) );
  XNOR U38894 ( .A(n13983), .B(n35925), .Z(n13985) );
  XNOR U38895 ( .A(q[2]), .B(DB[3138]), .Z(n35925) );
  XNOR U38896 ( .A(q[1]), .B(DB[3137]), .Z(n13983) );
  XOR U38897 ( .A(n35926), .B(n13948), .Z(n13911) );
  XOR U38898 ( .A(n35927), .B(n13936), .Z(n13948) );
  XNOR U38899 ( .A(q[6]), .B(DB[3149]), .Z(n13936) );
  IV U38900 ( .A(n13935), .Z(n35927) );
  XNOR U38901 ( .A(n13933), .B(n35928), .Z(n13935) );
  XNOR U38902 ( .A(q[5]), .B(DB[3148]), .Z(n35928) );
  XNOR U38903 ( .A(q[4]), .B(DB[3147]), .Z(n13933) );
  IV U38904 ( .A(n13947), .Z(n35926) );
  XOR U38905 ( .A(n35929), .B(n35930), .Z(n13947) );
  XNOR U38906 ( .A(n13943), .B(n13945), .Z(n35930) );
  XNOR U38907 ( .A(q[0]), .B(DB[3143]), .Z(n13945) );
  XNOR U38908 ( .A(q[3]), .B(DB[3146]), .Z(n13943) );
  IV U38909 ( .A(n13942), .Z(n35929) );
  XNOR U38910 ( .A(n13940), .B(n35931), .Z(n13942) );
  XNOR U38911 ( .A(q[2]), .B(DB[3145]), .Z(n35931) );
  XNOR U38912 ( .A(q[1]), .B(DB[3144]), .Z(n13940) );
  XOR U38913 ( .A(n35932), .B(n13905), .Z(n13868) );
  XOR U38914 ( .A(n35933), .B(n13893), .Z(n13905) );
  XNOR U38915 ( .A(q[6]), .B(DB[3156]), .Z(n13893) );
  IV U38916 ( .A(n13892), .Z(n35933) );
  XNOR U38917 ( .A(n13890), .B(n35934), .Z(n13892) );
  XNOR U38918 ( .A(q[5]), .B(DB[3155]), .Z(n35934) );
  XNOR U38919 ( .A(q[4]), .B(DB[3154]), .Z(n13890) );
  IV U38920 ( .A(n13904), .Z(n35932) );
  XOR U38921 ( .A(n35935), .B(n35936), .Z(n13904) );
  XNOR U38922 ( .A(n13900), .B(n13902), .Z(n35936) );
  XNOR U38923 ( .A(q[0]), .B(DB[3150]), .Z(n13902) );
  XNOR U38924 ( .A(q[3]), .B(DB[3153]), .Z(n13900) );
  IV U38925 ( .A(n13899), .Z(n35935) );
  XNOR U38926 ( .A(n13897), .B(n35937), .Z(n13899) );
  XNOR U38927 ( .A(q[2]), .B(DB[3152]), .Z(n35937) );
  XNOR U38928 ( .A(q[1]), .B(DB[3151]), .Z(n13897) );
  XOR U38929 ( .A(n35938), .B(n13862), .Z(n13825) );
  XOR U38930 ( .A(n35939), .B(n13850), .Z(n13862) );
  XNOR U38931 ( .A(q[6]), .B(DB[3163]), .Z(n13850) );
  IV U38932 ( .A(n13849), .Z(n35939) );
  XNOR U38933 ( .A(n13847), .B(n35940), .Z(n13849) );
  XNOR U38934 ( .A(q[5]), .B(DB[3162]), .Z(n35940) );
  XNOR U38935 ( .A(q[4]), .B(DB[3161]), .Z(n13847) );
  IV U38936 ( .A(n13861), .Z(n35938) );
  XOR U38937 ( .A(n35941), .B(n35942), .Z(n13861) );
  XNOR U38938 ( .A(n13857), .B(n13859), .Z(n35942) );
  XNOR U38939 ( .A(q[0]), .B(DB[3157]), .Z(n13859) );
  XNOR U38940 ( .A(q[3]), .B(DB[3160]), .Z(n13857) );
  IV U38941 ( .A(n13856), .Z(n35941) );
  XNOR U38942 ( .A(n13854), .B(n35943), .Z(n13856) );
  XNOR U38943 ( .A(q[2]), .B(DB[3159]), .Z(n35943) );
  XNOR U38944 ( .A(q[1]), .B(DB[3158]), .Z(n13854) );
  XOR U38945 ( .A(n35944), .B(n13819), .Z(n13782) );
  XOR U38946 ( .A(n35945), .B(n13807), .Z(n13819) );
  XNOR U38947 ( .A(q[6]), .B(DB[3170]), .Z(n13807) );
  IV U38948 ( .A(n13806), .Z(n35945) );
  XNOR U38949 ( .A(n13804), .B(n35946), .Z(n13806) );
  XNOR U38950 ( .A(q[5]), .B(DB[3169]), .Z(n35946) );
  XNOR U38951 ( .A(q[4]), .B(DB[3168]), .Z(n13804) );
  IV U38952 ( .A(n13818), .Z(n35944) );
  XOR U38953 ( .A(n35947), .B(n35948), .Z(n13818) );
  XNOR U38954 ( .A(n13814), .B(n13816), .Z(n35948) );
  XNOR U38955 ( .A(q[0]), .B(DB[3164]), .Z(n13816) );
  XNOR U38956 ( .A(q[3]), .B(DB[3167]), .Z(n13814) );
  IV U38957 ( .A(n13813), .Z(n35947) );
  XNOR U38958 ( .A(n13811), .B(n35949), .Z(n13813) );
  XNOR U38959 ( .A(q[2]), .B(DB[3166]), .Z(n35949) );
  XNOR U38960 ( .A(q[1]), .B(DB[3165]), .Z(n13811) );
  XOR U38961 ( .A(n35950), .B(n13776), .Z(n13739) );
  XOR U38962 ( .A(n35951), .B(n13764), .Z(n13776) );
  XNOR U38963 ( .A(q[6]), .B(DB[3177]), .Z(n13764) );
  IV U38964 ( .A(n13763), .Z(n35951) );
  XNOR U38965 ( .A(n13761), .B(n35952), .Z(n13763) );
  XNOR U38966 ( .A(q[5]), .B(DB[3176]), .Z(n35952) );
  XNOR U38967 ( .A(q[4]), .B(DB[3175]), .Z(n13761) );
  IV U38968 ( .A(n13775), .Z(n35950) );
  XOR U38969 ( .A(n35953), .B(n35954), .Z(n13775) );
  XNOR U38970 ( .A(n13771), .B(n13773), .Z(n35954) );
  XNOR U38971 ( .A(q[0]), .B(DB[3171]), .Z(n13773) );
  XNOR U38972 ( .A(q[3]), .B(DB[3174]), .Z(n13771) );
  IV U38973 ( .A(n13770), .Z(n35953) );
  XNOR U38974 ( .A(n13768), .B(n35955), .Z(n13770) );
  XNOR U38975 ( .A(q[2]), .B(DB[3173]), .Z(n35955) );
  XNOR U38976 ( .A(q[1]), .B(DB[3172]), .Z(n13768) );
  XOR U38977 ( .A(n35956), .B(n13733), .Z(n13696) );
  XOR U38978 ( .A(n35957), .B(n13721), .Z(n13733) );
  XNOR U38979 ( .A(q[6]), .B(DB[3184]), .Z(n13721) );
  IV U38980 ( .A(n13720), .Z(n35957) );
  XNOR U38981 ( .A(n13718), .B(n35958), .Z(n13720) );
  XNOR U38982 ( .A(q[5]), .B(DB[3183]), .Z(n35958) );
  XNOR U38983 ( .A(q[4]), .B(DB[3182]), .Z(n13718) );
  IV U38984 ( .A(n13732), .Z(n35956) );
  XOR U38985 ( .A(n35959), .B(n35960), .Z(n13732) );
  XNOR U38986 ( .A(n13728), .B(n13730), .Z(n35960) );
  XNOR U38987 ( .A(q[0]), .B(DB[3178]), .Z(n13730) );
  XNOR U38988 ( .A(q[3]), .B(DB[3181]), .Z(n13728) );
  IV U38989 ( .A(n13727), .Z(n35959) );
  XNOR U38990 ( .A(n13725), .B(n35961), .Z(n13727) );
  XNOR U38991 ( .A(q[2]), .B(DB[3180]), .Z(n35961) );
  XNOR U38992 ( .A(q[1]), .B(DB[3179]), .Z(n13725) );
  XOR U38993 ( .A(n35962), .B(n13690), .Z(n13653) );
  XOR U38994 ( .A(n35963), .B(n13678), .Z(n13690) );
  XNOR U38995 ( .A(q[6]), .B(DB[3191]), .Z(n13678) );
  IV U38996 ( .A(n13677), .Z(n35963) );
  XNOR U38997 ( .A(n13675), .B(n35964), .Z(n13677) );
  XNOR U38998 ( .A(q[5]), .B(DB[3190]), .Z(n35964) );
  XNOR U38999 ( .A(q[4]), .B(DB[3189]), .Z(n13675) );
  IV U39000 ( .A(n13689), .Z(n35962) );
  XOR U39001 ( .A(n35965), .B(n35966), .Z(n13689) );
  XNOR U39002 ( .A(n13685), .B(n13687), .Z(n35966) );
  XNOR U39003 ( .A(q[0]), .B(DB[3185]), .Z(n13687) );
  XNOR U39004 ( .A(q[3]), .B(DB[3188]), .Z(n13685) );
  IV U39005 ( .A(n13684), .Z(n35965) );
  XNOR U39006 ( .A(n13682), .B(n35967), .Z(n13684) );
  XNOR U39007 ( .A(q[2]), .B(DB[3187]), .Z(n35967) );
  XNOR U39008 ( .A(q[1]), .B(DB[3186]), .Z(n13682) );
  XOR U39009 ( .A(n35968), .B(n13647), .Z(n13610) );
  XOR U39010 ( .A(n35969), .B(n13635), .Z(n13647) );
  XNOR U39011 ( .A(q[6]), .B(DB[3198]), .Z(n13635) );
  IV U39012 ( .A(n13634), .Z(n35969) );
  XNOR U39013 ( .A(n13632), .B(n35970), .Z(n13634) );
  XNOR U39014 ( .A(q[5]), .B(DB[3197]), .Z(n35970) );
  XNOR U39015 ( .A(q[4]), .B(DB[3196]), .Z(n13632) );
  IV U39016 ( .A(n13646), .Z(n35968) );
  XOR U39017 ( .A(n35971), .B(n35972), .Z(n13646) );
  XNOR U39018 ( .A(n13642), .B(n13644), .Z(n35972) );
  XNOR U39019 ( .A(q[0]), .B(DB[3192]), .Z(n13644) );
  XNOR U39020 ( .A(q[3]), .B(DB[3195]), .Z(n13642) );
  IV U39021 ( .A(n13641), .Z(n35971) );
  XNOR U39022 ( .A(n13639), .B(n35973), .Z(n13641) );
  XNOR U39023 ( .A(q[2]), .B(DB[3194]), .Z(n35973) );
  XNOR U39024 ( .A(q[1]), .B(DB[3193]), .Z(n13639) );
  XOR U39025 ( .A(n35974), .B(n13604), .Z(n13567) );
  XOR U39026 ( .A(n35975), .B(n13592), .Z(n13604) );
  XNOR U39027 ( .A(q[6]), .B(DB[3205]), .Z(n13592) );
  IV U39028 ( .A(n13591), .Z(n35975) );
  XNOR U39029 ( .A(n13589), .B(n35976), .Z(n13591) );
  XNOR U39030 ( .A(q[5]), .B(DB[3204]), .Z(n35976) );
  XNOR U39031 ( .A(q[4]), .B(DB[3203]), .Z(n13589) );
  IV U39032 ( .A(n13603), .Z(n35974) );
  XOR U39033 ( .A(n35977), .B(n35978), .Z(n13603) );
  XNOR U39034 ( .A(n13599), .B(n13601), .Z(n35978) );
  XNOR U39035 ( .A(q[0]), .B(DB[3199]), .Z(n13601) );
  XNOR U39036 ( .A(q[3]), .B(DB[3202]), .Z(n13599) );
  IV U39037 ( .A(n13598), .Z(n35977) );
  XNOR U39038 ( .A(n13596), .B(n35979), .Z(n13598) );
  XNOR U39039 ( .A(q[2]), .B(DB[3201]), .Z(n35979) );
  XNOR U39040 ( .A(q[1]), .B(DB[3200]), .Z(n13596) );
  XOR U39041 ( .A(n35980), .B(n13561), .Z(n13524) );
  XOR U39042 ( .A(n35981), .B(n13549), .Z(n13561) );
  XNOR U39043 ( .A(q[6]), .B(DB[3212]), .Z(n13549) );
  IV U39044 ( .A(n13548), .Z(n35981) );
  XNOR U39045 ( .A(n13546), .B(n35982), .Z(n13548) );
  XNOR U39046 ( .A(q[5]), .B(DB[3211]), .Z(n35982) );
  XNOR U39047 ( .A(q[4]), .B(DB[3210]), .Z(n13546) );
  IV U39048 ( .A(n13560), .Z(n35980) );
  XOR U39049 ( .A(n35983), .B(n35984), .Z(n13560) );
  XNOR U39050 ( .A(n13556), .B(n13558), .Z(n35984) );
  XNOR U39051 ( .A(q[0]), .B(DB[3206]), .Z(n13558) );
  XNOR U39052 ( .A(q[3]), .B(DB[3209]), .Z(n13556) );
  IV U39053 ( .A(n13555), .Z(n35983) );
  XNOR U39054 ( .A(n13553), .B(n35985), .Z(n13555) );
  XNOR U39055 ( .A(q[2]), .B(DB[3208]), .Z(n35985) );
  XNOR U39056 ( .A(q[1]), .B(DB[3207]), .Z(n13553) );
  XOR U39057 ( .A(n35986), .B(n13518), .Z(n13481) );
  XOR U39058 ( .A(n35987), .B(n13506), .Z(n13518) );
  XNOR U39059 ( .A(q[6]), .B(DB[3219]), .Z(n13506) );
  IV U39060 ( .A(n13505), .Z(n35987) );
  XNOR U39061 ( .A(n13503), .B(n35988), .Z(n13505) );
  XNOR U39062 ( .A(q[5]), .B(DB[3218]), .Z(n35988) );
  XNOR U39063 ( .A(q[4]), .B(DB[3217]), .Z(n13503) );
  IV U39064 ( .A(n13517), .Z(n35986) );
  XOR U39065 ( .A(n35989), .B(n35990), .Z(n13517) );
  XNOR U39066 ( .A(n13513), .B(n13515), .Z(n35990) );
  XNOR U39067 ( .A(q[0]), .B(DB[3213]), .Z(n13515) );
  XNOR U39068 ( .A(q[3]), .B(DB[3216]), .Z(n13513) );
  IV U39069 ( .A(n13512), .Z(n35989) );
  XNOR U39070 ( .A(n13510), .B(n35991), .Z(n13512) );
  XNOR U39071 ( .A(q[2]), .B(DB[3215]), .Z(n35991) );
  XNOR U39072 ( .A(q[1]), .B(DB[3214]), .Z(n13510) );
  XOR U39073 ( .A(n35992), .B(n13475), .Z(n13438) );
  XOR U39074 ( .A(n35993), .B(n13463), .Z(n13475) );
  XNOR U39075 ( .A(q[6]), .B(DB[3226]), .Z(n13463) );
  IV U39076 ( .A(n13462), .Z(n35993) );
  XNOR U39077 ( .A(n13460), .B(n35994), .Z(n13462) );
  XNOR U39078 ( .A(q[5]), .B(DB[3225]), .Z(n35994) );
  XNOR U39079 ( .A(q[4]), .B(DB[3224]), .Z(n13460) );
  IV U39080 ( .A(n13474), .Z(n35992) );
  XOR U39081 ( .A(n35995), .B(n35996), .Z(n13474) );
  XNOR U39082 ( .A(n13470), .B(n13472), .Z(n35996) );
  XNOR U39083 ( .A(q[0]), .B(DB[3220]), .Z(n13472) );
  XNOR U39084 ( .A(q[3]), .B(DB[3223]), .Z(n13470) );
  IV U39085 ( .A(n13469), .Z(n35995) );
  XNOR U39086 ( .A(n13467), .B(n35997), .Z(n13469) );
  XNOR U39087 ( .A(q[2]), .B(DB[3222]), .Z(n35997) );
  XNOR U39088 ( .A(q[1]), .B(DB[3221]), .Z(n13467) );
  XOR U39089 ( .A(n35998), .B(n13432), .Z(n13395) );
  XOR U39090 ( .A(n35999), .B(n13420), .Z(n13432) );
  XNOR U39091 ( .A(q[6]), .B(DB[3233]), .Z(n13420) );
  IV U39092 ( .A(n13419), .Z(n35999) );
  XNOR U39093 ( .A(n13417), .B(n36000), .Z(n13419) );
  XNOR U39094 ( .A(q[5]), .B(DB[3232]), .Z(n36000) );
  XNOR U39095 ( .A(q[4]), .B(DB[3231]), .Z(n13417) );
  IV U39096 ( .A(n13431), .Z(n35998) );
  XOR U39097 ( .A(n36001), .B(n36002), .Z(n13431) );
  XNOR U39098 ( .A(n13427), .B(n13429), .Z(n36002) );
  XNOR U39099 ( .A(q[0]), .B(DB[3227]), .Z(n13429) );
  XNOR U39100 ( .A(q[3]), .B(DB[3230]), .Z(n13427) );
  IV U39101 ( .A(n13426), .Z(n36001) );
  XNOR U39102 ( .A(n13424), .B(n36003), .Z(n13426) );
  XNOR U39103 ( .A(q[2]), .B(DB[3229]), .Z(n36003) );
  XNOR U39104 ( .A(q[1]), .B(DB[3228]), .Z(n13424) );
  XOR U39105 ( .A(n36004), .B(n13389), .Z(n13352) );
  XOR U39106 ( .A(n36005), .B(n13377), .Z(n13389) );
  XNOR U39107 ( .A(q[6]), .B(DB[3240]), .Z(n13377) );
  IV U39108 ( .A(n13376), .Z(n36005) );
  XNOR U39109 ( .A(n13374), .B(n36006), .Z(n13376) );
  XNOR U39110 ( .A(q[5]), .B(DB[3239]), .Z(n36006) );
  XNOR U39111 ( .A(q[4]), .B(DB[3238]), .Z(n13374) );
  IV U39112 ( .A(n13388), .Z(n36004) );
  XOR U39113 ( .A(n36007), .B(n36008), .Z(n13388) );
  XNOR U39114 ( .A(n13384), .B(n13386), .Z(n36008) );
  XNOR U39115 ( .A(q[0]), .B(DB[3234]), .Z(n13386) );
  XNOR U39116 ( .A(q[3]), .B(DB[3237]), .Z(n13384) );
  IV U39117 ( .A(n13383), .Z(n36007) );
  XNOR U39118 ( .A(n13381), .B(n36009), .Z(n13383) );
  XNOR U39119 ( .A(q[2]), .B(DB[3236]), .Z(n36009) );
  XNOR U39120 ( .A(q[1]), .B(DB[3235]), .Z(n13381) );
  XOR U39121 ( .A(n36010), .B(n13346), .Z(n13309) );
  XOR U39122 ( .A(n36011), .B(n13334), .Z(n13346) );
  XNOR U39123 ( .A(q[6]), .B(DB[3247]), .Z(n13334) );
  IV U39124 ( .A(n13333), .Z(n36011) );
  XNOR U39125 ( .A(n13331), .B(n36012), .Z(n13333) );
  XNOR U39126 ( .A(q[5]), .B(DB[3246]), .Z(n36012) );
  XNOR U39127 ( .A(q[4]), .B(DB[3245]), .Z(n13331) );
  IV U39128 ( .A(n13345), .Z(n36010) );
  XOR U39129 ( .A(n36013), .B(n36014), .Z(n13345) );
  XNOR U39130 ( .A(n13341), .B(n13343), .Z(n36014) );
  XNOR U39131 ( .A(q[0]), .B(DB[3241]), .Z(n13343) );
  XNOR U39132 ( .A(q[3]), .B(DB[3244]), .Z(n13341) );
  IV U39133 ( .A(n13340), .Z(n36013) );
  XNOR U39134 ( .A(n13338), .B(n36015), .Z(n13340) );
  XNOR U39135 ( .A(q[2]), .B(DB[3243]), .Z(n36015) );
  XNOR U39136 ( .A(q[1]), .B(DB[3242]), .Z(n13338) );
  XOR U39137 ( .A(n36016), .B(n13303), .Z(n13266) );
  XOR U39138 ( .A(n36017), .B(n13291), .Z(n13303) );
  XNOR U39139 ( .A(q[6]), .B(DB[3254]), .Z(n13291) );
  IV U39140 ( .A(n13290), .Z(n36017) );
  XNOR U39141 ( .A(n13288), .B(n36018), .Z(n13290) );
  XNOR U39142 ( .A(q[5]), .B(DB[3253]), .Z(n36018) );
  XNOR U39143 ( .A(q[4]), .B(DB[3252]), .Z(n13288) );
  IV U39144 ( .A(n13302), .Z(n36016) );
  XOR U39145 ( .A(n36019), .B(n36020), .Z(n13302) );
  XNOR U39146 ( .A(n13298), .B(n13300), .Z(n36020) );
  XNOR U39147 ( .A(q[0]), .B(DB[3248]), .Z(n13300) );
  XNOR U39148 ( .A(q[3]), .B(DB[3251]), .Z(n13298) );
  IV U39149 ( .A(n13297), .Z(n36019) );
  XNOR U39150 ( .A(n13295), .B(n36021), .Z(n13297) );
  XNOR U39151 ( .A(q[2]), .B(DB[3250]), .Z(n36021) );
  XNOR U39152 ( .A(q[1]), .B(DB[3249]), .Z(n13295) );
  XOR U39153 ( .A(n36022), .B(n13260), .Z(n13223) );
  XOR U39154 ( .A(n36023), .B(n13248), .Z(n13260) );
  XNOR U39155 ( .A(q[6]), .B(DB[3261]), .Z(n13248) );
  IV U39156 ( .A(n13247), .Z(n36023) );
  XNOR U39157 ( .A(n13245), .B(n36024), .Z(n13247) );
  XNOR U39158 ( .A(q[5]), .B(DB[3260]), .Z(n36024) );
  XNOR U39159 ( .A(q[4]), .B(DB[3259]), .Z(n13245) );
  IV U39160 ( .A(n13259), .Z(n36022) );
  XOR U39161 ( .A(n36025), .B(n36026), .Z(n13259) );
  XNOR U39162 ( .A(n13255), .B(n13257), .Z(n36026) );
  XNOR U39163 ( .A(q[0]), .B(DB[3255]), .Z(n13257) );
  XNOR U39164 ( .A(q[3]), .B(DB[3258]), .Z(n13255) );
  IV U39165 ( .A(n13254), .Z(n36025) );
  XNOR U39166 ( .A(n13252), .B(n36027), .Z(n13254) );
  XNOR U39167 ( .A(q[2]), .B(DB[3257]), .Z(n36027) );
  XNOR U39168 ( .A(q[1]), .B(DB[3256]), .Z(n13252) );
  XOR U39169 ( .A(n36028), .B(n13217), .Z(n13180) );
  XOR U39170 ( .A(n36029), .B(n13205), .Z(n13217) );
  XNOR U39171 ( .A(q[6]), .B(DB[3268]), .Z(n13205) );
  IV U39172 ( .A(n13204), .Z(n36029) );
  XNOR U39173 ( .A(n13202), .B(n36030), .Z(n13204) );
  XNOR U39174 ( .A(q[5]), .B(DB[3267]), .Z(n36030) );
  XNOR U39175 ( .A(q[4]), .B(DB[3266]), .Z(n13202) );
  IV U39176 ( .A(n13216), .Z(n36028) );
  XOR U39177 ( .A(n36031), .B(n36032), .Z(n13216) );
  XNOR U39178 ( .A(n13212), .B(n13214), .Z(n36032) );
  XNOR U39179 ( .A(q[0]), .B(DB[3262]), .Z(n13214) );
  XNOR U39180 ( .A(q[3]), .B(DB[3265]), .Z(n13212) );
  IV U39181 ( .A(n13211), .Z(n36031) );
  XNOR U39182 ( .A(n13209), .B(n36033), .Z(n13211) );
  XNOR U39183 ( .A(q[2]), .B(DB[3264]), .Z(n36033) );
  XNOR U39184 ( .A(q[1]), .B(DB[3263]), .Z(n13209) );
  XOR U39185 ( .A(n36034), .B(n13174), .Z(n13137) );
  XOR U39186 ( .A(n36035), .B(n13162), .Z(n13174) );
  XNOR U39187 ( .A(q[6]), .B(DB[3275]), .Z(n13162) );
  IV U39188 ( .A(n13161), .Z(n36035) );
  XNOR U39189 ( .A(n13159), .B(n36036), .Z(n13161) );
  XNOR U39190 ( .A(q[5]), .B(DB[3274]), .Z(n36036) );
  XNOR U39191 ( .A(q[4]), .B(DB[3273]), .Z(n13159) );
  IV U39192 ( .A(n13173), .Z(n36034) );
  XOR U39193 ( .A(n36037), .B(n36038), .Z(n13173) );
  XNOR U39194 ( .A(n13169), .B(n13171), .Z(n36038) );
  XNOR U39195 ( .A(q[0]), .B(DB[3269]), .Z(n13171) );
  XNOR U39196 ( .A(q[3]), .B(DB[3272]), .Z(n13169) );
  IV U39197 ( .A(n13168), .Z(n36037) );
  XNOR U39198 ( .A(n13166), .B(n36039), .Z(n13168) );
  XNOR U39199 ( .A(q[2]), .B(DB[3271]), .Z(n36039) );
  XNOR U39200 ( .A(q[1]), .B(DB[3270]), .Z(n13166) );
  XOR U39201 ( .A(n36040), .B(n13131), .Z(n13094) );
  XOR U39202 ( .A(n36041), .B(n13119), .Z(n13131) );
  XNOR U39203 ( .A(q[6]), .B(DB[3282]), .Z(n13119) );
  IV U39204 ( .A(n13118), .Z(n36041) );
  XNOR U39205 ( .A(n13116), .B(n36042), .Z(n13118) );
  XNOR U39206 ( .A(q[5]), .B(DB[3281]), .Z(n36042) );
  XNOR U39207 ( .A(q[4]), .B(DB[3280]), .Z(n13116) );
  IV U39208 ( .A(n13130), .Z(n36040) );
  XOR U39209 ( .A(n36043), .B(n36044), .Z(n13130) );
  XNOR U39210 ( .A(n13126), .B(n13128), .Z(n36044) );
  XNOR U39211 ( .A(q[0]), .B(DB[3276]), .Z(n13128) );
  XNOR U39212 ( .A(q[3]), .B(DB[3279]), .Z(n13126) );
  IV U39213 ( .A(n13125), .Z(n36043) );
  XNOR U39214 ( .A(n13123), .B(n36045), .Z(n13125) );
  XNOR U39215 ( .A(q[2]), .B(DB[3278]), .Z(n36045) );
  XNOR U39216 ( .A(q[1]), .B(DB[3277]), .Z(n13123) );
  XOR U39217 ( .A(n36046), .B(n13088), .Z(n13051) );
  XOR U39218 ( .A(n36047), .B(n13076), .Z(n13088) );
  XNOR U39219 ( .A(q[6]), .B(DB[3289]), .Z(n13076) );
  IV U39220 ( .A(n13075), .Z(n36047) );
  XNOR U39221 ( .A(n13073), .B(n36048), .Z(n13075) );
  XNOR U39222 ( .A(q[5]), .B(DB[3288]), .Z(n36048) );
  XNOR U39223 ( .A(q[4]), .B(DB[3287]), .Z(n13073) );
  IV U39224 ( .A(n13087), .Z(n36046) );
  XOR U39225 ( .A(n36049), .B(n36050), .Z(n13087) );
  XNOR U39226 ( .A(n13083), .B(n13085), .Z(n36050) );
  XNOR U39227 ( .A(q[0]), .B(DB[3283]), .Z(n13085) );
  XNOR U39228 ( .A(q[3]), .B(DB[3286]), .Z(n13083) );
  IV U39229 ( .A(n13082), .Z(n36049) );
  XNOR U39230 ( .A(n13080), .B(n36051), .Z(n13082) );
  XNOR U39231 ( .A(q[2]), .B(DB[3285]), .Z(n36051) );
  XNOR U39232 ( .A(q[1]), .B(DB[3284]), .Z(n13080) );
  XOR U39233 ( .A(n36052), .B(n13045), .Z(n13008) );
  XOR U39234 ( .A(n36053), .B(n13033), .Z(n13045) );
  XNOR U39235 ( .A(q[6]), .B(DB[3296]), .Z(n13033) );
  IV U39236 ( .A(n13032), .Z(n36053) );
  XNOR U39237 ( .A(n13030), .B(n36054), .Z(n13032) );
  XNOR U39238 ( .A(q[5]), .B(DB[3295]), .Z(n36054) );
  XNOR U39239 ( .A(q[4]), .B(DB[3294]), .Z(n13030) );
  IV U39240 ( .A(n13044), .Z(n36052) );
  XOR U39241 ( .A(n36055), .B(n36056), .Z(n13044) );
  XNOR U39242 ( .A(n13040), .B(n13042), .Z(n36056) );
  XNOR U39243 ( .A(q[0]), .B(DB[3290]), .Z(n13042) );
  XNOR U39244 ( .A(q[3]), .B(DB[3293]), .Z(n13040) );
  IV U39245 ( .A(n13039), .Z(n36055) );
  XNOR U39246 ( .A(n13037), .B(n36057), .Z(n13039) );
  XNOR U39247 ( .A(q[2]), .B(DB[3292]), .Z(n36057) );
  XNOR U39248 ( .A(q[1]), .B(DB[3291]), .Z(n13037) );
  XOR U39249 ( .A(n36058), .B(n13002), .Z(n12965) );
  XOR U39250 ( .A(n36059), .B(n12990), .Z(n13002) );
  XNOR U39251 ( .A(q[6]), .B(DB[3303]), .Z(n12990) );
  IV U39252 ( .A(n12989), .Z(n36059) );
  XNOR U39253 ( .A(n12987), .B(n36060), .Z(n12989) );
  XNOR U39254 ( .A(q[5]), .B(DB[3302]), .Z(n36060) );
  XNOR U39255 ( .A(q[4]), .B(DB[3301]), .Z(n12987) );
  IV U39256 ( .A(n13001), .Z(n36058) );
  XOR U39257 ( .A(n36061), .B(n36062), .Z(n13001) );
  XNOR U39258 ( .A(n12997), .B(n12999), .Z(n36062) );
  XNOR U39259 ( .A(q[0]), .B(DB[3297]), .Z(n12999) );
  XNOR U39260 ( .A(q[3]), .B(DB[3300]), .Z(n12997) );
  IV U39261 ( .A(n12996), .Z(n36061) );
  XNOR U39262 ( .A(n12994), .B(n36063), .Z(n12996) );
  XNOR U39263 ( .A(q[2]), .B(DB[3299]), .Z(n36063) );
  XNOR U39264 ( .A(q[1]), .B(DB[3298]), .Z(n12994) );
  XOR U39265 ( .A(n36064), .B(n12959), .Z(n12922) );
  XOR U39266 ( .A(n36065), .B(n12947), .Z(n12959) );
  XNOR U39267 ( .A(q[6]), .B(DB[3310]), .Z(n12947) );
  IV U39268 ( .A(n12946), .Z(n36065) );
  XNOR U39269 ( .A(n12944), .B(n36066), .Z(n12946) );
  XNOR U39270 ( .A(q[5]), .B(DB[3309]), .Z(n36066) );
  XNOR U39271 ( .A(q[4]), .B(DB[3308]), .Z(n12944) );
  IV U39272 ( .A(n12958), .Z(n36064) );
  XOR U39273 ( .A(n36067), .B(n36068), .Z(n12958) );
  XNOR U39274 ( .A(n12954), .B(n12956), .Z(n36068) );
  XNOR U39275 ( .A(q[0]), .B(DB[3304]), .Z(n12956) );
  XNOR U39276 ( .A(q[3]), .B(DB[3307]), .Z(n12954) );
  IV U39277 ( .A(n12953), .Z(n36067) );
  XNOR U39278 ( .A(n12951), .B(n36069), .Z(n12953) );
  XNOR U39279 ( .A(q[2]), .B(DB[3306]), .Z(n36069) );
  XNOR U39280 ( .A(q[1]), .B(DB[3305]), .Z(n12951) );
  XOR U39281 ( .A(n36070), .B(n12916), .Z(n12879) );
  XOR U39282 ( .A(n36071), .B(n12904), .Z(n12916) );
  XNOR U39283 ( .A(q[6]), .B(DB[3317]), .Z(n12904) );
  IV U39284 ( .A(n12903), .Z(n36071) );
  XNOR U39285 ( .A(n12901), .B(n36072), .Z(n12903) );
  XNOR U39286 ( .A(q[5]), .B(DB[3316]), .Z(n36072) );
  XNOR U39287 ( .A(q[4]), .B(DB[3315]), .Z(n12901) );
  IV U39288 ( .A(n12915), .Z(n36070) );
  XOR U39289 ( .A(n36073), .B(n36074), .Z(n12915) );
  XNOR U39290 ( .A(n12911), .B(n12913), .Z(n36074) );
  XNOR U39291 ( .A(q[0]), .B(DB[3311]), .Z(n12913) );
  XNOR U39292 ( .A(q[3]), .B(DB[3314]), .Z(n12911) );
  IV U39293 ( .A(n12910), .Z(n36073) );
  XNOR U39294 ( .A(n12908), .B(n36075), .Z(n12910) );
  XNOR U39295 ( .A(q[2]), .B(DB[3313]), .Z(n36075) );
  XNOR U39296 ( .A(q[1]), .B(DB[3312]), .Z(n12908) );
  XOR U39297 ( .A(n36076), .B(n12873), .Z(n12836) );
  XOR U39298 ( .A(n36077), .B(n12861), .Z(n12873) );
  XNOR U39299 ( .A(q[6]), .B(DB[3324]), .Z(n12861) );
  IV U39300 ( .A(n12860), .Z(n36077) );
  XNOR U39301 ( .A(n12858), .B(n36078), .Z(n12860) );
  XNOR U39302 ( .A(q[5]), .B(DB[3323]), .Z(n36078) );
  XNOR U39303 ( .A(q[4]), .B(DB[3322]), .Z(n12858) );
  IV U39304 ( .A(n12872), .Z(n36076) );
  XOR U39305 ( .A(n36079), .B(n36080), .Z(n12872) );
  XNOR U39306 ( .A(n12868), .B(n12870), .Z(n36080) );
  XNOR U39307 ( .A(q[0]), .B(DB[3318]), .Z(n12870) );
  XNOR U39308 ( .A(q[3]), .B(DB[3321]), .Z(n12868) );
  IV U39309 ( .A(n12867), .Z(n36079) );
  XNOR U39310 ( .A(n12865), .B(n36081), .Z(n12867) );
  XNOR U39311 ( .A(q[2]), .B(DB[3320]), .Z(n36081) );
  XNOR U39312 ( .A(q[1]), .B(DB[3319]), .Z(n12865) );
  XOR U39313 ( .A(n36082), .B(n12830), .Z(n12793) );
  XOR U39314 ( .A(n36083), .B(n12818), .Z(n12830) );
  XNOR U39315 ( .A(q[6]), .B(DB[3331]), .Z(n12818) );
  IV U39316 ( .A(n12817), .Z(n36083) );
  XNOR U39317 ( .A(n12815), .B(n36084), .Z(n12817) );
  XNOR U39318 ( .A(q[5]), .B(DB[3330]), .Z(n36084) );
  XNOR U39319 ( .A(q[4]), .B(DB[3329]), .Z(n12815) );
  IV U39320 ( .A(n12829), .Z(n36082) );
  XOR U39321 ( .A(n36085), .B(n36086), .Z(n12829) );
  XNOR U39322 ( .A(n12825), .B(n12827), .Z(n36086) );
  XNOR U39323 ( .A(q[0]), .B(DB[3325]), .Z(n12827) );
  XNOR U39324 ( .A(q[3]), .B(DB[3328]), .Z(n12825) );
  IV U39325 ( .A(n12824), .Z(n36085) );
  XNOR U39326 ( .A(n12822), .B(n36087), .Z(n12824) );
  XNOR U39327 ( .A(q[2]), .B(DB[3327]), .Z(n36087) );
  XNOR U39328 ( .A(q[1]), .B(DB[3326]), .Z(n12822) );
  XOR U39329 ( .A(n36088), .B(n12787), .Z(n12750) );
  XOR U39330 ( .A(n36089), .B(n12775), .Z(n12787) );
  XNOR U39331 ( .A(q[6]), .B(DB[3338]), .Z(n12775) );
  IV U39332 ( .A(n12774), .Z(n36089) );
  XNOR U39333 ( .A(n12772), .B(n36090), .Z(n12774) );
  XNOR U39334 ( .A(q[5]), .B(DB[3337]), .Z(n36090) );
  XNOR U39335 ( .A(q[4]), .B(DB[3336]), .Z(n12772) );
  IV U39336 ( .A(n12786), .Z(n36088) );
  XOR U39337 ( .A(n36091), .B(n36092), .Z(n12786) );
  XNOR U39338 ( .A(n12782), .B(n12784), .Z(n36092) );
  XNOR U39339 ( .A(q[0]), .B(DB[3332]), .Z(n12784) );
  XNOR U39340 ( .A(q[3]), .B(DB[3335]), .Z(n12782) );
  IV U39341 ( .A(n12781), .Z(n36091) );
  XNOR U39342 ( .A(n12779), .B(n36093), .Z(n12781) );
  XNOR U39343 ( .A(q[2]), .B(DB[3334]), .Z(n36093) );
  XNOR U39344 ( .A(q[1]), .B(DB[3333]), .Z(n12779) );
  XOR U39345 ( .A(n36094), .B(n12744), .Z(n12707) );
  XOR U39346 ( .A(n36095), .B(n12732), .Z(n12744) );
  XNOR U39347 ( .A(q[6]), .B(DB[3345]), .Z(n12732) );
  IV U39348 ( .A(n12731), .Z(n36095) );
  XNOR U39349 ( .A(n12729), .B(n36096), .Z(n12731) );
  XNOR U39350 ( .A(q[5]), .B(DB[3344]), .Z(n36096) );
  XNOR U39351 ( .A(q[4]), .B(DB[3343]), .Z(n12729) );
  IV U39352 ( .A(n12743), .Z(n36094) );
  XOR U39353 ( .A(n36097), .B(n36098), .Z(n12743) );
  XNOR U39354 ( .A(n12739), .B(n12741), .Z(n36098) );
  XNOR U39355 ( .A(q[0]), .B(DB[3339]), .Z(n12741) );
  XNOR U39356 ( .A(q[3]), .B(DB[3342]), .Z(n12739) );
  IV U39357 ( .A(n12738), .Z(n36097) );
  XNOR U39358 ( .A(n12736), .B(n36099), .Z(n12738) );
  XNOR U39359 ( .A(q[2]), .B(DB[3341]), .Z(n36099) );
  XNOR U39360 ( .A(q[1]), .B(DB[3340]), .Z(n12736) );
  XOR U39361 ( .A(n36100), .B(n12701), .Z(n12664) );
  XOR U39362 ( .A(n36101), .B(n12689), .Z(n12701) );
  XNOR U39363 ( .A(q[6]), .B(DB[3352]), .Z(n12689) );
  IV U39364 ( .A(n12688), .Z(n36101) );
  XNOR U39365 ( .A(n12686), .B(n36102), .Z(n12688) );
  XNOR U39366 ( .A(q[5]), .B(DB[3351]), .Z(n36102) );
  XNOR U39367 ( .A(q[4]), .B(DB[3350]), .Z(n12686) );
  IV U39368 ( .A(n12700), .Z(n36100) );
  XOR U39369 ( .A(n36103), .B(n36104), .Z(n12700) );
  XNOR U39370 ( .A(n12696), .B(n12698), .Z(n36104) );
  XNOR U39371 ( .A(q[0]), .B(DB[3346]), .Z(n12698) );
  XNOR U39372 ( .A(q[3]), .B(DB[3349]), .Z(n12696) );
  IV U39373 ( .A(n12695), .Z(n36103) );
  XNOR U39374 ( .A(n12693), .B(n36105), .Z(n12695) );
  XNOR U39375 ( .A(q[2]), .B(DB[3348]), .Z(n36105) );
  XNOR U39376 ( .A(q[1]), .B(DB[3347]), .Z(n12693) );
  XOR U39377 ( .A(n36106), .B(n12658), .Z(n12621) );
  XOR U39378 ( .A(n36107), .B(n12646), .Z(n12658) );
  XNOR U39379 ( .A(q[6]), .B(DB[3359]), .Z(n12646) );
  IV U39380 ( .A(n12645), .Z(n36107) );
  XNOR U39381 ( .A(n12643), .B(n36108), .Z(n12645) );
  XNOR U39382 ( .A(q[5]), .B(DB[3358]), .Z(n36108) );
  XNOR U39383 ( .A(q[4]), .B(DB[3357]), .Z(n12643) );
  IV U39384 ( .A(n12657), .Z(n36106) );
  XOR U39385 ( .A(n36109), .B(n36110), .Z(n12657) );
  XNOR U39386 ( .A(n12653), .B(n12655), .Z(n36110) );
  XNOR U39387 ( .A(q[0]), .B(DB[3353]), .Z(n12655) );
  XNOR U39388 ( .A(q[3]), .B(DB[3356]), .Z(n12653) );
  IV U39389 ( .A(n12652), .Z(n36109) );
  XNOR U39390 ( .A(n12650), .B(n36111), .Z(n12652) );
  XNOR U39391 ( .A(q[2]), .B(DB[3355]), .Z(n36111) );
  XNOR U39392 ( .A(q[1]), .B(DB[3354]), .Z(n12650) );
  XOR U39393 ( .A(n36112), .B(n12615), .Z(n12578) );
  XOR U39394 ( .A(n36113), .B(n12603), .Z(n12615) );
  XNOR U39395 ( .A(q[6]), .B(DB[3366]), .Z(n12603) );
  IV U39396 ( .A(n12602), .Z(n36113) );
  XNOR U39397 ( .A(n12600), .B(n36114), .Z(n12602) );
  XNOR U39398 ( .A(q[5]), .B(DB[3365]), .Z(n36114) );
  XNOR U39399 ( .A(q[4]), .B(DB[3364]), .Z(n12600) );
  IV U39400 ( .A(n12614), .Z(n36112) );
  XOR U39401 ( .A(n36115), .B(n36116), .Z(n12614) );
  XNOR U39402 ( .A(n12610), .B(n12612), .Z(n36116) );
  XNOR U39403 ( .A(q[0]), .B(DB[3360]), .Z(n12612) );
  XNOR U39404 ( .A(q[3]), .B(DB[3363]), .Z(n12610) );
  IV U39405 ( .A(n12609), .Z(n36115) );
  XNOR U39406 ( .A(n12607), .B(n36117), .Z(n12609) );
  XNOR U39407 ( .A(q[2]), .B(DB[3362]), .Z(n36117) );
  XNOR U39408 ( .A(q[1]), .B(DB[3361]), .Z(n12607) );
  XOR U39409 ( .A(n36118), .B(n12572), .Z(n12535) );
  XOR U39410 ( .A(n36119), .B(n12560), .Z(n12572) );
  XNOR U39411 ( .A(q[6]), .B(DB[3373]), .Z(n12560) );
  IV U39412 ( .A(n12559), .Z(n36119) );
  XNOR U39413 ( .A(n12557), .B(n36120), .Z(n12559) );
  XNOR U39414 ( .A(q[5]), .B(DB[3372]), .Z(n36120) );
  XNOR U39415 ( .A(q[4]), .B(DB[3371]), .Z(n12557) );
  IV U39416 ( .A(n12571), .Z(n36118) );
  XOR U39417 ( .A(n36121), .B(n36122), .Z(n12571) );
  XNOR U39418 ( .A(n12567), .B(n12569), .Z(n36122) );
  XNOR U39419 ( .A(q[0]), .B(DB[3367]), .Z(n12569) );
  XNOR U39420 ( .A(q[3]), .B(DB[3370]), .Z(n12567) );
  IV U39421 ( .A(n12566), .Z(n36121) );
  XNOR U39422 ( .A(n12564), .B(n36123), .Z(n12566) );
  XNOR U39423 ( .A(q[2]), .B(DB[3369]), .Z(n36123) );
  XNOR U39424 ( .A(q[1]), .B(DB[3368]), .Z(n12564) );
  XOR U39425 ( .A(n36124), .B(n12529), .Z(n12492) );
  XOR U39426 ( .A(n36125), .B(n12517), .Z(n12529) );
  XNOR U39427 ( .A(q[6]), .B(DB[3380]), .Z(n12517) );
  IV U39428 ( .A(n12516), .Z(n36125) );
  XNOR U39429 ( .A(n12514), .B(n36126), .Z(n12516) );
  XNOR U39430 ( .A(q[5]), .B(DB[3379]), .Z(n36126) );
  XNOR U39431 ( .A(q[4]), .B(DB[3378]), .Z(n12514) );
  IV U39432 ( .A(n12528), .Z(n36124) );
  XOR U39433 ( .A(n36127), .B(n36128), .Z(n12528) );
  XNOR U39434 ( .A(n12524), .B(n12526), .Z(n36128) );
  XNOR U39435 ( .A(q[0]), .B(DB[3374]), .Z(n12526) );
  XNOR U39436 ( .A(q[3]), .B(DB[3377]), .Z(n12524) );
  IV U39437 ( .A(n12523), .Z(n36127) );
  XNOR U39438 ( .A(n12521), .B(n36129), .Z(n12523) );
  XNOR U39439 ( .A(q[2]), .B(DB[3376]), .Z(n36129) );
  XNOR U39440 ( .A(q[1]), .B(DB[3375]), .Z(n12521) );
  XOR U39441 ( .A(n36130), .B(n12486), .Z(n12449) );
  XOR U39442 ( .A(n36131), .B(n12474), .Z(n12486) );
  XNOR U39443 ( .A(q[6]), .B(DB[3387]), .Z(n12474) );
  IV U39444 ( .A(n12473), .Z(n36131) );
  XNOR U39445 ( .A(n12471), .B(n36132), .Z(n12473) );
  XNOR U39446 ( .A(q[5]), .B(DB[3386]), .Z(n36132) );
  XNOR U39447 ( .A(q[4]), .B(DB[3385]), .Z(n12471) );
  IV U39448 ( .A(n12485), .Z(n36130) );
  XOR U39449 ( .A(n36133), .B(n36134), .Z(n12485) );
  XNOR U39450 ( .A(n12481), .B(n12483), .Z(n36134) );
  XNOR U39451 ( .A(q[0]), .B(DB[3381]), .Z(n12483) );
  XNOR U39452 ( .A(q[3]), .B(DB[3384]), .Z(n12481) );
  IV U39453 ( .A(n12480), .Z(n36133) );
  XNOR U39454 ( .A(n12478), .B(n36135), .Z(n12480) );
  XNOR U39455 ( .A(q[2]), .B(DB[3383]), .Z(n36135) );
  XNOR U39456 ( .A(q[1]), .B(DB[3382]), .Z(n12478) );
  XOR U39457 ( .A(n36136), .B(n12443), .Z(n12406) );
  XOR U39458 ( .A(n36137), .B(n12431), .Z(n12443) );
  XNOR U39459 ( .A(q[6]), .B(DB[3394]), .Z(n12431) );
  IV U39460 ( .A(n12430), .Z(n36137) );
  XNOR U39461 ( .A(n12428), .B(n36138), .Z(n12430) );
  XNOR U39462 ( .A(q[5]), .B(DB[3393]), .Z(n36138) );
  XNOR U39463 ( .A(q[4]), .B(DB[3392]), .Z(n12428) );
  IV U39464 ( .A(n12442), .Z(n36136) );
  XOR U39465 ( .A(n36139), .B(n36140), .Z(n12442) );
  XNOR U39466 ( .A(n12438), .B(n12440), .Z(n36140) );
  XNOR U39467 ( .A(q[0]), .B(DB[3388]), .Z(n12440) );
  XNOR U39468 ( .A(q[3]), .B(DB[3391]), .Z(n12438) );
  IV U39469 ( .A(n12437), .Z(n36139) );
  XNOR U39470 ( .A(n12435), .B(n36141), .Z(n12437) );
  XNOR U39471 ( .A(q[2]), .B(DB[3390]), .Z(n36141) );
  XNOR U39472 ( .A(q[1]), .B(DB[3389]), .Z(n12435) );
  XOR U39473 ( .A(n36142), .B(n12400), .Z(n12363) );
  XOR U39474 ( .A(n36143), .B(n12388), .Z(n12400) );
  XNOR U39475 ( .A(q[6]), .B(DB[3401]), .Z(n12388) );
  IV U39476 ( .A(n12387), .Z(n36143) );
  XNOR U39477 ( .A(n12385), .B(n36144), .Z(n12387) );
  XNOR U39478 ( .A(q[5]), .B(DB[3400]), .Z(n36144) );
  XNOR U39479 ( .A(q[4]), .B(DB[3399]), .Z(n12385) );
  IV U39480 ( .A(n12399), .Z(n36142) );
  XOR U39481 ( .A(n36145), .B(n36146), .Z(n12399) );
  XNOR U39482 ( .A(n12395), .B(n12397), .Z(n36146) );
  XNOR U39483 ( .A(q[0]), .B(DB[3395]), .Z(n12397) );
  XNOR U39484 ( .A(q[3]), .B(DB[3398]), .Z(n12395) );
  IV U39485 ( .A(n12394), .Z(n36145) );
  XNOR U39486 ( .A(n12392), .B(n36147), .Z(n12394) );
  XNOR U39487 ( .A(q[2]), .B(DB[3397]), .Z(n36147) );
  XNOR U39488 ( .A(q[1]), .B(DB[3396]), .Z(n12392) );
  XOR U39489 ( .A(n36148), .B(n12357), .Z(n12320) );
  XOR U39490 ( .A(n36149), .B(n12345), .Z(n12357) );
  XNOR U39491 ( .A(q[6]), .B(DB[3408]), .Z(n12345) );
  IV U39492 ( .A(n12344), .Z(n36149) );
  XNOR U39493 ( .A(n12342), .B(n36150), .Z(n12344) );
  XNOR U39494 ( .A(q[5]), .B(DB[3407]), .Z(n36150) );
  XNOR U39495 ( .A(q[4]), .B(DB[3406]), .Z(n12342) );
  IV U39496 ( .A(n12356), .Z(n36148) );
  XOR U39497 ( .A(n36151), .B(n36152), .Z(n12356) );
  XNOR U39498 ( .A(n12352), .B(n12354), .Z(n36152) );
  XNOR U39499 ( .A(q[0]), .B(DB[3402]), .Z(n12354) );
  XNOR U39500 ( .A(q[3]), .B(DB[3405]), .Z(n12352) );
  IV U39501 ( .A(n12351), .Z(n36151) );
  XNOR U39502 ( .A(n12349), .B(n36153), .Z(n12351) );
  XNOR U39503 ( .A(q[2]), .B(DB[3404]), .Z(n36153) );
  XNOR U39504 ( .A(q[1]), .B(DB[3403]), .Z(n12349) );
  XOR U39505 ( .A(n36154), .B(n12314), .Z(n12277) );
  XOR U39506 ( .A(n36155), .B(n12302), .Z(n12314) );
  XNOR U39507 ( .A(q[6]), .B(DB[3415]), .Z(n12302) );
  IV U39508 ( .A(n12301), .Z(n36155) );
  XNOR U39509 ( .A(n12299), .B(n36156), .Z(n12301) );
  XNOR U39510 ( .A(q[5]), .B(DB[3414]), .Z(n36156) );
  XNOR U39511 ( .A(q[4]), .B(DB[3413]), .Z(n12299) );
  IV U39512 ( .A(n12313), .Z(n36154) );
  XOR U39513 ( .A(n36157), .B(n36158), .Z(n12313) );
  XNOR U39514 ( .A(n12309), .B(n12311), .Z(n36158) );
  XNOR U39515 ( .A(q[0]), .B(DB[3409]), .Z(n12311) );
  XNOR U39516 ( .A(q[3]), .B(DB[3412]), .Z(n12309) );
  IV U39517 ( .A(n12308), .Z(n36157) );
  XNOR U39518 ( .A(n12306), .B(n36159), .Z(n12308) );
  XNOR U39519 ( .A(q[2]), .B(DB[3411]), .Z(n36159) );
  XNOR U39520 ( .A(q[1]), .B(DB[3410]), .Z(n12306) );
  XOR U39521 ( .A(n36160), .B(n12271), .Z(n12234) );
  XOR U39522 ( .A(n36161), .B(n12259), .Z(n12271) );
  XNOR U39523 ( .A(q[6]), .B(DB[3422]), .Z(n12259) );
  IV U39524 ( .A(n12258), .Z(n36161) );
  XNOR U39525 ( .A(n12256), .B(n36162), .Z(n12258) );
  XNOR U39526 ( .A(q[5]), .B(DB[3421]), .Z(n36162) );
  XNOR U39527 ( .A(q[4]), .B(DB[3420]), .Z(n12256) );
  IV U39528 ( .A(n12270), .Z(n36160) );
  XOR U39529 ( .A(n36163), .B(n36164), .Z(n12270) );
  XNOR U39530 ( .A(n12266), .B(n12268), .Z(n36164) );
  XNOR U39531 ( .A(q[0]), .B(DB[3416]), .Z(n12268) );
  XNOR U39532 ( .A(q[3]), .B(DB[3419]), .Z(n12266) );
  IV U39533 ( .A(n12265), .Z(n36163) );
  XNOR U39534 ( .A(n12263), .B(n36165), .Z(n12265) );
  XNOR U39535 ( .A(q[2]), .B(DB[3418]), .Z(n36165) );
  XNOR U39536 ( .A(q[1]), .B(DB[3417]), .Z(n12263) );
  XOR U39537 ( .A(n36166), .B(n12228), .Z(n12191) );
  XOR U39538 ( .A(n36167), .B(n12216), .Z(n12228) );
  XNOR U39539 ( .A(q[6]), .B(DB[3429]), .Z(n12216) );
  IV U39540 ( .A(n12215), .Z(n36167) );
  XNOR U39541 ( .A(n12213), .B(n36168), .Z(n12215) );
  XNOR U39542 ( .A(q[5]), .B(DB[3428]), .Z(n36168) );
  XNOR U39543 ( .A(q[4]), .B(DB[3427]), .Z(n12213) );
  IV U39544 ( .A(n12227), .Z(n36166) );
  XOR U39545 ( .A(n36169), .B(n36170), .Z(n12227) );
  XNOR U39546 ( .A(n12223), .B(n12225), .Z(n36170) );
  XNOR U39547 ( .A(q[0]), .B(DB[3423]), .Z(n12225) );
  XNOR U39548 ( .A(q[3]), .B(DB[3426]), .Z(n12223) );
  IV U39549 ( .A(n12222), .Z(n36169) );
  XNOR U39550 ( .A(n12220), .B(n36171), .Z(n12222) );
  XNOR U39551 ( .A(q[2]), .B(DB[3425]), .Z(n36171) );
  XNOR U39552 ( .A(q[1]), .B(DB[3424]), .Z(n12220) );
  XOR U39553 ( .A(n36172), .B(n12185), .Z(n12148) );
  XOR U39554 ( .A(n36173), .B(n12173), .Z(n12185) );
  XNOR U39555 ( .A(q[6]), .B(DB[3436]), .Z(n12173) );
  IV U39556 ( .A(n12172), .Z(n36173) );
  XNOR U39557 ( .A(n12170), .B(n36174), .Z(n12172) );
  XNOR U39558 ( .A(q[5]), .B(DB[3435]), .Z(n36174) );
  XNOR U39559 ( .A(q[4]), .B(DB[3434]), .Z(n12170) );
  IV U39560 ( .A(n12184), .Z(n36172) );
  XOR U39561 ( .A(n36175), .B(n36176), .Z(n12184) );
  XNOR U39562 ( .A(n12180), .B(n12182), .Z(n36176) );
  XNOR U39563 ( .A(q[0]), .B(DB[3430]), .Z(n12182) );
  XNOR U39564 ( .A(q[3]), .B(DB[3433]), .Z(n12180) );
  IV U39565 ( .A(n12179), .Z(n36175) );
  XNOR U39566 ( .A(n12177), .B(n36177), .Z(n12179) );
  XNOR U39567 ( .A(q[2]), .B(DB[3432]), .Z(n36177) );
  XNOR U39568 ( .A(q[1]), .B(DB[3431]), .Z(n12177) );
  XOR U39569 ( .A(n36178), .B(n12142), .Z(n12105) );
  XOR U39570 ( .A(n36179), .B(n12130), .Z(n12142) );
  XNOR U39571 ( .A(q[6]), .B(DB[3443]), .Z(n12130) );
  IV U39572 ( .A(n12129), .Z(n36179) );
  XNOR U39573 ( .A(n12127), .B(n36180), .Z(n12129) );
  XNOR U39574 ( .A(q[5]), .B(DB[3442]), .Z(n36180) );
  XNOR U39575 ( .A(q[4]), .B(DB[3441]), .Z(n12127) );
  IV U39576 ( .A(n12141), .Z(n36178) );
  XOR U39577 ( .A(n36181), .B(n36182), .Z(n12141) );
  XNOR U39578 ( .A(n12137), .B(n12139), .Z(n36182) );
  XNOR U39579 ( .A(q[0]), .B(DB[3437]), .Z(n12139) );
  XNOR U39580 ( .A(q[3]), .B(DB[3440]), .Z(n12137) );
  IV U39581 ( .A(n12136), .Z(n36181) );
  XNOR U39582 ( .A(n12134), .B(n36183), .Z(n12136) );
  XNOR U39583 ( .A(q[2]), .B(DB[3439]), .Z(n36183) );
  XNOR U39584 ( .A(q[1]), .B(DB[3438]), .Z(n12134) );
  XOR U39585 ( .A(n36184), .B(n12099), .Z(n12062) );
  XOR U39586 ( .A(n36185), .B(n12087), .Z(n12099) );
  XNOR U39587 ( .A(q[6]), .B(DB[3450]), .Z(n12087) );
  IV U39588 ( .A(n12086), .Z(n36185) );
  XNOR U39589 ( .A(n12084), .B(n36186), .Z(n12086) );
  XNOR U39590 ( .A(q[5]), .B(DB[3449]), .Z(n36186) );
  XNOR U39591 ( .A(q[4]), .B(DB[3448]), .Z(n12084) );
  IV U39592 ( .A(n12098), .Z(n36184) );
  XOR U39593 ( .A(n36187), .B(n36188), .Z(n12098) );
  XNOR U39594 ( .A(n12094), .B(n12096), .Z(n36188) );
  XNOR U39595 ( .A(q[0]), .B(DB[3444]), .Z(n12096) );
  XNOR U39596 ( .A(q[3]), .B(DB[3447]), .Z(n12094) );
  IV U39597 ( .A(n12093), .Z(n36187) );
  XNOR U39598 ( .A(n12091), .B(n36189), .Z(n12093) );
  XNOR U39599 ( .A(q[2]), .B(DB[3446]), .Z(n36189) );
  XNOR U39600 ( .A(q[1]), .B(DB[3445]), .Z(n12091) );
  XOR U39601 ( .A(n36190), .B(n12056), .Z(n12019) );
  XOR U39602 ( .A(n36191), .B(n12044), .Z(n12056) );
  XNOR U39603 ( .A(q[6]), .B(DB[3457]), .Z(n12044) );
  IV U39604 ( .A(n12043), .Z(n36191) );
  XNOR U39605 ( .A(n12041), .B(n36192), .Z(n12043) );
  XNOR U39606 ( .A(q[5]), .B(DB[3456]), .Z(n36192) );
  XNOR U39607 ( .A(q[4]), .B(DB[3455]), .Z(n12041) );
  IV U39608 ( .A(n12055), .Z(n36190) );
  XOR U39609 ( .A(n36193), .B(n36194), .Z(n12055) );
  XNOR U39610 ( .A(n12051), .B(n12053), .Z(n36194) );
  XNOR U39611 ( .A(q[0]), .B(DB[3451]), .Z(n12053) );
  XNOR U39612 ( .A(q[3]), .B(DB[3454]), .Z(n12051) );
  IV U39613 ( .A(n12050), .Z(n36193) );
  XNOR U39614 ( .A(n12048), .B(n36195), .Z(n12050) );
  XNOR U39615 ( .A(q[2]), .B(DB[3453]), .Z(n36195) );
  XNOR U39616 ( .A(q[1]), .B(DB[3452]), .Z(n12048) );
  XOR U39617 ( .A(n36196), .B(n12013), .Z(n11976) );
  XOR U39618 ( .A(n36197), .B(n12001), .Z(n12013) );
  XNOR U39619 ( .A(q[6]), .B(DB[3464]), .Z(n12001) );
  IV U39620 ( .A(n12000), .Z(n36197) );
  XNOR U39621 ( .A(n11998), .B(n36198), .Z(n12000) );
  XNOR U39622 ( .A(q[5]), .B(DB[3463]), .Z(n36198) );
  XNOR U39623 ( .A(q[4]), .B(DB[3462]), .Z(n11998) );
  IV U39624 ( .A(n12012), .Z(n36196) );
  XOR U39625 ( .A(n36199), .B(n36200), .Z(n12012) );
  XNOR U39626 ( .A(n12008), .B(n12010), .Z(n36200) );
  XNOR U39627 ( .A(q[0]), .B(DB[3458]), .Z(n12010) );
  XNOR U39628 ( .A(q[3]), .B(DB[3461]), .Z(n12008) );
  IV U39629 ( .A(n12007), .Z(n36199) );
  XNOR U39630 ( .A(n12005), .B(n36201), .Z(n12007) );
  XNOR U39631 ( .A(q[2]), .B(DB[3460]), .Z(n36201) );
  XNOR U39632 ( .A(q[1]), .B(DB[3459]), .Z(n12005) );
  XOR U39633 ( .A(n36202), .B(n11970), .Z(n11933) );
  XOR U39634 ( .A(n36203), .B(n11958), .Z(n11970) );
  XNOR U39635 ( .A(q[6]), .B(DB[3471]), .Z(n11958) );
  IV U39636 ( .A(n11957), .Z(n36203) );
  XNOR U39637 ( .A(n11955), .B(n36204), .Z(n11957) );
  XNOR U39638 ( .A(q[5]), .B(DB[3470]), .Z(n36204) );
  XNOR U39639 ( .A(q[4]), .B(DB[3469]), .Z(n11955) );
  IV U39640 ( .A(n11969), .Z(n36202) );
  XOR U39641 ( .A(n36205), .B(n36206), .Z(n11969) );
  XNOR U39642 ( .A(n11965), .B(n11967), .Z(n36206) );
  XNOR U39643 ( .A(q[0]), .B(DB[3465]), .Z(n11967) );
  XNOR U39644 ( .A(q[3]), .B(DB[3468]), .Z(n11965) );
  IV U39645 ( .A(n11964), .Z(n36205) );
  XNOR U39646 ( .A(n11962), .B(n36207), .Z(n11964) );
  XNOR U39647 ( .A(q[2]), .B(DB[3467]), .Z(n36207) );
  XNOR U39648 ( .A(q[1]), .B(DB[3466]), .Z(n11962) );
  XOR U39649 ( .A(n36208), .B(n11927), .Z(n11890) );
  XOR U39650 ( .A(n36209), .B(n11915), .Z(n11927) );
  XNOR U39651 ( .A(q[6]), .B(DB[3478]), .Z(n11915) );
  IV U39652 ( .A(n11914), .Z(n36209) );
  XNOR U39653 ( .A(n11912), .B(n36210), .Z(n11914) );
  XNOR U39654 ( .A(q[5]), .B(DB[3477]), .Z(n36210) );
  XNOR U39655 ( .A(q[4]), .B(DB[3476]), .Z(n11912) );
  IV U39656 ( .A(n11926), .Z(n36208) );
  XOR U39657 ( .A(n36211), .B(n36212), .Z(n11926) );
  XNOR U39658 ( .A(n11922), .B(n11924), .Z(n36212) );
  XNOR U39659 ( .A(q[0]), .B(DB[3472]), .Z(n11924) );
  XNOR U39660 ( .A(q[3]), .B(DB[3475]), .Z(n11922) );
  IV U39661 ( .A(n11921), .Z(n36211) );
  XNOR U39662 ( .A(n11919), .B(n36213), .Z(n11921) );
  XNOR U39663 ( .A(q[2]), .B(DB[3474]), .Z(n36213) );
  XNOR U39664 ( .A(q[1]), .B(DB[3473]), .Z(n11919) );
  XOR U39665 ( .A(n36214), .B(n11884), .Z(n11847) );
  XOR U39666 ( .A(n36215), .B(n11872), .Z(n11884) );
  XNOR U39667 ( .A(q[6]), .B(DB[3485]), .Z(n11872) );
  IV U39668 ( .A(n11871), .Z(n36215) );
  XNOR U39669 ( .A(n11869), .B(n36216), .Z(n11871) );
  XNOR U39670 ( .A(q[5]), .B(DB[3484]), .Z(n36216) );
  XNOR U39671 ( .A(q[4]), .B(DB[3483]), .Z(n11869) );
  IV U39672 ( .A(n11883), .Z(n36214) );
  XOR U39673 ( .A(n36217), .B(n36218), .Z(n11883) );
  XNOR U39674 ( .A(n11879), .B(n11881), .Z(n36218) );
  XNOR U39675 ( .A(q[0]), .B(DB[3479]), .Z(n11881) );
  XNOR U39676 ( .A(q[3]), .B(DB[3482]), .Z(n11879) );
  IV U39677 ( .A(n11878), .Z(n36217) );
  XNOR U39678 ( .A(n11876), .B(n36219), .Z(n11878) );
  XNOR U39679 ( .A(q[2]), .B(DB[3481]), .Z(n36219) );
  XNOR U39680 ( .A(q[1]), .B(DB[3480]), .Z(n11876) );
  XOR U39681 ( .A(n36220), .B(n11841), .Z(n11804) );
  XOR U39682 ( .A(n36221), .B(n11829), .Z(n11841) );
  XNOR U39683 ( .A(q[6]), .B(DB[3492]), .Z(n11829) );
  IV U39684 ( .A(n11828), .Z(n36221) );
  XNOR U39685 ( .A(n11826), .B(n36222), .Z(n11828) );
  XNOR U39686 ( .A(q[5]), .B(DB[3491]), .Z(n36222) );
  XNOR U39687 ( .A(q[4]), .B(DB[3490]), .Z(n11826) );
  IV U39688 ( .A(n11840), .Z(n36220) );
  XOR U39689 ( .A(n36223), .B(n36224), .Z(n11840) );
  XNOR U39690 ( .A(n11836), .B(n11838), .Z(n36224) );
  XNOR U39691 ( .A(q[0]), .B(DB[3486]), .Z(n11838) );
  XNOR U39692 ( .A(q[3]), .B(DB[3489]), .Z(n11836) );
  IV U39693 ( .A(n11835), .Z(n36223) );
  XNOR U39694 ( .A(n11833), .B(n36225), .Z(n11835) );
  XNOR U39695 ( .A(q[2]), .B(DB[3488]), .Z(n36225) );
  XNOR U39696 ( .A(q[1]), .B(DB[3487]), .Z(n11833) );
  XOR U39697 ( .A(n36226), .B(n11798), .Z(n11761) );
  XOR U39698 ( .A(n36227), .B(n11786), .Z(n11798) );
  XNOR U39699 ( .A(q[6]), .B(DB[3499]), .Z(n11786) );
  IV U39700 ( .A(n11785), .Z(n36227) );
  XNOR U39701 ( .A(n11783), .B(n36228), .Z(n11785) );
  XNOR U39702 ( .A(q[5]), .B(DB[3498]), .Z(n36228) );
  XNOR U39703 ( .A(q[4]), .B(DB[3497]), .Z(n11783) );
  IV U39704 ( .A(n11797), .Z(n36226) );
  XOR U39705 ( .A(n36229), .B(n36230), .Z(n11797) );
  XNOR U39706 ( .A(n11793), .B(n11795), .Z(n36230) );
  XNOR U39707 ( .A(q[0]), .B(DB[3493]), .Z(n11795) );
  XNOR U39708 ( .A(q[3]), .B(DB[3496]), .Z(n11793) );
  IV U39709 ( .A(n11792), .Z(n36229) );
  XNOR U39710 ( .A(n11790), .B(n36231), .Z(n11792) );
  XNOR U39711 ( .A(q[2]), .B(DB[3495]), .Z(n36231) );
  XNOR U39712 ( .A(q[1]), .B(DB[3494]), .Z(n11790) );
  XOR U39713 ( .A(n36232), .B(n11755), .Z(n11718) );
  XOR U39714 ( .A(n36233), .B(n11743), .Z(n11755) );
  XNOR U39715 ( .A(q[6]), .B(DB[3506]), .Z(n11743) );
  IV U39716 ( .A(n11742), .Z(n36233) );
  XNOR U39717 ( .A(n11740), .B(n36234), .Z(n11742) );
  XNOR U39718 ( .A(q[5]), .B(DB[3505]), .Z(n36234) );
  XNOR U39719 ( .A(q[4]), .B(DB[3504]), .Z(n11740) );
  IV U39720 ( .A(n11754), .Z(n36232) );
  XOR U39721 ( .A(n36235), .B(n36236), .Z(n11754) );
  XNOR U39722 ( .A(n11750), .B(n11752), .Z(n36236) );
  XNOR U39723 ( .A(q[0]), .B(DB[3500]), .Z(n11752) );
  XNOR U39724 ( .A(q[3]), .B(DB[3503]), .Z(n11750) );
  IV U39725 ( .A(n11749), .Z(n36235) );
  XNOR U39726 ( .A(n11747), .B(n36237), .Z(n11749) );
  XNOR U39727 ( .A(q[2]), .B(DB[3502]), .Z(n36237) );
  XNOR U39728 ( .A(q[1]), .B(DB[3501]), .Z(n11747) );
  XOR U39729 ( .A(n36238), .B(n11712), .Z(n11675) );
  XOR U39730 ( .A(n36239), .B(n11700), .Z(n11712) );
  XNOR U39731 ( .A(q[6]), .B(DB[3513]), .Z(n11700) );
  IV U39732 ( .A(n11699), .Z(n36239) );
  XNOR U39733 ( .A(n11697), .B(n36240), .Z(n11699) );
  XNOR U39734 ( .A(q[5]), .B(DB[3512]), .Z(n36240) );
  XNOR U39735 ( .A(q[4]), .B(DB[3511]), .Z(n11697) );
  IV U39736 ( .A(n11711), .Z(n36238) );
  XOR U39737 ( .A(n36241), .B(n36242), .Z(n11711) );
  XNOR U39738 ( .A(n11707), .B(n11709), .Z(n36242) );
  XNOR U39739 ( .A(q[0]), .B(DB[3507]), .Z(n11709) );
  XNOR U39740 ( .A(q[3]), .B(DB[3510]), .Z(n11707) );
  IV U39741 ( .A(n11706), .Z(n36241) );
  XNOR U39742 ( .A(n11704), .B(n36243), .Z(n11706) );
  XNOR U39743 ( .A(q[2]), .B(DB[3509]), .Z(n36243) );
  XNOR U39744 ( .A(q[1]), .B(DB[3508]), .Z(n11704) );
  XOR U39745 ( .A(n36244), .B(n11669), .Z(n11632) );
  XOR U39746 ( .A(n36245), .B(n11657), .Z(n11669) );
  XNOR U39747 ( .A(q[6]), .B(DB[3520]), .Z(n11657) );
  IV U39748 ( .A(n11656), .Z(n36245) );
  XNOR U39749 ( .A(n11654), .B(n36246), .Z(n11656) );
  XNOR U39750 ( .A(q[5]), .B(DB[3519]), .Z(n36246) );
  XNOR U39751 ( .A(q[4]), .B(DB[3518]), .Z(n11654) );
  IV U39752 ( .A(n11668), .Z(n36244) );
  XOR U39753 ( .A(n36247), .B(n36248), .Z(n11668) );
  XNOR U39754 ( .A(n11664), .B(n11666), .Z(n36248) );
  XNOR U39755 ( .A(q[0]), .B(DB[3514]), .Z(n11666) );
  XNOR U39756 ( .A(q[3]), .B(DB[3517]), .Z(n11664) );
  IV U39757 ( .A(n11663), .Z(n36247) );
  XNOR U39758 ( .A(n11661), .B(n36249), .Z(n11663) );
  XNOR U39759 ( .A(q[2]), .B(DB[3516]), .Z(n36249) );
  XNOR U39760 ( .A(q[1]), .B(DB[3515]), .Z(n11661) );
  XOR U39761 ( .A(n36250), .B(n11626), .Z(n11589) );
  XOR U39762 ( .A(n36251), .B(n11614), .Z(n11626) );
  XNOR U39763 ( .A(q[6]), .B(DB[3527]), .Z(n11614) );
  IV U39764 ( .A(n11613), .Z(n36251) );
  XNOR U39765 ( .A(n11611), .B(n36252), .Z(n11613) );
  XNOR U39766 ( .A(q[5]), .B(DB[3526]), .Z(n36252) );
  XNOR U39767 ( .A(q[4]), .B(DB[3525]), .Z(n11611) );
  IV U39768 ( .A(n11625), .Z(n36250) );
  XOR U39769 ( .A(n36253), .B(n36254), .Z(n11625) );
  XNOR U39770 ( .A(n11621), .B(n11623), .Z(n36254) );
  XNOR U39771 ( .A(q[0]), .B(DB[3521]), .Z(n11623) );
  XNOR U39772 ( .A(q[3]), .B(DB[3524]), .Z(n11621) );
  IV U39773 ( .A(n11620), .Z(n36253) );
  XNOR U39774 ( .A(n11618), .B(n36255), .Z(n11620) );
  XNOR U39775 ( .A(q[2]), .B(DB[3523]), .Z(n36255) );
  XNOR U39776 ( .A(q[1]), .B(DB[3522]), .Z(n11618) );
  XOR U39777 ( .A(n36256), .B(n11583), .Z(n11546) );
  XOR U39778 ( .A(n36257), .B(n11571), .Z(n11583) );
  XNOR U39779 ( .A(q[6]), .B(DB[3534]), .Z(n11571) );
  IV U39780 ( .A(n11570), .Z(n36257) );
  XNOR U39781 ( .A(n11568), .B(n36258), .Z(n11570) );
  XNOR U39782 ( .A(q[5]), .B(DB[3533]), .Z(n36258) );
  XNOR U39783 ( .A(q[4]), .B(DB[3532]), .Z(n11568) );
  IV U39784 ( .A(n11582), .Z(n36256) );
  XOR U39785 ( .A(n36259), .B(n36260), .Z(n11582) );
  XNOR U39786 ( .A(n11578), .B(n11580), .Z(n36260) );
  XNOR U39787 ( .A(q[0]), .B(DB[3528]), .Z(n11580) );
  XNOR U39788 ( .A(q[3]), .B(DB[3531]), .Z(n11578) );
  IV U39789 ( .A(n11577), .Z(n36259) );
  XNOR U39790 ( .A(n11575), .B(n36261), .Z(n11577) );
  XNOR U39791 ( .A(q[2]), .B(DB[3530]), .Z(n36261) );
  XNOR U39792 ( .A(q[1]), .B(DB[3529]), .Z(n11575) );
  XOR U39793 ( .A(n36262), .B(n11540), .Z(n11503) );
  XOR U39794 ( .A(n36263), .B(n11528), .Z(n11540) );
  XNOR U39795 ( .A(q[6]), .B(DB[3541]), .Z(n11528) );
  IV U39796 ( .A(n11527), .Z(n36263) );
  XNOR U39797 ( .A(n11525), .B(n36264), .Z(n11527) );
  XNOR U39798 ( .A(q[5]), .B(DB[3540]), .Z(n36264) );
  XNOR U39799 ( .A(q[4]), .B(DB[3539]), .Z(n11525) );
  IV U39800 ( .A(n11539), .Z(n36262) );
  XOR U39801 ( .A(n36265), .B(n36266), .Z(n11539) );
  XNOR U39802 ( .A(n11535), .B(n11537), .Z(n36266) );
  XNOR U39803 ( .A(q[0]), .B(DB[3535]), .Z(n11537) );
  XNOR U39804 ( .A(q[3]), .B(DB[3538]), .Z(n11535) );
  IV U39805 ( .A(n11534), .Z(n36265) );
  XNOR U39806 ( .A(n11532), .B(n36267), .Z(n11534) );
  XNOR U39807 ( .A(q[2]), .B(DB[3537]), .Z(n36267) );
  XNOR U39808 ( .A(q[1]), .B(DB[3536]), .Z(n11532) );
  XOR U39809 ( .A(n36268), .B(n11497), .Z(n11460) );
  XOR U39810 ( .A(n36269), .B(n11485), .Z(n11497) );
  XNOR U39811 ( .A(q[6]), .B(DB[3548]), .Z(n11485) );
  IV U39812 ( .A(n11484), .Z(n36269) );
  XNOR U39813 ( .A(n11482), .B(n36270), .Z(n11484) );
  XNOR U39814 ( .A(q[5]), .B(DB[3547]), .Z(n36270) );
  XNOR U39815 ( .A(q[4]), .B(DB[3546]), .Z(n11482) );
  IV U39816 ( .A(n11496), .Z(n36268) );
  XOR U39817 ( .A(n36271), .B(n36272), .Z(n11496) );
  XNOR U39818 ( .A(n11492), .B(n11494), .Z(n36272) );
  XNOR U39819 ( .A(q[0]), .B(DB[3542]), .Z(n11494) );
  XNOR U39820 ( .A(q[3]), .B(DB[3545]), .Z(n11492) );
  IV U39821 ( .A(n11491), .Z(n36271) );
  XNOR U39822 ( .A(n11489), .B(n36273), .Z(n11491) );
  XNOR U39823 ( .A(q[2]), .B(DB[3544]), .Z(n36273) );
  XNOR U39824 ( .A(q[1]), .B(DB[3543]), .Z(n11489) );
  XOR U39825 ( .A(n36274), .B(n11454), .Z(n11417) );
  XOR U39826 ( .A(n36275), .B(n11442), .Z(n11454) );
  XNOR U39827 ( .A(q[6]), .B(DB[3555]), .Z(n11442) );
  IV U39828 ( .A(n11441), .Z(n36275) );
  XNOR U39829 ( .A(n11439), .B(n36276), .Z(n11441) );
  XNOR U39830 ( .A(q[5]), .B(DB[3554]), .Z(n36276) );
  XNOR U39831 ( .A(q[4]), .B(DB[3553]), .Z(n11439) );
  IV U39832 ( .A(n11453), .Z(n36274) );
  XOR U39833 ( .A(n36277), .B(n36278), .Z(n11453) );
  XNOR U39834 ( .A(n11449), .B(n11451), .Z(n36278) );
  XNOR U39835 ( .A(q[0]), .B(DB[3549]), .Z(n11451) );
  XNOR U39836 ( .A(q[3]), .B(DB[3552]), .Z(n11449) );
  IV U39837 ( .A(n11448), .Z(n36277) );
  XNOR U39838 ( .A(n11446), .B(n36279), .Z(n11448) );
  XNOR U39839 ( .A(q[2]), .B(DB[3551]), .Z(n36279) );
  XNOR U39840 ( .A(q[1]), .B(DB[3550]), .Z(n11446) );
  XOR U39841 ( .A(n36280), .B(n11411), .Z(n11374) );
  XOR U39842 ( .A(n36281), .B(n11399), .Z(n11411) );
  XNOR U39843 ( .A(q[6]), .B(DB[3562]), .Z(n11399) );
  IV U39844 ( .A(n11398), .Z(n36281) );
  XNOR U39845 ( .A(n11396), .B(n36282), .Z(n11398) );
  XNOR U39846 ( .A(q[5]), .B(DB[3561]), .Z(n36282) );
  XNOR U39847 ( .A(q[4]), .B(DB[3560]), .Z(n11396) );
  IV U39848 ( .A(n11410), .Z(n36280) );
  XOR U39849 ( .A(n36283), .B(n36284), .Z(n11410) );
  XNOR U39850 ( .A(n11406), .B(n11408), .Z(n36284) );
  XNOR U39851 ( .A(q[0]), .B(DB[3556]), .Z(n11408) );
  XNOR U39852 ( .A(q[3]), .B(DB[3559]), .Z(n11406) );
  IV U39853 ( .A(n11405), .Z(n36283) );
  XNOR U39854 ( .A(n11403), .B(n36285), .Z(n11405) );
  XNOR U39855 ( .A(q[2]), .B(DB[3558]), .Z(n36285) );
  XNOR U39856 ( .A(q[1]), .B(DB[3557]), .Z(n11403) );
  XOR U39857 ( .A(n36286), .B(n11368), .Z(n11331) );
  XOR U39858 ( .A(n36287), .B(n11356), .Z(n11368) );
  XNOR U39859 ( .A(q[6]), .B(DB[3569]), .Z(n11356) );
  IV U39860 ( .A(n11355), .Z(n36287) );
  XNOR U39861 ( .A(n11353), .B(n36288), .Z(n11355) );
  XNOR U39862 ( .A(q[5]), .B(DB[3568]), .Z(n36288) );
  XNOR U39863 ( .A(q[4]), .B(DB[3567]), .Z(n11353) );
  IV U39864 ( .A(n11367), .Z(n36286) );
  XOR U39865 ( .A(n36289), .B(n36290), .Z(n11367) );
  XNOR U39866 ( .A(n11363), .B(n11365), .Z(n36290) );
  XNOR U39867 ( .A(q[0]), .B(DB[3563]), .Z(n11365) );
  XNOR U39868 ( .A(q[3]), .B(DB[3566]), .Z(n11363) );
  IV U39869 ( .A(n11362), .Z(n36289) );
  XNOR U39870 ( .A(n11360), .B(n36291), .Z(n11362) );
  XNOR U39871 ( .A(q[2]), .B(DB[3565]), .Z(n36291) );
  XNOR U39872 ( .A(q[1]), .B(DB[3564]), .Z(n11360) );
  XOR U39873 ( .A(n36292), .B(n11325), .Z(n11287) );
  XOR U39874 ( .A(n36293), .B(n11313), .Z(n11325) );
  XNOR U39875 ( .A(q[6]), .B(DB[3576]), .Z(n11313) );
  IV U39876 ( .A(n11312), .Z(n36293) );
  XNOR U39877 ( .A(n11310), .B(n36294), .Z(n11312) );
  XNOR U39878 ( .A(q[5]), .B(DB[3575]), .Z(n36294) );
  XNOR U39879 ( .A(q[4]), .B(DB[3574]), .Z(n11310) );
  IV U39880 ( .A(n11324), .Z(n36292) );
  XOR U39881 ( .A(n36295), .B(n36296), .Z(n11324) );
  XNOR U39882 ( .A(n11320), .B(n11322), .Z(n36296) );
  XNOR U39883 ( .A(q[0]), .B(DB[3570]), .Z(n11322) );
  XNOR U39884 ( .A(q[3]), .B(DB[3573]), .Z(n11320) );
  IV U39885 ( .A(n11319), .Z(n36295) );
  XNOR U39886 ( .A(n11317), .B(n36297), .Z(n11319) );
  XNOR U39887 ( .A(q[2]), .B(DB[3572]), .Z(n36297) );
  XNOR U39888 ( .A(q[1]), .B(DB[3571]), .Z(n11317) );
endmodule

