
module hamming_N1600_CC32 ( clk, rst, x, y, o );
  input [49:0] x;
  input [49:0] y;
  output [10:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334;
  wire   [10:0] oglobal;

  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U53 ( .A(n220), .B(n222), .Z(n1) );
  XOR U54 ( .A(n220), .B(n222), .Z(n2) );
  NAND U55 ( .A(n2), .B(n221), .Z(n3) );
  NAND U56 ( .A(n1), .B(n3), .Z(n246) );
  XNOR U57 ( .A(n186), .B(n185), .Z(n214) );
  NAND U58 ( .A(n249), .B(n250), .Z(n4) );
  XOR U59 ( .A(n249), .B(n250), .Z(n5) );
  NANDN U60 ( .A(n248), .B(n5), .Z(n6) );
  NAND U61 ( .A(n4), .B(n6), .Z(n286) );
  NAND U62 ( .A(n294), .B(n296), .Z(n7) );
  XOR U63 ( .A(n294), .B(n296), .Z(n8) );
  NAND U64 ( .A(n8), .B(n295), .Z(n9) );
  NAND U65 ( .A(n7), .B(n9), .Z(n310) );
  NAND U66 ( .A(n299), .B(n300), .Z(n10) );
  XOR U67 ( .A(n299), .B(n300), .Z(n11) );
  NANDN U68 ( .A(n298), .B(n11), .Z(n12) );
  NAND U69 ( .A(n10), .B(n12), .Z(n315) );
  NAND U70 ( .A(n168), .B(n167), .Z(n13) );
  NAND U71 ( .A(n165), .B(n166), .Z(n14) );
  NAND U72 ( .A(n13), .B(n14), .Z(n272) );
  XOR U73 ( .A(n211), .B(n212), .Z(n15) );
  NANDN U74 ( .A(n213), .B(n15), .Z(n16) );
  NAND U75 ( .A(n211), .B(n212), .Z(n17) );
  AND U76 ( .A(n16), .B(n17), .Z(n245) );
  NAND U77 ( .A(n275), .B(n277), .Z(n18) );
  XOR U78 ( .A(n275), .B(n277), .Z(n19) );
  NAND U79 ( .A(n19), .B(n276), .Z(n20) );
  NAND U80 ( .A(n18), .B(n20), .Z(n300) );
  NAND U81 ( .A(n311), .B(n312), .Z(n21) );
  XOR U82 ( .A(n311), .B(n312), .Z(n22) );
  NAND U83 ( .A(n22), .B(n310), .Z(n23) );
  NAND U84 ( .A(n21), .B(n23), .Z(n324) );
  NAND U85 ( .A(n228), .B(n229), .Z(n24) );
  XOR U86 ( .A(n228), .B(n229), .Z(n25) );
  NANDN U87 ( .A(n227), .B(n25), .Z(n26) );
  NAND U88 ( .A(n24), .B(n26), .Z(n283) );
  NAND U89 ( .A(n317), .B(n318), .Z(n27) );
  XOR U90 ( .A(n317), .B(n318), .Z(n28) );
  NANDN U91 ( .A(n316), .B(n28), .Z(n29) );
  NAND U92 ( .A(n27), .B(n29), .Z(n320) );
  NAND U93 ( .A(n157), .B(n156), .Z(n30) );
  NAND U94 ( .A(n154), .B(n155), .Z(n31) );
  NAND U95 ( .A(n30), .B(n31), .Z(n271) );
  NAND U96 ( .A(n204), .B(n203), .Z(n32) );
  NAND U97 ( .A(n202), .B(oglobal[0]), .Z(n33) );
  NAND U98 ( .A(n32), .B(n33), .Z(n233) );
  NAND U99 ( .A(n138), .B(n137), .Z(n34) );
  NAND U100 ( .A(n135), .B(n136), .Z(n35) );
  AND U101 ( .A(n34), .B(n35), .Z(n238) );
  XNOR U102 ( .A(n192), .B(n191), .Z(n215) );
  NAND U103 ( .A(n263), .B(n264), .Z(n36) );
  XOR U104 ( .A(n263), .B(n264), .Z(n37) );
  NANDN U105 ( .A(n262), .B(n37), .Z(n38) );
  NAND U106 ( .A(n36), .B(n38), .Z(n291) );
  NAND U107 ( .A(n141), .B(n143), .Z(n39) );
  XOR U108 ( .A(n141), .B(n143), .Z(n40) );
  NAND U109 ( .A(n40), .B(n142), .Z(n41) );
  NAND U110 ( .A(n39), .B(n41), .Z(n276) );
  XOR U111 ( .A(n255), .B(n254), .Z(n42) );
  XNOR U112 ( .A(n257), .B(n42), .Z(n282) );
  NAND U113 ( .A(n302), .B(n304), .Z(n43) );
  XOR U114 ( .A(n302), .B(n304), .Z(n44) );
  NAND U115 ( .A(n44), .B(n303), .Z(n45) );
  NAND U116 ( .A(n43), .B(n45), .Z(n318) );
  XOR U117 ( .A(n315), .B(n313), .Z(n46) );
  NANDN U118 ( .A(n314), .B(n46), .Z(n47) );
  NAND U119 ( .A(n315), .B(n313), .Z(n48) );
  AND U120 ( .A(n47), .B(n48), .Z(n321) );
  XNOR U121 ( .A(n184), .B(n183), .Z(n185) );
  AND U122 ( .A(n231), .B(oglobal[1]), .Z(n290) );
  NAND U123 ( .A(n272), .B(n271), .Z(n49) );
  XOR U124 ( .A(n272), .B(n271), .Z(n50) );
  NANDN U125 ( .A(n273), .B(n50), .Z(n51) );
  NAND U126 ( .A(n49), .B(n51), .Z(n292) );
  NAND U127 ( .A(n245), .B(n247), .Z(n52) );
  XOR U128 ( .A(n245), .B(n247), .Z(n53) );
  NAND U129 ( .A(n53), .B(n246), .Z(n54) );
  NAND U130 ( .A(n52), .B(n54), .Z(n287) );
  XOR U131 ( .A(n280), .B(n278), .Z(n55) );
  NANDN U132 ( .A(n279), .B(n55), .Z(n56) );
  NAND U133 ( .A(n280), .B(n278), .Z(n57) );
  AND U134 ( .A(n56), .B(n57), .Z(n299) );
  NAND U135 ( .A(n252), .B(n253), .Z(n58) );
  XOR U136 ( .A(n252), .B(n253), .Z(n59) );
  NANDN U137 ( .A(n251), .B(n59), .Z(n60) );
  NAND U138 ( .A(n58), .B(n60), .Z(n303) );
  NAND U139 ( .A(n282), .B(n284), .Z(n61) );
  XOR U140 ( .A(n282), .B(n284), .Z(n62) );
  NANDN U141 ( .A(n283), .B(n62), .Z(n63) );
  NAND U142 ( .A(n61), .B(n63), .Z(n305) );
  NAND U143 ( .A(n320), .B(n322), .Z(n64) );
  XOR U144 ( .A(n320), .B(n322), .Z(n65) );
  NAND U145 ( .A(n65), .B(n321), .Z(n66) );
  NAND U146 ( .A(n64), .B(n66), .Z(n330) );
  NAND U147 ( .A(n130), .B(n129), .Z(n67) );
  NAND U148 ( .A(n127), .B(n128), .Z(n68) );
  NAND U149 ( .A(n67), .B(n68), .Z(n231) );
  XNOR U150 ( .A(n178), .B(n177), .Z(n179) );
  XNOR U151 ( .A(n190), .B(n189), .Z(n191) );
  NAND U152 ( .A(n208), .B(n207), .Z(n69) );
  NAND U153 ( .A(n205), .B(n206), .Z(n70) );
  AND U154 ( .A(n69), .B(n70), .Z(n232) );
  NAND U155 ( .A(n134), .B(n133), .Z(n71) );
  NAND U156 ( .A(n131), .B(n132), .Z(n72) );
  NAND U157 ( .A(n71), .B(n72), .Z(n239) );
  NAND U158 ( .A(n126), .B(n125), .Z(n73) );
  NANDN U159 ( .A(n124), .B(n123), .Z(n74) );
  NAND U160 ( .A(n73), .B(n74), .Z(n252) );
  NAND U161 ( .A(n291), .B(n293), .Z(n75) );
  XOR U162 ( .A(n291), .B(n293), .Z(n76) );
  NAND U163 ( .A(n76), .B(n292), .Z(n77) );
  NAND U164 ( .A(n75), .B(n77), .Z(n312) );
  NAND U165 ( .A(n144), .B(n146), .Z(n78) );
  XOR U166 ( .A(n144), .B(n146), .Z(n79) );
  NAND U167 ( .A(n79), .B(n145), .Z(n80) );
  NAND U168 ( .A(n78), .B(n80), .Z(n275) );
  XOR U169 ( .A(n226), .B(n224), .Z(n81) );
  NANDN U170 ( .A(n225), .B(n81), .Z(n82) );
  NAND U171 ( .A(n226), .B(n224), .Z(n83) );
  AND U172 ( .A(n82), .B(n83), .Z(n255) );
  OR U173 ( .A(n287), .B(n286), .Z(n84) );
  NAND U174 ( .A(n288), .B(n289), .Z(n85) );
  AND U175 ( .A(n84), .B(n85), .Z(n313) );
  NAND U176 ( .A(n306), .B(n307), .Z(n86) );
  XOR U177 ( .A(n306), .B(n307), .Z(n87) );
  NAND U178 ( .A(n87), .B(n305), .Z(n88) );
  NAND U179 ( .A(n86), .B(n88), .Z(n316) );
  XOR U180 ( .A(oglobal[5]), .B(n329), .Z(n89) );
  NANDN U181 ( .A(n330), .B(n89), .Z(n90) );
  NAND U182 ( .A(oglobal[5]), .B(n329), .Z(n91) );
  AND U183 ( .A(n90), .B(n91), .Z(n331) );
  NAND U184 ( .A(n334), .B(oglobal[9]), .Z(n92) );
  XNOR U185 ( .A(oglobal[10]), .B(n92), .Z(o[10]) );
  XOR U186 ( .A(x[5]), .B(y[5]), .Z(n183) );
  XNOR U187 ( .A(x[3]), .B(y[3]), .Z(n184) );
  XNOR U188 ( .A(x[7]), .B(y[7]), .Z(n186) );
  XOR U189 ( .A(x[2]), .B(y[2]), .Z(n177) );
  XNOR U190 ( .A(x[0]), .B(y[0]), .Z(n178) );
  XNOR U191 ( .A(x[1]), .B(y[1]), .Z(n180) );
  IV U192 ( .A(n180), .Z(n93) );
  XOR U193 ( .A(n179), .B(n93), .Z(n217) );
  XOR U194 ( .A(x[11]), .B(y[11]), .Z(n189) );
  XNOR U195 ( .A(x[9]), .B(y[9]), .Z(n190) );
  XNOR U196 ( .A(x[13]), .B(y[13]), .Z(n192) );
  XNOR U197 ( .A(n217), .B(n215), .Z(n94) );
  XOR U198 ( .A(n214), .B(n94), .Z(n226) );
  XOR U199 ( .A(x[28]), .B(y[28]), .Z(n150) );
  XOR U200 ( .A(x[32]), .B(y[32]), .Z(n148) );
  XNOR U201 ( .A(x[30]), .B(y[30]), .Z(n149) );
  XOR U202 ( .A(n148), .B(n149), .Z(n151) );
  XOR U203 ( .A(n150), .B(n151), .Z(n212) );
  XOR U204 ( .A(x[34]), .B(y[34]), .Z(n172) );
  XOR U205 ( .A(x[38]), .B(y[38]), .Z(n170) );
  XNOR U206 ( .A(x[36]), .B(y[36]), .Z(n171) );
  XOR U207 ( .A(n170), .B(n171), .Z(n173) );
  XNOR U208 ( .A(n172), .B(n173), .Z(n213) );
  XOR U209 ( .A(x[22]), .B(y[22]), .Z(n198) );
  XOR U210 ( .A(x[26]), .B(y[26]), .Z(n196) );
  XNOR U211 ( .A(x[24]), .B(y[24]), .Z(n197) );
  XOR U212 ( .A(n196), .B(n197), .Z(n199) );
  XOR U213 ( .A(n198), .B(n199), .Z(n211) );
  XOR U214 ( .A(n213), .B(n211), .Z(n95) );
  XOR U215 ( .A(n212), .B(n95), .Z(n225) );
  XOR U216 ( .A(x[33]), .B(y[33]), .Z(n134) );
  XOR U217 ( .A(x[47]), .B(y[47]), .Z(n132) );
  XOR U218 ( .A(x[31]), .B(y[31]), .Z(n131) );
  XOR U219 ( .A(n132), .B(n131), .Z(n133) );
  XOR U220 ( .A(n134), .B(n133), .Z(n141) );
  XOR U221 ( .A(x[29]), .B(y[29]), .Z(n118) );
  XOR U222 ( .A(x[49]), .B(y[49]), .Z(n116) );
  XOR U223 ( .A(x[27]), .B(y[27]), .Z(n115) );
  XOR U224 ( .A(n116), .B(n115), .Z(n117) );
  XOR U225 ( .A(n118), .B(n117), .Z(n143) );
  XOR U226 ( .A(x[37]), .B(y[37]), .Z(n130) );
  XOR U227 ( .A(x[45]), .B(y[45]), .Z(n128) );
  XOR U228 ( .A(x[35]), .B(y[35]), .Z(n127) );
  XOR U229 ( .A(n128), .B(n127), .Z(n129) );
  XOR U230 ( .A(n130), .B(n129), .Z(n142) );
  XNOR U231 ( .A(n143), .B(n142), .Z(n96) );
  XOR U232 ( .A(n141), .B(n96), .Z(n224) );
  XOR U233 ( .A(n225), .B(n224), .Z(n97) );
  XOR U234 ( .A(n226), .B(n97), .Z(n227) );
  XOR U235 ( .A(x[10]), .B(y[10]), .Z(n162) );
  XOR U236 ( .A(x[14]), .B(y[14]), .Z(n159) );
  XOR U237 ( .A(x[12]), .B(y[12]), .Z(n158) );
  XOR U238 ( .A(n159), .B(n158), .Z(n161) );
  XOR U239 ( .A(n162), .B(n161), .Z(n220) );
  XOR U240 ( .A(x[16]), .B(y[16]), .Z(n208) );
  XOR U241 ( .A(x[20]), .B(y[20]), .Z(n206) );
  XOR U242 ( .A(x[18]), .B(y[18]), .Z(n205) );
  XOR U243 ( .A(n206), .B(n205), .Z(n207) );
  XOR U244 ( .A(n208), .B(n207), .Z(n222) );
  XOR U245 ( .A(x[4]), .B(y[4]), .Z(n157) );
  XOR U246 ( .A(x[8]), .B(y[8]), .Z(n155) );
  XOR U247 ( .A(x[6]), .B(y[6]), .Z(n154) );
  XOR U248 ( .A(n155), .B(n154), .Z(n156) );
  XOR U249 ( .A(n157), .B(n156), .Z(n221) );
  XNOR U250 ( .A(n222), .B(n221), .Z(n98) );
  XOR U251 ( .A(n220), .B(n98), .Z(n125) );
  XOR U252 ( .A(x[44]), .B(y[44]), .Z(n168) );
  XOR U253 ( .A(x[48]), .B(y[48]), .Z(n166) );
  XOR U254 ( .A(x[46]), .B(y[46]), .Z(n165) );
  XOR U255 ( .A(n166), .B(n165), .Z(n167) );
  XOR U256 ( .A(n168), .B(n167), .Z(n124) );
  XOR U257 ( .A(x[40]), .B(y[40]), .Z(n204) );
  XOR U258 ( .A(x[42]), .B(y[42]), .Z(n202) );
  XOR U259 ( .A(oglobal[0]), .B(n202), .Z(n203) );
  XNOR U260 ( .A(n204), .B(n203), .Z(n123) );
  XNOR U261 ( .A(n124), .B(n123), .Z(n126) );
  XOR U262 ( .A(n125), .B(n126), .Z(n229) );
  XOR U263 ( .A(x[25]), .B(y[25]), .Z(n111) );
  XOR U264 ( .A(x[23]), .B(y[23]), .Z(n109) );
  XOR U265 ( .A(x[21]), .B(y[21]), .Z(n108) );
  XOR U266 ( .A(n109), .B(n108), .Z(n110) );
  XOR U267 ( .A(n111), .B(n110), .Z(n144) );
  XOR U268 ( .A(x[19]), .B(y[19]), .Z(n104) );
  XOR U269 ( .A(x[17]), .B(y[17]), .Z(n102) );
  XOR U270 ( .A(x[15]), .B(y[15]), .Z(n101) );
  XOR U271 ( .A(n102), .B(n101), .Z(n103) );
  XOR U272 ( .A(n104), .B(n103), .Z(n146) );
  XOR U273 ( .A(x[41]), .B(y[41]), .Z(n138) );
  XOR U274 ( .A(x[43]), .B(y[43]), .Z(n136) );
  XOR U275 ( .A(x[39]), .B(y[39]), .Z(n135) );
  XOR U276 ( .A(n136), .B(n135), .Z(n137) );
  XOR U277 ( .A(n138), .B(n137), .Z(n145) );
  XNOR U278 ( .A(n146), .B(n145), .Z(n99) );
  XOR U279 ( .A(n144), .B(n99), .Z(n228) );
  XOR U280 ( .A(n229), .B(n228), .Z(n100) );
  XOR U281 ( .A(n227), .B(n100), .Z(o[0]) );
  NAND U282 ( .A(n102), .B(n101), .Z(n107) );
  IV U283 ( .A(n103), .Z(n105) );
  NANDN U284 ( .A(n105), .B(n104), .Z(n106) );
  NAND U285 ( .A(n107), .B(n106), .Z(n264) );
  NAND U286 ( .A(n109), .B(n108), .Z(n114) );
  IV U287 ( .A(n110), .Z(n112) );
  NANDN U288 ( .A(n112), .B(n111), .Z(n113) );
  NAND U289 ( .A(n114), .B(n113), .Z(n263) );
  NAND U290 ( .A(n116), .B(n115), .Z(n121) );
  IV U291 ( .A(n117), .Z(n119) );
  NANDN U292 ( .A(n119), .B(n118), .Z(n120) );
  AND U293 ( .A(n121), .B(n120), .Z(n262) );
  XOR U294 ( .A(n263), .B(n262), .Z(n122) );
  XOR U295 ( .A(n264), .B(n122), .Z(n253) );
  XOR U296 ( .A(n231), .B(oglobal[1]), .Z(n240) );
  XOR U297 ( .A(n239), .B(n238), .Z(n139) );
  XNOR U298 ( .A(n240), .B(n139), .Z(n251) );
  XOR U299 ( .A(n252), .B(n251), .Z(n140) );
  XOR U300 ( .A(n253), .B(n140), .Z(n277) );
  XNOR U301 ( .A(n276), .B(n275), .Z(n147) );
  XNOR U302 ( .A(n277), .B(n147), .Z(n284) );
  NANDN U303 ( .A(n149), .B(n148), .Z(n153) );
  NANDN U304 ( .A(n151), .B(n150), .Z(n152) );
  NAND U305 ( .A(n153), .B(n152), .Z(n267) );
  IV U306 ( .A(n158), .Z(n160) );
  NANDN U307 ( .A(n160), .B(n159), .Z(n164) );
  NAND U308 ( .A(n162), .B(n161), .Z(n163) );
  AND U309 ( .A(n164), .B(n163), .Z(n273) );
  XOR U310 ( .A(n273), .B(n272), .Z(n169) );
  XNOR U311 ( .A(n271), .B(n169), .Z(n266) );
  NANDN U312 ( .A(n171), .B(n170), .Z(n175) );
  NANDN U313 ( .A(n173), .B(n172), .Z(n174) );
  AND U314 ( .A(n175), .B(n174), .Z(n265) );
  XOR U315 ( .A(n266), .B(n265), .Z(n176) );
  XOR U316 ( .A(n267), .B(n176), .Z(n280) );
  NANDN U317 ( .A(n178), .B(n177), .Z(n182) );
  NANDN U318 ( .A(n180), .B(n179), .Z(n181) );
  NAND U319 ( .A(n182), .B(n181), .Z(n250) );
  NANDN U320 ( .A(n184), .B(n183), .Z(n188) );
  NANDN U321 ( .A(n186), .B(n185), .Z(n187) );
  NAND U322 ( .A(n188), .B(n187), .Z(n249) );
  NANDN U323 ( .A(n190), .B(n189), .Z(n194) );
  NANDN U324 ( .A(n192), .B(n191), .Z(n193) );
  AND U325 ( .A(n194), .B(n193), .Z(n248) );
  XOR U326 ( .A(n249), .B(n248), .Z(n195) );
  XNOR U327 ( .A(n250), .B(n195), .Z(n279) );
  NANDN U328 ( .A(n197), .B(n196), .Z(n201) );
  NANDN U329 ( .A(n199), .B(n198), .Z(n200) );
  NAND U330 ( .A(n201), .B(n200), .Z(n234) );
  XOR U331 ( .A(n233), .B(n232), .Z(n209) );
  XOR U332 ( .A(n234), .B(n209), .Z(n278) );
  XOR U333 ( .A(n279), .B(n278), .Z(n210) );
  XOR U334 ( .A(n280), .B(n210), .Z(n257) );
  OR U335 ( .A(n215), .B(n214), .Z(n219) );
  AND U336 ( .A(n215), .B(n214), .Z(n216) );
  OR U337 ( .A(n217), .B(n216), .Z(n218) );
  AND U338 ( .A(n219), .B(n218), .Z(n247) );
  XOR U339 ( .A(n247), .B(n246), .Z(n223) );
  XOR U340 ( .A(n245), .B(n223), .Z(n256) );
  IV U341 ( .A(n256), .Z(n254) );
  XOR U342 ( .A(n282), .B(n283), .Z(n230) );
  XNOR U343 ( .A(n284), .B(n230), .Z(o[1]) );
  XOR U344 ( .A(oglobal[2]), .B(n290), .Z(n294) );
  NANDN U345 ( .A(n233), .B(n232), .Z(n237) );
  ANDN U346 ( .B(n233), .A(n232), .Z(n235) );
  OR U347 ( .A(n235), .B(n234), .Z(n236) );
  AND U348 ( .A(n237), .B(n236), .Z(n296) );
  NANDN U349 ( .A(n239), .B(n238), .Z(n243) );
  ANDN U350 ( .B(n239), .A(n238), .Z(n241) );
  OR U351 ( .A(n241), .B(n240), .Z(n242) );
  AND U352 ( .A(n243), .B(n242), .Z(n295) );
  XNOR U353 ( .A(n296), .B(n295), .Z(n244) );
  XOR U354 ( .A(n294), .B(n244), .Z(n288) );
  XOR U355 ( .A(n287), .B(n286), .Z(n289) );
  XOR U356 ( .A(n288), .B(n289), .Z(n304) );
  NANDN U357 ( .A(n254), .B(n255), .Z(n260) );
  NOR U358 ( .A(n256), .B(n255), .Z(n258) );
  NANDN U359 ( .A(n258), .B(n257), .Z(n259) );
  AND U360 ( .A(n260), .B(n259), .Z(n302) );
  XNOR U361 ( .A(n303), .B(n302), .Z(n261) );
  XOR U362 ( .A(n304), .B(n261), .Z(n307) );
  NANDN U363 ( .A(n266), .B(n265), .Z(n270) );
  ANDN U364 ( .B(n266), .A(n265), .Z(n268) );
  OR U365 ( .A(n268), .B(n267), .Z(n269) );
  AND U366 ( .A(n270), .B(n269), .Z(n293) );
  XNOR U367 ( .A(n293), .B(n292), .Z(n274) );
  XOR U368 ( .A(n291), .B(n274), .Z(n298) );
  XNOR U369 ( .A(n300), .B(n299), .Z(n281) );
  XOR U370 ( .A(n298), .B(n281), .Z(n306) );
  XNOR U371 ( .A(n306), .B(n305), .Z(n285) );
  XNOR U372 ( .A(n307), .B(n285), .Z(o[2]) );
  AND U373 ( .A(oglobal[2]), .B(n290), .Z(n309) );
  XOR U374 ( .A(n309), .B(oglobal[3]), .Z(n311) );
  XNOR U375 ( .A(n312), .B(n310), .Z(n297) );
  XOR U376 ( .A(n311), .B(n297), .Z(n314) );
  XOR U377 ( .A(n314), .B(n315), .Z(n301) );
  XOR U378 ( .A(n313), .B(n301), .Z(n317) );
  XNOR U379 ( .A(n318), .B(n316), .Z(n308) );
  XNOR U380 ( .A(n317), .B(n308), .Z(o[3]) );
  AND U381 ( .A(n309), .B(oglobal[3]), .Z(n323) );
  XOR U382 ( .A(oglobal[4]), .B(n323), .Z(n325) );
  XNOR U383 ( .A(n325), .B(n324), .Z(n322) );
  XOR U384 ( .A(n321), .B(n320), .Z(n319) );
  XNOR U385 ( .A(n322), .B(n319), .Z(o[4]) );
  NAND U386 ( .A(n323), .B(oglobal[4]), .Z(n327) );
  NAND U387 ( .A(n325), .B(n324), .Z(n326) );
  NAND U388 ( .A(n327), .B(n326), .Z(n329) );
  XOR U389 ( .A(n330), .B(n329), .Z(n328) );
  XNOR U390 ( .A(oglobal[5]), .B(n328), .Z(o[5]) );
  XNOR U391 ( .A(n331), .B(oglobal[6]), .Z(o[6]) );
  ANDN U392 ( .B(oglobal[6]), .A(n331), .Z(n332) );
  XOR U393 ( .A(n332), .B(oglobal[7]), .Z(o[7]) );
  AND U394 ( .A(n332), .B(oglobal[7]), .Z(n333) );
  XOR U395 ( .A(n333), .B(oglobal[8]), .Z(o[8]) );
  AND U396 ( .A(n333), .B(oglobal[8]), .Z(n334) );
  XOR U397 ( .A(oglobal[9]), .B(n334), .Z(o[9]) );
endmodule

