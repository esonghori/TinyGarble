
module Mult ( clk, rst, a, b, mult_func, c_mult );
  input [31:0] a;
  input [31:0] b;
  input [3:0] mult_func;
  output [31:0] c_mult;
  input clk, rst;
  wire   N118, N119, N120, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, \U3/U1/Z_0 ,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, \r60/A2[30] ,
         \r60/A2[31] , \r60/A2[32] , \r60/A2[33] , \r60/A2[34] , \r60/A2[35] ,
         \r60/A2[36] , \r60/A2[37] , \r60/A2[38] , \r60/A2[39] , \r60/A2[40] ,
         \r60/A2[41] , \r60/A2[42] , \r60/A2[43] , \r60/A2[44] , \r60/A2[45] ,
         \r60/A2[46] , \r60/A2[47] , \r60/A2[48] , \r60/A2[49] , \r60/A2[50] ,
         \r60/A2[51] , \r60/A2[52] , \r60/A2[53] , \r60/A2[54] , \r60/A2[55] ,
         \r60/A2[56] , \r60/A2[57] , \r60/A2[58] , \r60/A2[59] , \r60/A2[60] ,
         \r60/A2[61] , \r60/A1[30] , \r60/A1[31] , \r60/A1[32] , \r60/A1[33] ,
         \r60/A1[34] , \r60/A1[35] , \r60/A1[36] , \r60/A1[37] , \r60/A1[38] ,
         \r60/A1[39] , \r60/A1[40] , \r60/A1[41] , \r60/A1[42] , \r60/A1[43] ,
         \r60/A1[44] , \r60/A1[45] , \r60/A1[46] , \r60/A1[47] , \r60/A1[48] ,
         \r60/A1[49] , \r60/A1[50] , \r60/A1[51] , \r60/A1[52] , \r60/A1[53] ,
         \r60/A1[54] , \r60/A1[55] , \r60/A1[56] , \r60/A1[57] , \r60/A1[58] ,
         \r60/A1[59] , \r60/A1[60] , \r60/A1[61] , \r60/ZB , \r60/ZA ,
         \r60/QB , \r60/QA , \r60/SUMB[16][1] , \r60/SUMB[16][2] ,
         \r60/SUMB[16][3] , \r60/SUMB[16][4] , \r60/SUMB[16][5] ,
         \r60/SUMB[16][6] , \r60/SUMB[16][7] , \r60/SUMB[16][8] ,
         \r60/SUMB[16][9] , \r60/SUMB[16][10] , \r60/SUMB[16][11] ,
         \r60/SUMB[16][12] , \r60/SUMB[16][13] , \r60/SUMB[16][14] ,
         \r60/SUMB[16][15] , \r60/SUMB[16][16] , \r60/SUMB[16][17] ,
         \r60/SUMB[16][18] , \r60/SUMB[16][19] , \r60/SUMB[16][20] ,
         \r60/SUMB[16][21] , \r60/SUMB[16][22] , \r60/SUMB[16][23] ,
         \r60/SUMB[16][24] , \r60/SUMB[16][25] , \r60/SUMB[16][26] ,
         \r60/SUMB[16][27] , \r60/SUMB[16][28] , \r60/SUMB[16][29] ,
         \r60/SUMB[16][30] , \r60/SUMB[17][1] , \r60/SUMB[17][2] ,
         \r60/SUMB[17][3] , \r60/SUMB[17][4] , \r60/SUMB[17][5] ,
         \r60/SUMB[17][6] , \r60/SUMB[17][7] , \r60/SUMB[17][8] ,
         \r60/SUMB[17][9] , \r60/SUMB[17][10] , \r60/SUMB[17][11] ,
         \r60/SUMB[17][12] , \r60/SUMB[17][13] , \r60/SUMB[17][14] ,
         \r60/SUMB[17][15] , \r60/SUMB[17][16] , \r60/SUMB[17][17] ,
         \r60/SUMB[17][18] , \r60/SUMB[17][19] , \r60/SUMB[17][20] ,
         \r60/SUMB[17][21] , \r60/SUMB[17][22] , \r60/SUMB[17][23] ,
         \r60/SUMB[17][24] , \r60/SUMB[17][25] , \r60/SUMB[17][26] ,
         \r60/SUMB[17][27] , \r60/SUMB[17][28] , \r60/SUMB[17][29] ,
         \r60/SUMB[17][30] , \r60/SUMB[18][1] , \r60/SUMB[18][2] ,
         \r60/SUMB[18][3] , \r60/SUMB[18][4] , \r60/SUMB[18][5] ,
         \r60/SUMB[18][6] , \r60/SUMB[18][7] , \r60/SUMB[18][8] ,
         \r60/SUMB[18][9] , \r60/SUMB[18][10] , \r60/SUMB[18][11] ,
         \r60/SUMB[18][12] , \r60/SUMB[18][13] , \r60/SUMB[18][14] ,
         \r60/SUMB[18][15] , \r60/SUMB[18][16] , \r60/SUMB[18][17] ,
         \r60/SUMB[18][18] , \r60/SUMB[18][19] , \r60/SUMB[18][20] ,
         \r60/SUMB[18][21] , \r60/SUMB[18][22] , \r60/SUMB[18][23] ,
         \r60/SUMB[18][24] , \r60/SUMB[18][25] , \r60/SUMB[18][26] ,
         \r60/SUMB[18][27] , \r60/SUMB[18][28] , \r60/SUMB[18][29] ,
         \r60/SUMB[18][30] , \r60/SUMB[19][1] , \r60/SUMB[19][2] ,
         \r60/SUMB[19][3] , \r60/SUMB[19][4] , \r60/SUMB[19][5] ,
         \r60/SUMB[19][6] , \r60/SUMB[19][7] , \r60/SUMB[19][8] ,
         \r60/SUMB[19][9] , \r60/SUMB[19][10] , \r60/SUMB[19][11] ,
         \r60/SUMB[19][12] , \r60/SUMB[19][13] , \r60/SUMB[19][14] ,
         \r60/SUMB[19][15] , \r60/SUMB[19][16] , \r60/SUMB[19][17] ,
         \r60/SUMB[19][18] , \r60/SUMB[19][19] , \r60/SUMB[19][20] ,
         \r60/SUMB[19][21] , \r60/SUMB[19][22] , \r60/SUMB[19][23] ,
         \r60/SUMB[19][24] , \r60/SUMB[19][25] , \r60/SUMB[19][26] ,
         \r60/SUMB[19][27] , \r60/SUMB[19][28] , \r60/SUMB[19][29] ,
         \r60/SUMB[19][30] , \r60/SUMB[20][1] , \r60/SUMB[20][2] ,
         \r60/SUMB[20][3] , \r60/SUMB[20][4] , \r60/SUMB[20][5] ,
         \r60/SUMB[20][6] , \r60/SUMB[20][7] , \r60/SUMB[20][8] ,
         \r60/SUMB[20][9] , \r60/SUMB[20][10] , \r60/SUMB[20][11] ,
         \r60/SUMB[20][12] , \r60/SUMB[20][13] , \r60/SUMB[20][14] ,
         \r60/SUMB[20][15] , \r60/SUMB[20][16] , \r60/SUMB[20][17] ,
         \r60/SUMB[20][18] , \r60/SUMB[20][19] , \r60/SUMB[20][20] ,
         \r60/SUMB[20][21] , \r60/SUMB[20][22] , \r60/SUMB[20][23] ,
         \r60/SUMB[20][24] , \r60/SUMB[20][25] , \r60/SUMB[20][26] ,
         \r60/SUMB[20][27] , \r60/SUMB[20][28] , \r60/SUMB[20][29] ,
         \r60/SUMB[20][30] , \r60/SUMB[21][1] , \r60/SUMB[21][2] ,
         \r60/SUMB[21][3] , \r60/SUMB[21][4] , \r60/SUMB[21][5] ,
         \r60/SUMB[21][6] , \r60/SUMB[21][7] , \r60/SUMB[21][8] ,
         \r60/SUMB[21][9] , \r60/SUMB[21][10] , \r60/SUMB[21][11] ,
         \r60/SUMB[21][12] , \r60/SUMB[21][13] , \r60/SUMB[21][14] ,
         \r60/SUMB[21][15] , \r60/SUMB[21][16] , \r60/SUMB[21][17] ,
         \r60/SUMB[21][18] , \r60/SUMB[21][19] , \r60/SUMB[21][20] ,
         \r60/SUMB[21][21] , \r60/SUMB[21][22] , \r60/SUMB[21][23] ,
         \r60/SUMB[21][24] , \r60/SUMB[21][25] , \r60/SUMB[21][26] ,
         \r60/SUMB[21][27] , \r60/SUMB[21][28] , \r60/SUMB[21][29] ,
         \r60/SUMB[21][30] , \r60/SUMB[22][1] , \r60/SUMB[22][2] ,
         \r60/SUMB[22][3] , \r60/SUMB[22][4] , \r60/SUMB[22][5] ,
         \r60/SUMB[22][6] , \r60/SUMB[22][7] , \r60/SUMB[22][8] ,
         \r60/SUMB[22][9] , \r60/SUMB[22][10] , \r60/SUMB[22][11] ,
         \r60/SUMB[22][12] , \r60/SUMB[22][13] , \r60/SUMB[22][14] ,
         \r60/SUMB[22][15] , \r60/SUMB[22][16] , \r60/SUMB[22][17] ,
         \r60/SUMB[22][18] , \r60/SUMB[22][19] , \r60/SUMB[22][20] ,
         \r60/SUMB[22][21] , \r60/SUMB[22][22] , \r60/SUMB[22][23] ,
         \r60/SUMB[22][24] , \r60/SUMB[22][25] , \r60/SUMB[22][26] ,
         \r60/SUMB[22][27] , \r60/SUMB[22][28] , \r60/SUMB[22][29] ,
         \r60/SUMB[22][30] , \r60/SUMB[23][1] , \r60/SUMB[23][2] ,
         \r60/SUMB[23][3] , \r60/SUMB[23][4] , \r60/SUMB[23][5] ,
         \r60/SUMB[23][6] , \r60/SUMB[23][7] , \r60/SUMB[23][8] ,
         \r60/SUMB[23][9] , \r60/SUMB[23][10] , \r60/SUMB[23][11] ,
         \r60/SUMB[23][12] , \r60/SUMB[23][13] , \r60/SUMB[23][14] ,
         \r60/SUMB[23][15] , \r60/SUMB[23][16] , \r60/SUMB[23][17] ,
         \r60/SUMB[23][18] , \r60/SUMB[23][19] , \r60/SUMB[23][20] ,
         \r60/SUMB[23][21] , \r60/SUMB[23][22] , \r60/SUMB[23][23] ,
         \r60/SUMB[23][24] , \r60/SUMB[23][25] , \r60/SUMB[23][26] ,
         \r60/SUMB[23][27] , \r60/SUMB[23][28] , \r60/SUMB[23][29] ,
         \r60/SUMB[23][30] , \r60/SUMB[24][1] , \r60/SUMB[24][2] ,
         \r60/SUMB[24][3] , \r60/SUMB[24][4] , \r60/SUMB[24][5] ,
         \r60/SUMB[24][6] , \r60/SUMB[24][7] , \r60/SUMB[24][8] ,
         \r60/SUMB[24][9] , \r60/SUMB[24][10] , \r60/SUMB[24][11] ,
         \r60/SUMB[24][12] , \r60/SUMB[24][13] , \r60/SUMB[24][14] ,
         \r60/SUMB[24][15] , \r60/SUMB[24][16] , \r60/SUMB[24][17] ,
         \r60/SUMB[24][18] , \r60/SUMB[24][19] , \r60/SUMB[24][20] ,
         \r60/SUMB[24][21] , \r60/SUMB[24][22] , \r60/SUMB[24][23] ,
         \r60/SUMB[24][24] , \r60/SUMB[24][25] , \r60/SUMB[24][26] ,
         \r60/SUMB[24][27] , \r60/SUMB[24][28] , \r60/SUMB[24][29] ,
         \r60/SUMB[24][30] , \r60/SUMB[25][1] , \r60/SUMB[25][2] ,
         \r60/SUMB[25][3] , \r60/SUMB[25][4] , \r60/SUMB[25][5] ,
         \r60/SUMB[25][6] , \r60/SUMB[25][7] , \r60/SUMB[25][8] ,
         \r60/SUMB[25][9] , \r60/SUMB[25][10] , \r60/SUMB[25][11] ,
         \r60/SUMB[25][12] , \r60/SUMB[25][13] , \r60/SUMB[25][14] ,
         \r60/SUMB[25][15] , \r60/SUMB[25][16] , \r60/SUMB[25][17] ,
         \r60/SUMB[25][18] , \r60/SUMB[25][19] , \r60/SUMB[25][20] ,
         \r60/SUMB[25][21] , \r60/SUMB[25][22] , \r60/SUMB[25][23] ,
         \r60/SUMB[25][24] , \r60/SUMB[25][25] , \r60/SUMB[25][26] ,
         \r60/SUMB[25][27] , \r60/SUMB[25][28] , \r60/SUMB[25][29] ,
         \r60/SUMB[25][30] , \r60/SUMB[26][1] , \r60/SUMB[26][2] ,
         \r60/SUMB[26][3] , \r60/SUMB[26][4] , \r60/SUMB[26][5] ,
         \r60/SUMB[26][6] , \r60/SUMB[26][7] , \r60/SUMB[26][8] ,
         \r60/SUMB[26][9] , \r60/SUMB[26][10] , \r60/SUMB[26][11] ,
         \r60/SUMB[26][12] , \r60/SUMB[26][13] , \r60/SUMB[26][14] ,
         \r60/SUMB[26][15] , \r60/SUMB[26][16] , \r60/SUMB[26][17] ,
         \r60/SUMB[26][18] , \r60/SUMB[26][19] , \r60/SUMB[26][20] ,
         \r60/SUMB[26][21] , \r60/SUMB[26][22] , \r60/SUMB[26][23] ,
         \r60/SUMB[26][24] , \r60/SUMB[26][25] , \r60/SUMB[26][26] ,
         \r60/SUMB[26][27] , \r60/SUMB[26][28] , \r60/SUMB[26][29] ,
         \r60/SUMB[26][30] , \r60/SUMB[27][1] , \r60/SUMB[27][2] ,
         \r60/SUMB[27][3] , \r60/SUMB[27][4] , \r60/SUMB[27][5] ,
         \r60/SUMB[27][6] , \r60/SUMB[27][7] , \r60/SUMB[27][8] ,
         \r60/SUMB[27][9] , \r60/SUMB[27][10] , \r60/SUMB[27][11] ,
         \r60/SUMB[27][12] , \r60/SUMB[27][13] , \r60/SUMB[27][14] ,
         \r60/SUMB[27][15] , \r60/SUMB[27][16] , \r60/SUMB[27][17] ,
         \r60/SUMB[27][18] , \r60/SUMB[27][19] , \r60/SUMB[27][20] ,
         \r60/SUMB[27][21] , \r60/SUMB[27][22] , \r60/SUMB[27][23] ,
         \r60/SUMB[27][24] , \r60/SUMB[27][25] , \r60/SUMB[27][26] ,
         \r60/SUMB[27][27] , \r60/SUMB[27][28] , \r60/SUMB[27][29] ,
         \r60/SUMB[27][30] , \r60/SUMB[28][1] , \r60/SUMB[28][2] ,
         \r60/SUMB[28][3] , \r60/SUMB[28][4] , \r60/SUMB[28][5] ,
         \r60/SUMB[28][6] , \r60/SUMB[28][7] , \r60/SUMB[28][8] ,
         \r60/SUMB[28][9] , \r60/SUMB[28][10] , \r60/SUMB[28][11] ,
         \r60/SUMB[28][12] , \r60/SUMB[28][13] , \r60/SUMB[28][14] ,
         \r60/SUMB[28][15] , \r60/SUMB[28][16] , \r60/SUMB[28][17] ,
         \r60/SUMB[28][18] , \r60/SUMB[28][19] , \r60/SUMB[28][20] ,
         \r60/SUMB[28][21] , \r60/SUMB[28][22] , \r60/SUMB[28][23] ,
         \r60/SUMB[28][24] , \r60/SUMB[28][25] , \r60/SUMB[28][26] ,
         \r60/SUMB[28][27] , \r60/SUMB[28][28] , \r60/SUMB[28][29] ,
         \r60/SUMB[28][30] , \r60/SUMB[29][1] , \r60/SUMB[29][2] ,
         \r60/SUMB[29][3] , \r60/SUMB[29][4] , \r60/SUMB[29][5] ,
         \r60/SUMB[29][6] , \r60/SUMB[29][7] , \r60/SUMB[29][8] ,
         \r60/SUMB[29][9] , \r60/SUMB[29][10] , \r60/SUMB[29][11] ,
         \r60/SUMB[29][12] , \r60/SUMB[29][13] , \r60/SUMB[29][14] ,
         \r60/SUMB[29][15] , \r60/SUMB[29][16] , \r60/SUMB[29][17] ,
         \r60/SUMB[29][18] , \r60/SUMB[29][19] , \r60/SUMB[29][20] ,
         \r60/SUMB[29][21] , \r60/SUMB[29][22] , \r60/SUMB[29][23] ,
         \r60/SUMB[29][24] , \r60/SUMB[29][25] , \r60/SUMB[29][26] ,
         \r60/SUMB[29][27] , \r60/SUMB[29][28] , \r60/SUMB[29][29] ,
         \r60/SUMB[29][30] , \r60/SUMB[30][1] , \r60/SUMB[30][2] ,
         \r60/SUMB[30][3] , \r60/SUMB[30][4] , \r60/SUMB[30][5] ,
         \r60/SUMB[30][6] , \r60/SUMB[30][7] , \r60/SUMB[30][8] ,
         \r60/SUMB[30][9] , \r60/SUMB[30][10] , \r60/SUMB[30][11] ,
         \r60/SUMB[30][12] , \r60/SUMB[30][13] , \r60/SUMB[30][14] ,
         \r60/SUMB[30][15] , \r60/SUMB[30][16] , \r60/SUMB[30][17] ,
         \r60/SUMB[30][18] , \r60/SUMB[30][19] , \r60/SUMB[30][20] ,
         \r60/SUMB[30][21] , \r60/SUMB[30][22] , \r60/SUMB[30][23] ,
         \r60/SUMB[30][24] , \r60/SUMB[30][25] , \r60/SUMB[30][26] ,
         \r60/SUMB[30][27] , \r60/SUMB[30][28] , \r60/SUMB[30][29] ,
         \r60/SUMB[30][30] , \r60/SUMB[31][0] , \r60/SUMB[31][1] ,
         \r60/SUMB[31][2] , \r60/SUMB[31][3] , \r60/SUMB[31][4] ,
         \r60/SUMB[31][5] , \r60/SUMB[31][6] , \r60/SUMB[31][7] ,
         \r60/SUMB[31][8] , \r60/SUMB[31][9] , \r60/SUMB[31][10] ,
         \r60/SUMB[31][11] , \r60/SUMB[31][12] , \r60/SUMB[31][13] ,
         \r60/SUMB[31][14] , \r60/SUMB[31][15] , \r60/SUMB[31][16] ,
         \r60/SUMB[31][17] , \r60/SUMB[31][18] , \r60/SUMB[31][19] ,
         \r60/SUMB[31][20] , \r60/SUMB[31][21] , \r60/SUMB[31][22] ,
         \r60/SUMB[31][23] , \r60/SUMB[31][24] , \r60/SUMB[31][25] ,
         \r60/SUMB[31][26] , \r60/SUMB[31][27] , \r60/SUMB[31][28] ,
         \r60/SUMB[31][29] , \r60/SUMB[31][30] , \r60/SUMB[31][31] ,
         \r60/CARRYB[16][0] , \r60/CARRYB[16][1] , \r60/CARRYB[16][2] ,
         \r60/CARRYB[16][3] , \r60/CARRYB[16][4] , \r60/CARRYB[16][5] ,
         \r60/CARRYB[16][6] , \r60/CARRYB[16][7] , \r60/CARRYB[16][8] ,
         \r60/CARRYB[16][9] , \r60/CARRYB[16][10] , \r60/CARRYB[16][11] ,
         \r60/CARRYB[16][12] , \r60/CARRYB[16][13] , \r60/CARRYB[16][14] ,
         \r60/CARRYB[16][15] , \r60/CARRYB[16][16] , \r60/CARRYB[16][17] ,
         \r60/CARRYB[16][18] , \r60/CARRYB[16][19] , \r60/CARRYB[16][20] ,
         \r60/CARRYB[16][21] , \r60/CARRYB[16][22] , \r60/CARRYB[16][23] ,
         \r60/CARRYB[16][24] , \r60/CARRYB[16][25] , \r60/CARRYB[16][26] ,
         \r60/CARRYB[16][27] , \r60/CARRYB[16][28] , \r60/CARRYB[16][29] ,
         \r60/CARRYB[16][30] , \r60/CARRYB[17][0] , \r60/CARRYB[17][1] ,
         \r60/CARRYB[17][2] , \r60/CARRYB[17][3] , \r60/CARRYB[17][4] ,
         \r60/CARRYB[17][5] , \r60/CARRYB[17][6] , \r60/CARRYB[17][7] ,
         \r60/CARRYB[17][8] , \r60/CARRYB[17][9] , \r60/CARRYB[17][10] ,
         \r60/CARRYB[17][11] , \r60/CARRYB[17][12] , \r60/CARRYB[17][13] ,
         \r60/CARRYB[17][14] , \r60/CARRYB[17][15] , \r60/CARRYB[17][16] ,
         \r60/CARRYB[17][17] , \r60/CARRYB[17][18] , \r60/CARRYB[17][19] ,
         \r60/CARRYB[17][20] , \r60/CARRYB[17][21] , \r60/CARRYB[17][22] ,
         \r60/CARRYB[17][23] , \r60/CARRYB[17][24] , \r60/CARRYB[17][25] ,
         \r60/CARRYB[17][26] , \r60/CARRYB[17][27] , \r60/CARRYB[17][28] ,
         \r60/CARRYB[17][29] , \r60/CARRYB[17][30] , \r60/CARRYB[18][0] ,
         \r60/CARRYB[18][1] , \r60/CARRYB[18][2] , \r60/CARRYB[18][3] ,
         \r60/CARRYB[18][4] , \r60/CARRYB[18][5] , \r60/CARRYB[18][6] ,
         \r60/CARRYB[18][7] , \r60/CARRYB[18][8] , \r60/CARRYB[18][9] ,
         \r60/CARRYB[18][10] , \r60/CARRYB[18][11] , \r60/CARRYB[18][12] ,
         \r60/CARRYB[18][13] , \r60/CARRYB[18][14] , \r60/CARRYB[18][15] ,
         \r60/CARRYB[18][16] , \r60/CARRYB[18][17] , \r60/CARRYB[18][18] ,
         \r60/CARRYB[18][19] , \r60/CARRYB[18][20] , \r60/CARRYB[18][21] ,
         \r60/CARRYB[18][22] , \r60/CARRYB[18][23] , \r60/CARRYB[18][24] ,
         \r60/CARRYB[18][25] , \r60/CARRYB[18][26] , \r60/CARRYB[18][27] ,
         \r60/CARRYB[18][28] , \r60/CARRYB[18][29] , \r60/CARRYB[18][30] ,
         \r60/CARRYB[19][0] , \r60/CARRYB[19][1] , \r60/CARRYB[19][2] ,
         \r60/CARRYB[19][3] , \r60/CARRYB[19][4] , \r60/CARRYB[19][5] ,
         \r60/CARRYB[19][6] , \r60/CARRYB[19][7] , \r60/CARRYB[19][8] ,
         \r60/CARRYB[19][9] , \r60/CARRYB[19][10] , \r60/CARRYB[19][11] ,
         \r60/CARRYB[19][12] , \r60/CARRYB[19][13] , \r60/CARRYB[19][14] ,
         \r60/CARRYB[19][15] , \r60/CARRYB[19][16] , \r60/CARRYB[19][17] ,
         \r60/CARRYB[19][18] , \r60/CARRYB[19][19] , \r60/CARRYB[19][20] ,
         \r60/CARRYB[19][21] , \r60/CARRYB[19][22] , \r60/CARRYB[19][23] ,
         \r60/CARRYB[19][24] , \r60/CARRYB[19][25] , \r60/CARRYB[19][26] ,
         \r60/CARRYB[19][27] , \r60/CARRYB[19][28] , \r60/CARRYB[19][29] ,
         \r60/CARRYB[19][30] , \r60/CARRYB[20][0] , \r60/CARRYB[20][1] ,
         \r60/CARRYB[20][2] , \r60/CARRYB[20][3] , \r60/CARRYB[20][4] ,
         \r60/CARRYB[20][5] , \r60/CARRYB[20][6] , \r60/CARRYB[20][7] ,
         \r60/CARRYB[20][8] , \r60/CARRYB[20][9] , \r60/CARRYB[20][10] ,
         \r60/CARRYB[20][11] , \r60/CARRYB[20][12] , \r60/CARRYB[20][13] ,
         \r60/CARRYB[20][14] , \r60/CARRYB[20][15] , \r60/CARRYB[20][16] ,
         \r60/CARRYB[20][17] , \r60/CARRYB[20][18] , \r60/CARRYB[20][19] ,
         \r60/CARRYB[20][20] , \r60/CARRYB[20][21] , \r60/CARRYB[20][22] ,
         \r60/CARRYB[20][23] , \r60/CARRYB[20][24] , \r60/CARRYB[20][25] ,
         \r60/CARRYB[20][26] , \r60/CARRYB[20][27] , \r60/CARRYB[20][28] ,
         \r60/CARRYB[20][29] , \r60/CARRYB[20][30] , \r60/CARRYB[21][0] ,
         \r60/CARRYB[21][1] , \r60/CARRYB[21][2] , \r60/CARRYB[21][3] ,
         \r60/CARRYB[21][4] , \r60/CARRYB[21][5] , \r60/CARRYB[21][6] ,
         \r60/CARRYB[21][7] , \r60/CARRYB[21][8] , \r60/CARRYB[21][9] ,
         \r60/CARRYB[21][10] , \r60/CARRYB[21][11] , \r60/CARRYB[21][12] ,
         \r60/CARRYB[21][13] , \r60/CARRYB[21][14] , \r60/CARRYB[21][15] ,
         \r60/CARRYB[21][16] , \r60/CARRYB[21][17] , \r60/CARRYB[21][18] ,
         \r60/CARRYB[21][19] , \r60/CARRYB[21][20] , \r60/CARRYB[21][21] ,
         \r60/CARRYB[21][22] , \r60/CARRYB[21][23] , \r60/CARRYB[21][24] ,
         \r60/CARRYB[21][25] , \r60/CARRYB[21][26] , \r60/CARRYB[21][27] ,
         \r60/CARRYB[21][28] , \r60/CARRYB[21][29] , \r60/CARRYB[21][30] ,
         \r60/CARRYB[22][0] , \r60/CARRYB[22][1] , \r60/CARRYB[22][2] ,
         \r60/CARRYB[22][3] , \r60/CARRYB[22][4] , \r60/CARRYB[22][5] ,
         \r60/CARRYB[22][6] , \r60/CARRYB[22][7] , \r60/CARRYB[22][8] ,
         \r60/CARRYB[22][9] , \r60/CARRYB[22][10] , \r60/CARRYB[22][11] ,
         \r60/CARRYB[22][12] , \r60/CARRYB[22][13] , \r60/CARRYB[22][14] ,
         \r60/CARRYB[22][15] , \r60/CARRYB[22][16] , \r60/CARRYB[22][17] ,
         \r60/CARRYB[22][18] , \r60/CARRYB[22][19] , \r60/CARRYB[22][20] ,
         \r60/CARRYB[22][21] , \r60/CARRYB[22][22] , \r60/CARRYB[22][23] ,
         \r60/CARRYB[22][24] , \r60/CARRYB[22][25] , \r60/CARRYB[22][26] ,
         \r60/CARRYB[22][27] , \r60/CARRYB[22][28] , \r60/CARRYB[22][29] ,
         \r60/CARRYB[22][30] , \r60/CARRYB[23][0] , \r60/CARRYB[23][1] ,
         \r60/CARRYB[23][2] , \r60/CARRYB[23][3] , \r60/CARRYB[23][4] ,
         \r60/CARRYB[23][5] , \r60/CARRYB[23][6] , \r60/CARRYB[23][7] ,
         \r60/CARRYB[23][8] , \r60/CARRYB[23][9] , \r60/CARRYB[23][10] ,
         \r60/CARRYB[23][11] , \r60/CARRYB[23][12] , \r60/CARRYB[23][13] ,
         \r60/CARRYB[23][14] , \r60/CARRYB[23][15] , \r60/CARRYB[23][16] ,
         \r60/CARRYB[23][17] , \r60/CARRYB[23][18] , \r60/CARRYB[23][19] ,
         \r60/CARRYB[23][20] , \r60/CARRYB[23][21] , \r60/CARRYB[23][22] ,
         \r60/CARRYB[23][23] , \r60/CARRYB[23][24] , \r60/CARRYB[23][25] ,
         \r60/CARRYB[23][26] , \r60/CARRYB[23][27] , \r60/CARRYB[23][28] ,
         \r60/CARRYB[23][29] , \r60/CARRYB[23][30] , \r60/CARRYB[24][0] ,
         \r60/CARRYB[24][1] , \r60/CARRYB[24][2] , \r60/CARRYB[24][3] ,
         \r60/CARRYB[24][4] , \r60/CARRYB[24][5] , \r60/CARRYB[24][6] ,
         \r60/CARRYB[24][7] , \r60/CARRYB[24][8] , \r60/CARRYB[24][9] ,
         \r60/CARRYB[24][10] , \r60/CARRYB[24][11] , \r60/CARRYB[24][12] ,
         \r60/CARRYB[24][13] , \r60/CARRYB[24][14] , \r60/CARRYB[24][15] ,
         \r60/CARRYB[24][16] , \r60/CARRYB[24][17] , \r60/CARRYB[24][18] ,
         \r60/CARRYB[24][19] , \r60/CARRYB[24][20] , \r60/CARRYB[24][21] ,
         \r60/CARRYB[24][22] , \r60/CARRYB[24][23] , \r60/CARRYB[24][24] ,
         \r60/CARRYB[24][25] , \r60/CARRYB[24][26] , \r60/CARRYB[24][27] ,
         \r60/CARRYB[24][28] , \r60/CARRYB[24][29] , \r60/CARRYB[24][30] ,
         \r60/CARRYB[25][0] , \r60/CARRYB[25][1] , \r60/CARRYB[25][2] ,
         \r60/CARRYB[25][3] , \r60/CARRYB[25][4] , \r60/CARRYB[25][5] ,
         \r60/CARRYB[25][6] , \r60/CARRYB[25][7] , \r60/CARRYB[25][8] ,
         \r60/CARRYB[25][9] , \r60/CARRYB[25][10] , \r60/CARRYB[25][11] ,
         \r60/CARRYB[25][12] , \r60/CARRYB[25][13] , \r60/CARRYB[25][14] ,
         \r60/CARRYB[25][15] , \r60/CARRYB[25][16] , \r60/CARRYB[25][17] ,
         \r60/CARRYB[25][18] , \r60/CARRYB[25][19] , \r60/CARRYB[25][20] ,
         \r60/CARRYB[25][21] , \r60/CARRYB[25][22] , \r60/CARRYB[25][23] ,
         \r60/CARRYB[25][24] , \r60/CARRYB[25][25] , \r60/CARRYB[25][26] ,
         \r60/CARRYB[25][27] , \r60/CARRYB[25][28] , \r60/CARRYB[25][29] ,
         \r60/CARRYB[25][30] , \r60/CARRYB[26][0] , \r60/CARRYB[26][1] ,
         \r60/CARRYB[26][2] , \r60/CARRYB[26][3] , \r60/CARRYB[26][4] ,
         \r60/CARRYB[26][5] , \r60/CARRYB[26][6] , \r60/CARRYB[26][7] ,
         \r60/CARRYB[26][8] , \r60/CARRYB[26][9] , \r60/CARRYB[26][10] ,
         \r60/CARRYB[26][11] , \r60/CARRYB[26][12] , \r60/CARRYB[26][13] ,
         \r60/CARRYB[26][14] , \r60/CARRYB[26][15] , \r60/CARRYB[26][16] ,
         \r60/CARRYB[26][17] , \r60/CARRYB[26][18] , \r60/CARRYB[26][19] ,
         \r60/CARRYB[26][20] , \r60/CARRYB[26][21] , \r60/CARRYB[26][22] ,
         \r60/CARRYB[26][23] , \r60/CARRYB[26][24] , \r60/CARRYB[26][25] ,
         \r60/CARRYB[26][26] , \r60/CARRYB[26][27] , \r60/CARRYB[26][28] ,
         \r60/CARRYB[26][29] , \r60/CARRYB[26][30] , \r60/CARRYB[27][0] ,
         \r60/CARRYB[27][1] , \r60/CARRYB[27][2] , \r60/CARRYB[27][3] ,
         \r60/CARRYB[27][4] , \r60/CARRYB[27][5] , \r60/CARRYB[27][6] ,
         \r60/CARRYB[27][7] , \r60/CARRYB[27][8] , \r60/CARRYB[27][9] ,
         \r60/CARRYB[27][10] , \r60/CARRYB[27][11] , \r60/CARRYB[27][12] ,
         \r60/CARRYB[27][13] , \r60/CARRYB[27][14] , \r60/CARRYB[27][15] ,
         \r60/CARRYB[27][16] , \r60/CARRYB[27][17] , \r60/CARRYB[27][18] ,
         \r60/CARRYB[27][19] , \r60/CARRYB[27][20] , \r60/CARRYB[27][21] ,
         \r60/CARRYB[27][22] , \r60/CARRYB[27][23] , \r60/CARRYB[27][24] ,
         \r60/CARRYB[27][25] , \r60/CARRYB[27][26] , \r60/CARRYB[27][27] ,
         \r60/CARRYB[27][28] , \r60/CARRYB[27][29] , \r60/CARRYB[27][30] ,
         \r60/CARRYB[28][0] , \r60/CARRYB[28][1] , \r60/CARRYB[28][2] ,
         \r60/CARRYB[28][3] , \r60/CARRYB[28][4] , \r60/CARRYB[28][5] ,
         \r60/CARRYB[28][6] , \r60/CARRYB[28][7] , \r60/CARRYB[28][8] ,
         \r60/CARRYB[28][9] , \r60/CARRYB[28][10] , \r60/CARRYB[28][11] ,
         \r60/CARRYB[28][12] , \r60/CARRYB[28][13] , \r60/CARRYB[28][14] ,
         \r60/CARRYB[28][15] , \r60/CARRYB[28][16] , \r60/CARRYB[28][17] ,
         \r60/CARRYB[28][18] , \r60/CARRYB[28][19] , \r60/CARRYB[28][20] ,
         \r60/CARRYB[28][21] , \r60/CARRYB[28][22] , \r60/CARRYB[28][23] ,
         \r60/CARRYB[28][24] , \r60/CARRYB[28][25] , \r60/CARRYB[28][26] ,
         \r60/CARRYB[28][27] , \r60/CARRYB[28][28] , \r60/CARRYB[28][29] ,
         \r60/CARRYB[28][30] , \r60/CARRYB[29][0] , \r60/CARRYB[29][1] ,
         \r60/CARRYB[29][2] , \r60/CARRYB[29][3] , \r60/CARRYB[29][4] ,
         \r60/CARRYB[29][5] , \r60/CARRYB[29][6] , \r60/CARRYB[29][7] ,
         \r60/CARRYB[29][8] , \r60/CARRYB[29][9] , \r60/CARRYB[29][10] ,
         \r60/CARRYB[29][11] , \r60/CARRYB[29][12] , \r60/CARRYB[29][13] ,
         \r60/CARRYB[29][14] , \r60/CARRYB[29][15] , \r60/CARRYB[29][16] ,
         \r60/CARRYB[29][17] , \r60/CARRYB[29][18] , \r60/CARRYB[29][19] ,
         \r60/CARRYB[29][20] , \r60/CARRYB[29][21] , \r60/CARRYB[29][22] ,
         \r60/CARRYB[29][23] , \r60/CARRYB[29][24] , \r60/CARRYB[29][25] ,
         \r60/CARRYB[29][26] , \r60/CARRYB[29][27] , \r60/CARRYB[29][28] ,
         \r60/CARRYB[29][29] , \r60/CARRYB[29][30] , \r60/CARRYB[30][0] ,
         \r60/CARRYB[30][1] , \r60/CARRYB[30][2] , \r60/CARRYB[30][3] ,
         \r60/CARRYB[30][4] , \r60/CARRYB[30][5] , \r60/CARRYB[30][6] ,
         \r60/CARRYB[30][7] , \r60/CARRYB[30][8] , \r60/CARRYB[30][9] ,
         \r60/CARRYB[30][10] , \r60/CARRYB[30][11] , \r60/CARRYB[30][12] ,
         \r60/CARRYB[30][13] , \r60/CARRYB[30][14] , \r60/CARRYB[30][15] ,
         \r60/CARRYB[30][16] , \r60/CARRYB[30][17] , \r60/CARRYB[30][18] ,
         \r60/CARRYB[30][19] , \r60/CARRYB[30][20] , \r60/CARRYB[30][21] ,
         \r60/CARRYB[30][22] , \r60/CARRYB[30][23] , \r60/CARRYB[30][24] ,
         \r60/CARRYB[30][25] , \r60/CARRYB[30][26] , \r60/CARRYB[30][27] ,
         \r60/CARRYB[30][28] , \r60/CARRYB[30][29] , \r60/CARRYB[30][30] ,
         \r60/CARRYB[31][0] , \r60/CARRYB[31][1] , \r60/CARRYB[31][2] ,
         \r60/CARRYB[31][3] , \r60/CARRYB[31][4] , \r60/CARRYB[31][5] ,
         \r60/CARRYB[31][6] , \r60/CARRYB[31][7] , \r60/CARRYB[31][8] ,
         \r60/CARRYB[31][9] , \r60/CARRYB[31][10] , \r60/CARRYB[31][11] ,
         \r60/CARRYB[31][12] , \r60/CARRYB[31][13] , \r60/CARRYB[31][14] ,
         \r60/CARRYB[31][15] , \r60/CARRYB[31][16] , \r60/CARRYB[31][17] ,
         \r60/CARRYB[31][18] , \r60/CARRYB[31][19] , \r60/CARRYB[31][20] ,
         \r60/CARRYB[31][21] , \r60/CARRYB[31][22] , \r60/CARRYB[31][23] ,
         \r60/CARRYB[31][24] , \r60/CARRYB[31][25] , \r60/CARRYB[31][26] ,
         \r60/CARRYB[31][27] , \r60/CARRYB[31][28] , \r60/CARRYB[31][29] ,
         \r60/CARRYB[31][30] , \r60/CARRYB[31][31] , \r60/SUMB[1][1] ,
         \r60/SUMB[1][2] , \r60/SUMB[1][3] , \r60/SUMB[1][4] ,
         \r60/SUMB[1][5] , \r60/SUMB[1][6] , \r60/SUMB[1][7] ,
         \r60/SUMB[1][8] , \r60/SUMB[1][9] , \r60/SUMB[1][10] ,
         \r60/SUMB[1][11] , \r60/SUMB[1][12] , \r60/SUMB[1][13] ,
         \r60/SUMB[1][14] , \r60/SUMB[1][15] , \r60/SUMB[1][16] ,
         \r60/SUMB[1][17] , \r60/SUMB[1][18] , \r60/SUMB[1][19] ,
         \r60/SUMB[1][20] , \r60/SUMB[1][21] , \r60/SUMB[1][22] ,
         \r60/SUMB[1][23] , \r60/SUMB[1][24] , \r60/SUMB[1][25] ,
         \r60/SUMB[1][26] , \r60/SUMB[1][27] , \r60/SUMB[1][28] ,
         \r60/SUMB[1][29] , \r60/SUMB[1][30] , \r60/SUMB[2][1] ,
         \r60/SUMB[2][2] , \r60/SUMB[2][3] , \r60/SUMB[2][4] ,
         \r60/SUMB[2][5] , \r60/SUMB[2][6] , \r60/SUMB[2][7] ,
         \r60/SUMB[2][8] , \r60/SUMB[2][9] , \r60/SUMB[2][10] ,
         \r60/SUMB[2][11] , \r60/SUMB[2][12] , \r60/SUMB[2][13] ,
         \r60/SUMB[2][14] , \r60/SUMB[2][15] , \r60/SUMB[2][16] ,
         \r60/SUMB[2][17] , \r60/SUMB[2][18] , \r60/SUMB[2][19] ,
         \r60/SUMB[2][20] , \r60/SUMB[2][21] , \r60/SUMB[2][22] ,
         \r60/SUMB[2][23] , \r60/SUMB[2][24] , \r60/SUMB[2][25] ,
         \r60/SUMB[2][26] , \r60/SUMB[2][27] , \r60/SUMB[2][28] ,
         \r60/SUMB[2][29] , \r60/SUMB[2][30] , \r60/SUMB[3][1] ,
         \r60/SUMB[3][2] , \r60/SUMB[3][3] , \r60/SUMB[3][4] ,
         \r60/SUMB[3][5] , \r60/SUMB[3][6] , \r60/SUMB[3][7] ,
         \r60/SUMB[3][8] , \r60/SUMB[3][9] , \r60/SUMB[3][10] ,
         \r60/SUMB[3][11] , \r60/SUMB[3][12] , \r60/SUMB[3][13] ,
         \r60/SUMB[3][14] , \r60/SUMB[3][15] , \r60/SUMB[3][16] ,
         \r60/SUMB[3][17] , \r60/SUMB[3][18] , \r60/SUMB[3][19] ,
         \r60/SUMB[3][20] , \r60/SUMB[3][21] , \r60/SUMB[3][22] ,
         \r60/SUMB[3][23] , \r60/SUMB[3][24] , \r60/SUMB[3][25] ,
         \r60/SUMB[3][26] , \r60/SUMB[3][27] , \r60/SUMB[3][28] ,
         \r60/SUMB[3][29] , \r60/SUMB[3][30] , \r60/SUMB[4][1] ,
         \r60/SUMB[4][2] , \r60/SUMB[4][3] , \r60/SUMB[4][4] ,
         \r60/SUMB[4][5] , \r60/SUMB[4][6] , \r60/SUMB[4][7] ,
         \r60/SUMB[4][8] , \r60/SUMB[4][9] , \r60/SUMB[4][10] ,
         \r60/SUMB[4][11] , \r60/SUMB[4][12] , \r60/SUMB[4][13] ,
         \r60/SUMB[4][14] , \r60/SUMB[4][15] , \r60/SUMB[4][16] ,
         \r60/SUMB[4][17] , \r60/SUMB[4][18] , \r60/SUMB[4][19] ,
         \r60/SUMB[4][20] , \r60/SUMB[4][21] , \r60/SUMB[4][22] ,
         \r60/SUMB[4][23] , \r60/SUMB[4][24] , \r60/SUMB[4][25] ,
         \r60/SUMB[4][26] , \r60/SUMB[4][27] , \r60/SUMB[4][28] ,
         \r60/SUMB[4][29] , \r60/SUMB[4][30] , \r60/SUMB[5][1] ,
         \r60/SUMB[5][2] , \r60/SUMB[5][3] , \r60/SUMB[5][4] ,
         \r60/SUMB[5][5] , \r60/SUMB[5][6] , \r60/SUMB[5][7] ,
         \r60/SUMB[5][8] , \r60/SUMB[5][9] , \r60/SUMB[5][10] ,
         \r60/SUMB[5][11] , \r60/SUMB[5][12] , \r60/SUMB[5][13] ,
         \r60/SUMB[5][14] , \r60/SUMB[5][15] , \r60/SUMB[5][16] ,
         \r60/SUMB[5][17] , \r60/SUMB[5][18] , \r60/SUMB[5][19] ,
         \r60/SUMB[5][20] , \r60/SUMB[5][21] , \r60/SUMB[5][22] ,
         \r60/SUMB[5][23] , \r60/SUMB[5][24] , \r60/SUMB[5][25] ,
         \r60/SUMB[5][26] , \r60/SUMB[5][27] , \r60/SUMB[5][28] ,
         \r60/SUMB[5][29] , \r60/SUMB[5][30] , \r60/SUMB[6][1] ,
         \r60/SUMB[6][2] , \r60/SUMB[6][3] , \r60/SUMB[6][4] ,
         \r60/SUMB[6][5] , \r60/SUMB[6][6] , \r60/SUMB[6][7] ,
         \r60/SUMB[6][8] , \r60/SUMB[6][9] , \r60/SUMB[6][10] ,
         \r60/SUMB[6][11] , \r60/SUMB[6][12] , \r60/SUMB[6][13] ,
         \r60/SUMB[6][14] , \r60/SUMB[6][15] , \r60/SUMB[6][16] ,
         \r60/SUMB[6][17] , \r60/SUMB[6][18] , \r60/SUMB[6][19] ,
         \r60/SUMB[6][20] , \r60/SUMB[6][21] , \r60/SUMB[6][22] ,
         \r60/SUMB[6][23] , \r60/SUMB[6][24] , \r60/SUMB[6][25] ,
         \r60/SUMB[6][26] , \r60/SUMB[6][27] , \r60/SUMB[6][28] ,
         \r60/SUMB[6][29] , \r60/SUMB[6][30] , \r60/SUMB[7][1] ,
         \r60/SUMB[7][2] , \r60/SUMB[7][3] , \r60/SUMB[7][4] ,
         \r60/SUMB[7][5] , \r60/SUMB[7][6] , \r60/SUMB[7][7] ,
         \r60/SUMB[7][8] , \r60/SUMB[7][9] , \r60/SUMB[7][10] ,
         \r60/SUMB[7][11] , \r60/SUMB[7][12] , \r60/SUMB[7][13] ,
         \r60/SUMB[7][14] , \r60/SUMB[7][15] , \r60/SUMB[7][16] ,
         \r60/SUMB[7][17] , \r60/SUMB[7][18] , \r60/SUMB[7][19] ,
         \r60/SUMB[7][20] , \r60/SUMB[7][21] , \r60/SUMB[7][22] ,
         \r60/SUMB[7][23] , \r60/SUMB[7][24] , \r60/SUMB[7][25] ,
         \r60/SUMB[7][26] , \r60/SUMB[7][27] , \r60/SUMB[7][28] ,
         \r60/SUMB[7][29] , \r60/SUMB[7][30] , \r60/SUMB[8][1] ,
         \r60/SUMB[8][2] , \r60/SUMB[8][3] , \r60/SUMB[8][4] ,
         \r60/SUMB[8][5] , \r60/SUMB[8][6] , \r60/SUMB[8][7] ,
         \r60/SUMB[8][8] , \r60/SUMB[8][9] , \r60/SUMB[8][10] ,
         \r60/SUMB[8][11] , \r60/SUMB[8][12] , \r60/SUMB[8][13] ,
         \r60/SUMB[8][14] , \r60/SUMB[8][15] , \r60/SUMB[8][16] ,
         \r60/SUMB[8][17] , \r60/SUMB[8][18] , \r60/SUMB[8][19] ,
         \r60/SUMB[8][20] , \r60/SUMB[8][21] , \r60/SUMB[8][22] ,
         \r60/SUMB[8][23] , \r60/SUMB[8][24] , \r60/SUMB[8][25] ,
         \r60/SUMB[8][26] , \r60/SUMB[8][27] , \r60/SUMB[8][28] ,
         \r60/SUMB[8][29] , \r60/SUMB[8][30] , \r60/SUMB[9][1] ,
         \r60/SUMB[9][2] , \r60/SUMB[9][3] , \r60/SUMB[9][4] ,
         \r60/SUMB[9][5] , \r60/SUMB[9][6] , \r60/SUMB[9][7] ,
         \r60/SUMB[9][8] , \r60/SUMB[9][9] , \r60/SUMB[9][10] ,
         \r60/SUMB[9][11] , \r60/SUMB[9][12] , \r60/SUMB[9][13] ,
         \r60/SUMB[9][14] , \r60/SUMB[9][15] , \r60/SUMB[9][16] ,
         \r60/SUMB[9][17] , \r60/SUMB[9][18] , \r60/SUMB[9][19] ,
         \r60/SUMB[9][20] , \r60/SUMB[9][21] , \r60/SUMB[9][22] ,
         \r60/SUMB[9][23] , \r60/SUMB[9][24] , \r60/SUMB[9][25] ,
         \r60/SUMB[9][26] , \r60/SUMB[9][27] , \r60/SUMB[9][28] ,
         \r60/SUMB[9][29] , \r60/SUMB[9][30] , \r60/SUMB[10][1] ,
         \r60/SUMB[10][2] , \r60/SUMB[10][3] , \r60/SUMB[10][4] ,
         \r60/SUMB[10][5] , \r60/SUMB[10][6] , \r60/SUMB[10][7] ,
         \r60/SUMB[10][8] , \r60/SUMB[10][9] , \r60/SUMB[10][10] ,
         \r60/SUMB[10][11] , \r60/SUMB[10][12] , \r60/SUMB[10][13] ,
         \r60/SUMB[10][14] , \r60/SUMB[10][15] , \r60/SUMB[10][16] ,
         \r60/SUMB[10][17] , \r60/SUMB[10][18] , \r60/SUMB[10][19] ,
         \r60/SUMB[10][20] , \r60/SUMB[10][21] , \r60/SUMB[10][22] ,
         \r60/SUMB[10][23] , \r60/SUMB[10][24] , \r60/SUMB[10][25] ,
         \r60/SUMB[10][26] , \r60/SUMB[10][27] , \r60/SUMB[10][28] ,
         \r60/SUMB[10][29] , \r60/SUMB[10][30] , \r60/SUMB[11][1] ,
         \r60/SUMB[11][2] , \r60/SUMB[11][3] , \r60/SUMB[11][4] ,
         \r60/SUMB[11][5] , \r60/SUMB[11][6] , \r60/SUMB[11][7] ,
         \r60/SUMB[11][8] , \r60/SUMB[11][9] , \r60/SUMB[11][10] ,
         \r60/SUMB[11][11] , \r60/SUMB[11][12] , \r60/SUMB[11][13] ,
         \r60/SUMB[11][14] , \r60/SUMB[11][15] , \r60/SUMB[11][16] ,
         \r60/SUMB[11][17] , \r60/SUMB[11][18] , \r60/SUMB[11][19] ,
         \r60/SUMB[11][20] , \r60/SUMB[11][21] , \r60/SUMB[11][22] ,
         \r60/SUMB[11][23] , \r60/SUMB[11][24] , \r60/SUMB[11][25] ,
         \r60/SUMB[11][26] , \r60/SUMB[11][27] , \r60/SUMB[11][28] ,
         \r60/SUMB[11][29] , \r60/SUMB[11][30] , \r60/SUMB[12][1] ,
         \r60/SUMB[12][2] , \r60/SUMB[12][3] , \r60/SUMB[12][4] ,
         \r60/SUMB[12][5] , \r60/SUMB[12][6] , \r60/SUMB[12][7] ,
         \r60/SUMB[12][8] , \r60/SUMB[12][9] , \r60/SUMB[12][10] ,
         \r60/SUMB[12][11] , \r60/SUMB[12][12] , \r60/SUMB[12][13] ,
         \r60/SUMB[12][14] , \r60/SUMB[12][15] , \r60/SUMB[12][16] ,
         \r60/SUMB[12][17] , \r60/SUMB[12][18] , \r60/SUMB[12][19] ,
         \r60/SUMB[12][20] , \r60/SUMB[12][21] , \r60/SUMB[12][22] ,
         \r60/SUMB[12][23] , \r60/SUMB[12][24] , \r60/SUMB[12][25] ,
         \r60/SUMB[12][26] , \r60/SUMB[12][27] , \r60/SUMB[12][28] ,
         \r60/SUMB[12][29] , \r60/SUMB[12][30] , \r60/SUMB[13][1] ,
         \r60/SUMB[13][2] , \r60/SUMB[13][3] , \r60/SUMB[13][4] ,
         \r60/SUMB[13][5] , \r60/SUMB[13][6] , \r60/SUMB[13][7] ,
         \r60/SUMB[13][8] , \r60/SUMB[13][9] , \r60/SUMB[13][10] ,
         \r60/SUMB[13][11] , \r60/SUMB[13][12] , \r60/SUMB[13][13] ,
         \r60/SUMB[13][14] , \r60/SUMB[13][15] , \r60/SUMB[13][16] ,
         \r60/SUMB[13][17] , \r60/SUMB[13][18] , \r60/SUMB[13][19] ,
         \r60/SUMB[13][20] , \r60/SUMB[13][21] , \r60/SUMB[13][22] ,
         \r60/SUMB[13][23] , \r60/SUMB[13][24] , \r60/SUMB[13][25] ,
         \r60/SUMB[13][26] , \r60/SUMB[13][27] , \r60/SUMB[13][28] ,
         \r60/SUMB[13][29] , \r60/SUMB[13][30] , \r60/SUMB[14][1] ,
         \r60/SUMB[14][2] , \r60/SUMB[14][3] , \r60/SUMB[14][4] ,
         \r60/SUMB[14][5] , \r60/SUMB[14][6] , \r60/SUMB[14][7] ,
         \r60/SUMB[14][8] , \r60/SUMB[14][9] , \r60/SUMB[14][10] ,
         \r60/SUMB[14][11] , \r60/SUMB[14][12] , \r60/SUMB[14][13] ,
         \r60/SUMB[14][14] , \r60/SUMB[14][15] , \r60/SUMB[14][16] ,
         \r60/SUMB[14][17] , \r60/SUMB[14][18] , \r60/SUMB[14][19] ,
         \r60/SUMB[14][20] , \r60/SUMB[14][21] , \r60/SUMB[14][22] ,
         \r60/SUMB[14][23] , \r60/SUMB[14][24] , \r60/SUMB[14][25] ,
         \r60/SUMB[14][26] , \r60/SUMB[14][27] , \r60/SUMB[14][28] ,
         \r60/SUMB[14][29] , \r60/SUMB[14][30] , \r60/SUMB[15][1] ,
         \r60/SUMB[15][2] , \r60/SUMB[15][3] , \r60/SUMB[15][4] ,
         \r60/SUMB[15][5] , \r60/SUMB[15][6] , \r60/SUMB[15][7] ,
         \r60/SUMB[15][8] , \r60/SUMB[15][9] , \r60/SUMB[15][10] ,
         \r60/SUMB[15][11] , \r60/SUMB[15][12] , \r60/SUMB[15][13] ,
         \r60/SUMB[15][14] , \r60/SUMB[15][15] , \r60/SUMB[15][16] ,
         \r60/SUMB[15][17] , \r60/SUMB[15][18] , \r60/SUMB[15][19] ,
         \r60/SUMB[15][20] , \r60/SUMB[15][21] , \r60/SUMB[15][22] ,
         \r60/SUMB[15][23] , \r60/SUMB[15][24] , \r60/SUMB[15][25] ,
         \r60/SUMB[15][26] , \r60/SUMB[15][27] , \r60/SUMB[15][28] ,
         \r60/SUMB[15][29] , \r60/SUMB[15][30] , \r60/CARRYB[1][0] ,
         \r60/CARRYB[1][1] , \r60/CARRYB[1][2] , \r60/CARRYB[1][3] ,
         \r60/CARRYB[1][4] , \r60/CARRYB[1][5] , \r60/CARRYB[1][6] ,
         \r60/CARRYB[1][7] , \r60/CARRYB[1][8] , \r60/CARRYB[1][9] ,
         \r60/CARRYB[1][10] , \r60/CARRYB[1][11] , \r60/CARRYB[1][12] ,
         \r60/CARRYB[1][13] , \r60/CARRYB[1][14] , \r60/CARRYB[1][15] ,
         \r60/CARRYB[1][16] , \r60/CARRYB[1][17] , \r60/CARRYB[1][18] ,
         \r60/CARRYB[1][19] , \r60/CARRYB[1][20] , \r60/CARRYB[1][21] ,
         \r60/CARRYB[1][22] , \r60/CARRYB[1][23] , \r60/CARRYB[1][24] ,
         \r60/CARRYB[1][25] , \r60/CARRYB[1][26] , \r60/CARRYB[1][27] ,
         \r60/CARRYB[1][28] , \r60/CARRYB[1][29] , \r60/CARRYB[1][30] ,
         \r60/CARRYB[2][0] , \r60/CARRYB[2][1] , \r60/CARRYB[2][2] ,
         \r60/CARRYB[2][3] , \r60/CARRYB[2][4] , \r60/CARRYB[2][5] ,
         \r60/CARRYB[2][6] , \r60/CARRYB[2][7] , \r60/CARRYB[2][8] ,
         \r60/CARRYB[2][9] , \r60/CARRYB[2][10] , \r60/CARRYB[2][11] ,
         \r60/CARRYB[2][12] , \r60/CARRYB[2][13] , \r60/CARRYB[2][14] ,
         \r60/CARRYB[2][15] , \r60/CARRYB[2][16] , \r60/CARRYB[2][17] ,
         \r60/CARRYB[2][18] , \r60/CARRYB[2][19] , \r60/CARRYB[2][20] ,
         \r60/CARRYB[2][21] , \r60/CARRYB[2][22] , \r60/CARRYB[2][23] ,
         \r60/CARRYB[2][24] , \r60/CARRYB[2][25] , \r60/CARRYB[2][26] ,
         \r60/CARRYB[2][27] , \r60/CARRYB[2][28] , \r60/CARRYB[2][29] ,
         \r60/CARRYB[2][30] , \r60/CARRYB[3][0] , \r60/CARRYB[3][1] ,
         \r60/CARRYB[3][2] , \r60/CARRYB[3][3] , \r60/CARRYB[3][4] ,
         \r60/CARRYB[3][5] , \r60/CARRYB[3][6] , \r60/CARRYB[3][7] ,
         \r60/CARRYB[3][8] , \r60/CARRYB[3][9] , \r60/CARRYB[3][10] ,
         \r60/CARRYB[3][11] , \r60/CARRYB[3][12] , \r60/CARRYB[3][13] ,
         \r60/CARRYB[3][14] , \r60/CARRYB[3][15] , \r60/CARRYB[3][16] ,
         \r60/CARRYB[3][17] , \r60/CARRYB[3][18] , \r60/CARRYB[3][19] ,
         \r60/CARRYB[3][20] , \r60/CARRYB[3][21] , \r60/CARRYB[3][22] ,
         \r60/CARRYB[3][23] , \r60/CARRYB[3][24] , \r60/CARRYB[3][25] ,
         \r60/CARRYB[3][26] , \r60/CARRYB[3][27] , \r60/CARRYB[3][28] ,
         \r60/CARRYB[3][29] , \r60/CARRYB[3][30] , \r60/CARRYB[4][0] ,
         \r60/CARRYB[4][1] , \r60/CARRYB[4][2] , \r60/CARRYB[4][3] ,
         \r60/CARRYB[4][4] , \r60/CARRYB[4][5] , \r60/CARRYB[4][6] ,
         \r60/CARRYB[4][7] , \r60/CARRYB[4][8] , \r60/CARRYB[4][9] ,
         \r60/CARRYB[4][10] , \r60/CARRYB[4][11] , \r60/CARRYB[4][12] ,
         \r60/CARRYB[4][13] , \r60/CARRYB[4][14] , \r60/CARRYB[4][15] ,
         \r60/CARRYB[4][16] , \r60/CARRYB[4][17] , \r60/CARRYB[4][18] ,
         \r60/CARRYB[4][19] , \r60/CARRYB[4][20] , \r60/CARRYB[4][21] ,
         \r60/CARRYB[4][22] , \r60/CARRYB[4][23] , \r60/CARRYB[4][24] ,
         \r60/CARRYB[4][25] , \r60/CARRYB[4][26] , \r60/CARRYB[4][27] ,
         \r60/CARRYB[4][28] , \r60/CARRYB[4][29] , \r60/CARRYB[4][30] ,
         \r60/CARRYB[5][0] , \r60/CARRYB[5][1] , \r60/CARRYB[5][2] ,
         \r60/CARRYB[5][3] , \r60/CARRYB[5][4] , \r60/CARRYB[5][5] ,
         \r60/CARRYB[5][6] , \r60/CARRYB[5][7] , \r60/CARRYB[5][8] ,
         \r60/CARRYB[5][9] , \r60/CARRYB[5][10] , \r60/CARRYB[5][11] ,
         \r60/CARRYB[5][12] , \r60/CARRYB[5][13] , \r60/CARRYB[5][14] ,
         \r60/CARRYB[5][15] , \r60/CARRYB[5][16] , \r60/CARRYB[5][17] ,
         \r60/CARRYB[5][18] , \r60/CARRYB[5][19] , \r60/CARRYB[5][20] ,
         \r60/CARRYB[5][21] , \r60/CARRYB[5][22] , \r60/CARRYB[5][23] ,
         \r60/CARRYB[5][24] , \r60/CARRYB[5][25] , \r60/CARRYB[5][26] ,
         \r60/CARRYB[5][27] , \r60/CARRYB[5][28] , \r60/CARRYB[5][29] ,
         \r60/CARRYB[5][30] , \r60/CARRYB[6][0] , \r60/CARRYB[6][1] ,
         \r60/CARRYB[6][2] , \r60/CARRYB[6][3] , \r60/CARRYB[6][4] ,
         \r60/CARRYB[6][5] , \r60/CARRYB[6][6] , \r60/CARRYB[6][7] ,
         \r60/CARRYB[6][8] , \r60/CARRYB[6][9] , \r60/CARRYB[6][10] ,
         \r60/CARRYB[6][11] , \r60/CARRYB[6][12] , \r60/CARRYB[6][13] ,
         \r60/CARRYB[6][14] , \r60/CARRYB[6][15] , \r60/CARRYB[6][16] ,
         \r60/CARRYB[6][17] , \r60/CARRYB[6][18] , \r60/CARRYB[6][19] ,
         \r60/CARRYB[6][20] , \r60/CARRYB[6][21] , \r60/CARRYB[6][22] ,
         \r60/CARRYB[6][23] , \r60/CARRYB[6][24] , \r60/CARRYB[6][25] ,
         \r60/CARRYB[6][26] , \r60/CARRYB[6][27] , \r60/CARRYB[6][28] ,
         \r60/CARRYB[6][29] , \r60/CARRYB[6][30] , \r60/CARRYB[7][0] ,
         \r60/CARRYB[7][1] , \r60/CARRYB[7][2] , \r60/CARRYB[7][3] ,
         \r60/CARRYB[7][4] , \r60/CARRYB[7][5] , \r60/CARRYB[7][6] ,
         \r60/CARRYB[7][7] , \r60/CARRYB[7][8] , \r60/CARRYB[7][9] ,
         \r60/CARRYB[7][10] , \r60/CARRYB[7][11] , \r60/CARRYB[7][12] ,
         \r60/CARRYB[7][13] , \r60/CARRYB[7][14] , \r60/CARRYB[7][15] ,
         \r60/CARRYB[7][16] , \r60/CARRYB[7][17] , \r60/CARRYB[7][18] ,
         \r60/CARRYB[7][19] , \r60/CARRYB[7][20] , \r60/CARRYB[7][21] ,
         \r60/CARRYB[7][22] , \r60/CARRYB[7][23] , \r60/CARRYB[7][24] ,
         \r60/CARRYB[7][25] , \r60/CARRYB[7][26] , \r60/CARRYB[7][27] ,
         \r60/CARRYB[7][28] , \r60/CARRYB[7][29] , \r60/CARRYB[7][30] ,
         \r60/CARRYB[8][0] , \r60/CARRYB[8][1] , \r60/CARRYB[8][2] ,
         \r60/CARRYB[8][3] , \r60/CARRYB[8][4] , \r60/CARRYB[8][5] ,
         \r60/CARRYB[8][6] , \r60/CARRYB[8][7] , \r60/CARRYB[8][8] ,
         \r60/CARRYB[8][9] , \r60/CARRYB[8][10] , \r60/CARRYB[8][11] ,
         \r60/CARRYB[8][12] , \r60/CARRYB[8][13] , \r60/CARRYB[8][14] ,
         \r60/CARRYB[8][15] , \r60/CARRYB[8][16] , \r60/CARRYB[8][17] ,
         \r60/CARRYB[8][18] , \r60/CARRYB[8][19] , \r60/CARRYB[8][20] ,
         \r60/CARRYB[8][21] , \r60/CARRYB[8][22] , \r60/CARRYB[8][23] ,
         \r60/CARRYB[8][24] , \r60/CARRYB[8][25] , \r60/CARRYB[8][26] ,
         \r60/CARRYB[8][27] , \r60/CARRYB[8][28] , \r60/CARRYB[8][29] ,
         \r60/CARRYB[8][30] , \r60/CARRYB[9][0] , \r60/CARRYB[9][1] ,
         \r60/CARRYB[9][2] , \r60/CARRYB[9][3] , \r60/CARRYB[9][4] ,
         \r60/CARRYB[9][5] , \r60/CARRYB[9][6] , \r60/CARRYB[9][7] ,
         \r60/CARRYB[9][8] , \r60/CARRYB[9][9] , \r60/CARRYB[9][10] ,
         \r60/CARRYB[9][11] , \r60/CARRYB[9][12] , \r60/CARRYB[9][13] ,
         \r60/CARRYB[9][14] , \r60/CARRYB[9][15] , \r60/CARRYB[9][16] ,
         \r60/CARRYB[9][17] , \r60/CARRYB[9][18] , \r60/CARRYB[9][19] ,
         \r60/CARRYB[9][20] , \r60/CARRYB[9][21] , \r60/CARRYB[9][22] ,
         \r60/CARRYB[9][23] , \r60/CARRYB[9][24] , \r60/CARRYB[9][25] ,
         \r60/CARRYB[9][26] , \r60/CARRYB[9][27] , \r60/CARRYB[9][28] ,
         \r60/CARRYB[9][29] , \r60/CARRYB[9][30] , \r60/CARRYB[10][0] ,
         \r60/CARRYB[10][1] , \r60/CARRYB[10][2] , \r60/CARRYB[10][3] ,
         \r60/CARRYB[10][4] , \r60/CARRYB[10][5] , \r60/CARRYB[10][6] ,
         \r60/CARRYB[10][7] , \r60/CARRYB[10][8] , \r60/CARRYB[10][9] ,
         \r60/CARRYB[10][10] , \r60/CARRYB[10][11] , \r60/CARRYB[10][12] ,
         \r60/CARRYB[10][13] , \r60/CARRYB[10][14] , \r60/CARRYB[10][15] ,
         \r60/CARRYB[10][16] , \r60/CARRYB[10][17] , \r60/CARRYB[10][18] ,
         \r60/CARRYB[10][19] , \r60/CARRYB[10][20] , \r60/CARRYB[10][21] ,
         \r60/CARRYB[10][22] , \r60/CARRYB[10][23] , \r60/CARRYB[10][24] ,
         \r60/CARRYB[10][25] , \r60/CARRYB[10][26] , \r60/CARRYB[10][27] ,
         \r60/CARRYB[10][28] , \r60/CARRYB[10][29] , \r60/CARRYB[10][30] ,
         \r60/CARRYB[11][0] , \r60/CARRYB[11][1] , \r60/CARRYB[11][2] ,
         \r60/CARRYB[11][3] , \r60/CARRYB[11][4] , \r60/CARRYB[11][5] ,
         \r60/CARRYB[11][6] , \r60/CARRYB[11][7] , \r60/CARRYB[11][8] ,
         \r60/CARRYB[11][9] , \r60/CARRYB[11][10] , \r60/CARRYB[11][11] ,
         \r60/CARRYB[11][12] , \r60/CARRYB[11][13] , \r60/CARRYB[11][14] ,
         \r60/CARRYB[11][15] , \r60/CARRYB[11][16] , \r60/CARRYB[11][17] ,
         \r60/CARRYB[11][18] , \r60/CARRYB[11][19] , \r60/CARRYB[11][20] ,
         \r60/CARRYB[11][21] , \r60/CARRYB[11][22] , \r60/CARRYB[11][23] ,
         \r60/CARRYB[11][24] , \r60/CARRYB[11][25] , \r60/CARRYB[11][26] ,
         \r60/CARRYB[11][27] , \r60/CARRYB[11][28] , \r60/CARRYB[11][29] ,
         \r60/CARRYB[11][30] , \r60/CARRYB[12][0] , \r60/CARRYB[12][1] ,
         \r60/CARRYB[12][2] , \r60/CARRYB[12][3] , \r60/CARRYB[12][4] ,
         \r60/CARRYB[12][5] , \r60/CARRYB[12][6] , \r60/CARRYB[12][7] ,
         \r60/CARRYB[12][8] , \r60/CARRYB[12][9] , \r60/CARRYB[12][10] ,
         \r60/CARRYB[12][11] , \r60/CARRYB[12][12] , \r60/CARRYB[12][13] ,
         \r60/CARRYB[12][14] , \r60/CARRYB[12][15] , \r60/CARRYB[12][16] ,
         \r60/CARRYB[12][17] , \r60/CARRYB[12][18] , \r60/CARRYB[12][19] ,
         \r60/CARRYB[12][20] , \r60/CARRYB[12][21] , \r60/CARRYB[12][22] ,
         \r60/CARRYB[12][23] , \r60/CARRYB[12][24] , \r60/CARRYB[12][25] ,
         \r60/CARRYB[12][26] , \r60/CARRYB[12][27] , \r60/CARRYB[12][28] ,
         \r60/CARRYB[12][29] , \r60/CARRYB[12][30] , \r60/CARRYB[13][0] ,
         \r60/CARRYB[13][1] , \r60/CARRYB[13][2] , \r60/CARRYB[13][3] ,
         \r60/CARRYB[13][4] , \r60/CARRYB[13][5] , \r60/CARRYB[13][6] ,
         \r60/CARRYB[13][7] , \r60/CARRYB[13][8] , \r60/CARRYB[13][9] ,
         \r60/CARRYB[13][10] , \r60/CARRYB[13][11] , \r60/CARRYB[13][12] ,
         \r60/CARRYB[13][13] , \r60/CARRYB[13][14] , \r60/CARRYB[13][15] ,
         \r60/CARRYB[13][16] , \r60/CARRYB[13][17] , \r60/CARRYB[13][18] ,
         \r60/CARRYB[13][19] , \r60/CARRYB[13][20] , \r60/CARRYB[13][21] ,
         \r60/CARRYB[13][22] , \r60/CARRYB[13][23] , \r60/CARRYB[13][24] ,
         \r60/CARRYB[13][25] , \r60/CARRYB[13][26] , \r60/CARRYB[13][27] ,
         \r60/CARRYB[13][28] , \r60/CARRYB[13][29] , \r60/CARRYB[13][30] ,
         \r60/CARRYB[14][0] , \r60/CARRYB[14][1] , \r60/CARRYB[14][2] ,
         \r60/CARRYB[14][3] , \r60/CARRYB[14][4] , \r60/CARRYB[14][5] ,
         \r60/CARRYB[14][6] , \r60/CARRYB[14][7] , \r60/CARRYB[14][8] ,
         \r60/CARRYB[14][9] , \r60/CARRYB[14][10] , \r60/CARRYB[14][11] ,
         \r60/CARRYB[14][12] , \r60/CARRYB[14][13] , \r60/CARRYB[14][14] ,
         \r60/CARRYB[14][15] , \r60/CARRYB[14][16] , \r60/CARRYB[14][17] ,
         \r60/CARRYB[14][18] , \r60/CARRYB[14][19] , \r60/CARRYB[14][20] ,
         \r60/CARRYB[14][21] , \r60/CARRYB[14][22] , \r60/CARRYB[14][23] ,
         \r60/CARRYB[14][24] , \r60/CARRYB[14][25] , \r60/CARRYB[14][26] ,
         \r60/CARRYB[14][27] , \r60/CARRYB[14][28] , \r60/CARRYB[14][29] ,
         \r60/CARRYB[14][30] , \r60/CARRYB[15][0] , \r60/CARRYB[15][1] ,
         \r60/CARRYB[15][2] , \r60/CARRYB[15][3] , \r60/CARRYB[15][4] ,
         \r60/CARRYB[15][5] , \r60/CARRYB[15][6] , \r60/CARRYB[15][7] ,
         \r60/CARRYB[15][8] , \r60/CARRYB[15][9] , \r60/CARRYB[15][10] ,
         \r60/CARRYB[15][11] , \r60/CARRYB[15][12] , \r60/CARRYB[15][13] ,
         \r60/CARRYB[15][14] , \r60/CARRYB[15][15] , \r60/CARRYB[15][16] ,
         \r60/CARRYB[15][17] , \r60/CARRYB[15][18] , \r60/CARRYB[15][19] ,
         \r60/CARRYB[15][20] , \r60/CARRYB[15][21] , \r60/CARRYB[15][22] ,
         \r60/CARRYB[15][23] , \r60/CARRYB[15][24] , \r60/CARRYB[15][25] ,
         \r60/CARRYB[15][26] , \r60/CARRYB[15][27] , \r60/CARRYB[15][28] ,
         \r60/CARRYB[15][29] , \r60/CARRYB[15][30] , \r60/ab[0][1] ,
         \r60/ab[0][2] , \r60/ab[0][3] , \r60/ab[0][4] , \r60/ab[0][5] ,
         \r60/ab[0][6] , \r60/ab[0][7] , \r60/ab[0][8] , \r60/ab[0][9] ,
         \r60/ab[0][10] , \r60/ab[0][11] , \r60/ab[0][12] , \r60/ab[0][13] ,
         \r60/ab[0][14] , \r60/ab[0][15] , \r60/ab[0][16] , \r60/ab[0][17] ,
         \r60/ab[0][18] , \r60/ab[0][19] , \r60/ab[0][20] , \r60/ab[0][21] ,
         \r60/ab[0][22] , \r60/ab[0][23] , \r60/ab[0][24] , \r60/ab[0][25] ,
         \r60/ab[0][26] , \r60/ab[0][27] , \r60/ab[0][28] , \r60/ab[0][29] ,
         \r60/ab[0][30] , \r60/ab[0][31] , \r60/ab[1][0] , \r60/ab[1][1] ,
         \r60/ab[1][2] , \r60/ab[1][3] , \r60/ab[1][4] , \r60/ab[1][5] ,
         \r60/ab[1][6] , \r60/ab[1][7] , \r60/ab[1][8] , \r60/ab[1][9] ,
         \r60/ab[1][10] , \r60/ab[1][11] , \r60/ab[1][12] , \r60/ab[1][13] ,
         \r60/ab[1][14] , \r60/ab[1][15] , \r60/ab[1][16] , \r60/ab[1][17] ,
         \r60/ab[1][18] , \r60/ab[1][19] , \r60/ab[1][20] , \r60/ab[1][21] ,
         \r60/ab[1][22] , \r60/ab[1][23] , \r60/ab[1][24] , \r60/ab[1][25] ,
         \r60/ab[1][26] , \r60/ab[1][27] , \r60/ab[1][28] , \r60/ab[1][29] ,
         \r60/ab[1][30] , \r60/ab[1][31] , \r60/ab[2][0] , \r60/ab[2][1] ,
         \r60/ab[2][2] , \r60/ab[2][3] , \r60/ab[2][4] , \r60/ab[2][5] ,
         \r60/ab[2][6] , \r60/ab[2][7] , \r60/ab[2][8] , \r60/ab[2][9] ,
         \r60/ab[2][10] , \r60/ab[2][11] , \r60/ab[2][12] , \r60/ab[2][13] ,
         \r60/ab[2][14] , \r60/ab[2][15] , \r60/ab[2][16] , \r60/ab[2][17] ,
         \r60/ab[2][18] , \r60/ab[2][19] , \r60/ab[2][20] , \r60/ab[2][21] ,
         \r60/ab[2][22] , \r60/ab[2][23] , \r60/ab[2][24] , \r60/ab[2][25] ,
         \r60/ab[2][26] , \r60/ab[2][27] , \r60/ab[2][28] , \r60/ab[2][29] ,
         \r60/ab[2][30] , \r60/ab[2][31] , \r60/ab[3][0] , \r60/ab[3][1] ,
         \r60/ab[3][2] , \r60/ab[3][3] , \r60/ab[3][4] , \r60/ab[3][5] ,
         \r60/ab[3][6] , \r60/ab[3][7] , \r60/ab[3][8] , \r60/ab[3][9] ,
         \r60/ab[3][10] , \r60/ab[3][11] , \r60/ab[3][12] , \r60/ab[3][13] ,
         \r60/ab[3][14] , \r60/ab[3][15] , \r60/ab[3][16] , \r60/ab[3][17] ,
         \r60/ab[3][18] , \r60/ab[3][19] , \r60/ab[3][20] , \r60/ab[3][21] ,
         \r60/ab[3][22] , \r60/ab[3][23] , \r60/ab[3][24] , \r60/ab[3][25] ,
         \r60/ab[3][26] , \r60/ab[3][27] , \r60/ab[3][28] , \r60/ab[3][29] ,
         \r60/ab[3][30] , \r60/ab[3][31] , \r60/ab[4][0] , \r60/ab[4][1] ,
         \r60/ab[4][2] , \r60/ab[4][3] , \r60/ab[4][4] , \r60/ab[4][5] ,
         \r60/ab[4][6] , \r60/ab[4][7] , \r60/ab[4][8] , \r60/ab[4][9] ,
         \r60/ab[4][10] , \r60/ab[4][11] , \r60/ab[4][12] , \r60/ab[4][13] ,
         \r60/ab[4][14] , \r60/ab[4][15] , \r60/ab[4][16] , \r60/ab[4][17] ,
         \r60/ab[4][18] , \r60/ab[4][19] , \r60/ab[4][20] , \r60/ab[4][21] ,
         \r60/ab[4][22] , \r60/ab[4][23] , \r60/ab[4][24] , \r60/ab[4][25] ,
         \r60/ab[4][26] , \r60/ab[4][27] , \r60/ab[4][28] , \r60/ab[4][29] ,
         \r60/ab[4][30] , \r60/ab[4][31] , \r60/ab[5][0] , \r60/ab[5][1] ,
         \r60/ab[5][2] , \r60/ab[5][3] , \r60/ab[5][4] , \r60/ab[5][5] ,
         \r60/ab[5][6] , \r60/ab[5][7] , \r60/ab[5][8] , \r60/ab[5][9] ,
         \r60/ab[5][10] , \r60/ab[5][11] , \r60/ab[5][12] , \r60/ab[5][13] ,
         \r60/ab[5][14] , \r60/ab[5][15] , \r60/ab[5][16] , \r60/ab[5][17] ,
         \r60/ab[5][18] , \r60/ab[5][19] , \r60/ab[5][20] , \r60/ab[5][21] ,
         \r60/ab[5][22] , \r60/ab[5][23] , \r60/ab[5][24] , \r60/ab[5][25] ,
         \r60/ab[5][26] , \r60/ab[5][27] , \r60/ab[5][28] , \r60/ab[5][29] ,
         \r60/ab[5][30] , \r60/ab[5][31] , \r60/ab[6][0] , \r60/ab[6][1] ,
         \r60/ab[6][2] , \r60/ab[6][3] , \r60/ab[6][4] , \r60/ab[6][5] ,
         \r60/ab[6][6] , \r60/ab[6][7] , \r60/ab[6][8] , \r60/ab[6][9] ,
         \r60/ab[6][10] , \r60/ab[6][11] , \r60/ab[6][12] , \r60/ab[6][13] ,
         \r60/ab[6][14] , \r60/ab[6][15] , \r60/ab[6][16] , \r60/ab[6][17] ,
         \r60/ab[6][18] , \r60/ab[6][19] , \r60/ab[6][20] , \r60/ab[6][21] ,
         \r60/ab[6][22] , \r60/ab[6][23] , \r60/ab[6][24] , \r60/ab[6][25] ,
         \r60/ab[6][26] , \r60/ab[6][27] , \r60/ab[6][28] , \r60/ab[6][29] ,
         \r60/ab[6][30] , \r60/ab[6][31] , \r60/ab[7][0] , \r60/ab[7][1] ,
         \r60/ab[7][2] , \r60/ab[7][3] , \r60/ab[7][4] , \r60/ab[7][5] ,
         \r60/ab[7][6] , \r60/ab[7][7] , \r60/ab[7][8] , \r60/ab[7][9] ,
         \r60/ab[7][10] , \r60/ab[7][11] , \r60/ab[7][12] , \r60/ab[7][13] ,
         \r60/ab[7][14] , \r60/ab[7][15] , \r60/ab[7][16] , \r60/ab[7][17] ,
         \r60/ab[7][18] , \r60/ab[7][19] , \r60/ab[7][20] , \r60/ab[7][21] ,
         \r60/ab[7][22] , \r60/ab[7][23] , \r60/ab[7][24] , \r60/ab[7][25] ,
         \r60/ab[7][26] , \r60/ab[7][27] , \r60/ab[7][28] , \r60/ab[7][29] ,
         \r60/ab[7][30] , \r60/ab[7][31] , \r60/ab[8][0] , \r60/ab[8][1] ,
         \r60/ab[8][2] , \r60/ab[8][3] , \r60/ab[8][4] , \r60/ab[8][5] ,
         \r60/ab[8][6] , \r60/ab[8][7] , \r60/ab[8][8] , \r60/ab[8][9] ,
         \r60/ab[8][10] , \r60/ab[8][11] , \r60/ab[8][12] , \r60/ab[8][13] ,
         \r60/ab[8][14] , \r60/ab[8][15] , \r60/ab[8][16] , \r60/ab[8][17] ,
         \r60/ab[8][18] , \r60/ab[8][19] , \r60/ab[8][20] , \r60/ab[8][21] ,
         \r60/ab[8][22] , \r60/ab[8][23] , \r60/ab[8][24] , \r60/ab[8][25] ,
         \r60/ab[8][26] , \r60/ab[8][27] , \r60/ab[8][28] , \r60/ab[8][29] ,
         \r60/ab[8][30] , \r60/ab[8][31] , \r60/ab[9][0] , \r60/ab[9][1] ,
         \r60/ab[9][2] , \r60/ab[9][3] , \r60/ab[9][4] , \r60/ab[9][5] ,
         \r60/ab[9][6] , \r60/ab[9][7] , \r60/ab[9][8] , \r60/ab[9][9] ,
         \r60/ab[9][10] , \r60/ab[9][11] , \r60/ab[9][12] , \r60/ab[9][13] ,
         \r60/ab[9][14] , \r60/ab[9][15] , \r60/ab[9][16] , \r60/ab[9][17] ,
         \r60/ab[9][18] , \r60/ab[9][19] , \r60/ab[9][20] , \r60/ab[9][21] ,
         \r60/ab[9][22] , \r60/ab[9][23] , \r60/ab[9][24] , \r60/ab[9][25] ,
         \r60/ab[9][26] , \r60/ab[9][27] , \r60/ab[9][28] , \r60/ab[9][29] ,
         \r60/ab[9][30] , \r60/ab[9][31] , \r60/ab[10][0] , \r60/ab[10][1] ,
         \r60/ab[10][2] , \r60/ab[10][3] , \r60/ab[10][4] , \r60/ab[10][5] ,
         \r60/ab[10][6] , \r60/ab[10][7] , \r60/ab[10][8] , \r60/ab[10][9] ,
         \r60/ab[10][10] , \r60/ab[10][11] , \r60/ab[10][12] ,
         \r60/ab[10][13] , \r60/ab[10][14] , \r60/ab[10][15] ,
         \r60/ab[10][16] , \r60/ab[10][17] , \r60/ab[10][18] ,
         \r60/ab[10][19] , \r60/ab[10][20] , \r60/ab[10][21] ,
         \r60/ab[10][22] , \r60/ab[10][23] , \r60/ab[10][24] ,
         \r60/ab[10][25] , \r60/ab[10][26] , \r60/ab[10][27] ,
         \r60/ab[10][28] , \r60/ab[10][29] , \r60/ab[10][30] ,
         \r60/ab[10][31] , \r60/ab[11][0] , \r60/ab[11][1] , \r60/ab[11][2] ,
         \r60/ab[11][3] , \r60/ab[11][4] , \r60/ab[11][5] , \r60/ab[11][6] ,
         \r60/ab[11][7] , \r60/ab[11][8] , \r60/ab[11][9] , \r60/ab[11][10] ,
         \r60/ab[11][11] , \r60/ab[11][12] , \r60/ab[11][13] ,
         \r60/ab[11][14] , \r60/ab[11][15] , \r60/ab[11][16] ,
         \r60/ab[11][17] , \r60/ab[11][18] , \r60/ab[11][19] ,
         \r60/ab[11][20] , \r60/ab[11][21] , \r60/ab[11][22] ,
         \r60/ab[11][23] , \r60/ab[11][24] , \r60/ab[11][25] ,
         \r60/ab[11][26] , \r60/ab[11][27] , \r60/ab[11][28] ,
         \r60/ab[11][29] , \r60/ab[11][30] , \r60/ab[11][31] , \r60/ab[12][0] ,
         \r60/ab[12][1] , \r60/ab[12][2] , \r60/ab[12][3] , \r60/ab[12][4] ,
         \r60/ab[12][5] , \r60/ab[12][6] , \r60/ab[12][7] , \r60/ab[12][8] ,
         \r60/ab[12][9] , \r60/ab[12][10] , \r60/ab[12][11] , \r60/ab[12][12] ,
         \r60/ab[12][13] , \r60/ab[12][14] , \r60/ab[12][15] ,
         \r60/ab[12][16] , \r60/ab[12][17] , \r60/ab[12][18] ,
         \r60/ab[12][19] , \r60/ab[12][20] , \r60/ab[12][21] ,
         \r60/ab[12][22] , \r60/ab[12][23] , \r60/ab[12][24] ,
         \r60/ab[12][25] , \r60/ab[12][26] , \r60/ab[12][27] ,
         \r60/ab[12][28] , \r60/ab[12][29] , \r60/ab[12][30] ,
         \r60/ab[12][31] , \r60/ab[13][0] , \r60/ab[13][1] , \r60/ab[13][2] ,
         \r60/ab[13][3] , \r60/ab[13][4] , \r60/ab[13][5] , \r60/ab[13][6] ,
         \r60/ab[13][7] , \r60/ab[13][8] , \r60/ab[13][9] , \r60/ab[13][10] ,
         \r60/ab[13][11] , \r60/ab[13][12] , \r60/ab[13][13] ,
         \r60/ab[13][14] , \r60/ab[13][15] , \r60/ab[13][16] ,
         \r60/ab[13][17] , \r60/ab[13][18] , \r60/ab[13][19] ,
         \r60/ab[13][20] , \r60/ab[13][21] , \r60/ab[13][22] ,
         \r60/ab[13][23] , \r60/ab[13][24] , \r60/ab[13][25] ,
         \r60/ab[13][26] , \r60/ab[13][27] , \r60/ab[13][28] ,
         \r60/ab[13][29] , \r60/ab[13][30] , \r60/ab[13][31] , \r60/ab[14][0] ,
         \r60/ab[14][1] , \r60/ab[14][2] , \r60/ab[14][3] , \r60/ab[14][4] ,
         \r60/ab[14][5] , \r60/ab[14][6] , \r60/ab[14][7] , \r60/ab[14][8] ,
         \r60/ab[14][9] , \r60/ab[14][10] , \r60/ab[14][11] , \r60/ab[14][12] ,
         \r60/ab[14][13] , \r60/ab[14][14] , \r60/ab[14][15] ,
         \r60/ab[14][16] , \r60/ab[14][17] , \r60/ab[14][18] ,
         \r60/ab[14][19] , \r60/ab[14][20] , \r60/ab[14][21] ,
         \r60/ab[14][22] , \r60/ab[14][23] , \r60/ab[14][24] ,
         \r60/ab[14][25] , \r60/ab[14][26] , \r60/ab[14][27] ,
         \r60/ab[14][28] , \r60/ab[14][29] , \r60/ab[14][30] ,
         \r60/ab[14][31] , \r60/ab[15][0] , \r60/ab[15][1] , \r60/ab[15][2] ,
         \r60/ab[15][3] , \r60/ab[15][4] , \r60/ab[15][5] , \r60/ab[15][6] ,
         \r60/ab[15][7] , \r60/ab[15][8] , \r60/ab[15][9] , \r60/ab[15][10] ,
         \r60/ab[15][11] , \r60/ab[15][12] , \r60/ab[15][13] ,
         \r60/ab[15][14] , \r60/ab[15][15] , \r60/ab[15][16] ,
         \r60/ab[15][17] , \r60/ab[15][18] , \r60/ab[15][19] ,
         \r60/ab[15][20] , \r60/ab[15][21] , \r60/ab[15][22] ,
         \r60/ab[15][23] , \r60/ab[15][24] , \r60/ab[15][25] ,
         \r60/ab[15][26] , \r60/ab[15][27] , \r60/ab[15][28] ,
         \r60/ab[15][29] , \r60/ab[15][30] , \r60/ab[15][31] , \r60/ab[16][0] ,
         \r60/ab[16][1] , \r60/ab[16][2] , \r60/ab[16][3] , \r60/ab[16][4] ,
         \r60/ab[16][5] , \r60/ab[16][6] , \r60/ab[16][7] , \r60/ab[16][8] ,
         \r60/ab[16][9] , \r60/ab[16][10] , \r60/ab[16][11] , \r60/ab[16][12] ,
         \r60/ab[16][13] , \r60/ab[16][14] , \r60/ab[16][15] ,
         \r60/ab[16][16] , \r60/ab[16][17] , \r60/ab[16][18] ,
         \r60/ab[16][19] , \r60/ab[16][20] , \r60/ab[16][21] ,
         \r60/ab[16][22] , \r60/ab[16][23] , \r60/ab[16][24] ,
         \r60/ab[16][25] , \r60/ab[16][26] , \r60/ab[16][27] ,
         \r60/ab[16][28] , \r60/ab[16][29] , \r60/ab[16][30] ,
         \r60/ab[16][31] , \r60/ab[17][0] , \r60/ab[17][1] , \r60/ab[17][2] ,
         \r60/ab[17][3] , \r60/ab[17][4] , \r60/ab[17][5] , \r60/ab[17][6] ,
         \r60/ab[17][7] , \r60/ab[17][8] , \r60/ab[17][9] , \r60/ab[17][10] ,
         \r60/ab[17][11] , \r60/ab[17][12] , \r60/ab[17][13] ,
         \r60/ab[17][14] , \r60/ab[17][15] , \r60/ab[17][16] ,
         \r60/ab[17][17] , \r60/ab[17][18] , \r60/ab[17][19] ,
         \r60/ab[17][20] , \r60/ab[17][21] , \r60/ab[17][22] ,
         \r60/ab[17][23] , \r60/ab[17][24] , \r60/ab[17][25] ,
         \r60/ab[17][26] , \r60/ab[17][27] , \r60/ab[17][28] ,
         \r60/ab[17][29] , \r60/ab[17][30] , \r60/ab[17][31] , \r60/ab[18][0] ,
         \r60/ab[18][1] , \r60/ab[18][2] , \r60/ab[18][3] , \r60/ab[18][4] ,
         \r60/ab[18][5] , \r60/ab[18][6] , \r60/ab[18][7] , \r60/ab[18][8] ,
         \r60/ab[18][9] , \r60/ab[18][10] , \r60/ab[18][11] , \r60/ab[18][12] ,
         \r60/ab[18][13] , \r60/ab[18][14] , \r60/ab[18][15] ,
         \r60/ab[18][16] , \r60/ab[18][17] , \r60/ab[18][18] ,
         \r60/ab[18][19] , \r60/ab[18][20] , \r60/ab[18][21] ,
         \r60/ab[18][22] , \r60/ab[18][23] , \r60/ab[18][24] ,
         \r60/ab[18][25] , \r60/ab[18][26] , \r60/ab[18][27] ,
         \r60/ab[18][28] , \r60/ab[18][29] , \r60/ab[18][30] ,
         \r60/ab[18][31] , \r60/ab[19][0] , \r60/ab[19][1] , \r60/ab[19][2] ,
         \r60/ab[19][3] , \r60/ab[19][4] , \r60/ab[19][5] , \r60/ab[19][6] ,
         \r60/ab[19][7] , \r60/ab[19][8] , \r60/ab[19][9] , \r60/ab[19][10] ,
         \r60/ab[19][11] , \r60/ab[19][12] , \r60/ab[19][13] ,
         \r60/ab[19][14] , \r60/ab[19][15] , \r60/ab[19][16] ,
         \r60/ab[19][17] , \r60/ab[19][18] , \r60/ab[19][19] ,
         \r60/ab[19][20] , \r60/ab[19][21] , \r60/ab[19][22] ,
         \r60/ab[19][23] , \r60/ab[19][24] , \r60/ab[19][25] ,
         \r60/ab[19][26] , \r60/ab[19][27] , \r60/ab[19][28] ,
         \r60/ab[19][29] , \r60/ab[19][30] , \r60/ab[19][31] , \r60/ab[20][0] ,
         \r60/ab[20][1] , \r60/ab[20][2] , \r60/ab[20][3] , \r60/ab[20][4] ,
         \r60/ab[20][5] , \r60/ab[20][6] , \r60/ab[20][7] , \r60/ab[20][8] ,
         \r60/ab[20][9] , \r60/ab[20][10] , \r60/ab[20][11] , \r60/ab[20][12] ,
         \r60/ab[20][13] , \r60/ab[20][14] , \r60/ab[20][15] ,
         \r60/ab[20][16] , \r60/ab[20][17] , \r60/ab[20][18] ,
         \r60/ab[20][19] , \r60/ab[20][20] , \r60/ab[20][21] ,
         \r60/ab[20][22] , \r60/ab[20][23] , \r60/ab[20][24] ,
         \r60/ab[20][25] , \r60/ab[20][26] , \r60/ab[20][27] ,
         \r60/ab[20][28] , \r60/ab[20][29] , \r60/ab[20][30] ,
         \r60/ab[20][31] , \r60/ab[21][0] , \r60/ab[21][1] , \r60/ab[21][2] ,
         \r60/ab[21][3] , \r60/ab[21][4] , \r60/ab[21][5] , \r60/ab[21][6] ,
         \r60/ab[21][7] , \r60/ab[21][8] , \r60/ab[21][9] , \r60/ab[21][10] ,
         \r60/ab[21][11] , \r60/ab[21][12] , \r60/ab[21][13] ,
         \r60/ab[21][14] , \r60/ab[21][15] , \r60/ab[21][16] ,
         \r60/ab[21][17] , \r60/ab[21][18] , \r60/ab[21][19] ,
         \r60/ab[21][20] , \r60/ab[21][21] , \r60/ab[21][22] ,
         \r60/ab[21][23] , \r60/ab[21][24] , \r60/ab[21][25] ,
         \r60/ab[21][26] , \r60/ab[21][27] , \r60/ab[21][28] ,
         \r60/ab[21][29] , \r60/ab[21][30] , \r60/ab[21][31] , \r60/ab[22][0] ,
         \r60/ab[22][1] , \r60/ab[22][2] , \r60/ab[22][3] , \r60/ab[22][4] ,
         \r60/ab[22][5] , \r60/ab[22][6] , \r60/ab[22][7] , \r60/ab[22][8] ,
         \r60/ab[22][9] , \r60/ab[22][10] , \r60/ab[22][11] , \r60/ab[22][12] ,
         \r60/ab[22][13] , \r60/ab[22][14] , \r60/ab[22][15] ,
         \r60/ab[22][16] , \r60/ab[22][17] , \r60/ab[22][18] ,
         \r60/ab[22][19] , \r60/ab[22][20] , \r60/ab[22][21] ,
         \r60/ab[22][22] , \r60/ab[22][23] , \r60/ab[22][24] ,
         \r60/ab[22][25] , \r60/ab[22][26] , \r60/ab[22][27] ,
         \r60/ab[22][28] , \r60/ab[22][29] , \r60/ab[22][30] ,
         \r60/ab[22][31] , \r60/ab[23][0] , \r60/ab[23][1] , \r60/ab[23][2] ,
         \r60/ab[23][3] , \r60/ab[23][4] , \r60/ab[23][5] , \r60/ab[23][6] ,
         \r60/ab[23][7] , \r60/ab[23][8] , \r60/ab[23][9] , \r60/ab[23][10] ,
         \r60/ab[23][11] , \r60/ab[23][12] , \r60/ab[23][13] ,
         \r60/ab[23][14] , \r60/ab[23][15] , \r60/ab[23][16] ,
         \r60/ab[23][17] , \r60/ab[23][18] , \r60/ab[23][19] ,
         \r60/ab[23][20] , \r60/ab[23][21] , \r60/ab[23][22] ,
         \r60/ab[23][23] , \r60/ab[23][24] , \r60/ab[23][25] ,
         \r60/ab[23][26] , \r60/ab[23][27] , \r60/ab[23][28] ,
         \r60/ab[23][29] , \r60/ab[23][30] , \r60/ab[23][31] , \r60/ab[24][0] ,
         \r60/ab[24][1] , \r60/ab[24][2] , \r60/ab[24][3] , \r60/ab[24][4] ,
         \r60/ab[24][5] , \r60/ab[24][6] , \r60/ab[24][7] , \r60/ab[24][8] ,
         \r60/ab[24][9] , \r60/ab[24][10] , \r60/ab[24][11] , \r60/ab[24][12] ,
         \r60/ab[24][13] , \r60/ab[24][14] , \r60/ab[24][15] ,
         \r60/ab[24][16] , \r60/ab[24][17] , \r60/ab[24][18] ,
         \r60/ab[24][19] , \r60/ab[24][20] , \r60/ab[24][21] ,
         \r60/ab[24][22] , \r60/ab[24][23] , \r60/ab[24][24] ,
         \r60/ab[24][25] , \r60/ab[24][26] , \r60/ab[24][27] ,
         \r60/ab[24][28] , \r60/ab[24][29] , \r60/ab[24][30] ,
         \r60/ab[24][31] , \r60/ab[25][0] , \r60/ab[25][1] , \r60/ab[25][2] ,
         \r60/ab[25][3] , \r60/ab[25][4] , \r60/ab[25][5] , \r60/ab[25][6] ,
         \r60/ab[25][7] , \r60/ab[25][8] , \r60/ab[25][9] , \r60/ab[25][10] ,
         \r60/ab[25][11] , \r60/ab[25][12] , \r60/ab[25][13] ,
         \r60/ab[25][14] , \r60/ab[25][15] , \r60/ab[25][16] ,
         \r60/ab[25][17] , \r60/ab[25][18] , \r60/ab[25][19] ,
         \r60/ab[25][20] , \r60/ab[25][21] , \r60/ab[25][22] ,
         \r60/ab[25][23] , \r60/ab[25][24] , \r60/ab[25][25] ,
         \r60/ab[25][26] , \r60/ab[25][27] , \r60/ab[25][28] ,
         \r60/ab[25][29] , \r60/ab[25][30] , \r60/ab[25][31] , \r60/ab[26][0] ,
         \r60/ab[26][1] , \r60/ab[26][2] , \r60/ab[26][3] , \r60/ab[26][4] ,
         \r60/ab[26][5] , \r60/ab[26][6] , \r60/ab[26][7] , \r60/ab[26][8] ,
         \r60/ab[26][9] , \r60/ab[26][10] , \r60/ab[26][11] , \r60/ab[26][12] ,
         \r60/ab[26][13] , \r60/ab[26][14] , \r60/ab[26][15] ,
         \r60/ab[26][16] , \r60/ab[26][17] , \r60/ab[26][18] ,
         \r60/ab[26][19] , \r60/ab[26][20] , \r60/ab[26][21] ,
         \r60/ab[26][22] , \r60/ab[26][23] , \r60/ab[26][24] ,
         \r60/ab[26][25] , \r60/ab[26][26] , \r60/ab[26][27] ,
         \r60/ab[26][28] , \r60/ab[26][29] , \r60/ab[26][30] ,
         \r60/ab[26][31] , \r60/ab[27][0] , \r60/ab[27][1] , \r60/ab[27][2] ,
         \r60/ab[27][3] , \r60/ab[27][4] , \r60/ab[27][5] , \r60/ab[27][6] ,
         \r60/ab[27][7] , \r60/ab[27][8] , \r60/ab[27][9] , \r60/ab[27][10] ,
         \r60/ab[27][11] , \r60/ab[27][12] , \r60/ab[27][13] ,
         \r60/ab[27][14] , \r60/ab[27][15] , \r60/ab[27][16] ,
         \r60/ab[27][17] , \r60/ab[27][18] , \r60/ab[27][19] ,
         \r60/ab[27][20] , \r60/ab[27][21] , \r60/ab[27][22] ,
         \r60/ab[27][23] , \r60/ab[27][24] , \r60/ab[27][25] ,
         \r60/ab[27][26] , \r60/ab[27][27] , \r60/ab[27][28] ,
         \r60/ab[27][29] , \r60/ab[27][30] , \r60/ab[27][31] , \r60/ab[28][0] ,
         \r60/ab[28][1] , \r60/ab[28][2] , \r60/ab[28][3] , \r60/ab[28][4] ,
         \r60/ab[28][5] , \r60/ab[28][6] , \r60/ab[28][7] , \r60/ab[28][8] ,
         \r60/ab[28][9] , \r60/ab[28][10] , \r60/ab[28][11] , \r60/ab[28][12] ,
         \r60/ab[28][13] , \r60/ab[28][14] , \r60/ab[28][15] ,
         \r60/ab[28][16] , \r60/ab[28][17] , \r60/ab[28][18] ,
         \r60/ab[28][19] , \r60/ab[28][20] , \r60/ab[28][21] ,
         \r60/ab[28][22] , \r60/ab[28][23] , \r60/ab[28][24] ,
         \r60/ab[28][25] , \r60/ab[28][26] , \r60/ab[28][27] ,
         \r60/ab[28][28] , \r60/ab[28][29] , \r60/ab[28][30] ,
         \r60/ab[28][31] , \r60/ab[29][0] , \r60/ab[29][1] , \r60/ab[29][2] ,
         \r60/ab[29][3] , \r60/ab[29][4] , \r60/ab[29][5] , \r60/ab[29][6] ,
         \r60/ab[29][7] , \r60/ab[29][8] , \r60/ab[29][9] , \r60/ab[29][10] ,
         \r60/ab[29][11] , \r60/ab[29][12] , \r60/ab[29][13] ,
         \r60/ab[29][14] , \r60/ab[29][15] , \r60/ab[29][16] ,
         \r60/ab[29][17] , \r60/ab[29][18] , \r60/ab[29][19] ,
         \r60/ab[29][20] , \r60/ab[29][21] , \r60/ab[29][22] ,
         \r60/ab[29][23] , \r60/ab[29][24] , \r60/ab[29][25] ,
         \r60/ab[29][26] , \r60/ab[29][27] , \r60/ab[29][28] ,
         \r60/ab[29][29] , \r60/ab[29][30] , \r60/ab[29][31] , \r60/ab[30][0] ,
         \r60/ab[30][1] , \r60/ab[30][2] , \r60/ab[30][3] , \r60/ab[30][4] ,
         \r60/ab[30][5] , \r60/ab[30][6] , \r60/ab[30][7] , \r60/ab[30][8] ,
         \r60/ab[30][9] , \r60/ab[30][10] , \r60/ab[30][11] , \r60/ab[30][12] ,
         \r60/ab[30][13] , \r60/ab[30][14] , \r60/ab[30][15] ,
         \r60/ab[30][16] , \r60/ab[30][17] , \r60/ab[30][18] ,
         \r60/ab[30][19] , \r60/ab[30][20] , \r60/ab[30][21] ,
         \r60/ab[30][22] , \r60/ab[30][23] , \r60/ab[30][24] ,
         \r60/ab[30][25] , \r60/ab[30][26] , \r60/ab[30][27] ,
         \r60/ab[30][28] , \r60/ab[30][29] , \r60/ab[30][30] ,
         \r60/ab[30][31] , \r60/ab[31][0] , \r60/ab[31][1] , \r60/ab[31][2] ,
         \r60/ab[31][3] , \r60/ab[31][4] , \r60/ab[31][5] , \r60/ab[31][6] ,
         \r60/ab[31][7] , \r60/ab[31][8] , \r60/ab[31][9] , \r60/ab[31][10] ,
         \r60/ab[31][11] , \r60/ab[31][12] , \r60/ab[31][13] ,
         \r60/ab[31][14] , \r60/ab[31][15] , \r60/ab[31][16] ,
         \r60/ab[31][17] , \r60/ab[31][18] , \r60/ab[31][19] ,
         \r60/ab[31][20] , \r60/ab[31][21] , \r60/ab[31][22] ,
         \r60/ab[31][23] , \r60/ab[31][24] , \r60/ab[31][25] ,
         \r60/ab[31][26] , \r60/ab[31][27] , \r60/ab[31][28] ,
         \r60/ab[31][29] , \r60/ab[31][30] , \r60/ab[31][31] , n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325;
  wire   [31:0] Lo;
  wire   [31:0] Hi;

  DFF \Hi_reg[31]  ( .D(n679), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[31]) );
  DFF \Hi_reg[30]  ( .D(n678), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[30]) );
  DFF \Hi_reg[29]  ( .D(n677), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[29]) );
  DFF \Hi_reg[28]  ( .D(n676), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[28]) );
  DFF \Hi_reg[27]  ( .D(n675), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[27]) );
  DFF \Hi_reg[26]  ( .D(n674), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[26]) );
  DFF \Hi_reg[25]  ( .D(n673), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[25]) );
  DFF \Hi_reg[24]  ( .D(n672), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[24]) );
  DFF \Hi_reg[23]  ( .D(n671), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[23]) );
  DFF \Hi_reg[22]  ( .D(n670), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[22]) );
  DFF \Hi_reg[21]  ( .D(n669), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[21]) );
  DFF \Hi_reg[20]  ( .D(n668), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[20]) );
  DFF \Hi_reg[19]  ( .D(n667), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[19]) );
  DFF \Hi_reg[18]  ( .D(n666), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[18]) );
  DFF \Hi_reg[17]  ( .D(n665), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[17]) );
  DFF \Hi_reg[16]  ( .D(n664), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[16]) );
  DFF \Hi_reg[15]  ( .D(n663), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[15]) );
  DFF \Hi_reg[14]  ( .D(n662), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[14]) );
  DFF \Hi_reg[13]  ( .D(n661), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[13]) );
  DFF \Hi_reg[12]  ( .D(n660), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[12]) );
  DFF \Hi_reg[11]  ( .D(n659), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[11]) );
  DFF \Hi_reg[10]  ( .D(n658), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[10]) );
  DFF \Hi_reg[9]  ( .D(n657), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[9]) );
  DFF \Hi_reg[8]  ( .D(n656), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[8]) );
  DFF \Hi_reg[7]  ( .D(n655), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[7]) );
  DFF \Hi_reg[6]  ( .D(n654), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[6]) );
  DFF \Hi_reg[5]  ( .D(n653), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[5]) );
  DFF \Hi_reg[4]  ( .D(n652), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[4]) );
  DFF \Hi_reg[3]  ( .D(n651), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[3]) );
  DFF \Hi_reg[2]  ( .D(n650), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[2]) );
  DFF \Hi_reg[1]  ( .D(n649), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[1]) );
  DFF \Hi_reg[0]  ( .D(n648), .CLK(clk), .RST(rst), .I(1'b0), .Q(Hi[0]) );
  DFF \Lo_reg[31]  ( .D(n647), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[31]) );
  DFF \Lo_reg[30]  ( .D(n646), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[30]) );
  DFF \Lo_reg[29]  ( .D(n645), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[29]) );
  DFF \Lo_reg[28]  ( .D(n644), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[28]) );
  DFF \Lo_reg[27]  ( .D(n643), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[27]) );
  DFF \Lo_reg[26]  ( .D(n642), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[26]) );
  DFF \Lo_reg[25]  ( .D(n641), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[25]) );
  DFF \Lo_reg[24]  ( .D(n640), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[24]) );
  DFF \Lo_reg[23]  ( .D(n639), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[23]) );
  DFF \Lo_reg[22]  ( .D(n638), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[22]) );
  DFF \Lo_reg[21]  ( .D(n637), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[21]) );
  DFF \Lo_reg[20]  ( .D(n636), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[20]) );
  DFF \Lo_reg[19]  ( .D(n635), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[19]) );
  DFF \Lo_reg[18]  ( .D(n634), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[18]) );
  DFF \Lo_reg[17]  ( .D(n633), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[17]) );
  DFF \Lo_reg[16]  ( .D(n632), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[16]) );
  DFF \Lo_reg[15]  ( .D(n631), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[15]) );
  DFF \Lo_reg[14]  ( .D(n630), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[14]) );
  DFF \Lo_reg[13]  ( .D(n629), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[13]) );
  DFF \Lo_reg[12]  ( .D(n628), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[12]) );
  DFF \Lo_reg[11]  ( .D(n627), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[11]) );
  DFF \Lo_reg[10]  ( .D(n626), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[10]) );
  DFF \Lo_reg[9]  ( .D(n625), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[9]) );
  DFF \Lo_reg[8]  ( .D(n624), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[8]) );
  DFF \Lo_reg[7]  ( .D(n623), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[7]) );
  DFF \Lo_reg[6]  ( .D(n622), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[6]) );
  DFF \Lo_reg[5]  ( .D(n621), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[5]) );
  DFF \Lo_reg[4]  ( .D(n620), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[4]) );
  DFF \Lo_reg[3]  ( .D(n619), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[3]) );
  DFF \Lo_reg[2]  ( .D(n618), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[2]) );
  DFF \Lo_reg[1]  ( .D(n617), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[1]) );
  DFF \Lo_reg[0]  ( .D(n616), .CLK(clk), .RST(rst), .I(1'b0), .Q(Lo[0]) );
  FADDER \r60/S3_2_30  ( .CIN(\r60/ab[2][30] ), .IN0(\r60/CARRYB[1][30] ), 
        .IN1(\r60/ab[1][31] ), .COUT(\r60/CARRYB[2][30] ), .SUM(
        \r60/SUMB[2][30] ) );
  FADDER \r60/S2_2_29  ( .CIN(\r60/ab[2][29] ), .IN0(\r60/CARRYB[1][29] ), 
        .IN1(\r60/SUMB[1][30] ), .COUT(\r60/CARRYB[2][29] ), .SUM(
        \r60/SUMB[2][29] ) );
  FADDER \r60/S2_2_28  ( .CIN(\r60/ab[2][28] ), .IN0(\r60/CARRYB[1][28] ), 
        .IN1(\r60/SUMB[1][29] ), .COUT(\r60/CARRYB[2][28] ), .SUM(
        \r60/SUMB[2][28] ) );
  FADDER \r60/S2_2_27  ( .CIN(\r60/ab[2][27] ), .IN0(\r60/CARRYB[1][27] ), 
        .IN1(\r60/SUMB[1][28] ), .COUT(\r60/CARRYB[2][27] ), .SUM(
        \r60/SUMB[2][27] ) );
  FADDER \r60/S2_2_26  ( .CIN(\r60/ab[2][26] ), .IN0(\r60/CARRYB[1][26] ), 
        .IN1(\r60/SUMB[1][27] ), .COUT(\r60/CARRYB[2][26] ), .SUM(
        \r60/SUMB[2][26] ) );
  FADDER \r60/S2_2_25  ( .CIN(\r60/ab[2][25] ), .IN0(\r60/CARRYB[1][25] ), 
        .IN1(\r60/SUMB[1][26] ), .COUT(\r60/CARRYB[2][25] ), .SUM(
        \r60/SUMB[2][25] ) );
  FADDER \r60/S2_2_24  ( .CIN(\r60/ab[2][24] ), .IN0(\r60/CARRYB[1][24] ), 
        .IN1(\r60/SUMB[1][25] ), .COUT(\r60/CARRYB[2][24] ), .SUM(
        \r60/SUMB[2][24] ) );
  FADDER \r60/S2_2_23  ( .CIN(\r60/ab[2][23] ), .IN0(\r60/CARRYB[1][23] ), 
        .IN1(\r60/SUMB[1][24] ), .COUT(\r60/CARRYB[2][23] ), .SUM(
        \r60/SUMB[2][23] ) );
  FADDER \r60/S2_2_22  ( .CIN(\r60/ab[2][22] ), .IN0(\r60/CARRYB[1][22] ), 
        .IN1(\r60/SUMB[1][23] ), .COUT(\r60/CARRYB[2][22] ), .SUM(
        \r60/SUMB[2][22] ) );
  FADDER \r60/S2_2_21  ( .CIN(\r60/ab[2][21] ), .IN0(\r60/CARRYB[1][21] ), 
        .IN1(\r60/SUMB[1][22] ), .COUT(\r60/CARRYB[2][21] ), .SUM(
        \r60/SUMB[2][21] ) );
  FADDER \r60/S2_2_20  ( .CIN(\r60/ab[2][20] ), .IN0(\r60/CARRYB[1][20] ), 
        .IN1(\r60/SUMB[1][21] ), .COUT(\r60/CARRYB[2][20] ), .SUM(
        \r60/SUMB[2][20] ) );
  FADDER \r60/S2_2_19  ( .CIN(\r60/ab[2][19] ), .IN0(\r60/CARRYB[1][19] ), 
        .IN1(\r60/SUMB[1][20] ), .COUT(\r60/CARRYB[2][19] ), .SUM(
        \r60/SUMB[2][19] ) );
  FADDER \r60/S2_2_18  ( .CIN(\r60/ab[2][18] ), .IN0(\r60/CARRYB[1][18] ), 
        .IN1(\r60/SUMB[1][19] ), .COUT(\r60/CARRYB[2][18] ), .SUM(
        \r60/SUMB[2][18] ) );
  FADDER \r60/S2_2_17  ( .CIN(\r60/ab[2][17] ), .IN0(\r60/CARRYB[1][17] ), 
        .IN1(\r60/SUMB[1][18] ), .COUT(\r60/CARRYB[2][17] ), .SUM(
        \r60/SUMB[2][17] ) );
  FADDER \r60/S2_2_16  ( .CIN(\r60/ab[2][16] ), .IN0(\r60/CARRYB[1][16] ), 
        .IN1(\r60/SUMB[1][17] ), .COUT(\r60/CARRYB[2][16] ), .SUM(
        \r60/SUMB[2][16] ) );
  FADDER \r60/S2_2_15  ( .CIN(\r60/ab[2][15] ), .IN0(\r60/CARRYB[1][15] ), 
        .IN1(\r60/SUMB[1][16] ), .COUT(\r60/CARRYB[2][15] ), .SUM(
        \r60/SUMB[2][15] ) );
  FADDER \r60/S2_2_14  ( .CIN(\r60/ab[2][14] ), .IN0(\r60/CARRYB[1][14] ), 
        .IN1(\r60/SUMB[1][15] ), .COUT(\r60/CARRYB[2][14] ), .SUM(
        \r60/SUMB[2][14] ) );
  FADDER \r60/S2_2_13  ( .CIN(\r60/ab[2][13] ), .IN0(\r60/CARRYB[1][13] ), 
        .IN1(\r60/SUMB[1][14] ), .COUT(\r60/CARRYB[2][13] ), .SUM(
        \r60/SUMB[2][13] ) );
  FADDER \r60/S2_2_12  ( .CIN(\r60/ab[2][12] ), .IN0(\r60/CARRYB[1][12] ), 
        .IN1(\r60/SUMB[1][13] ), .COUT(\r60/CARRYB[2][12] ), .SUM(
        \r60/SUMB[2][12] ) );
  FADDER \r60/S2_2_11  ( .CIN(\r60/ab[2][11] ), .IN0(\r60/CARRYB[1][11] ), 
        .IN1(\r60/SUMB[1][12] ), .COUT(\r60/CARRYB[2][11] ), .SUM(
        \r60/SUMB[2][11] ) );
  FADDER \r60/S2_2_10  ( .CIN(\r60/ab[2][10] ), .IN0(\r60/CARRYB[1][10] ), 
        .IN1(\r60/SUMB[1][11] ), .COUT(\r60/CARRYB[2][10] ), .SUM(
        \r60/SUMB[2][10] ) );
  FADDER \r60/S2_2_9  ( .CIN(\r60/ab[2][9] ), .IN0(\r60/CARRYB[1][9] ), .IN1(
        \r60/SUMB[1][10] ), .COUT(\r60/CARRYB[2][9] ), .SUM(\r60/SUMB[2][9] )
         );
  FADDER \r60/S2_2_8  ( .CIN(\r60/ab[2][8] ), .IN0(\r60/CARRYB[1][8] ), .IN1(
        \r60/SUMB[1][9] ), .COUT(\r60/CARRYB[2][8] ), .SUM(\r60/SUMB[2][8] )
         );
  FADDER \r60/S2_2_7  ( .CIN(\r60/ab[2][7] ), .IN0(\r60/CARRYB[1][7] ), .IN1(
        \r60/SUMB[1][8] ), .COUT(\r60/CARRYB[2][7] ), .SUM(\r60/SUMB[2][7] )
         );
  FADDER \r60/S2_2_6  ( .CIN(\r60/ab[2][6] ), .IN0(\r60/CARRYB[1][6] ), .IN1(
        \r60/SUMB[1][7] ), .COUT(\r60/CARRYB[2][6] ), .SUM(\r60/SUMB[2][6] )
         );
  FADDER \r60/S2_2_5  ( .CIN(\r60/ab[2][5] ), .IN0(\r60/CARRYB[1][5] ), .IN1(
        \r60/SUMB[1][6] ), .COUT(\r60/CARRYB[2][5] ), .SUM(\r60/SUMB[2][5] )
         );
  FADDER \r60/S2_2_4  ( .CIN(\r60/ab[2][4] ), .IN0(\r60/CARRYB[1][4] ), .IN1(
        \r60/SUMB[1][5] ), .COUT(\r60/CARRYB[2][4] ), .SUM(\r60/SUMB[2][4] )
         );
  FADDER \r60/S2_2_3  ( .CIN(\r60/ab[2][3] ), .IN0(\r60/CARRYB[1][3] ), .IN1(
        \r60/SUMB[1][4] ), .COUT(\r60/CARRYB[2][3] ), .SUM(\r60/SUMB[2][3] )
         );
  FADDER \r60/S2_2_2  ( .CIN(\r60/ab[2][2] ), .IN0(\r60/CARRYB[1][2] ), .IN1(
        \r60/SUMB[1][3] ), .COUT(\r60/CARRYB[2][2] ), .SUM(\r60/SUMB[2][2] )
         );
  FADDER \r60/S2_2_1  ( .CIN(\r60/ab[2][1] ), .IN0(\r60/CARRYB[1][1] ), .IN1(
        \r60/SUMB[1][2] ), .COUT(\r60/CARRYB[2][1] ), .SUM(\r60/SUMB[2][1] )
         );
  FADDER \r60/S1_2_0  ( .CIN(\r60/ab[2][0] ), .IN0(\r60/CARRYB[1][0] ), .IN1(
        \r60/SUMB[1][1] ), .COUT(\r60/CARRYB[2][0] ), .SUM(N119) );
  FADDER \r60/S3_3_30  ( .CIN(\r60/ab[3][30] ), .IN0(\r60/CARRYB[2][30] ), 
        .IN1(\r60/ab[2][31] ), .COUT(\r60/CARRYB[3][30] ), .SUM(
        \r60/SUMB[3][30] ) );
  FADDER \r60/S2_3_29  ( .CIN(\r60/ab[3][29] ), .IN0(\r60/CARRYB[2][29] ), 
        .IN1(\r60/SUMB[2][30] ), .COUT(\r60/CARRYB[3][29] ), .SUM(
        \r60/SUMB[3][29] ) );
  FADDER \r60/S2_3_28  ( .CIN(\r60/ab[3][28] ), .IN0(\r60/CARRYB[2][28] ), 
        .IN1(\r60/SUMB[2][29] ), .COUT(\r60/CARRYB[3][28] ), .SUM(
        \r60/SUMB[3][28] ) );
  FADDER \r60/S2_3_27  ( .CIN(\r60/ab[3][27] ), .IN0(\r60/CARRYB[2][27] ), 
        .IN1(\r60/SUMB[2][28] ), .COUT(\r60/CARRYB[3][27] ), .SUM(
        \r60/SUMB[3][27] ) );
  FADDER \r60/S2_3_26  ( .CIN(\r60/ab[3][26] ), .IN0(\r60/CARRYB[2][26] ), 
        .IN1(\r60/SUMB[2][27] ), .COUT(\r60/CARRYB[3][26] ), .SUM(
        \r60/SUMB[3][26] ) );
  FADDER \r60/S2_3_25  ( .CIN(\r60/ab[3][25] ), .IN0(\r60/CARRYB[2][25] ), 
        .IN1(\r60/SUMB[2][26] ), .COUT(\r60/CARRYB[3][25] ), .SUM(
        \r60/SUMB[3][25] ) );
  FADDER \r60/S2_3_24  ( .CIN(\r60/ab[3][24] ), .IN0(\r60/CARRYB[2][24] ), 
        .IN1(\r60/SUMB[2][25] ), .COUT(\r60/CARRYB[3][24] ), .SUM(
        \r60/SUMB[3][24] ) );
  FADDER \r60/S2_3_23  ( .CIN(\r60/ab[3][23] ), .IN0(\r60/CARRYB[2][23] ), 
        .IN1(\r60/SUMB[2][24] ), .COUT(\r60/CARRYB[3][23] ), .SUM(
        \r60/SUMB[3][23] ) );
  FADDER \r60/S2_3_22  ( .CIN(\r60/ab[3][22] ), .IN0(\r60/CARRYB[2][22] ), 
        .IN1(\r60/SUMB[2][23] ), .COUT(\r60/CARRYB[3][22] ), .SUM(
        \r60/SUMB[3][22] ) );
  FADDER \r60/S2_3_21  ( .CIN(\r60/ab[3][21] ), .IN0(\r60/CARRYB[2][21] ), 
        .IN1(\r60/SUMB[2][22] ), .COUT(\r60/CARRYB[3][21] ), .SUM(
        \r60/SUMB[3][21] ) );
  FADDER \r60/S2_3_20  ( .CIN(\r60/ab[3][20] ), .IN0(\r60/CARRYB[2][20] ), 
        .IN1(\r60/SUMB[2][21] ), .COUT(\r60/CARRYB[3][20] ), .SUM(
        \r60/SUMB[3][20] ) );
  FADDER \r60/S2_3_19  ( .CIN(\r60/ab[3][19] ), .IN0(\r60/CARRYB[2][19] ), 
        .IN1(\r60/SUMB[2][20] ), .COUT(\r60/CARRYB[3][19] ), .SUM(
        \r60/SUMB[3][19] ) );
  FADDER \r60/S2_3_18  ( .CIN(\r60/ab[3][18] ), .IN0(\r60/CARRYB[2][18] ), 
        .IN1(\r60/SUMB[2][19] ), .COUT(\r60/CARRYB[3][18] ), .SUM(
        \r60/SUMB[3][18] ) );
  FADDER \r60/S2_3_17  ( .CIN(\r60/ab[3][17] ), .IN0(\r60/CARRYB[2][17] ), 
        .IN1(\r60/SUMB[2][18] ), .COUT(\r60/CARRYB[3][17] ), .SUM(
        \r60/SUMB[3][17] ) );
  FADDER \r60/S2_3_16  ( .CIN(\r60/ab[3][16] ), .IN0(\r60/CARRYB[2][16] ), 
        .IN1(\r60/SUMB[2][17] ), .COUT(\r60/CARRYB[3][16] ), .SUM(
        \r60/SUMB[3][16] ) );
  FADDER \r60/S2_3_15  ( .CIN(\r60/ab[3][15] ), .IN0(\r60/CARRYB[2][15] ), 
        .IN1(\r60/SUMB[2][16] ), .COUT(\r60/CARRYB[3][15] ), .SUM(
        \r60/SUMB[3][15] ) );
  FADDER \r60/S2_3_14  ( .CIN(\r60/ab[3][14] ), .IN0(\r60/CARRYB[2][14] ), 
        .IN1(\r60/SUMB[2][15] ), .COUT(\r60/CARRYB[3][14] ), .SUM(
        \r60/SUMB[3][14] ) );
  FADDER \r60/S2_3_13  ( .CIN(\r60/ab[3][13] ), .IN0(\r60/CARRYB[2][13] ), 
        .IN1(\r60/SUMB[2][14] ), .COUT(\r60/CARRYB[3][13] ), .SUM(
        \r60/SUMB[3][13] ) );
  FADDER \r60/S2_3_12  ( .CIN(\r60/ab[3][12] ), .IN0(\r60/CARRYB[2][12] ), 
        .IN1(\r60/SUMB[2][13] ), .COUT(\r60/CARRYB[3][12] ), .SUM(
        \r60/SUMB[3][12] ) );
  FADDER \r60/S2_3_11  ( .CIN(\r60/ab[3][11] ), .IN0(\r60/CARRYB[2][11] ), 
        .IN1(\r60/SUMB[2][12] ), .COUT(\r60/CARRYB[3][11] ), .SUM(
        \r60/SUMB[3][11] ) );
  FADDER \r60/S2_3_10  ( .CIN(\r60/ab[3][10] ), .IN0(\r60/CARRYB[2][10] ), 
        .IN1(\r60/SUMB[2][11] ), .COUT(\r60/CARRYB[3][10] ), .SUM(
        \r60/SUMB[3][10] ) );
  FADDER \r60/S2_3_9  ( .CIN(\r60/ab[3][9] ), .IN0(\r60/CARRYB[2][9] ), .IN1(
        \r60/SUMB[2][10] ), .COUT(\r60/CARRYB[3][9] ), .SUM(\r60/SUMB[3][9] )
         );
  FADDER \r60/S2_3_8  ( .CIN(\r60/ab[3][8] ), .IN0(\r60/CARRYB[2][8] ), .IN1(
        \r60/SUMB[2][9] ), .COUT(\r60/CARRYB[3][8] ), .SUM(\r60/SUMB[3][8] )
         );
  FADDER \r60/S2_3_7  ( .CIN(\r60/ab[3][7] ), .IN0(\r60/CARRYB[2][7] ), .IN1(
        \r60/SUMB[2][8] ), .COUT(\r60/CARRYB[3][7] ), .SUM(\r60/SUMB[3][7] )
         );
  FADDER \r60/S2_3_6  ( .CIN(\r60/ab[3][6] ), .IN0(\r60/CARRYB[2][6] ), .IN1(
        \r60/SUMB[2][7] ), .COUT(\r60/CARRYB[3][6] ), .SUM(\r60/SUMB[3][6] )
         );
  FADDER \r60/S2_3_5  ( .CIN(\r60/ab[3][5] ), .IN0(\r60/CARRYB[2][5] ), .IN1(
        \r60/SUMB[2][6] ), .COUT(\r60/CARRYB[3][5] ), .SUM(\r60/SUMB[3][5] )
         );
  FADDER \r60/S2_3_4  ( .CIN(\r60/ab[3][4] ), .IN0(\r60/CARRYB[2][4] ), .IN1(
        \r60/SUMB[2][5] ), .COUT(\r60/CARRYB[3][4] ), .SUM(\r60/SUMB[3][4] )
         );
  FADDER \r60/S2_3_3  ( .CIN(\r60/ab[3][3] ), .IN0(\r60/CARRYB[2][3] ), .IN1(
        \r60/SUMB[2][4] ), .COUT(\r60/CARRYB[3][3] ), .SUM(\r60/SUMB[3][3] )
         );
  FADDER \r60/S2_3_2  ( .CIN(\r60/ab[3][2] ), .IN0(\r60/CARRYB[2][2] ), .IN1(
        \r60/SUMB[2][3] ), .COUT(\r60/CARRYB[3][2] ), .SUM(\r60/SUMB[3][2] )
         );
  FADDER \r60/S2_3_1  ( .CIN(\r60/ab[3][1] ), .IN0(\r60/CARRYB[2][1] ), .IN1(
        \r60/SUMB[2][2] ), .COUT(\r60/CARRYB[3][1] ), .SUM(\r60/SUMB[3][1] )
         );
  FADDER \r60/S1_3_0  ( .CIN(\r60/ab[3][0] ), .IN0(\r60/CARRYB[2][0] ), .IN1(
        \r60/SUMB[2][1] ), .COUT(\r60/CARRYB[3][0] ), .SUM(N120) );
  FADDER \r60/S3_4_30  ( .CIN(\r60/ab[4][30] ), .IN0(\r60/CARRYB[3][30] ), 
        .IN1(\r60/ab[3][31] ), .COUT(\r60/CARRYB[4][30] ), .SUM(
        \r60/SUMB[4][30] ) );
  FADDER \r60/S2_4_29  ( .CIN(\r60/ab[4][29] ), .IN0(\r60/CARRYB[3][29] ), 
        .IN1(\r60/SUMB[3][30] ), .COUT(\r60/CARRYB[4][29] ), .SUM(
        \r60/SUMB[4][29] ) );
  FADDER \r60/S2_4_28  ( .CIN(\r60/ab[4][28] ), .IN0(\r60/CARRYB[3][28] ), 
        .IN1(\r60/SUMB[3][29] ), .COUT(\r60/CARRYB[4][28] ), .SUM(
        \r60/SUMB[4][28] ) );
  FADDER \r60/S2_4_27  ( .CIN(\r60/ab[4][27] ), .IN0(\r60/CARRYB[3][27] ), 
        .IN1(\r60/SUMB[3][28] ), .COUT(\r60/CARRYB[4][27] ), .SUM(
        \r60/SUMB[4][27] ) );
  FADDER \r60/S2_4_26  ( .CIN(\r60/ab[4][26] ), .IN0(\r60/CARRYB[3][26] ), 
        .IN1(\r60/SUMB[3][27] ), .COUT(\r60/CARRYB[4][26] ), .SUM(
        \r60/SUMB[4][26] ) );
  FADDER \r60/S2_4_25  ( .CIN(\r60/ab[4][25] ), .IN0(\r60/CARRYB[3][25] ), 
        .IN1(\r60/SUMB[3][26] ), .COUT(\r60/CARRYB[4][25] ), .SUM(
        \r60/SUMB[4][25] ) );
  FADDER \r60/S2_4_24  ( .CIN(\r60/ab[4][24] ), .IN0(\r60/CARRYB[3][24] ), 
        .IN1(\r60/SUMB[3][25] ), .COUT(\r60/CARRYB[4][24] ), .SUM(
        \r60/SUMB[4][24] ) );
  FADDER \r60/S2_4_23  ( .CIN(\r60/ab[4][23] ), .IN0(\r60/CARRYB[3][23] ), 
        .IN1(\r60/SUMB[3][24] ), .COUT(\r60/CARRYB[4][23] ), .SUM(
        \r60/SUMB[4][23] ) );
  FADDER \r60/S2_4_22  ( .CIN(\r60/ab[4][22] ), .IN0(\r60/CARRYB[3][22] ), 
        .IN1(\r60/SUMB[3][23] ), .COUT(\r60/CARRYB[4][22] ), .SUM(
        \r60/SUMB[4][22] ) );
  FADDER \r60/S2_4_21  ( .CIN(\r60/ab[4][21] ), .IN0(\r60/CARRYB[3][21] ), 
        .IN1(\r60/SUMB[3][22] ), .COUT(\r60/CARRYB[4][21] ), .SUM(
        \r60/SUMB[4][21] ) );
  FADDER \r60/S2_4_20  ( .CIN(\r60/ab[4][20] ), .IN0(\r60/CARRYB[3][20] ), 
        .IN1(\r60/SUMB[3][21] ), .COUT(\r60/CARRYB[4][20] ), .SUM(
        \r60/SUMB[4][20] ) );
  FADDER \r60/S2_4_19  ( .CIN(\r60/ab[4][19] ), .IN0(\r60/CARRYB[3][19] ), 
        .IN1(\r60/SUMB[3][20] ), .COUT(\r60/CARRYB[4][19] ), .SUM(
        \r60/SUMB[4][19] ) );
  FADDER \r60/S2_4_18  ( .CIN(\r60/ab[4][18] ), .IN0(\r60/CARRYB[3][18] ), 
        .IN1(\r60/SUMB[3][19] ), .COUT(\r60/CARRYB[4][18] ), .SUM(
        \r60/SUMB[4][18] ) );
  FADDER \r60/S2_4_17  ( .CIN(\r60/ab[4][17] ), .IN0(\r60/CARRYB[3][17] ), 
        .IN1(\r60/SUMB[3][18] ), .COUT(\r60/CARRYB[4][17] ), .SUM(
        \r60/SUMB[4][17] ) );
  FADDER \r60/S2_4_16  ( .CIN(\r60/ab[4][16] ), .IN0(\r60/CARRYB[3][16] ), 
        .IN1(\r60/SUMB[3][17] ), .COUT(\r60/CARRYB[4][16] ), .SUM(
        \r60/SUMB[4][16] ) );
  FADDER \r60/S2_4_15  ( .CIN(\r60/ab[4][15] ), .IN0(\r60/CARRYB[3][15] ), 
        .IN1(\r60/SUMB[3][16] ), .COUT(\r60/CARRYB[4][15] ), .SUM(
        \r60/SUMB[4][15] ) );
  FADDER \r60/S2_4_14  ( .CIN(\r60/ab[4][14] ), .IN0(\r60/CARRYB[3][14] ), 
        .IN1(\r60/SUMB[3][15] ), .COUT(\r60/CARRYB[4][14] ), .SUM(
        \r60/SUMB[4][14] ) );
  FADDER \r60/S2_4_13  ( .CIN(\r60/ab[4][13] ), .IN0(\r60/CARRYB[3][13] ), 
        .IN1(\r60/SUMB[3][14] ), .COUT(\r60/CARRYB[4][13] ), .SUM(
        \r60/SUMB[4][13] ) );
  FADDER \r60/S2_4_12  ( .CIN(\r60/ab[4][12] ), .IN0(\r60/CARRYB[3][12] ), 
        .IN1(\r60/SUMB[3][13] ), .COUT(\r60/CARRYB[4][12] ), .SUM(
        \r60/SUMB[4][12] ) );
  FADDER \r60/S2_4_11  ( .CIN(\r60/ab[4][11] ), .IN0(\r60/CARRYB[3][11] ), 
        .IN1(\r60/SUMB[3][12] ), .COUT(\r60/CARRYB[4][11] ), .SUM(
        \r60/SUMB[4][11] ) );
  FADDER \r60/S2_4_10  ( .CIN(\r60/ab[4][10] ), .IN0(\r60/CARRYB[3][10] ), 
        .IN1(\r60/SUMB[3][11] ), .COUT(\r60/CARRYB[4][10] ), .SUM(
        \r60/SUMB[4][10] ) );
  FADDER \r60/S2_4_9  ( .CIN(\r60/ab[4][9] ), .IN0(\r60/CARRYB[3][9] ), .IN1(
        \r60/SUMB[3][10] ), .COUT(\r60/CARRYB[4][9] ), .SUM(\r60/SUMB[4][9] )
         );
  FADDER \r60/S2_4_8  ( .CIN(\r60/ab[4][8] ), .IN0(\r60/CARRYB[3][8] ), .IN1(
        \r60/SUMB[3][9] ), .COUT(\r60/CARRYB[4][8] ), .SUM(\r60/SUMB[4][8] )
         );
  FADDER \r60/S2_4_7  ( .CIN(\r60/ab[4][7] ), .IN0(\r60/CARRYB[3][7] ), .IN1(
        \r60/SUMB[3][8] ), .COUT(\r60/CARRYB[4][7] ), .SUM(\r60/SUMB[4][7] )
         );
  FADDER \r60/S2_4_6  ( .CIN(\r60/ab[4][6] ), .IN0(\r60/CARRYB[3][6] ), .IN1(
        \r60/SUMB[3][7] ), .COUT(\r60/CARRYB[4][6] ), .SUM(\r60/SUMB[4][6] )
         );
  FADDER \r60/S2_4_5  ( .CIN(\r60/ab[4][5] ), .IN0(\r60/CARRYB[3][5] ), .IN1(
        \r60/SUMB[3][6] ), .COUT(\r60/CARRYB[4][5] ), .SUM(\r60/SUMB[4][5] )
         );
  FADDER \r60/S2_4_4  ( .CIN(\r60/ab[4][4] ), .IN0(\r60/CARRYB[3][4] ), .IN1(
        \r60/SUMB[3][5] ), .COUT(\r60/CARRYB[4][4] ), .SUM(\r60/SUMB[4][4] )
         );
  FADDER \r60/S2_4_3  ( .CIN(\r60/ab[4][3] ), .IN0(\r60/CARRYB[3][3] ), .IN1(
        \r60/SUMB[3][4] ), .COUT(\r60/CARRYB[4][3] ), .SUM(\r60/SUMB[4][3] )
         );
  FADDER \r60/S2_4_2  ( .CIN(\r60/ab[4][2] ), .IN0(\r60/CARRYB[3][2] ), .IN1(
        \r60/SUMB[3][3] ), .COUT(\r60/CARRYB[4][2] ), .SUM(\r60/SUMB[4][2] )
         );
  FADDER \r60/S2_4_1  ( .CIN(\r60/ab[4][1] ), .IN0(\r60/CARRYB[3][1] ), .IN1(
        \r60/SUMB[3][2] ), .COUT(\r60/CARRYB[4][1] ), .SUM(\r60/SUMB[4][1] )
         );
  FADDER \r60/S1_4_0  ( .CIN(\r60/ab[4][0] ), .IN0(\r60/CARRYB[3][0] ), .IN1(
        \r60/SUMB[3][1] ), .COUT(\r60/CARRYB[4][0] ), .SUM(N121) );
  FADDER \r60/S3_5_30  ( .CIN(\r60/ab[5][30] ), .IN0(\r60/CARRYB[4][30] ), 
        .IN1(\r60/ab[4][31] ), .COUT(\r60/CARRYB[5][30] ), .SUM(
        \r60/SUMB[5][30] ) );
  FADDER \r60/S2_5_29  ( .CIN(\r60/ab[5][29] ), .IN0(\r60/CARRYB[4][29] ), 
        .IN1(\r60/SUMB[4][30] ), .COUT(\r60/CARRYB[5][29] ), .SUM(
        \r60/SUMB[5][29] ) );
  FADDER \r60/S2_5_28  ( .CIN(\r60/ab[5][28] ), .IN0(\r60/CARRYB[4][28] ), 
        .IN1(\r60/SUMB[4][29] ), .COUT(\r60/CARRYB[5][28] ), .SUM(
        \r60/SUMB[5][28] ) );
  FADDER \r60/S2_5_27  ( .CIN(\r60/ab[5][27] ), .IN0(\r60/CARRYB[4][27] ), 
        .IN1(\r60/SUMB[4][28] ), .COUT(\r60/CARRYB[5][27] ), .SUM(
        \r60/SUMB[5][27] ) );
  FADDER \r60/S2_5_26  ( .CIN(\r60/ab[5][26] ), .IN0(\r60/CARRYB[4][26] ), 
        .IN1(\r60/SUMB[4][27] ), .COUT(\r60/CARRYB[5][26] ), .SUM(
        \r60/SUMB[5][26] ) );
  FADDER \r60/S2_5_25  ( .CIN(\r60/ab[5][25] ), .IN0(\r60/CARRYB[4][25] ), 
        .IN1(\r60/SUMB[4][26] ), .COUT(\r60/CARRYB[5][25] ), .SUM(
        \r60/SUMB[5][25] ) );
  FADDER \r60/S2_5_24  ( .CIN(\r60/ab[5][24] ), .IN0(\r60/CARRYB[4][24] ), 
        .IN1(\r60/SUMB[4][25] ), .COUT(\r60/CARRYB[5][24] ), .SUM(
        \r60/SUMB[5][24] ) );
  FADDER \r60/S2_5_23  ( .CIN(\r60/ab[5][23] ), .IN0(\r60/CARRYB[4][23] ), 
        .IN1(\r60/SUMB[4][24] ), .COUT(\r60/CARRYB[5][23] ), .SUM(
        \r60/SUMB[5][23] ) );
  FADDER \r60/S2_5_22  ( .CIN(\r60/ab[5][22] ), .IN0(\r60/CARRYB[4][22] ), 
        .IN1(\r60/SUMB[4][23] ), .COUT(\r60/CARRYB[5][22] ), .SUM(
        \r60/SUMB[5][22] ) );
  FADDER \r60/S2_5_21  ( .CIN(\r60/ab[5][21] ), .IN0(\r60/CARRYB[4][21] ), 
        .IN1(\r60/SUMB[4][22] ), .COUT(\r60/CARRYB[5][21] ), .SUM(
        \r60/SUMB[5][21] ) );
  FADDER \r60/S2_5_20  ( .CIN(\r60/ab[5][20] ), .IN0(\r60/CARRYB[4][20] ), 
        .IN1(\r60/SUMB[4][21] ), .COUT(\r60/CARRYB[5][20] ), .SUM(
        \r60/SUMB[5][20] ) );
  FADDER \r60/S2_5_19  ( .CIN(\r60/ab[5][19] ), .IN0(\r60/CARRYB[4][19] ), 
        .IN1(\r60/SUMB[4][20] ), .COUT(\r60/CARRYB[5][19] ), .SUM(
        \r60/SUMB[5][19] ) );
  FADDER \r60/S2_5_18  ( .CIN(\r60/ab[5][18] ), .IN0(\r60/CARRYB[4][18] ), 
        .IN1(\r60/SUMB[4][19] ), .COUT(\r60/CARRYB[5][18] ), .SUM(
        \r60/SUMB[5][18] ) );
  FADDER \r60/S2_5_17  ( .CIN(\r60/ab[5][17] ), .IN0(\r60/CARRYB[4][17] ), 
        .IN1(\r60/SUMB[4][18] ), .COUT(\r60/CARRYB[5][17] ), .SUM(
        \r60/SUMB[5][17] ) );
  FADDER \r60/S2_5_16  ( .CIN(\r60/ab[5][16] ), .IN0(\r60/CARRYB[4][16] ), 
        .IN1(\r60/SUMB[4][17] ), .COUT(\r60/CARRYB[5][16] ), .SUM(
        \r60/SUMB[5][16] ) );
  FADDER \r60/S2_5_15  ( .CIN(\r60/ab[5][15] ), .IN0(\r60/CARRYB[4][15] ), 
        .IN1(\r60/SUMB[4][16] ), .COUT(\r60/CARRYB[5][15] ), .SUM(
        \r60/SUMB[5][15] ) );
  FADDER \r60/S2_5_14  ( .CIN(\r60/ab[5][14] ), .IN0(\r60/CARRYB[4][14] ), 
        .IN1(\r60/SUMB[4][15] ), .COUT(\r60/CARRYB[5][14] ), .SUM(
        \r60/SUMB[5][14] ) );
  FADDER \r60/S2_5_13  ( .CIN(\r60/ab[5][13] ), .IN0(\r60/CARRYB[4][13] ), 
        .IN1(\r60/SUMB[4][14] ), .COUT(\r60/CARRYB[5][13] ), .SUM(
        \r60/SUMB[5][13] ) );
  FADDER \r60/S2_5_12  ( .CIN(\r60/ab[5][12] ), .IN0(\r60/CARRYB[4][12] ), 
        .IN1(\r60/SUMB[4][13] ), .COUT(\r60/CARRYB[5][12] ), .SUM(
        \r60/SUMB[5][12] ) );
  FADDER \r60/S2_5_11  ( .CIN(\r60/ab[5][11] ), .IN0(\r60/CARRYB[4][11] ), 
        .IN1(\r60/SUMB[4][12] ), .COUT(\r60/CARRYB[5][11] ), .SUM(
        \r60/SUMB[5][11] ) );
  FADDER \r60/S2_5_10  ( .CIN(\r60/ab[5][10] ), .IN0(\r60/CARRYB[4][10] ), 
        .IN1(\r60/SUMB[4][11] ), .COUT(\r60/CARRYB[5][10] ), .SUM(
        \r60/SUMB[5][10] ) );
  FADDER \r60/S2_5_9  ( .CIN(\r60/ab[5][9] ), .IN0(\r60/CARRYB[4][9] ), .IN1(
        \r60/SUMB[4][10] ), .COUT(\r60/CARRYB[5][9] ), .SUM(\r60/SUMB[5][9] )
         );
  FADDER \r60/S2_5_8  ( .CIN(\r60/ab[5][8] ), .IN0(\r60/CARRYB[4][8] ), .IN1(
        \r60/SUMB[4][9] ), .COUT(\r60/CARRYB[5][8] ), .SUM(\r60/SUMB[5][8] )
         );
  FADDER \r60/S2_5_7  ( .CIN(\r60/ab[5][7] ), .IN0(\r60/CARRYB[4][7] ), .IN1(
        \r60/SUMB[4][8] ), .COUT(\r60/CARRYB[5][7] ), .SUM(\r60/SUMB[5][7] )
         );
  FADDER \r60/S2_5_6  ( .CIN(\r60/ab[5][6] ), .IN0(\r60/CARRYB[4][6] ), .IN1(
        \r60/SUMB[4][7] ), .COUT(\r60/CARRYB[5][6] ), .SUM(\r60/SUMB[5][6] )
         );
  FADDER \r60/S2_5_5  ( .CIN(\r60/ab[5][5] ), .IN0(\r60/CARRYB[4][5] ), .IN1(
        \r60/SUMB[4][6] ), .COUT(\r60/CARRYB[5][5] ), .SUM(\r60/SUMB[5][5] )
         );
  FADDER \r60/S2_5_4  ( .CIN(\r60/ab[5][4] ), .IN0(\r60/CARRYB[4][4] ), .IN1(
        \r60/SUMB[4][5] ), .COUT(\r60/CARRYB[5][4] ), .SUM(\r60/SUMB[5][4] )
         );
  FADDER \r60/S2_5_3  ( .CIN(\r60/ab[5][3] ), .IN0(\r60/CARRYB[4][3] ), .IN1(
        \r60/SUMB[4][4] ), .COUT(\r60/CARRYB[5][3] ), .SUM(\r60/SUMB[5][3] )
         );
  FADDER \r60/S2_5_2  ( .CIN(\r60/ab[5][2] ), .IN0(\r60/CARRYB[4][2] ), .IN1(
        \r60/SUMB[4][3] ), .COUT(\r60/CARRYB[5][2] ), .SUM(\r60/SUMB[5][2] )
         );
  FADDER \r60/S2_5_1  ( .CIN(\r60/ab[5][1] ), .IN0(\r60/CARRYB[4][1] ), .IN1(
        \r60/SUMB[4][2] ), .COUT(\r60/CARRYB[5][1] ), .SUM(\r60/SUMB[5][1] )
         );
  FADDER \r60/S1_5_0  ( .CIN(\r60/ab[5][0] ), .IN0(\r60/CARRYB[4][0] ), .IN1(
        \r60/SUMB[4][1] ), .COUT(\r60/CARRYB[5][0] ), .SUM(N122) );
  FADDER \r60/S3_6_30  ( .CIN(\r60/ab[6][30] ), .IN0(\r60/CARRYB[5][30] ), 
        .IN1(\r60/ab[5][31] ), .COUT(\r60/CARRYB[6][30] ), .SUM(
        \r60/SUMB[6][30] ) );
  FADDER \r60/S2_6_29  ( .CIN(\r60/ab[6][29] ), .IN0(\r60/CARRYB[5][29] ), 
        .IN1(\r60/SUMB[5][30] ), .COUT(\r60/CARRYB[6][29] ), .SUM(
        \r60/SUMB[6][29] ) );
  FADDER \r60/S2_6_28  ( .CIN(\r60/ab[6][28] ), .IN0(\r60/CARRYB[5][28] ), 
        .IN1(\r60/SUMB[5][29] ), .COUT(\r60/CARRYB[6][28] ), .SUM(
        \r60/SUMB[6][28] ) );
  FADDER \r60/S2_6_27  ( .CIN(\r60/ab[6][27] ), .IN0(\r60/CARRYB[5][27] ), 
        .IN1(\r60/SUMB[5][28] ), .COUT(\r60/CARRYB[6][27] ), .SUM(
        \r60/SUMB[6][27] ) );
  FADDER \r60/S2_6_26  ( .CIN(\r60/ab[6][26] ), .IN0(\r60/CARRYB[5][26] ), 
        .IN1(\r60/SUMB[5][27] ), .COUT(\r60/CARRYB[6][26] ), .SUM(
        \r60/SUMB[6][26] ) );
  FADDER \r60/S2_6_25  ( .CIN(\r60/ab[6][25] ), .IN0(\r60/CARRYB[5][25] ), 
        .IN1(\r60/SUMB[5][26] ), .COUT(\r60/CARRYB[6][25] ), .SUM(
        \r60/SUMB[6][25] ) );
  FADDER \r60/S2_6_24  ( .CIN(\r60/ab[6][24] ), .IN0(\r60/CARRYB[5][24] ), 
        .IN1(\r60/SUMB[5][25] ), .COUT(\r60/CARRYB[6][24] ), .SUM(
        \r60/SUMB[6][24] ) );
  FADDER \r60/S2_6_23  ( .CIN(\r60/ab[6][23] ), .IN0(\r60/CARRYB[5][23] ), 
        .IN1(\r60/SUMB[5][24] ), .COUT(\r60/CARRYB[6][23] ), .SUM(
        \r60/SUMB[6][23] ) );
  FADDER \r60/S2_6_22  ( .CIN(\r60/ab[6][22] ), .IN0(\r60/CARRYB[5][22] ), 
        .IN1(\r60/SUMB[5][23] ), .COUT(\r60/CARRYB[6][22] ), .SUM(
        \r60/SUMB[6][22] ) );
  FADDER \r60/S2_6_21  ( .CIN(\r60/ab[6][21] ), .IN0(\r60/CARRYB[5][21] ), 
        .IN1(\r60/SUMB[5][22] ), .COUT(\r60/CARRYB[6][21] ), .SUM(
        \r60/SUMB[6][21] ) );
  FADDER \r60/S2_6_20  ( .CIN(\r60/ab[6][20] ), .IN0(\r60/CARRYB[5][20] ), 
        .IN1(\r60/SUMB[5][21] ), .COUT(\r60/CARRYB[6][20] ), .SUM(
        \r60/SUMB[6][20] ) );
  FADDER \r60/S2_6_19  ( .CIN(\r60/ab[6][19] ), .IN0(\r60/CARRYB[5][19] ), 
        .IN1(\r60/SUMB[5][20] ), .COUT(\r60/CARRYB[6][19] ), .SUM(
        \r60/SUMB[6][19] ) );
  FADDER \r60/S2_6_18  ( .CIN(\r60/ab[6][18] ), .IN0(\r60/CARRYB[5][18] ), 
        .IN1(\r60/SUMB[5][19] ), .COUT(\r60/CARRYB[6][18] ), .SUM(
        \r60/SUMB[6][18] ) );
  FADDER \r60/S2_6_17  ( .CIN(\r60/ab[6][17] ), .IN0(\r60/CARRYB[5][17] ), 
        .IN1(\r60/SUMB[5][18] ), .COUT(\r60/CARRYB[6][17] ), .SUM(
        \r60/SUMB[6][17] ) );
  FADDER \r60/S2_6_16  ( .CIN(\r60/ab[6][16] ), .IN0(\r60/CARRYB[5][16] ), 
        .IN1(\r60/SUMB[5][17] ), .COUT(\r60/CARRYB[6][16] ), .SUM(
        \r60/SUMB[6][16] ) );
  FADDER \r60/S2_6_15  ( .CIN(\r60/ab[6][15] ), .IN0(\r60/CARRYB[5][15] ), 
        .IN1(\r60/SUMB[5][16] ), .COUT(\r60/CARRYB[6][15] ), .SUM(
        \r60/SUMB[6][15] ) );
  FADDER \r60/S2_6_14  ( .CIN(\r60/ab[6][14] ), .IN0(\r60/CARRYB[5][14] ), 
        .IN1(\r60/SUMB[5][15] ), .COUT(\r60/CARRYB[6][14] ), .SUM(
        \r60/SUMB[6][14] ) );
  FADDER \r60/S2_6_13  ( .CIN(\r60/ab[6][13] ), .IN0(\r60/CARRYB[5][13] ), 
        .IN1(\r60/SUMB[5][14] ), .COUT(\r60/CARRYB[6][13] ), .SUM(
        \r60/SUMB[6][13] ) );
  FADDER \r60/S2_6_12  ( .CIN(\r60/ab[6][12] ), .IN0(\r60/CARRYB[5][12] ), 
        .IN1(\r60/SUMB[5][13] ), .COUT(\r60/CARRYB[6][12] ), .SUM(
        \r60/SUMB[6][12] ) );
  FADDER \r60/S2_6_11  ( .CIN(\r60/ab[6][11] ), .IN0(\r60/CARRYB[5][11] ), 
        .IN1(\r60/SUMB[5][12] ), .COUT(\r60/CARRYB[6][11] ), .SUM(
        \r60/SUMB[6][11] ) );
  FADDER \r60/S2_6_10  ( .CIN(\r60/ab[6][10] ), .IN0(\r60/CARRYB[5][10] ), 
        .IN1(\r60/SUMB[5][11] ), .COUT(\r60/CARRYB[6][10] ), .SUM(
        \r60/SUMB[6][10] ) );
  FADDER \r60/S2_6_9  ( .CIN(\r60/ab[6][9] ), .IN0(\r60/CARRYB[5][9] ), .IN1(
        \r60/SUMB[5][10] ), .COUT(\r60/CARRYB[6][9] ), .SUM(\r60/SUMB[6][9] )
         );
  FADDER \r60/S2_6_8  ( .CIN(\r60/ab[6][8] ), .IN0(\r60/CARRYB[5][8] ), .IN1(
        \r60/SUMB[5][9] ), .COUT(\r60/CARRYB[6][8] ), .SUM(\r60/SUMB[6][8] )
         );
  FADDER \r60/S2_6_7  ( .CIN(\r60/ab[6][7] ), .IN0(\r60/CARRYB[5][7] ), .IN1(
        \r60/SUMB[5][8] ), .COUT(\r60/CARRYB[6][7] ), .SUM(\r60/SUMB[6][7] )
         );
  FADDER \r60/S2_6_6  ( .CIN(\r60/ab[6][6] ), .IN0(\r60/CARRYB[5][6] ), .IN1(
        \r60/SUMB[5][7] ), .COUT(\r60/CARRYB[6][6] ), .SUM(\r60/SUMB[6][6] )
         );
  FADDER \r60/S2_6_5  ( .CIN(\r60/ab[6][5] ), .IN0(\r60/CARRYB[5][5] ), .IN1(
        \r60/SUMB[5][6] ), .COUT(\r60/CARRYB[6][5] ), .SUM(\r60/SUMB[6][5] )
         );
  FADDER \r60/S2_6_4  ( .CIN(\r60/ab[6][4] ), .IN0(\r60/CARRYB[5][4] ), .IN1(
        \r60/SUMB[5][5] ), .COUT(\r60/CARRYB[6][4] ), .SUM(\r60/SUMB[6][4] )
         );
  FADDER \r60/S2_6_3  ( .CIN(\r60/ab[6][3] ), .IN0(\r60/CARRYB[5][3] ), .IN1(
        \r60/SUMB[5][4] ), .COUT(\r60/CARRYB[6][3] ), .SUM(\r60/SUMB[6][3] )
         );
  FADDER \r60/S2_6_2  ( .CIN(\r60/ab[6][2] ), .IN0(\r60/CARRYB[5][2] ), .IN1(
        \r60/SUMB[5][3] ), .COUT(\r60/CARRYB[6][2] ), .SUM(\r60/SUMB[6][2] )
         );
  FADDER \r60/S2_6_1  ( .CIN(\r60/ab[6][1] ), .IN0(\r60/CARRYB[5][1] ), .IN1(
        \r60/SUMB[5][2] ), .COUT(\r60/CARRYB[6][1] ), .SUM(\r60/SUMB[6][1] )
         );
  FADDER \r60/S1_6_0  ( .CIN(\r60/ab[6][0] ), .IN0(\r60/CARRYB[5][0] ), .IN1(
        \r60/SUMB[5][1] ), .COUT(\r60/CARRYB[6][0] ), .SUM(N123) );
  FADDER \r60/S3_7_30  ( .CIN(\r60/ab[7][30] ), .IN0(\r60/CARRYB[6][30] ), 
        .IN1(\r60/ab[6][31] ), .COUT(\r60/CARRYB[7][30] ), .SUM(
        \r60/SUMB[7][30] ) );
  FADDER \r60/S2_7_29  ( .CIN(\r60/ab[7][29] ), .IN0(\r60/CARRYB[6][29] ), 
        .IN1(\r60/SUMB[6][30] ), .COUT(\r60/CARRYB[7][29] ), .SUM(
        \r60/SUMB[7][29] ) );
  FADDER \r60/S2_7_28  ( .CIN(\r60/ab[7][28] ), .IN0(\r60/CARRYB[6][28] ), 
        .IN1(\r60/SUMB[6][29] ), .COUT(\r60/CARRYB[7][28] ), .SUM(
        \r60/SUMB[7][28] ) );
  FADDER \r60/S2_7_27  ( .CIN(\r60/ab[7][27] ), .IN0(\r60/CARRYB[6][27] ), 
        .IN1(\r60/SUMB[6][28] ), .COUT(\r60/CARRYB[7][27] ), .SUM(
        \r60/SUMB[7][27] ) );
  FADDER \r60/S2_7_26  ( .CIN(\r60/ab[7][26] ), .IN0(\r60/CARRYB[6][26] ), 
        .IN1(\r60/SUMB[6][27] ), .COUT(\r60/CARRYB[7][26] ), .SUM(
        \r60/SUMB[7][26] ) );
  FADDER \r60/S2_7_25  ( .CIN(\r60/ab[7][25] ), .IN0(\r60/CARRYB[6][25] ), 
        .IN1(\r60/SUMB[6][26] ), .COUT(\r60/CARRYB[7][25] ), .SUM(
        \r60/SUMB[7][25] ) );
  FADDER \r60/S2_7_24  ( .CIN(\r60/ab[7][24] ), .IN0(\r60/CARRYB[6][24] ), 
        .IN1(\r60/SUMB[6][25] ), .COUT(\r60/CARRYB[7][24] ), .SUM(
        \r60/SUMB[7][24] ) );
  FADDER \r60/S2_7_23  ( .CIN(\r60/ab[7][23] ), .IN0(\r60/CARRYB[6][23] ), 
        .IN1(\r60/SUMB[6][24] ), .COUT(\r60/CARRYB[7][23] ), .SUM(
        \r60/SUMB[7][23] ) );
  FADDER \r60/S2_7_22  ( .CIN(\r60/ab[7][22] ), .IN0(\r60/CARRYB[6][22] ), 
        .IN1(\r60/SUMB[6][23] ), .COUT(\r60/CARRYB[7][22] ), .SUM(
        \r60/SUMB[7][22] ) );
  FADDER \r60/S2_7_21  ( .CIN(\r60/ab[7][21] ), .IN0(\r60/CARRYB[6][21] ), 
        .IN1(\r60/SUMB[6][22] ), .COUT(\r60/CARRYB[7][21] ), .SUM(
        \r60/SUMB[7][21] ) );
  FADDER \r60/S2_7_20  ( .CIN(\r60/ab[7][20] ), .IN0(\r60/CARRYB[6][20] ), 
        .IN1(\r60/SUMB[6][21] ), .COUT(\r60/CARRYB[7][20] ), .SUM(
        \r60/SUMB[7][20] ) );
  FADDER \r60/S2_7_19  ( .CIN(\r60/ab[7][19] ), .IN0(\r60/CARRYB[6][19] ), 
        .IN1(\r60/SUMB[6][20] ), .COUT(\r60/CARRYB[7][19] ), .SUM(
        \r60/SUMB[7][19] ) );
  FADDER \r60/S2_7_18  ( .CIN(\r60/ab[7][18] ), .IN0(\r60/CARRYB[6][18] ), 
        .IN1(\r60/SUMB[6][19] ), .COUT(\r60/CARRYB[7][18] ), .SUM(
        \r60/SUMB[7][18] ) );
  FADDER \r60/S2_7_17  ( .CIN(\r60/ab[7][17] ), .IN0(\r60/CARRYB[6][17] ), 
        .IN1(\r60/SUMB[6][18] ), .COUT(\r60/CARRYB[7][17] ), .SUM(
        \r60/SUMB[7][17] ) );
  FADDER \r60/S2_7_16  ( .CIN(\r60/ab[7][16] ), .IN0(\r60/CARRYB[6][16] ), 
        .IN1(\r60/SUMB[6][17] ), .COUT(\r60/CARRYB[7][16] ), .SUM(
        \r60/SUMB[7][16] ) );
  FADDER \r60/S2_7_15  ( .CIN(\r60/ab[7][15] ), .IN0(\r60/CARRYB[6][15] ), 
        .IN1(\r60/SUMB[6][16] ), .COUT(\r60/CARRYB[7][15] ), .SUM(
        \r60/SUMB[7][15] ) );
  FADDER \r60/S2_7_14  ( .CIN(\r60/ab[7][14] ), .IN0(\r60/CARRYB[6][14] ), 
        .IN1(\r60/SUMB[6][15] ), .COUT(\r60/CARRYB[7][14] ), .SUM(
        \r60/SUMB[7][14] ) );
  FADDER \r60/S2_7_13  ( .CIN(\r60/ab[7][13] ), .IN0(\r60/CARRYB[6][13] ), 
        .IN1(\r60/SUMB[6][14] ), .COUT(\r60/CARRYB[7][13] ), .SUM(
        \r60/SUMB[7][13] ) );
  FADDER \r60/S2_7_12  ( .CIN(\r60/ab[7][12] ), .IN0(\r60/CARRYB[6][12] ), 
        .IN1(\r60/SUMB[6][13] ), .COUT(\r60/CARRYB[7][12] ), .SUM(
        \r60/SUMB[7][12] ) );
  FADDER \r60/S2_7_11  ( .CIN(\r60/ab[7][11] ), .IN0(\r60/CARRYB[6][11] ), 
        .IN1(\r60/SUMB[6][12] ), .COUT(\r60/CARRYB[7][11] ), .SUM(
        \r60/SUMB[7][11] ) );
  FADDER \r60/S2_7_10  ( .CIN(\r60/ab[7][10] ), .IN0(\r60/CARRYB[6][10] ), 
        .IN1(\r60/SUMB[6][11] ), .COUT(\r60/CARRYB[7][10] ), .SUM(
        \r60/SUMB[7][10] ) );
  FADDER \r60/S2_7_9  ( .CIN(\r60/ab[7][9] ), .IN0(\r60/CARRYB[6][9] ), .IN1(
        \r60/SUMB[6][10] ), .COUT(\r60/CARRYB[7][9] ), .SUM(\r60/SUMB[7][9] )
         );
  FADDER \r60/S2_7_8  ( .CIN(\r60/ab[7][8] ), .IN0(\r60/CARRYB[6][8] ), .IN1(
        \r60/SUMB[6][9] ), .COUT(\r60/CARRYB[7][8] ), .SUM(\r60/SUMB[7][8] )
         );
  FADDER \r60/S2_7_7  ( .CIN(\r60/ab[7][7] ), .IN0(\r60/CARRYB[6][7] ), .IN1(
        \r60/SUMB[6][8] ), .COUT(\r60/CARRYB[7][7] ), .SUM(\r60/SUMB[7][7] )
         );
  FADDER \r60/S2_7_6  ( .CIN(\r60/ab[7][6] ), .IN0(\r60/CARRYB[6][6] ), .IN1(
        \r60/SUMB[6][7] ), .COUT(\r60/CARRYB[7][6] ), .SUM(\r60/SUMB[7][6] )
         );
  FADDER \r60/S2_7_5  ( .CIN(\r60/ab[7][5] ), .IN0(\r60/CARRYB[6][5] ), .IN1(
        \r60/SUMB[6][6] ), .COUT(\r60/CARRYB[7][5] ), .SUM(\r60/SUMB[7][5] )
         );
  FADDER \r60/S2_7_4  ( .CIN(\r60/ab[7][4] ), .IN0(\r60/CARRYB[6][4] ), .IN1(
        \r60/SUMB[6][5] ), .COUT(\r60/CARRYB[7][4] ), .SUM(\r60/SUMB[7][4] )
         );
  FADDER \r60/S2_7_3  ( .CIN(\r60/ab[7][3] ), .IN0(\r60/CARRYB[6][3] ), .IN1(
        \r60/SUMB[6][4] ), .COUT(\r60/CARRYB[7][3] ), .SUM(\r60/SUMB[7][3] )
         );
  FADDER \r60/S2_7_2  ( .CIN(\r60/ab[7][2] ), .IN0(\r60/CARRYB[6][2] ), .IN1(
        \r60/SUMB[6][3] ), .COUT(\r60/CARRYB[7][2] ), .SUM(\r60/SUMB[7][2] )
         );
  FADDER \r60/S2_7_1  ( .CIN(\r60/ab[7][1] ), .IN0(\r60/CARRYB[6][1] ), .IN1(
        \r60/SUMB[6][2] ), .COUT(\r60/CARRYB[7][1] ), .SUM(\r60/SUMB[7][1] )
         );
  FADDER \r60/S1_7_0  ( .CIN(\r60/ab[7][0] ), .IN0(\r60/CARRYB[6][0] ), .IN1(
        \r60/SUMB[6][1] ), .COUT(\r60/CARRYB[7][0] ), .SUM(N124) );
  FADDER \r60/S3_8_30  ( .CIN(\r60/ab[8][30] ), .IN0(\r60/CARRYB[7][30] ), 
        .IN1(\r60/ab[7][31] ), .COUT(\r60/CARRYB[8][30] ), .SUM(
        \r60/SUMB[8][30] ) );
  FADDER \r60/S2_8_29  ( .CIN(\r60/ab[8][29] ), .IN0(\r60/CARRYB[7][29] ), 
        .IN1(\r60/SUMB[7][30] ), .COUT(\r60/CARRYB[8][29] ), .SUM(
        \r60/SUMB[8][29] ) );
  FADDER \r60/S2_8_28  ( .CIN(\r60/ab[8][28] ), .IN0(\r60/CARRYB[7][28] ), 
        .IN1(\r60/SUMB[7][29] ), .COUT(\r60/CARRYB[8][28] ), .SUM(
        \r60/SUMB[8][28] ) );
  FADDER \r60/S2_8_27  ( .CIN(\r60/ab[8][27] ), .IN0(\r60/CARRYB[7][27] ), 
        .IN1(\r60/SUMB[7][28] ), .COUT(\r60/CARRYB[8][27] ), .SUM(
        \r60/SUMB[8][27] ) );
  FADDER \r60/S2_8_26  ( .CIN(\r60/ab[8][26] ), .IN0(\r60/CARRYB[7][26] ), 
        .IN1(\r60/SUMB[7][27] ), .COUT(\r60/CARRYB[8][26] ), .SUM(
        \r60/SUMB[8][26] ) );
  FADDER \r60/S2_8_25  ( .CIN(\r60/ab[8][25] ), .IN0(\r60/CARRYB[7][25] ), 
        .IN1(\r60/SUMB[7][26] ), .COUT(\r60/CARRYB[8][25] ), .SUM(
        \r60/SUMB[8][25] ) );
  FADDER \r60/S2_8_24  ( .CIN(\r60/ab[8][24] ), .IN0(\r60/CARRYB[7][24] ), 
        .IN1(\r60/SUMB[7][25] ), .COUT(\r60/CARRYB[8][24] ), .SUM(
        \r60/SUMB[8][24] ) );
  FADDER \r60/S2_8_23  ( .CIN(\r60/ab[8][23] ), .IN0(\r60/CARRYB[7][23] ), 
        .IN1(\r60/SUMB[7][24] ), .COUT(\r60/CARRYB[8][23] ), .SUM(
        \r60/SUMB[8][23] ) );
  FADDER \r60/S2_8_22  ( .CIN(\r60/ab[8][22] ), .IN0(\r60/CARRYB[7][22] ), 
        .IN1(\r60/SUMB[7][23] ), .COUT(\r60/CARRYB[8][22] ), .SUM(
        \r60/SUMB[8][22] ) );
  FADDER \r60/S2_8_21  ( .CIN(\r60/ab[8][21] ), .IN0(\r60/CARRYB[7][21] ), 
        .IN1(\r60/SUMB[7][22] ), .COUT(\r60/CARRYB[8][21] ), .SUM(
        \r60/SUMB[8][21] ) );
  FADDER \r60/S2_8_20  ( .CIN(\r60/ab[8][20] ), .IN0(\r60/CARRYB[7][20] ), 
        .IN1(\r60/SUMB[7][21] ), .COUT(\r60/CARRYB[8][20] ), .SUM(
        \r60/SUMB[8][20] ) );
  FADDER \r60/S2_8_19  ( .CIN(\r60/ab[8][19] ), .IN0(\r60/CARRYB[7][19] ), 
        .IN1(\r60/SUMB[7][20] ), .COUT(\r60/CARRYB[8][19] ), .SUM(
        \r60/SUMB[8][19] ) );
  FADDER \r60/S2_8_18  ( .CIN(\r60/ab[8][18] ), .IN0(\r60/CARRYB[7][18] ), 
        .IN1(\r60/SUMB[7][19] ), .COUT(\r60/CARRYB[8][18] ), .SUM(
        \r60/SUMB[8][18] ) );
  FADDER \r60/S2_8_17  ( .CIN(\r60/ab[8][17] ), .IN0(\r60/CARRYB[7][17] ), 
        .IN1(\r60/SUMB[7][18] ), .COUT(\r60/CARRYB[8][17] ), .SUM(
        \r60/SUMB[8][17] ) );
  FADDER \r60/S2_8_16  ( .CIN(\r60/ab[8][16] ), .IN0(\r60/CARRYB[7][16] ), 
        .IN1(\r60/SUMB[7][17] ), .COUT(\r60/CARRYB[8][16] ), .SUM(
        \r60/SUMB[8][16] ) );
  FADDER \r60/S2_8_15  ( .CIN(\r60/ab[8][15] ), .IN0(\r60/CARRYB[7][15] ), 
        .IN1(\r60/SUMB[7][16] ), .COUT(\r60/CARRYB[8][15] ), .SUM(
        \r60/SUMB[8][15] ) );
  FADDER \r60/S2_8_14  ( .CIN(\r60/ab[8][14] ), .IN0(\r60/CARRYB[7][14] ), 
        .IN1(\r60/SUMB[7][15] ), .COUT(\r60/CARRYB[8][14] ), .SUM(
        \r60/SUMB[8][14] ) );
  FADDER \r60/S2_8_13  ( .CIN(\r60/ab[8][13] ), .IN0(\r60/CARRYB[7][13] ), 
        .IN1(\r60/SUMB[7][14] ), .COUT(\r60/CARRYB[8][13] ), .SUM(
        \r60/SUMB[8][13] ) );
  FADDER \r60/S2_8_12  ( .CIN(\r60/ab[8][12] ), .IN0(\r60/CARRYB[7][12] ), 
        .IN1(\r60/SUMB[7][13] ), .COUT(\r60/CARRYB[8][12] ), .SUM(
        \r60/SUMB[8][12] ) );
  FADDER \r60/S2_8_11  ( .CIN(\r60/ab[8][11] ), .IN0(\r60/CARRYB[7][11] ), 
        .IN1(\r60/SUMB[7][12] ), .COUT(\r60/CARRYB[8][11] ), .SUM(
        \r60/SUMB[8][11] ) );
  FADDER \r60/S2_8_10  ( .CIN(\r60/ab[8][10] ), .IN0(\r60/CARRYB[7][10] ), 
        .IN1(\r60/SUMB[7][11] ), .COUT(\r60/CARRYB[8][10] ), .SUM(
        \r60/SUMB[8][10] ) );
  FADDER \r60/S2_8_9  ( .CIN(\r60/ab[8][9] ), .IN0(\r60/CARRYB[7][9] ), .IN1(
        \r60/SUMB[7][10] ), .COUT(\r60/CARRYB[8][9] ), .SUM(\r60/SUMB[8][9] )
         );
  FADDER \r60/S2_8_8  ( .CIN(\r60/ab[8][8] ), .IN0(\r60/CARRYB[7][8] ), .IN1(
        \r60/SUMB[7][9] ), .COUT(\r60/CARRYB[8][8] ), .SUM(\r60/SUMB[8][8] )
         );
  FADDER \r60/S2_8_7  ( .CIN(\r60/ab[8][7] ), .IN0(\r60/CARRYB[7][7] ), .IN1(
        \r60/SUMB[7][8] ), .COUT(\r60/CARRYB[8][7] ), .SUM(\r60/SUMB[8][7] )
         );
  FADDER \r60/S2_8_6  ( .CIN(\r60/ab[8][6] ), .IN0(\r60/CARRYB[7][6] ), .IN1(
        \r60/SUMB[7][7] ), .COUT(\r60/CARRYB[8][6] ), .SUM(\r60/SUMB[8][6] )
         );
  FADDER \r60/S2_8_5  ( .CIN(\r60/ab[8][5] ), .IN0(\r60/CARRYB[7][5] ), .IN1(
        \r60/SUMB[7][6] ), .COUT(\r60/CARRYB[8][5] ), .SUM(\r60/SUMB[8][5] )
         );
  FADDER \r60/S2_8_4  ( .CIN(\r60/ab[8][4] ), .IN0(\r60/CARRYB[7][4] ), .IN1(
        \r60/SUMB[7][5] ), .COUT(\r60/CARRYB[8][4] ), .SUM(\r60/SUMB[8][4] )
         );
  FADDER \r60/S2_8_3  ( .CIN(\r60/ab[8][3] ), .IN0(\r60/CARRYB[7][3] ), .IN1(
        \r60/SUMB[7][4] ), .COUT(\r60/CARRYB[8][3] ), .SUM(\r60/SUMB[8][3] )
         );
  FADDER \r60/S2_8_2  ( .CIN(\r60/ab[8][2] ), .IN0(\r60/CARRYB[7][2] ), .IN1(
        \r60/SUMB[7][3] ), .COUT(\r60/CARRYB[8][2] ), .SUM(\r60/SUMB[8][2] )
         );
  FADDER \r60/S2_8_1  ( .CIN(\r60/ab[8][1] ), .IN0(\r60/CARRYB[7][1] ), .IN1(
        \r60/SUMB[7][2] ), .COUT(\r60/CARRYB[8][1] ), .SUM(\r60/SUMB[8][1] )
         );
  FADDER \r60/S1_8_0  ( .CIN(\r60/ab[8][0] ), .IN0(\r60/CARRYB[7][0] ), .IN1(
        \r60/SUMB[7][1] ), .COUT(\r60/CARRYB[8][0] ), .SUM(N125) );
  FADDER \r60/S3_9_30  ( .CIN(\r60/ab[9][30] ), .IN0(\r60/CARRYB[8][30] ), 
        .IN1(\r60/ab[8][31] ), .COUT(\r60/CARRYB[9][30] ), .SUM(
        \r60/SUMB[9][30] ) );
  FADDER \r60/S2_9_29  ( .CIN(\r60/ab[9][29] ), .IN0(\r60/CARRYB[8][29] ), 
        .IN1(\r60/SUMB[8][30] ), .COUT(\r60/CARRYB[9][29] ), .SUM(
        \r60/SUMB[9][29] ) );
  FADDER \r60/S2_9_28  ( .CIN(\r60/ab[9][28] ), .IN0(\r60/CARRYB[8][28] ), 
        .IN1(\r60/SUMB[8][29] ), .COUT(\r60/CARRYB[9][28] ), .SUM(
        \r60/SUMB[9][28] ) );
  FADDER \r60/S2_9_27  ( .CIN(\r60/ab[9][27] ), .IN0(\r60/CARRYB[8][27] ), 
        .IN1(\r60/SUMB[8][28] ), .COUT(\r60/CARRYB[9][27] ), .SUM(
        \r60/SUMB[9][27] ) );
  FADDER \r60/S2_9_26  ( .CIN(\r60/ab[9][26] ), .IN0(\r60/CARRYB[8][26] ), 
        .IN1(\r60/SUMB[8][27] ), .COUT(\r60/CARRYB[9][26] ), .SUM(
        \r60/SUMB[9][26] ) );
  FADDER \r60/S2_9_25  ( .CIN(\r60/ab[9][25] ), .IN0(\r60/CARRYB[8][25] ), 
        .IN1(\r60/SUMB[8][26] ), .COUT(\r60/CARRYB[9][25] ), .SUM(
        \r60/SUMB[9][25] ) );
  FADDER \r60/S2_9_24  ( .CIN(\r60/ab[9][24] ), .IN0(\r60/CARRYB[8][24] ), 
        .IN1(\r60/SUMB[8][25] ), .COUT(\r60/CARRYB[9][24] ), .SUM(
        \r60/SUMB[9][24] ) );
  FADDER \r60/S2_9_23  ( .CIN(\r60/ab[9][23] ), .IN0(\r60/CARRYB[8][23] ), 
        .IN1(\r60/SUMB[8][24] ), .COUT(\r60/CARRYB[9][23] ), .SUM(
        \r60/SUMB[9][23] ) );
  FADDER \r60/S2_9_22  ( .CIN(\r60/ab[9][22] ), .IN0(\r60/CARRYB[8][22] ), 
        .IN1(\r60/SUMB[8][23] ), .COUT(\r60/CARRYB[9][22] ), .SUM(
        \r60/SUMB[9][22] ) );
  FADDER \r60/S2_9_21  ( .CIN(\r60/ab[9][21] ), .IN0(\r60/CARRYB[8][21] ), 
        .IN1(\r60/SUMB[8][22] ), .COUT(\r60/CARRYB[9][21] ), .SUM(
        \r60/SUMB[9][21] ) );
  FADDER \r60/S2_9_20  ( .CIN(\r60/ab[9][20] ), .IN0(\r60/CARRYB[8][20] ), 
        .IN1(\r60/SUMB[8][21] ), .COUT(\r60/CARRYB[9][20] ), .SUM(
        \r60/SUMB[9][20] ) );
  FADDER \r60/S2_9_19  ( .CIN(\r60/ab[9][19] ), .IN0(\r60/CARRYB[8][19] ), 
        .IN1(\r60/SUMB[8][20] ), .COUT(\r60/CARRYB[9][19] ), .SUM(
        \r60/SUMB[9][19] ) );
  FADDER \r60/S2_9_18  ( .CIN(\r60/ab[9][18] ), .IN0(\r60/CARRYB[8][18] ), 
        .IN1(\r60/SUMB[8][19] ), .COUT(\r60/CARRYB[9][18] ), .SUM(
        \r60/SUMB[9][18] ) );
  FADDER \r60/S2_9_17  ( .CIN(\r60/ab[9][17] ), .IN0(\r60/CARRYB[8][17] ), 
        .IN1(\r60/SUMB[8][18] ), .COUT(\r60/CARRYB[9][17] ), .SUM(
        \r60/SUMB[9][17] ) );
  FADDER \r60/S2_9_16  ( .CIN(\r60/ab[9][16] ), .IN0(\r60/CARRYB[8][16] ), 
        .IN1(\r60/SUMB[8][17] ), .COUT(\r60/CARRYB[9][16] ), .SUM(
        \r60/SUMB[9][16] ) );
  FADDER \r60/S2_9_15  ( .CIN(\r60/ab[9][15] ), .IN0(\r60/CARRYB[8][15] ), 
        .IN1(\r60/SUMB[8][16] ), .COUT(\r60/CARRYB[9][15] ), .SUM(
        \r60/SUMB[9][15] ) );
  FADDER \r60/S2_9_14  ( .CIN(\r60/ab[9][14] ), .IN0(\r60/CARRYB[8][14] ), 
        .IN1(\r60/SUMB[8][15] ), .COUT(\r60/CARRYB[9][14] ), .SUM(
        \r60/SUMB[9][14] ) );
  FADDER \r60/S2_9_13  ( .CIN(\r60/ab[9][13] ), .IN0(\r60/CARRYB[8][13] ), 
        .IN1(\r60/SUMB[8][14] ), .COUT(\r60/CARRYB[9][13] ), .SUM(
        \r60/SUMB[9][13] ) );
  FADDER \r60/S2_9_12  ( .CIN(\r60/ab[9][12] ), .IN0(\r60/CARRYB[8][12] ), 
        .IN1(\r60/SUMB[8][13] ), .COUT(\r60/CARRYB[9][12] ), .SUM(
        \r60/SUMB[9][12] ) );
  FADDER \r60/S2_9_11  ( .CIN(\r60/ab[9][11] ), .IN0(\r60/CARRYB[8][11] ), 
        .IN1(\r60/SUMB[8][12] ), .COUT(\r60/CARRYB[9][11] ), .SUM(
        \r60/SUMB[9][11] ) );
  FADDER \r60/S2_9_10  ( .CIN(\r60/ab[9][10] ), .IN0(\r60/CARRYB[8][10] ), 
        .IN1(\r60/SUMB[8][11] ), .COUT(\r60/CARRYB[9][10] ), .SUM(
        \r60/SUMB[9][10] ) );
  FADDER \r60/S2_9_9  ( .CIN(\r60/ab[9][9] ), .IN0(\r60/CARRYB[8][9] ), .IN1(
        \r60/SUMB[8][10] ), .COUT(\r60/CARRYB[9][9] ), .SUM(\r60/SUMB[9][9] )
         );
  FADDER \r60/S2_9_8  ( .CIN(\r60/ab[9][8] ), .IN0(\r60/CARRYB[8][8] ), .IN1(
        \r60/SUMB[8][9] ), .COUT(\r60/CARRYB[9][8] ), .SUM(\r60/SUMB[9][8] )
         );
  FADDER \r60/S2_9_7  ( .CIN(\r60/ab[9][7] ), .IN0(\r60/CARRYB[8][7] ), .IN1(
        \r60/SUMB[8][8] ), .COUT(\r60/CARRYB[9][7] ), .SUM(\r60/SUMB[9][7] )
         );
  FADDER \r60/S2_9_6  ( .CIN(\r60/ab[9][6] ), .IN0(\r60/CARRYB[8][6] ), .IN1(
        \r60/SUMB[8][7] ), .COUT(\r60/CARRYB[9][6] ), .SUM(\r60/SUMB[9][6] )
         );
  FADDER \r60/S2_9_5  ( .CIN(\r60/ab[9][5] ), .IN0(\r60/CARRYB[8][5] ), .IN1(
        \r60/SUMB[8][6] ), .COUT(\r60/CARRYB[9][5] ), .SUM(\r60/SUMB[9][5] )
         );
  FADDER \r60/S2_9_4  ( .CIN(\r60/ab[9][4] ), .IN0(\r60/CARRYB[8][4] ), .IN1(
        \r60/SUMB[8][5] ), .COUT(\r60/CARRYB[9][4] ), .SUM(\r60/SUMB[9][4] )
         );
  FADDER \r60/S2_9_3  ( .CIN(\r60/ab[9][3] ), .IN0(\r60/CARRYB[8][3] ), .IN1(
        \r60/SUMB[8][4] ), .COUT(\r60/CARRYB[9][3] ), .SUM(\r60/SUMB[9][3] )
         );
  FADDER \r60/S2_9_2  ( .CIN(\r60/ab[9][2] ), .IN0(\r60/CARRYB[8][2] ), .IN1(
        \r60/SUMB[8][3] ), .COUT(\r60/CARRYB[9][2] ), .SUM(\r60/SUMB[9][2] )
         );
  FADDER \r60/S2_9_1  ( .CIN(\r60/ab[9][1] ), .IN0(\r60/CARRYB[8][1] ), .IN1(
        \r60/SUMB[8][2] ), .COUT(\r60/CARRYB[9][1] ), .SUM(\r60/SUMB[9][1] )
         );
  FADDER \r60/S1_9_0  ( .CIN(\r60/ab[9][0] ), .IN0(\r60/CARRYB[8][0] ), .IN1(
        \r60/SUMB[8][1] ), .COUT(\r60/CARRYB[9][0] ), .SUM(N126) );
  FADDER \r60/S3_10_30  ( .CIN(\r60/ab[10][30] ), .IN0(\r60/CARRYB[9][30] ), 
        .IN1(\r60/ab[9][31] ), .COUT(\r60/CARRYB[10][30] ), .SUM(
        \r60/SUMB[10][30] ) );
  FADDER \r60/S2_10_29  ( .CIN(\r60/ab[10][29] ), .IN0(\r60/CARRYB[9][29] ), 
        .IN1(\r60/SUMB[9][30] ), .COUT(\r60/CARRYB[10][29] ), .SUM(
        \r60/SUMB[10][29] ) );
  FADDER \r60/S2_10_28  ( .CIN(\r60/ab[10][28] ), .IN0(\r60/CARRYB[9][28] ), 
        .IN1(\r60/SUMB[9][29] ), .COUT(\r60/CARRYB[10][28] ), .SUM(
        \r60/SUMB[10][28] ) );
  FADDER \r60/S2_10_27  ( .CIN(\r60/ab[10][27] ), .IN0(\r60/CARRYB[9][27] ), 
        .IN1(\r60/SUMB[9][28] ), .COUT(\r60/CARRYB[10][27] ), .SUM(
        \r60/SUMB[10][27] ) );
  FADDER \r60/S2_10_26  ( .CIN(\r60/ab[10][26] ), .IN0(\r60/CARRYB[9][26] ), 
        .IN1(\r60/SUMB[9][27] ), .COUT(\r60/CARRYB[10][26] ), .SUM(
        \r60/SUMB[10][26] ) );
  FADDER \r60/S2_10_25  ( .CIN(\r60/ab[10][25] ), .IN0(\r60/CARRYB[9][25] ), 
        .IN1(\r60/SUMB[9][26] ), .COUT(\r60/CARRYB[10][25] ), .SUM(
        \r60/SUMB[10][25] ) );
  FADDER \r60/S2_10_24  ( .CIN(\r60/ab[10][24] ), .IN0(\r60/CARRYB[9][24] ), 
        .IN1(\r60/SUMB[9][25] ), .COUT(\r60/CARRYB[10][24] ), .SUM(
        \r60/SUMB[10][24] ) );
  FADDER \r60/S2_10_23  ( .CIN(\r60/ab[10][23] ), .IN0(\r60/CARRYB[9][23] ), 
        .IN1(\r60/SUMB[9][24] ), .COUT(\r60/CARRYB[10][23] ), .SUM(
        \r60/SUMB[10][23] ) );
  FADDER \r60/S2_10_22  ( .CIN(\r60/ab[10][22] ), .IN0(\r60/CARRYB[9][22] ), 
        .IN1(\r60/SUMB[9][23] ), .COUT(\r60/CARRYB[10][22] ), .SUM(
        \r60/SUMB[10][22] ) );
  FADDER \r60/S2_10_21  ( .CIN(\r60/ab[10][21] ), .IN0(\r60/CARRYB[9][21] ), 
        .IN1(\r60/SUMB[9][22] ), .COUT(\r60/CARRYB[10][21] ), .SUM(
        \r60/SUMB[10][21] ) );
  FADDER \r60/S2_10_20  ( .CIN(\r60/ab[10][20] ), .IN0(\r60/CARRYB[9][20] ), 
        .IN1(\r60/SUMB[9][21] ), .COUT(\r60/CARRYB[10][20] ), .SUM(
        \r60/SUMB[10][20] ) );
  FADDER \r60/S2_10_19  ( .CIN(\r60/ab[10][19] ), .IN0(\r60/CARRYB[9][19] ), 
        .IN1(\r60/SUMB[9][20] ), .COUT(\r60/CARRYB[10][19] ), .SUM(
        \r60/SUMB[10][19] ) );
  FADDER \r60/S2_10_18  ( .CIN(\r60/ab[10][18] ), .IN0(\r60/CARRYB[9][18] ), 
        .IN1(\r60/SUMB[9][19] ), .COUT(\r60/CARRYB[10][18] ), .SUM(
        \r60/SUMB[10][18] ) );
  FADDER \r60/S2_10_17  ( .CIN(\r60/ab[10][17] ), .IN0(\r60/CARRYB[9][17] ), 
        .IN1(\r60/SUMB[9][18] ), .COUT(\r60/CARRYB[10][17] ), .SUM(
        \r60/SUMB[10][17] ) );
  FADDER \r60/S2_10_16  ( .CIN(\r60/ab[10][16] ), .IN0(\r60/CARRYB[9][16] ), 
        .IN1(\r60/SUMB[9][17] ), .COUT(\r60/CARRYB[10][16] ), .SUM(
        \r60/SUMB[10][16] ) );
  FADDER \r60/S2_10_15  ( .CIN(\r60/ab[10][15] ), .IN0(\r60/CARRYB[9][15] ), 
        .IN1(\r60/SUMB[9][16] ), .COUT(\r60/CARRYB[10][15] ), .SUM(
        \r60/SUMB[10][15] ) );
  FADDER \r60/S2_10_14  ( .CIN(\r60/ab[10][14] ), .IN0(\r60/CARRYB[9][14] ), 
        .IN1(\r60/SUMB[9][15] ), .COUT(\r60/CARRYB[10][14] ), .SUM(
        \r60/SUMB[10][14] ) );
  FADDER \r60/S2_10_13  ( .CIN(\r60/ab[10][13] ), .IN0(\r60/CARRYB[9][13] ), 
        .IN1(\r60/SUMB[9][14] ), .COUT(\r60/CARRYB[10][13] ), .SUM(
        \r60/SUMB[10][13] ) );
  FADDER \r60/S2_10_12  ( .CIN(\r60/ab[10][12] ), .IN0(\r60/CARRYB[9][12] ), 
        .IN1(\r60/SUMB[9][13] ), .COUT(\r60/CARRYB[10][12] ), .SUM(
        \r60/SUMB[10][12] ) );
  FADDER \r60/S2_10_11  ( .CIN(\r60/ab[10][11] ), .IN0(\r60/CARRYB[9][11] ), 
        .IN1(\r60/SUMB[9][12] ), .COUT(\r60/CARRYB[10][11] ), .SUM(
        \r60/SUMB[10][11] ) );
  FADDER \r60/S2_10_10  ( .CIN(\r60/ab[10][10] ), .IN0(\r60/CARRYB[9][10] ), 
        .IN1(\r60/SUMB[9][11] ), .COUT(\r60/CARRYB[10][10] ), .SUM(
        \r60/SUMB[10][10] ) );
  FADDER \r60/S2_10_9  ( .CIN(\r60/ab[10][9] ), .IN0(\r60/CARRYB[9][9] ), 
        .IN1(\r60/SUMB[9][10] ), .COUT(\r60/CARRYB[10][9] ), .SUM(
        \r60/SUMB[10][9] ) );
  FADDER \r60/S2_10_8  ( .CIN(\r60/ab[10][8] ), .IN0(\r60/CARRYB[9][8] ), 
        .IN1(\r60/SUMB[9][9] ), .COUT(\r60/CARRYB[10][8] ), .SUM(
        \r60/SUMB[10][8] ) );
  FADDER \r60/S2_10_7  ( .CIN(\r60/ab[10][7] ), .IN0(\r60/CARRYB[9][7] ), 
        .IN1(\r60/SUMB[9][8] ), .COUT(\r60/CARRYB[10][7] ), .SUM(
        \r60/SUMB[10][7] ) );
  FADDER \r60/S2_10_6  ( .CIN(\r60/ab[10][6] ), .IN0(\r60/CARRYB[9][6] ), 
        .IN1(\r60/SUMB[9][7] ), .COUT(\r60/CARRYB[10][6] ), .SUM(
        \r60/SUMB[10][6] ) );
  FADDER \r60/S2_10_5  ( .CIN(\r60/ab[10][5] ), .IN0(\r60/CARRYB[9][5] ), 
        .IN1(\r60/SUMB[9][6] ), .COUT(\r60/CARRYB[10][5] ), .SUM(
        \r60/SUMB[10][5] ) );
  FADDER \r60/S2_10_4  ( .CIN(\r60/ab[10][4] ), .IN0(\r60/CARRYB[9][4] ), 
        .IN1(\r60/SUMB[9][5] ), .COUT(\r60/CARRYB[10][4] ), .SUM(
        \r60/SUMB[10][4] ) );
  FADDER \r60/S2_10_3  ( .CIN(\r60/ab[10][3] ), .IN0(\r60/CARRYB[9][3] ), 
        .IN1(\r60/SUMB[9][4] ), .COUT(\r60/CARRYB[10][3] ), .SUM(
        \r60/SUMB[10][3] ) );
  FADDER \r60/S2_10_2  ( .CIN(\r60/ab[10][2] ), .IN0(\r60/CARRYB[9][2] ), 
        .IN1(\r60/SUMB[9][3] ), .COUT(\r60/CARRYB[10][2] ), .SUM(
        \r60/SUMB[10][2] ) );
  FADDER \r60/S2_10_1  ( .CIN(\r60/ab[10][1] ), .IN0(\r60/CARRYB[9][1] ), 
        .IN1(\r60/SUMB[9][2] ), .COUT(\r60/CARRYB[10][1] ), .SUM(
        \r60/SUMB[10][1] ) );
  FADDER \r60/S1_10_0  ( .CIN(\r60/ab[10][0] ), .IN0(\r60/CARRYB[9][0] ), 
        .IN1(\r60/SUMB[9][1] ), .COUT(\r60/CARRYB[10][0] ), .SUM(N127) );
  FADDER \r60/S3_11_30  ( .CIN(\r60/ab[11][30] ), .IN0(\r60/CARRYB[10][30] ), 
        .IN1(\r60/ab[10][31] ), .COUT(\r60/CARRYB[11][30] ), .SUM(
        \r60/SUMB[11][30] ) );
  FADDER \r60/S2_11_29  ( .CIN(\r60/ab[11][29] ), .IN0(\r60/CARRYB[10][29] ), 
        .IN1(\r60/SUMB[10][30] ), .COUT(\r60/CARRYB[11][29] ), .SUM(
        \r60/SUMB[11][29] ) );
  FADDER \r60/S2_11_28  ( .CIN(\r60/ab[11][28] ), .IN0(\r60/CARRYB[10][28] ), 
        .IN1(\r60/SUMB[10][29] ), .COUT(\r60/CARRYB[11][28] ), .SUM(
        \r60/SUMB[11][28] ) );
  FADDER \r60/S2_11_27  ( .CIN(\r60/ab[11][27] ), .IN0(\r60/CARRYB[10][27] ), 
        .IN1(\r60/SUMB[10][28] ), .COUT(\r60/CARRYB[11][27] ), .SUM(
        \r60/SUMB[11][27] ) );
  FADDER \r60/S2_11_26  ( .CIN(\r60/ab[11][26] ), .IN0(\r60/CARRYB[10][26] ), 
        .IN1(\r60/SUMB[10][27] ), .COUT(\r60/CARRYB[11][26] ), .SUM(
        \r60/SUMB[11][26] ) );
  FADDER \r60/S2_11_25  ( .CIN(\r60/ab[11][25] ), .IN0(\r60/CARRYB[10][25] ), 
        .IN1(\r60/SUMB[10][26] ), .COUT(\r60/CARRYB[11][25] ), .SUM(
        \r60/SUMB[11][25] ) );
  FADDER \r60/S2_11_24  ( .CIN(\r60/ab[11][24] ), .IN0(\r60/CARRYB[10][24] ), 
        .IN1(\r60/SUMB[10][25] ), .COUT(\r60/CARRYB[11][24] ), .SUM(
        \r60/SUMB[11][24] ) );
  FADDER \r60/S2_11_23  ( .CIN(\r60/ab[11][23] ), .IN0(\r60/CARRYB[10][23] ), 
        .IN1(\r60/SUMB[10][24] ), .COUT(\r60/CARRYB[11][23] ), .SUM(
        \r60/SUMB[11][23] ) );
  FADDER \r60/S2_11_22  ( .CIN(\r60/ab[11][22] ), .IN0(\r60/CARRYB[10][22] ), 
        .IN1(\r60/SUMB[10][23] ), .COUT(\r60/CARRYB[11][22] ), .SUM(
        \r60/SUMB[11][22] ) );
  FADDER \r60/S2_11_21  ( .CIN(\r60/ab[11][21] ), .IN0(\r60/CARRYB[10][21] ), 
        .IN1(\r60/SUMB[10][22] ), .COUT(\r60/CARRYB[11][21] ), .SUM(
        \r60/SUMB[11][21] ) );
  FADDER \r60/S2_11_20  ( .CIN(\r60/ab[11][20] ), .IN0(\r60/CARRYB[10][20] ), 
        .IN1(\r60/SUMB[10][21] ), .COUT(\r60/CARRYB[11][20] ), .SUM(
        \r60/SUMB[11][20] ) );
  FADDER \r60/S2_11_19  ( .CIN(\r60/ab[11][19] ), .IN0(\r60/CARRYB[10][19] ), 
        .IN1(\r60/SUMB[10][20] ), .COUT(\r60/CARRYB[11][19] ), .SUM(
        \r60/SUMB[11][19] ) );
  FADDER \r60/S2_11_18  ( .CIN(\r60/ab[11][18] ), .IN0(\r60/CARRYB[10][18] ), 
        .IN1(\r60/SUMB[10][19] ), .COUT(\r60/CARRYB[11][18] ), .SUM(
        \r60/SUMB[11][18] ) );
  FADDER \r60/S2_11_17  ( .CIN(\r60/ab[11][17] ), .IN0(\r60/CARRYB[10][17] ), 
        .IN1(\r60/SUMB[10][18] ), .COUT(\r60/CARRYB[11][17] ), .SUM(
        \r60/SUMB[11][17] ) );
  FADDER \r60/S2_11_16  ( .CIN(\r60/ab[11][16] ), .IN0(\r60/CARRYB[10][16] ), 
        .IN1(\r60/SUMB[10][17] ), .COUT(\r60/CARRYB[11][16] ), .SUM(
        \r60/SUMB[11][16] ) );
  FADDER \r60/S2_11_15  ( .CIN(\r60/ab[11][15] ), .IN0(\r60/CARRYB[10][15] ), 
        .IN1(\r60/SUMB[10][16] ), .COUT(\r60/CARRYB[11][15] ), .SUM(
        \r60/SUMB[11][15] ) );
  FADDER \r60/S2_11_14  ( .CIN(\r60/ab[11][14] ), .IN0(\r60/CARRYB[10][14] ), 
        .IN1(\r60/SUMB[10][15] ), .COUT(\r60/CARRYB[11][14] ), .SUM(
        \r60/SUMB[11][14] ) );
  FADDER \r60/S2_11_13  ( .CIN(\r60/ab[11][13] ), .IN0(\r60/CARRYB[10][13] ), 
        .IN1(\r60/SUMB[10][14] ), .COUT(\r60/CARRYB[11][13] ), .SUM(
        \r60/SUMB[11][13] ) );
  FADDER \r60/S2_11_12  ( .CIN(\r60/ab[11][12] ), .IN0(\r60/CARRYB[10][12] ), 
        .IN1(\r60/SUMB[10][13] ), .COUT(\r60/CARRYB[11][12] ), .SUM(
        \r60/SUMB[11][12] ) );
  FADDER \r60/S2_11_11  ( .CIN(\r60/ab[11][11] ), .IN0(\r60/CARRYB[10][11] ), 
        .IN1(\r60/SUMB[10][12] ), .COUT(\r60/CARRYB[11][11] ), .SUM(
        \r60/SUMB[11][11] ) );
  FADDER \r60/S2_11_10  ( .CIN(\r60/ab[11][10] ), .IN0(\r60/CARRYB[10][10] ), 
        .IN1(\r60/SUMB[10][11] ), .COUT(\r60/CARRYB[11][10] ), .SUM(
        \r60/SUMB[11][10] ) );
  FADDER \r60/S2_11_9  ( .CIN(\r60/ab[11][9] ), .IN0(\r60/CARRYB[10][9] ), 
        .IN1(\r60/SUMB[10][10] ), .COUT(\r60/CARRYB[11][9] ), .SUM(
        \r60/SUMB[11][9] ) );
  FADDER \r60/S2_11_8  ( .CIN(\r60/ab[11][8] ), .IN0(\r60/CARRYB[10][8] ), 
        .IN1(\r60/SUMB[10][9] ), .COUT(\r60/CARRYB[11][8] ), .SUM(
        \r60/SUMB[11][8] ) );
  FADDER \r60/S2_11_7  ( .CIN(\r60/ab[11][7] ), .IN0(\r60/CARRYB[10][7] ), 
        .IN1(\r60/SUMB[10][8] ), .COUT(\r60/CARRYB[11][7] ), .SUM(
        \r60/SUMB[11][7] ) );
  FADDER \r60/S2_11_6  ( .CIN(\r60/ab[11][6] ), .IN0(\r60/CARRYB[10][6] ), 
        .IN1(\r60/SUMB[10][7] ), .COUT(\r60/CARRYB[11][6] ), .SUM(
        \r60/SUMB[11][6] ) );
  FADDER \r60/S2_11_5  ( .CIN(\r60/ab[11][5] ), .IN0(\r60/CARRYB[10][5] ), 
        .IN1(\r60/SUMB[10][6] ), .COUT(\r60/CARRYB[11][5] ), .SUM(
        \r60/SUMB[11][5] ) );
  FADDER \r60/S2_11_4  ( .CIN(\r60/ab[11][4] ), .IN0(\r60/CARRYB[10][4] ), 
        .IN1(\r60/SUMB[10][5] ), .COUT(\r60/CARRYB[11][4] ), .SUM(
        \r60/SUMB[11][4] ) );
  FADDER \r60/S2_11_3  ( .CIN(\r60/ab[11][3] ), .IN0(\r60/CARRYB[10][3] ), 
        .IN1(\r60/SUMB[10][4] ), .COUT(\r60/CARRYB[11][3] ), .SUM(
        \r60/SUMB[11][3] ) );
  FADDER \r60/S2_11_2  ( .CIN(\r60/ab[11][2] ), .IN0(\r60/CARRYB[10][2] ), 
        .IN1(\r60/SUMB[10][3] ), .COUT(\r60/CARRYB[11][2] ), .SUM(
        \r60/SUMB[11][2] ) );
  FADDER \r60/S2_11_1  ( .CIN(\r60/ab[11][1] ), .IN0(\r60/CARRYB[10][1] ), 
        .IN1(\r60/SUMB[10][2] ), .COUT(\r60/CARRYB[11][1] ), .SUM(
        \r60/SUMB[11][1] ) );
  FADDER \r60/S1_11_0  ( .CIN(\r60/ab[11][0] ), .IN0(\r60/CARRYB[10][0] ), 
        .IN1(\r60/SUMB[10][1] ), .COUT(\r60/CARRYB[11][0] ), .SUM(N128) );
  FADDER \r60/S3_12_30  ( .CIN(\r60/ab[12][30] ), .IN0(\r60/CARRYB[11][30] ), 
        .IN1(\r60/ab[11][31] ), .COUT(\r60/CARRYB[12][30] ), .SUM(
        \r60/SUMB[12][30] ) );
  FADDER \r60/S2_12_29  ( .CIN(\r60/ab[12][29] ), .IN0(\r60/CARRYB[11][29] ), 
        .IN1(\r60/SUMB[11][30] ), .COUT(\r60/CARRYB[12][29] ), .SUM(
        \r60/SUMB[12][29] ) );
  FADDER \r60/S2_12_28  ( .CIN(\r60/ab[12][28] ), .IN0(\r60/CARRYB[11][28] ), 
        .IN1(\r60/SUMB[11][29] ), .COUT(\r60/CARRYB[12][28] ), .SUM(
        \r60/SUMB[12][28] ) );
  FADDER \r60/S2_12_27  ( .CIN(\r60/ab[12][27] ), .IN0(\r60/CARRYB[11][27] ), 
        .IN1(\r60/SUMB[11][28] ), .COUT(\r60/CARRYB[12][27] ), .SUM(
        \r60/SUMB[12][27] ) );
  FADDER \r60/S2_12_26  ( .CIN(\r60/ab[12][26] ), .IN0(\r60/CARRYB[11][26] ), 
        .IN1(\r60/SUMB[11][27] ), .COUT(\r60/CARRYB[12][26] ), .SUM(
        \r60/SUMB[12][26] ) );
  FADDER \r60/S2_12_25  ( .CIN(\r60/ab[12][25] ), .IN0(\r60/CARRYB[11][25] ), 
        .IN1(\r60/SUMB[11][26] ), .COUT(\r60/CARRYB[12][25] ), .SUM(
        \r60/SUMB[12][25] ) );
  FADDER \r60/S2_12_24  ( .CIN(\r60/ab[12][24] ), .IN0(\r60/CARRYB[11][24] ), 
        .IN1(\r60/SUMB[11][25] ), .COUT(\r60/CARRYB[12][24] ), .SUM(
        \r60/SUMB[12][24] ) );
  FADDER \r60/S2_12_23  ( .CIN(\r60/ab[12][23] ), .IN0(\r60/CARRYB[11][23] ), 
        .IN1(\r60/SUMB[11][24] ), .COUT(\r60/CARRYB[12][23] ), .SUM(
        \r60/SUMB[12][23] ) );
  FADDER \r60/S2_12_22  ( .CIN(\r60/ab[12][22] ), .IN0(\r60/CARRYB[11][22] ), 
        .IN1(\r60/SUMB[11][23] ), .COUT(\r60/CARRYB[12][22] ), .SUM(
        \r60/SUMB[12][22] ) );
  FADDER \r60/S2_12_21  ( .CIN(\r60/ab[12][21] ), .IN0(\r60/CARRYB[11][21] ), 
        .IN1(\r60/SUMB[11][22] ), .COUT(\r60/CARRYB[12][21] ), .SUM(
        \r60/SUMB[12][21] ) );
  FADDER \r60/S2_12_20  ( .CIN(\r60/ab[12][20] ), .IN0(\r60/CARRYB[11][20] ), 
        .IN1(\r60/SUMB[11][21] ), .COUT(\r60/CARRYB[12][20] ), .SUM(
        \r60/SUMB[12][20] ) );
  FADDER \r60/S2_12_19  ( .CIN(\r60/ab[12][19] ), .IN0(\r60/CARRYB[11][19] ), 
        .IN1(\r60/SUMB[11][20] ), .COUT(\r60/CARRYB[12][19] ), .SUM(
        \r60/SUMB[12][19] ) );
  FADDER \r60/S2_12_18  ( .CIN(\r60/ab[12][18] ), .IN0(\r60/CARRYB[11][18] ), 
        .IN1(\r60/SUMB[11][19] ), .COUT(\r60/CARRYB[12][18] ), .SUM(
        \r60/SUMB[12][18] ) );
  FADDER \r60/S2_12_17  ( .CIN(\r60/ab[12][17] ), .IN0(\r60/CARRYB[11][17] ), 
        .IN1(\r60/SUMB[11][18] ), .COUT(\r60/CARRYB[12][17] ), .SUM(
        \r60/SUMB[12][17] ) );
  FADDER \r60/S2_12_16  ( .CIN(\r60/ab[12][16] ), .IN0(\r60/CARRYB[11][16] ), 
        .IN1(\r60/SUMB[11][17] ), .COUT(\r60/CARRYB[12][16] ), .SUM(
        \r60/SUMB[12][16] ) );
  FADDER \r60/S2_12_15  ( .CIN(\r60/ab[12][15] ), .IN0(\r60/CARRYB[11][15] ), 
        .IN1(\r60/SUMB[11][16] ), .COUT(\r60/CARRYB[12][15] ), .SUM(
        \r60/SUMB[12][15] ) );
  FADDER \r60/S2_12_14  ( .CIN(\r60/ab[12][14] ), .IN0(\r60/CARRYB[11][14] ), 
        .IN1(\r60/SUMB[11][15] ), .COUT(\r60/CARRYB[12][14] ), .SUM(
        \r60/SUMB[12][14] ) );
  FADDER \r60/S2_12_13  ( .CIN(\r60/ab[12][13] ), .IN0(\r60/CARRYB[11][13] ), 
        .IN1(\r60/SUMB[11][14] ), .COUT(\r60/CARRYB[12][13] ), .SUM(
        \r60/SUMB[12][13] ) );
  FADDER \r60/S2_12_12  ( .CIN(\r60/ab[12][12] ), .IN0(\r60/CARRYB[11][12] ), 
        .IN1(\r60/SUMB[11][13] ), .COUT(\r60/CARRYB[12][12] ), .SUM(
        \r60/SUMB[12][12] ) );
  FADDER \r60/S2_12_11  ( .CIN(\r60/ab[12][11] ), .IN0(\r60/CARRYB[11][11] ), 
        .IN1(\r60/SUMB[11][12] ), .COUT(\r60/CARRYB[12][11] ), .SUM(
        \r60/SUMB[12][11] ) );
  FADDER \r60/S2_12_10  ( .CIN(\r60/ab[12][10] ), .IN0(\r60/CARRYB[11][10] ), 
        .IN1(\r60/SUMB[11][11] ), .COUT(\r60/CARRYB[12][10] ), .SUM(
        \r60/SUMB[12][10] ) );
  FADDER \r60/S2_12_9  ( .CIN(\r60/ab[12][9] ), .IN0(\r60/CARRYB[11][9] ), 
        .IN1(\r60/SUMB[11][10] ), .COUT(\r60/CARRYB[12][9] ), .SUM(
        \r60/SUMB[12][9] ) );
  FADDER \r60/S2_12_8  ( .CIN(\r60/ab[12][8] ), .IN0(\r60/CARRYB[11][8] ), 
        .IN1(\r60/SUMB[11][9] ), .COUT(\r60/CARRYB[12][8] ), .SUM(
        \r60/SUMB[12][8] ) );
  FADDER \r60/S2_12_7  ( .CIN(\r60/ab[12][7] ), .IN0(\r60/CARRYB[11][7] ), 
        .IN1(\r60/SUMB[11][8] ), .COUT(\r60/CARRYB[12][7] ), .SUM(
        \r60/SUMB[12][7] ) );
  FADDER \r60/S2_12_6  ( .CIN(\r60/ab[12][6] ), .IN0(\r60/CARRYB[11][6] ), 
        .IN1(\r60/SUMB[11][7] ), .COUT(\r60/CARRYB[12][6] ), .SUM(
        \r60/SUMB[12][6] ) );
  FADDER \r60/S2_12_5  ( .CIN(\r60/ab[12][5] ), .IN0(\r60/CARRYB[11][5] ), 
        .IN1(\r60/SUMB[11][6] ), .COUT(\r60/CARRYB[12][5] ), .SUM(
        \r60/SUMB[12][5] ) );
  FADDER \r60/S2_12_4  ( .CIN(\r60/ab[12][4] ), .IN0(\r60/CARRYB[11][4] ), 
        .IN1(\r60/SUMB[11][5] ), .COUT(\r60/CARRYB[12][4] ), .SUM(
        \r60/SUMB[12][4] ) );
  FADDER \r60/S2_12_3  ( .CIN(\r60/ab[12][3] ), .IN0(\r60/CARRYB[11][3] ), 
        .IN1(\r60/SUMB[11][4] ), .COUT(\r60/CARRYB[12][3] ), .SUM(
        \r60/SUMB[12][3] ) );
  FADDER \r60/S2_12_2  ( .CIN(\r60/ab[12][2] ), .IN0(\r60/CARRYB[11][2] ), 
        .IN1(\r60/SUMB[11][3] ), .COUT(\r60/CARRYB[12][2] ), .SUM(
        \r60/SUMB[12][2] ) );
  FADDER \r60/S2_12_1  ( .CIN(\r60/ab[12][1] ), .IN0(\r60/CARRYB[11][1] ), 
        .IN1(\r60/SUMB[11][2] ), .COUT(\r60/CARRYB[12][1] ), .SUM(
        \r60/SUMB[12][1] ) );
  FADDER \r60/S1_12_0  ( .CIN(\r60/ab[12][0] ), .IN0(\r60/CARRYB[11][0] ), 
        .IN1(\r60/SUMB[11][1] ), .COUT(\r60/CARRYB[12][0] ), .SUM(N129) );
  FADDER \r60/S3_13_30  ( .CIN(\r60/ab[13][30] ), .IN0(\r60/CARRYB[12][30] ), 
        .IN1(\r60/ab[12][31] ), .COUT(\r60/CARRYB[13][30] ), .SUM(
        \r60/SUMB[13][30] ) );
  FADDER \r60/S2_13_29  ( .CIN(\r60/ab[13][29] ), .IN0(\r60/CARRYB[12][29] ), 
        .IN1(\r60/SUMB[12][30] ), .COUT(\r60/CARRYB[13][29] ), .SUM(
        \r60/SUMB[13][29] ) );
  FADDER \r60/S2_13_28  ( .CIN(\r60/ab[13][28] ), .IN0(\r60/CARRYB[12][28] ), 
        .IN1(\r60/SUMB[12][29] ), .COUT(\r60/CARRYB[13][28] ), .SUM(
        \r60/SUMB[13][28] ) );
  FADDER \r60/S2_13_27  ( .CIN(\r60/ab[13][27] ), .IN0(\r60/CARRYB[12][27] ), 
        .IN1(\r60/SUMB[12][28] ), .COUT(\r60/CARRYB[13][27] ), .SUM(
        \r60/SUMB[13][27] ) );
  FADDER \r60/S2_13_26  ( .CIN(\r60/ab[13][26] ), .IN0(\r60/CARRYB[12][26] ), 
        .IN1(\r60/SUMB[12][27] ), .COUT(\r60/CARRYB[13][26] ), .SUM(
        \r60/SUMB[13][26] ) );
  FADDER \r60/S2_13_25  ( .CIN(\r60/ab[13][25] ), .IN0(\r60/CARRYB[12][25] ), 
        .IN1(\r60/SUMB[12][26] ), .COUT(\r60/CARRYB[13][25] ), .SUM(
        \r60/SUMB[13][25] ) );
  FADDER \r60/S2_13_24  ( .CIN(\r60/ab[13][24] ), .IN0(\r60/CARRYB[12][24] ), 
        .IN1(\r60/SUMB[12][25] ), .COUT(\r60/CARRYB[13][24] ), .SUM(
        \r60/SUMB[13][24] ) );
  FADDER \r60/S2_13_23  ( .CIN(\r60/ab[13][23] ), .IN0(\r60/CARRYB[12][23] ), 
        .IN1(\r60/SUMB[12][24] ), .COUT(\r60/CARRYB[13][23] ), .SUM(
        \r60/SUMB[13][23] ) );
  FADDER \r60/S2_13_22  ( .CIN(\r60/ab[13][22] ), .IN0(\r60/CARRYB[12][22] ), 
        .IN1(\r60/SUMB[12][23] ), .COUT(\r60/CARRYB[13][22] ), .SUM(
        \r60/SUMB[13][22] ) );
  FADDER \r60/S2_13_21  ( .CIN(\r60/ab[13][21] ), .IN0(\r60/CARRYB[12][21] ), 
        .IN1(\r60/SUMB[12][22] ), .COUT(\r60/CARRYB[13][21] ), .SUM(
        \r60/SUMB[13][21] ) );
  FADDER \r60/S2_13_20  ( .CIN(\r60/ab[13][20] ), .IN0(\r60/CARRYB[12][20] ), 
        .IN1(\r60/SUMB[12][21] ), .COUT(\r60/CARRYB[13][20] ), .SUM(
        \r60/SUMB[13][20] ) );
  FADDER \r60/S2_13_19  ( .CIN(\r60/ab[13][19] ), .IN0(\r60/CARRYB[12][19] ), 
        .IN1(\r60/SUMB[12][20] ), .COUT(\r60/CARRYB[13][19] ), .SUM(
        \r60/SUMB[13][19] ) );
  FADDER \r60/S2_13_18  ( .CIN(\r60/ab[13][18] ), .IN0(\r60/CARRYB[12][18] ), 
        .IN1(\r60/SUMB[12][19] ), .COUT(\r60/CARRYB[13][18] ), .SUM(
        \r60/SUMB[13][18] ) );
  FADDER \r60/S2_13_17  ( .CIN(\r60/ab[13][17] ), .IN0(\r60/CARRYB[12][17] ), 
        .IN1(\r60/SUMB[12][18] ), .COUT(\r60/CARRYB[13][17] ), .SUM(
        \r60/SUMB[13][17] ) );
  FADDER \r60/S2_13_16  ( .CIN(\r60/ab[13][16] ), .IN0(\r60/CARRYB[12][16] ), 
        .IN1(\r60/SUMB[12][17] ), .COUT(\r60/CARRYB[13][16] ), .SUM(
        \r60/SUMB[13][16] ) );
  FADDER \r60/S2_13_15  ( .CIN(\r60/ab[13][15] ), .IN0(\r60/CARRYB[12][15] ), 
        .IN1(\r60/SUMB[12][16] ), .COUT(\r60/CARRYB[13][15] ), .SUM(
        \r60/SUMB[13][15] ) );
  FADDER \r60/S2_13_14  ( .CIN(\r60/ab[13][14] ), .IN0(\r60/CARRYB[12][14] ), 
        .IN1(\r60/SUMB[12][15] ), .COUT(\r60/CARRYB[13][14] ), .SUM(
        \r60/SUMB[13][14] ) );
  FADDER \r60/S2_13_13  ( .CIN(\r60/ab[13][13] ), .IN0(\r60/CARRYB[12][13] ), 
        .IN1(\r60/SUMB[12][14] ), .COUT(\r60/CARRYB[13][13] ), .SUM(
        \r60/SUMB[13][13] ) );
  FADDER \r60/S2_13_12  ( .CIN(\r60/ab[13][12] ), .IN0(\r60/CARRYB[12][12] ), 
        .IN1(\r60/SUMB[12][13] ), .COUT(\r60/CARRYB[13][12] ), .SUM(
        \r60/SUMB[13][12] ) );
  FADDER \r60/S2_13_11  ( .CIN(\r60/ab[13][11] ), .IN0(\r60/CARRYB[12][11] ), 
        .IN1(\r60/SUMB[12][12] ), .COUT(\r60/CARRYB[13][11] ), .SUM(
        \r60/SUMB[13][11] ) );
  FADDER \r60/S2_13_10  ( .CIN(\r60/ab[13][10] ), .IN0(\r60/CARRYB[12][10] ), 
        .IN1(\r60/SUMB[12][11] ), .COUT(\r60/CARRYB[13][10] ), .SUM(
        \r60/SUMB[13][10] ) );
  FADDER \r60/S2_13_9  ( .CIN(\r60/ab[13][9] ), .IN0(\r60/CARRYB[12][9] ), 
        .IN1(\r60/SUMB[12][10] ), .COUT(\r60/CARRYB[13][9] ), .SUM(
        \r60/SUMB[13][9] ) );
  FADDER \r60/S2_13_8  ( .CIN(\r60/ab[13][8] ), .IN0(\r60/CARRYB[12][8] ), 
        .IN1(\r60/SUMB[12][9] ), .COUT(\r60/CARRYB[13][8] ), .SUM(
        \r60/SUMB[13][8] ) );
  FADDER \r60/S2_13_7  ( .CIN(\r60/ab[13][7] ), .IN0(\r60/CARRYB[12][7] ), 
        .IN1(\r60/SUMB[12][8] ), .COUT(\r60/CARRYB[13][7] ), .SUM(
        \r60/SUMB[13][7] ) );
  FADDER \r60/S2_13_6  ( .CIN(\r60/ab[13][6] ), .IN0(\r60/CARRYB[12][6] ), 
        .IN1(\r60/SUMB[12][7] ), .COUT(\r60/CARRYB[13][6] ), .SUM(
        \r60/SUMB[13][6] ) );
  FADDER \r60/S2_13_5  ( .CIN(\r60/ab[13][5] ), .IN0(\r60/CARRYB[12][5] ), 
        .IN1(\r60/SUMB[12][6] ), .COUT(\r60/CARRYB[13][5] ), .SUM(
        \r60/SUMB[13][5] ) );
  FADDER \r60/S2_13_4  ( .CIN(\r60/ab[13][4] ), .IN0(\r60/CARRYB[12][4] ), 
        .IN1(\r60/SUMB[12][5] ), .COUT(\r60/CARRYB[13][4] ), .SUM(
        \r60/SUMB[13][4] ) );
  FADDER \r60/S2_13_3  ( .CIN(\r60/ab[13][3] ), .IN0(\r60/CARRYB[12][3] ), 
        .IN1(\r60/SUMB[12][4] ), .COUT(\r60/CARRYB[13][3] ), .SUM(
        \r60/SUMB[13][3] ) );
  FADDER \r60/S2_13_2  ( .CIN(\r60/ab[13][2] ), .IN0(\r60/CARRYB[12][2] ), 
        .IN1(\r60/SUMB[12][3] ), .COUT(\r60/CARRYB[13][2] ), .SUM(
        \r60/SUMB[13][2] ) );
  FADDER \r60/S2_13_1  ( .CIN(\r60/ab[13][1] ), .IN0(\r60/CARRYB[12][1] ), 
        .IN1(\r60/SUMB[12][2] ), .COUT(\r60/CARRYB[13][1] ), .SUM(
        \r60/SUMB[13][1] ) );
  FADDER \r60/S1_13_0  ( .CIN(\r60/ab[13][0] ), .IN0(\r60/CARRYB[12][0] ), 
        .IN1(\r60/SUMB[12][1] ), .COUT(\r60/CARRYB[13][0] ), .SUM(N130) );
  FADDER \r60/S3_14_30  ( .CIN(\r60/ab[14][30] ), .IN0(\r60/CARRYB[13][30] ), 
        .IN1(\r60/ab[13][31] ), .COUT(\r60/CARRYB[14][30] ), .SUM(
        \r60/SUMB[14][30] ) );
  FADDER \r60/S2_14_29  ( .CIN(\r60/ab[14][29] ), .IN0(\r60/CARRYB[13][29] ), 
        .IN1(\r60/SUMB[13][30] ), .COUT(\r60/CARRYB[14][29] ), .SUM(
        \r60/SUMB[14][29] ) );
  FADDER \r60/S2_14_28  ( .CIN(\r60/ab[14][28] ), .IN0(\r60/CARRYB[13][28] ), 
        .IN1(\r60/SUMB[13][29] ), .COUT(\r60/CARRYB[14][28] ), .SUM(
        \r60/SUMB[14][28] ) );
  FADDER \r60/S2_14_27  ( .CIN(\r60/ab[14][27] ), .IN0(\r60/CARRYB[13][27] ), 
        .IN1(\r60/SUMB[13][28] ), .COUT(\r60/CARRYB[14][27] ), .SUM(
        \r60/SUMB[14][27] ) );
  FADDER \r60/S2_14_26  ( .CIN(\r60/ab[14][26] ), .IN0(\r60/CARRYB[13][26] ), 
        .IN1(\r60/SUMB[13][27] ), .COUT(\r60/CARRYB[14][26] ), .SUM(
        \r60/SUMB[14][26] ) );
  FADDER \r60/S2_14_25  ( .CIN(\r60/ab[14][25] ), .IN0(\r60/CARRYB[13][25] ), 
        .IN1(\r60/SUMB[13][26] ), .COUT(\r60/CARRYB[14][25] ), .SUM(
        \r60/SUMB[14][25] ) );
  FADDER \r60/S2_14_24  ( .CIN(\r60/ab[14][24] ), .IN0(\r60/CARRYB[13][24] ), 
        .IN1(\r60/SUMB[13][25] ), .COUT(\r60/CARRYB[14][24] ), .SUM(
        \r60/SUMB[14][24] ) );
  FADDER \r60/S2_14_23  ( .CIN(\r60/ab[14][23] ), .IN0(\r60/CARRYB[13][23] ), 
        .IN1(\r60/SUMB[13][24] ), .COUT(\r60/CARRYB[14][23] ), .SUM(
        \r60/SUMB[14][23] ) );
  FADDER \r60/S2_14_22  ( .CIN(\r60/ab[14][22] ), .IN0(\r60/CARRYB[13][22] ), 
        .IN1(\r60/SUMB[13][23] ), .COUT(\r60/CARRYB[14][22] ), .SUM(
        \r60/SUMB[14][22] ) );
  FADDER \r60/S2_14_21  ( .CIN(\r60/ab[14][21] ), .IN0(\r60/CARRYB[13][21] ), 
        .IN1(\r60/SUMB[13][22] ), .COUT(\r60/CARRYB[14][21] ), .SUM(
        \r60/SUMB[14][21] ) );
  FADDER \r60/S2_14_20  ( .CIN(\r60/ab[14][20] ), .IN0(\r60/CARRYB[13][20] ), 
        .IN1(\r60/SUMB[13][21] ), .COUT(\r60/CARRYB[14][20] ), .SUM(
        \r60/SUMB[14][20] ) );
  FADDER \r60/S2_14_19  ( .CIN(\r60/ab[14][19] ), .IN0(\r60/CARRYB[13][19] ), 
        .IN1(\r60/SUMB[13][20] ), .COUT(\r60/CARRYB[14][19] ), .SUM(
        \r60/SUMB[14][19] ) );
  FADDER \r60/S2_14_18  ( .CIN(\r60/ab[14][18] ), .IN0(\r60/CARRYB[13][18] ), 
        .IN1(\r60/SUMB[13][19] ), .COUT(\r60/CARRYB[14][18] ), .SUM(
        \r60/SUMB[14][18] ) );
  FADDER \r60/S2_14_17  ( .CIN(\r60/ab[14][17] ), .IN0(\r60/CARRYB[13][17] ), 
        .IN1(\r60/SUMB[13][18] ), .COUT(\r60/CARRYB[14][17] ), .SUM(
        \r60/SUMB[14][17] ) );
  FADDER \r60/S2_14_16  ( .CIN(\r60/ab[14][16] ), .IN0(\r60/CARRYB[13][16] ), 
        .IN1(\r60/SUMB[13][17] ), .COUT(\r60/CARRYB[14][16] ), .SUM(
        \r60/SUMB[14][16] ) );
  FADDER \r60/S2_14_15  ( .CIN(\r60/ab[14][15] ), .IN0(\r60/CARRYB[13][15] ), 
        .IN1(\r60/SUMB[13][16] ), .COUT(\r60/CARRYB[14][15] ), .SUM(
        \r60/SUMB[14][15] ) );
  FADDER \r60/S2_14_14  ( .CIN(\r60/ab[14][14] ), .IN0(\r60/CARRYB[13][14] ), 
        .IN1(\r60/SUMB[13][15] ), .COUT(\r60/CARRYB[14][14] ), .SUM(
        \r60/SUMB[14][14] ) );
  FADDER \r60/S2_14_13  ( .CIN(\r60/ab[14][13] ), .IN0(\r60/CARRYB[13][13] ), 
        .IN1(\r60/SUMB[13][14] ), .COUT(\r60/CARRYB[14][13] ), .SUM(
        \r60/SUMB[14][13] ) );
  FADDER \r60/S2_14_12  ( .CIN(\r60/ab[14][12] ), .IN0(\r60/CARRYB[13][12] ), 
        .IN1(\r60/SUMB[13][13] ), .COUT(\r60/CARRYB[14][12] ), .SUM(
        \r60/SUMB[14][12] ) );
  FADDER \r60/S2_14_11  ( .CIN(\r60/ab[14][11] ), .IN0(\r60/CARRYB[13][11] ), 
        .IN1(\r60/SUMB[13][12] ), .COUT(\r60/CARRYB[14][11] ), .SUM(
        \r60/SUMB[14][11] ) );
  FADDER \r60/S2_14_10  ( .CIN(\r60/ab[14][10] ), .IN0(\r60/CARRYB[13][10] ), 
        .IN1(\r60/SUMB[13][11] ), .COUT(\r60/CARRYB[14][10] ), .SUM(
        \r60/SUMB[14][10] ) );
  FADDER \r60/S2_14_9  ( .CIN(\r60/ab[14][9] ), .IN0(\r60/CARRYB[13][9] ), 
        .IN1(\r60/SUMB[13][10] ), .COUT(\r60/CARRYB[14][9] ), .SUM(
        \r60/SUMB[14][9] ) );
  FADDER \r60/S2_14_8  ( .CIN(\r60/ab[14][8] ), .IN0(\r60/CARRYB[13][8] ), 
        .IN1(\r60/SUMB[13][9] ), .COUT(\r60/CARRYB[14][8] ), .SUM(
        \r60/SUMB[14][8] ) );
  FADDER \r60/S2_14_7  ( .CIN(\r60/ab[14][7] ), .IN0(\r60/CARRYB[13][7] ), 
        .IN1(\r60/SUMB[13][8] ), .COUT(\r60/CARRYB[14][7] ), .SUM(
        \r60/SUMB[14][7] ) );
  FADDER \r60/S2_14_6  ( .CIN(\r60/ab[14][6] ), .IN0(\r60/CARRYB[13][6] ), 
        .IN1(\r60/SUMB[13][7] ), .COUT(\r60/CARRYB[14][6] ), .SUM(
        \r60/SUMB[14][6] ) );
  FADDER \r60/S2_14_5  ( .CIN(\r60/ab[14][5] ), .IN0(\r60/CARRYB[13][5] ), 
        .IN1(\r60/SUMB[13][6] ), .COUT(\r60/CARRYB[14][5] ), .SUM(
        \r60/SUMB[14][5] ) );
  FADDER \r60/S2_14_4  ( .CIN(\r60/ab[14][4] ), .IN0(\r60/CARRYB[13][4] ), 
        .IN1(\r60/SUMB[13][5] ), .COUT(\r60/CARRYB[14][4] ), .SUM(
        \r60/SUMB[14][4] ) );
  FADDER \r60/S2_14_3  ( .CIN(\r60/ab[14][3] ), .IN0(\r60/CARRYB[13][3] ), 
        .IN1(\r60/SUMB[13][4] ), .COUT(\r60/CARRYB[14][3] ), .SUM(
        \r60/SUMB[14][3] ) );
  FADDER \r60/S2_14_2  ( .CIN(\r60/ab[14][2] ), .IN0(\r60/CARRYB[13][2] ), 
        .IN1(\r60/SUMB[13][3] ), .COUT(\r60/CARRYB[14][2] ), .SUM(
        \r60/SUMB[14][2] ) );
  FADDER \r60/S2_14_1  ( .CIN(\r60/ab[14][1] ), .IN0(\r60/CARRYB[13][1] ), 
        .IN1(\r60/SUMB[13][2] ), .COUT(\r60/CARRYB[14][1] ), .SUM(
        \r60/SUMB[14][1] ) );
  FADDER \r60/S1_14_0  ( .CIN(\r60/ab[14][0] ), .IN0(\r60/CARRYB[13][0] ), 
        .IN1(\r60/SUMB[13][1] ), .COUT(\r60/CARRYB[14][0] ), .SUM(N131) );
  FADDER \r60/S3_15_30  ( .CIN(\r60/ab[15][30] ), .IN0(\r60/CARRYB[14][30] ), 
        .IN1(\r60/ab[14][31] ), .COUT(\r60/CARRYB[15][30] ), .SUM(
        \r60/SUMB[15][30] ) );
  FADDER \r60/S2_15_29  ( .CIN(\r60/ab[15][29] ), .IN0(\r60/CARRYB[14][29] ), 
        .IN1(\r60/SUMB[14][30] ), .COUT(\r60/CARRYB[15][29] ), .SUM(
        \r60/SUMB[15][29] ) );
  FADDER \r60/S2_15_28  ( .CIN(\r60/ab[15][28] ), .IN0(\r60/CARRYB[14][28] ), 
        .IN1(\r60/SUMB[14][29] ), .COUT(\r60/CARRYB[15][28] ), .SUM(
        \r60/SUMB[15][28] ) );
  FADDER \r60/S2_15_27  ( .CIN(\r60/ab[15][27] ), .IN0(\r60/CARRYB[14][27] ), 
        .IN1(\r60/SUMB[14][28] ), .COUT(\r60/CARRYB[15][27] ), .SUM(
        \r60/SUMB[15][27] ) );
  FADDER \r60/S2_15_26  ( .CIN(\r60/ab[15][26] ), .IN0(\r60/CARRYB[14][26] ), 
        .IN1(\r60/SUMB[14][27] ), .COUT(\r60/CARRYB[15][26] ), .SUM(
        \r60/SUMB[15][26] ) );
  FADDER \r60/S2_15_25  ( .CIN(\r60/ab[15][25] ), .IN0(\r60/CARRYB[14][25] ), 
        .IN1(\r60/SUMB[14][26] ), .COUT(\r60/CARRYB[15][25] ), .SUM(
        \r60/SUMB[15][25] ) );
  FADDER \r60/S2_15_24  ( .CIN(\r60/ab[15][24] ), .IN0(\r60/CARRYB[14][24] ), 
        .IN1(\r60/SUMB[14][25] ), .COUT(\r60/CARRYB[15][24] ), .SUM(
        \r60/SUMB[15][24] ) );
  FADDER \r60/S2_15_23  ( .CIN(\r60/ab[15][23] ), .IN0(\r60/CARRYB[14][23] ), 
        .IN1(\r60/SUMB[14][24] ), .COUT(\r60/CARRYB[15][23] ), .SUM(
        \r60/SUMB[15][23] ) );
  FADDER \r60/S2_15_22  ( .CIN(\r60/ab[15][22] ), .IN0(\r60/CARRYB[14][22] ), 
        .IN1(\r60/SUMB[14][23] ), .COUT(\r60/CARRYB[15][22] ), .SUM(
        \r60/SUMB[15][22] ) );
  FADDER \r60/S2_15_21  ( .CIN(\r60/ab[15][21] ), .IN0(\r60/CARRYB[14][21] ), 
        .IN1(\r60/SUMB[14][22] ), .COUT(\r60/CARRYB[15][21] ), .SUM(
        \r60/SUMB[15][21] ) );
  FADDER \r60/S2_15_20  ( .CIN(\r60/ab[15][20] ), .IN0(\r60/CARRYB[14][20] ), 
        .IN1(\r60/SUMB[14][21] ), .COUT(\r60/CARRYB[15][20] ), .SUM(
        \r60/SUMB[15][20] ) );
  FADDER \r60/S2_15_19  ( .CIN(\r60/ab[15][19] ), .IN0(\r60/CARRYB[14][19] ), 
        .IN1(\r60/SUMB[14][20] ), .COUT(\r60/CARRYB[15][19] ), .SUM(
        \r60/SUMB[15][19] ) );
  FADDER \r60/S2_15_18  ( .CIN(\r60/ab[15][18] ), .IN0(\r60/CARRYB[14][18] ), 
        .IN1(\r60/SUMB[14][19] ), .COUT(\r60/CARRYB[15][18] ), .SUM(
        \r60/SUMB[15][18] ) );
  FADDER \r60/S2_15_17  ( .CIN(\r60/ab[15][17] ), .IN0(\r60/CARRYB[14][17] ), 
        .IN1(\r60/SUMB[14][18] ), .COUT(\r60/CARRYB[15][17] ), .SUM(
        \r60/SUMB[15][17] ) );
  FADDER \r60/S2_15_16  ( .CIN(\r60/ab[15][16] ), .IN0(\r60/CARRYB[14][16] ), 
        .IN1(\r60/SUMB[14][17] ), .COUT(\r60/CARRYB[15][16] ), .SUM(
        \r60/SUMB[15][16] ) );
  FADDER \r60/S2_15_15  ( .CIN(\r60/ab[15][15] ), .IN0(\r60/CARRYB[14][15] ), 
        .IN1(\r60/SUMB[14][16] ), .COUT(\r60/CARRYB[15][15] ), .SUM(
        \r60/SUMB[15][15] ) );
  FADDER \r60/S2_15_14  ( .CIN(\r60/ab[15][14] ), .IN0(\r60/CARRYB[14][14] ), 
        .IN1(\r60/SUMB[14][15] ), .COUT(\r60/CARRYB[15][14] ), .SUM(
        \r60/SUMB[15][14] ) );
  FADDER \r60/S2_15_13  ( .CIN(\r60/ab[15][13] ), .IN0(\r60/CARRYB[14][13] ), 
        .IN1(\r60/SUMB[14][14] ), .COUT(\r60/CARRYB[15][13] ), .SUM(
        \r60/SUMB[15][13] ) );
  FADDER \r60/S2_15_12  ( .CIN(\r60/ab[15][12] ), .IN0(\r60/CARRYB[14][12] ), 
        .IN1(\r60/SUMB[14][13] ), .COUT(\r60/CARRYB[15][12] ), .SUM(
        \r60/SUMB[15][12] ) );
  FADDER \r60/S2_15_11  ( .CIN(\r60/ab[15][11] ), .IN0(\r60/CARRYB[14][11] ), 
        .IN1(\r60/SUMB[14][12] ), .COUT(\r60/CARRYB[15][11] ), .SUM(
        \r60/SUMB[15][11] ) );
  FADDER \r60/S2_15_10  ( .CIN(\r60/ab[15][10] ), .IN0(\r60/CARRYB[14][10] ), 
        .IN1(\r60/SUMB[14][11] ), .COUT(\r60/CARRYB[15][10] ), .SUM(
        \r60/SUMB[15][10] ) );
  FADDER \r60/S2_15_9  ( .CIN(\r60/ab[15][9] ), .IN0(\r60/CARRYB[14][9] ), 
        .IN1(\r60/SUMB[14][10] ), .COUT(\r60/CARRYB[15][9] ), .SUM(
        \r60/SUMB[15][9] ) );
  FADDER \r60/S2_15_8  ( .CIN(\r60/ab[15][8] ), .IN0(\r60/CARRYB[14][8] ), 
        .IN1(\r60/SUMB[14][9] ), .COUT(\r60/CARRYB[15][8] ), .SUM(
        \r60/SUMB[15][8] ) );
  FADDER \r60/S2_15_7  ( .CIN(\r60/ab[15][7] ), .IN0(\r60/CARRYB[14][7] ), 
        .IN1(\r60/SUMB[14][8] ), .COUT(\r60/CARRYB[15][7] ), .SUM(
        \r60/SUMB[15][7] ) );
  FADDER \r60/S2_15_6  ( .CIN(\r60/ab[15][6] ), .IN0(\r60/CARRYB[14][6] ), 
        .IN1(\r60/SUMB[14][7] ), .COUT(\r60/CARRYB[15][6] ), .SUM(
        \r60/SUMB[15][6] ) );
  FADDER \r60/S2_15_5  ( .CIN(\r60/ab[15][5] ), .IN0(\r60/CARRYB[14][5] ), 
        .IN1(\r60/SUMB[14][6] ), .COUT(\r60/CARRYB[15][5] ), .SUM(
        \r60/SUMB[15][5] ) );
  FADDER \r60/S2_15_4  ( .CIN(\r60/ab[15][4] ), .IN0(\r60/CARRYB[14][4] ), 
        .IN1(\r60/SUMB[14][5] ), .COUT(\r60/CARRYB[15][4] ), .SUM(
        \r60/SUMB[15][4] ) );
  FADDER \r60/S2_15_3  ( .CIN(\r60/ab[15][3] ), .IN0(\r60/CARRYB[14][3] ), 
        .IN1(\r60/SUMB[14][4] ), .COUT(\r60/CARRYB[15][3] ), .SUM(
        \r60/SUMB[15][3] ) );
  FADDER \r60/S2_15_2  ( .CIN(\r60/ab[15][2] ), .IN0(\r60/CARRYB[14][2] ), 
        .IN1(\r60/SUMB[14][3] ), .COUT(\r60/CARRYB[15][2] ), .SUM(
        \r60/SUMB[15][2] ) );
  FADDER \r60/S2_15_1  ( .CIN(\r60/ab[15][1] ), .IN0(\r60/CARRYB[14][1] ), 
        .IN1(\r60/SUMB[14][2] ), .COUT(\r60/CARRYB[15][1] ), .SUM(
        \r60/SUMB[15][1] ) );
  FADDER \r60/S1_15_0  ( .CIN(\r60/ab[15][0] ), .IN0(\r60/CARRYB[14][0] ), 
        .IN1(\r60/SUMB[14][1] ), .COUT(\r60/CARRYB[15][0] ), .SUM(N132) );
  FADDER \r60/S3_16_30  ( .CIN(\r60/ab[16][30] ), .IN0(\r60/CARRYB[15][30] ), 
        .IN1(\r60/ab[15][31] ), .COUT(\r60/CARRYB[16][30] ), .SUM(
        \r60/SUMB[16][30] ) );
  FADDER \r60/S2_16_29  ( .CIN(\r60/ab[16][29] ), .IN0(\r60/CARRYB[15][29] ), 
        .IN1(\r60/SUMB[15][30] ), .COUT(\r60/CARRYB[16][29] ), .SUM(
        \r60/SUMB[16][29] ) );
  FADDER \r60/S2_16_28  ( .CIN(\r60/ab[16][28] ), .IN0(\r60/CARRYB[15][28] ), 
        .IN1(\r60/SUMB[15][29] ), .COUT(\r60/CARRYB[16][28] ), .SUM(
        \r60/SUMB[16][28] ) );
  FADDER \r60/S2_16_27  ( .CIN(\r60/ab[16][27] ), .IN0(\r60/CARRYB[15][27] ), 
        .IN1(\r60/SUMB[15][28] ), .COUT(\r60/CARRYB[16][27] ), .SUM(
        \r60/SUMB[16][27] ) );
  FADDER \r60/S2_16_26  ( .CIN(\r60/ab[16][26] ), .IN0(\r60/CARRYB[15][26] ), 
        .IN1(\r60/SUMB[15][27] ), .COUT(\r60/CARRYB[16][26] ), .SUM(
        \r60/SUMB[16][26] ) );
  FADDER \r60/S2_16_25  ( .CIN(\r60/ab[16][25] ), .IN0(\r60/CARRYB[15][25] ), 
        .IN1(\r60/SUMB[15][26] ), .COUT(\r60/CARRYB[16][25] ), .SUM(
        \r60/SUMB[16][25] ) );
  FADDER \r60/S2_16_24  ( .CIN(\r60/ab[16][24] ), .IN0(\r60/CARRYB[15][24] ), 
        .IN1(\r60/SUMB[15][25] ), .COUT(\r60/CARRYB[16][24] ), .SUM(
        \r60/SUMB[16][24] ) );
  FADDER \r60/S2_16_23  ( .CIN(\r60/ab[16][23] ), .IN0(\r60/CARRYB[15][23] ), 
        .IN1(\r60/SUMB[15][24] ), .COUT(\r60/CARRYB[16][23] ), .SUM(
        \r60/SUMB[16][23] ) );
  FADDER \r60/S2_16_22  ( .CIN(\r60/ab[16][22] ), .IN0(\r60/CARRYB[15][22] ), 
        .IN1(\r60/SUMB[15][23] ), .COUT(\r60/CARRYB[16][22] ), .SUM(
        \r60/SUMB[16][22] ) );
  FADDER \r60/S2_16_21  ( .CIN(\r60/ab[16][21] ), .IN0(\r60/CARRYB[15][21] ), 
        .IN1(\r60/SUMB[15][22] ), .COUT(\r60/CARRYB[16][21] ), .SUM(
        \r60/SUMB[16][21] ) );
  FADDER \r60/S2_16_20  ( .CIN(\r60/ab[16][20] ), .IN0(\r60/CARRYB[15][20] ), 
        .IN1(\r60/SUMB[15][21] ), .COUT(\r60/CARRYB[16][20] ), .SUM(
        \r60/SUMB[16][20] ) );
  FADDER \r60/S2_16_19  ( .CIN(\r60/ab[16][19] ), .IN0(\r60/CARRYB[15][19] ), 
        .IN1(\r60/SUMB[15][20] ), .COUT(\r60/CARRYB[16][19] ), .SUM(
        \r60/SUMB[16][19] ) );
  FADDER \r60/S2_16_18  ( .CIN(\r60/ab[16][18] ), .IN0(\r60/CARRYB[15][18] ), 
        .IN1(\r60/SUMB[15][19] ), .COUT(\r60/CARRYB[16][18] ), .SUM(
        \r60/SUMB[16][18] ) );
  FADDER \r60/S2_16_17  ( .CIN(\r60/ab[16][17] ), .IN0(\r60/CARRYB[15][17] ), 
        .IN1(\r60/SUMB[15][18] ), .COUT(\r60/CARRYB[16][17] ), .SUM(
        \r60/SUMB[16][17] ) );
  FADDER \r60/S2_16_16  ( .CIN(\r60/ab[16][16] ), .IN0(\r60/CARRYB[15][16] ), 
        .IN1(\r60/SUMB[15][17] ), .COUT(\r60/CARRYB[16][16] ), .SUM(
        \r60/SUMB[16][16] ) );
  FADDER \r60/S2_16_15  ( .CIN(\r60/ab[16][15] ), .IN0(\r60/CARRYB[15][15] ), 
        .IN1(\r60/SUMB[15][16] ), .COUT(\r60/CARRYB[16][15] ), .SUM(
        \r60/SUMB[16][15] ) );
  FADDER \r60/S2_16_14  ( .CIN(\r60/ab[16][14] ), .IN0(\r60/CARRYB[15][14] ), 
        .IN1(\r60/SUMB[15][15] ), .COUT(\r60/CARRYB[16][14] ), .SUM(
        \r60/SUMB[16][14] ) );
  FADDER \r60/S2_16_13  ( .CIN(\r60/ab[16][13] ), .IN0(\r60/CARRYB[15][13] ), 
        .IN1(\r60/SUMB[15][14] ), .COUT(\r60/CARRYB[16][13] ), .SUM(
        \r60/SUMB[16][13] ) );
  FADDER \r60/S2_16_12  ( .CIN(\r60/ab[16][12] ), .IN0(\r60/CARRYB[15][12] ), 
        .IN1(\r60/SUMB[15][13] ), .COUT(\r60/CARRYB[16][12] ), .SUM(
        \r60/SUMB[16][12] ) );
  FADDER \r60/S2_16_11  ( .CIN(\r60/ab[16][11] ), .IN0(\r60/CARRYB[15][11] ), 
        .IN1(\r60/SUMB[15][12] ), .COUT(\r60/CARRYB[16][11] ), .SUM(
        \r60/SUMB[16][11] ) );
  FADDER \r60/S2_16_10  ( .CIN(\r60/ab[16][10] ), .IN0(\r60/CARRYB[15][10] ), 
        .IN1(\r60/SUMB[15][11] ), .COUT(\r60/CARRYB[16][10] ), .SUM(
        \r60/SUMB[16][10] ) );
  FADDER \r60/S2_16_9  ( .CIN(\r60/ab[16][9] ), .IN0(\r60/CARRYB[15][9] ), 
        .IN1(\r60/SUMB[15][10] ), .COUT(\r60/CARRYB[16][9] ), .SUM(
        \r60/SUMB[16][9] ) );
  FADDER \r60/S2_16_8  ( .CIN(\r60/ab[16][8] ), .IN0(\r60/CARRYB[15][8] ), 
        .IN1(\r60/SUMB[15][9] ), .COUT(\r60/CARRYB[16][8] ), .SUM(
        \r60/SUMB[16][8] ) );
  FADDER \r60/S2_16_7  ( .CIN(\r60/ab[16][7] ), .IN0(\r60/CARRYB[15][7] ), 
        .IN1(\r60/SUMB[15][8] ), .COUT(\r60/CARRYB[16][7] ), .SUM(
        \r60/SUMB[16][7] ) );
  FADDER \r60/S2_16_6  ( .CIN(\r60/ab[16][6] ), .IN0(\r60/CARRYB[15][6] ), 
        .IN1(\r60/SUMB[15][7] ), .COUT(\r60/CARRYB[16][6] ), .SUM(
        \r60/SUMB[16][6] ) );
  FADDER \r60/S2_16_5  ( .CIN(\r60/ab[16][5] ), .IN0(\r60/CARRYB[15][5] ), 
        .IN1(\r60/SUMB[15][6] ), .COUT(\r60/CARRYB[16][5] ), .SUM(
        \r60/SUMB[16][5] ) );
  FADDER \r60/S2_16_4  ( .CIN(\r60/ab[16][4] ), .IN0(\r60/CARRYB[15][4] ), 
        .IN1(\r60/SUMB[15][5] ), .COUT(\r60/CARRYB[16][4] ), .SUM(
        \r60/SUMB[16][4] ) );
  FADDER \r60/S2_16_3  ( .CIN(\r60/ab[16][3] ), .IN0(\r60/CARRYB[15][3] ), 
        .IN1(\r60/SUMB[15][4] ), .COUT(\r60/CARRYB[16][3] ), .SUM(
        \r60/SUMB[16][3] ) );
  FADDER \r60/S2_16_2  ( .CIN(\r60/ab[16][2] ), .IN0(\r60/CARRYB[15][2] ), 
        .IN1(\r60/SUMB[15][3] ), .COUT(\r60/CARRYB[16][2] ), .SUM(
        \r60/SUMB[16][2] ) );
  FADDER \r60/S2_16_1  ( .CIN(\r60/ab[16][1] ), .IN0(\r60/CARRYB[15][1] ), 
        .IN1(\r60/SUMB[15][2] ), .COUT(\r60/CARRYB[16][1] ), .SUM(
        \r60/SUMB[16][1] ) );
  FADDER \r60/S1_16_0  ( .CIN(\r60/ab[16][0] ), .IN0(\r60/CARRYB[15][0] ), 
        .IN1(\r60/SUMB[15][1] ), .COUT(\r60/CARRYB[16][0] ), .SUM(N133) );
  FADDER \r60/S3_17_30  ( .CIN(\r60/ab[17][30] ), .IN0(\r60/CARRYB[16][30] ), 
        .IN1(\r60/ab[16][31] ), .COUT(\r60/CARRYB[17][30] ), .SUM(
        \r60/SUMB[17][30] ) );
  FADDER \r60/S2_17_29  ( .CIN(\r60/ab[17][29] ), .IN0(\r60/CARRYB[16][29] ), 
        .IN1(\r60/SUMB[16][30] ), .COUT(\r60/CARRYB[17][29] ), .SUM(
        \r60/SUMB[17][29] ) );
  FADDER \r60/S2_17_28  ( .CIN(\r60/ab[17][28] ), .IN0(\r60/CARRYB[16][28] ), 
        .IN1(\r60/SUMB[16][29] ), .COUT(\r60/CARRYB[17][28] ), .SUM(
        \r60/SUMB[17][28] ) );
  FADDER \r60/S2_17_27  ( .CIN(\r60/ab[17][27] ), .IN0(\r60/CARRYB[16][27] ), 
        .IN1(\r60/SUMB[16][28] ), .COUT(\r60/CARRYB[17][27] ), .SUM(
        \r60/SUMB[17][27] ) );
  FADDER \r60/S2_17_26  ( .CIN(\r60/ab[17][26] ), .IN0(\r60/CARRYB[16][26] ), 
        .IN1(\r60/SUMB[16][27] ), .COUT(\r60/CARRYB[17][26] ), .SUM(
        \r60/SUMB[17][26] ) );
  FADDER \r60/S2_17_25  ( .CIN(\r60/ab[17][25] ), .IN0(\r60/CARRYB[16][25] ), 
        .IN1(\r60/SUMB[16][26] ), .COUT(\r60/CARRYB[17][25] ), .SUM(
        \r60/SUMB[17][25] ) );
  FADDER \r60/S2_17_24  ( .CIN(\r60/ab[17][24] ), .IN0(\r60/CARRYB[16][24] ), 
        .IN1(\r60/SUMB[16][25] ), .COUT(\r60/CARRYB[17][24] ), .SUM(
        \r60/SUMB[17][24] ) );
  FADDER \r60/S2_17_23  ( .CIN(\r60/ab[17][23] ), .IN0(\r60/CARRYB[16][23] ), 
        .IN1(\r60/SUMB[16][24] ), .COUT(\r60/CARRYB[17][23] ), .SUM(
        \r60/SUMB[17][23] ) );
  FADDER \r60/S2_17_22  ( .CIN(\r60/ab[17][22] ), .IN0(\r60/CARRYB[16][22] ), 
        .IN1(\r60/SUMB[16][23] ), .COUT(\r60/CARRYB[17][22] ), .SUM(
        \r60/SUMB[17][22] ) );
  FADDER \r60/S2_17_21  ( .CIN(\r60/ab[17][21] ), .IN0(\r60/CARRYB[16][21] ), 
        .IN1(\r60/SUMB[16][22] ), .COUT(\r60/CARRYB[17][21] ), .SUM(
        \r60/SUMB[17][21] ) );
  FADDER \r60/S2_17_20  ( .CIN(\r60/ab[17][20] ), .IN0(\r60/CARRYB[16][20] ), 
        .IN1(\r60/SUMB[16][21] ), .COUT(\r60/CARRYB[17][20] ), .SUM(
        \r60/SUMB[17][20] ) );
  FADDER \r60/S2_17_19  ( .CIN(\r60/ab[17][19] ), .IN0(\r60/CARRYB[16][19] ), 
        .IN1(\r60/SUMB[16][20] ), .COUT(\r60/CARRYB[17][19] ), .SUM(
        \r60/SUMB[17][19] ) );
  FADDER \r60/S2_17_18  ( .CIN(\r60/ab[17][18] ), .IN0(\r60/CARRYB[16][18] ), 
        .IN1(\r60/SUMB[16][19] ), .COUT(\r60/CARRYB[17][18] ), .SUM(
        \r60/SUMB[17][18] ) );
  FADDER \r60/S2_17_17  ( .CIN(\r60/ab[17][17] ), .IN0(\r60/CARRYB[16][17] ), 
        .IN1(\r60/SUMB[16][18] ), .COUT(\r60/CARRYB[17][17] ), .SUM(
        \r60/SUMB[17][17] ) );
  FADDER \r60/S2_17_16  ( .CIN(\r60/ab[17][16] ), .IN0(\r60/CARRYB[16][16] ), 
        .IN1(\r60/SUMB[16][17] ), .COUT(\r60/CARRYB[17][16] ), .SUM(
        \r60/SUMB[17][16] ) );
  FADDER \r60/S2_17_15  ( .CIN(\r60/ab[17][15] ), .IN0(\r60/CARRYB[16][15] ), 
        .IN1(\r60/SUMB[16][16] ), .COUT(\r60/CARRYB[17][15] ), .SUM(
        \r60/SUMB[17][15] ) );
  FADDER \r60/S2_17_14  ( .CIN(\r60/ab[17][14] ), .IN0(\r60/CARRYB[16][14] ), 
        .IN1(\r60/SUMB[16][15] ), .COUT(\r60/CARRYB[17][14] ), .SUM(
        \r60/SUMB[17][14] ) );
  FADDER \r60/S2_17_13  ( .CIN(\r60/ab[17][13] ), .IN0(\r60/CARRYB[16][13] ), 
        .IN1(\r60/SUMB[16][14] ), .COUT(\r60/CARRYB[17][13] ), .SUM(
        \r60/SUMB[17][13] ) );
  FADDER \r60/S2_17_12  ( .CIN(\r60/ab[17][12] ), .IN0(\r60/CARRYB[16][12] ), 
        .IN1(\r60/SUMB[16][13] ), .COUT(\r60/CARRYB[17][12] ), .SUM(
        \r60/SUMB[17][12] ) );
  FADDER \r60/S2_17_11  ( .CIN(\r60/ab[17][11] ), .IN0(\r60/CARRYB[16][11] ), 
        .IN1(\r60/SUMB[16][12] ), .COUT(\r60/CARRYB[17][11] ), .SUM(
        \r60/SUMB[17][11] ) );
  FADDER \r60/S2_17_10  ( .CIN(\r60/ab[17][10] ), .IN0(\r60/CARRYB[16][10] ), 
        .IN1(\r60/SUMB[16][11] ), .COUT(\r60/CARRYB[17][10] ), .SUM(
        \r60/SUMB[17][10] ) );
  FADDER \r60/S2_17_9  ( .CIN(\r60/ab[17][9] ), .IN0(\r60/CARRYB[16][9] ), 
        .IN1(\r60/SUMB[16][10] ), .COUT(\r60/CARRYB[17][9] ), .SUM(
        \r60/SUMB[17][9] ) );
  FADDER \r60/S2_17_8  ( .CIN(\r60/ab[17][8] ), .IN0(\r60/CARRYB[16][8] ), 
        .IN1(\r60/SUMB[16][9] ), .COUT(\r60/CARRYB[17][8] ), .SUM(
        \r60/SUMB[17][8] ) );
  FADDER \r60/S2_17_7  ( .CIN(\r60/ab[17][7] ), .IN0(\r60/CARRYB[16][7] ), 
        .IN1(\r60/SUMB[16][8] ), .COUT(\r60/CARRYB[17][7] ), .SUM(
        \r60/SUMB[17][7] ) );
  FADDER \r60/S2_17_6  ( .CIN(\r60/ab[17][6] ), .IN0(\r60/CARRYB[16][6] ), 
        .IN1(\r60/SUMB[16][7] ), .COUT(\r60/CARRYB[17][6] ), .SUM(
        \r60/SUMB[17][6] ) );
  FADDER \r60/S2_17_5  ( .CIN(\r60/ab[17][5] ), .IN0(\r60/CARRYB[16][5] ), 
        .IN1(\r60/SUMB[16][6] ), .COUT(\r60/CARRYB[17][5] ), .SUM(
        \r60/SUMB[17][5] ) );
  FADDER \r60/S2_17_4  ( .CIN(\r60/ab[17][4] ), .IN0(\r60/CARRYB[16][4] ), 
        .IN1(\r60/SUMB[16][5] ), .COUT(\r60/CARRYB[17][4] ), .SUM(
        \r60/SUMB[17][4] ) );
  FADDER \r60/S2_17_3  ( .CIN(\r60/ab[17][3] ), .IN0(\r60/CARRYB[16][3] ), 
        .IN1(\r60/SUMB[16][4] ), .COUT(\r60/CARRYB[17][3] ), .SUM(
        \r60/SUMB[17][3] ) );
  FADDER \r60/S2_17_2  ( .CIN(\r60/ab[17][2] ), .IN0(\r60/CARRYB[16][2] ), 
        .IN1(\r60/SUMB[16][3] ), .COUT(\r60/CARRYB[17][2] ), .SUM(
        \r60/SUMB[17][2] ) );
  FADDER \r60/S2_17_1  ( .CIN(\r60/ab[17][1] ), .IN0(\r60/CARRYB[16][1] ), 
        .IN1(\r60/SUMB[16][2] ), .COUT(\r60/CARRYB[17][1] ), .SUM(
        \r60/SUMB[17][1] ) );
  FADDER \r60/S1_17_0  ( .CIN(\r60/ab[17][0] ), .IN0(\r60/CARRYB[16][0] ), 
        .IN1(\r60/SUMB[16][1] ), .COUT(\r60/CARRYB[17][0] ), .SUM(N134) );
  FADDER \r60/S3_18_30  ( .CIN(\r60/ab[18][30] ), .IN0(\r60/CARRYB[17][30] ), 
        .IN1(\r60/ab[17][31] ), .COUT(\r60/CARRYB[18][30] ), .SUM(
        \r60/SUMB[18][30] ) );
  FADDER \r60/S2_18_29  ( .CIN(\r60/ab[18][29] ), .IN0(\r60/CARRYB[17][29] ), 
        .IN1(\r60/SUMB[17][30] ), .COUT(\r60/CARRYB[18][29] ), .SUM(
        \r60/SUMB[18][29] ) );
  FADDER \r60/S2_18_28  ( .CIN(\r60/ab[18][28] ), .IN0(\r60/CARRYB[17][28] ), 
        .IN1(\r60/SUMB[17][29] ), .COUT(\r60/CARRYB[18][28] ), .SUM(
        \r60/SUMB[18][28] ) );
  FADDER \r60/S2_18_27  ( .CIN(\r60/ab[18][27] ), .IN0(\r60/CARRYB[17][27] ), 
        .IN1(\r60/SUMB[17][28] ), .COUT(\r60/CARRYB[18][27] ), .SUM(
        \r60/SUMB[18][27] ) );
  FADDER \r60/S2_18_26  ( .CIN(\r60/ab[18][26] ), .IN0(\r60/CARRYB[17][26] ), 
        .IN1(\r60/SUMB[17][27] ), .COUT(\r60/CARRYB[18][26] ), .SUM(
        \r60/SUMB[18][26] ) );
  FADDER \r60/S2_18_25  ( .CIN(\r60/ab[18][25] ), .IN0(\r60/CARRYB[17][25] ), 
        .IN1(\r60/SUMB[17][26] ), .COUT(\r60/CARRYB[18][25] ), .SUM(
        \r60/SUMB[18][25] ) );
  FADDER \r60/S2_18_24  ( .CIN(\r60/ab[18][24] ), .IN0(\r60/CARRYB[17][24] ), 
        .IN1(\r60/SUMB[17][25] ), .COUT(\r60/CARRYB[18][24] ), .SUM(
        \r60/SUMB[18][24] ) );
  FADDER \r60/S2_18_23  ( .CIN(\r60/ab[18][23] ), .IN0(\r60/CARRYB[17][23] ), 
        .IN1(\r60/SUMB[17][24] ), .COUT(\r60/CARRYB[18][23] ), .SUM(
        \r60/SUMB[18][23] ) );
  FADDER \r60/S2_18_22  ( .CIN(\r60/ab[18][22] ), .IN0(\r60/CARRYB[17][22] ), 
        .IN1(\r60/SUMB[17][23] ), .COUT(\r60/CARRYB[18][22] ), .SUM(
        \r60/SUMB[18][22] ) );
  FADDER \r60/S2_18_21  ( .CIN(\r60/ab[18][21] ), .IN0(\r60/CARRYB[17][21] ), 
        .IN1(\r60/SUMB[17][22] ), .COUT(\r60/CARRYB[18][21] ), .SUM(
        \r60/SUMB[18][21] ) );
  FADDER \r60/S2_18_20  ( .CIN(\r60/ab[18][20] ), .IN0(\r60/CARRYB[17][20] ), 
        .IN1(\r60/SUMB[17][21] ), .COUT(\r60/CARRYB[18][20] ), .SUM(
        \r60/SUMB[18][20] ) );
  FADDER \r60/S2_18_19  ( .CIN(\r60/ab[18][19] ), .IN0(\r60/CARRYB[17][19] ), 
        .IN1(\r60/SUMB[17][20] ), .COUT(\r60/CARRYB[18][19] ), .SUM(
        \r60/SUMB[18][19] ) );
  FADDER \r60/S2_18_18  ( .CIN(\r60/ab[18][18] ), .IN0(\r60/CARRYB[17][18] ), 
        .IN1(\r60/SUMB[17][19] ), .COUT(\r60/CARRYB[18][18] ), .SUM(
        \r60/SUMB[18][18] ) );
  FADDER \r60/S2_18_17  ( .CIN(\r60/ab[18][17] ), .IN0(\r60/CARRYB[17][17] ), 
        .IN1(\r60/SUMB[17][18] ), .COUT(\r60/CARRYB[18][17] ), .SUM(
        \r60/SUMB[18][17] ) );
  FADDER \r60/S2_18_16  ( .CIN(\r60/ab[18][16] ), .IN0(\r60/CARRYB[17][16] ), 
        .IN1(\r60/SUMB[17][17] ), .COUT(\r60/CARRYB[18][16] ), .SUM(
        \r60/SUMB[18][16] ) );
  FADDER \r60/S2_18_15  ( .CIN(\r60/ab[18][15] ), .IN0(\r60/CARRYB[17][15] ), 
        .IN1(\r60/SUMB[17][16] ), .COUT(\r60/CARRYB[18][15] ), .SUM(
        \r60/SUMB[18][15] ) );
  FADDER \r60/S2_18_14  ( .CIN(\r60/ab[18][14] ), .IN0(\r60/CARRYB[17][14] ), 
        .IN1(\r60/SUMB[17][15] ), .COUT(\r60/CARRYB[18][14] ), .SUM(
        \r60/SUMB[18][14] ) );
  FADDER \r60/S2_18_13  ( .CIN(\r60/ab[18][13] ), .IN0(\r60/CARRYB[17][13] ), 
        .IN1(\r60/SUMB[17][14] ), .COUT(\r60/CARRYB[18][13] ), .SUM(
        \r60/SUMB[18][13] ) );
  FADDER \r60/S2_18_12  ( .CIN(\r60/ab[18][12] ), .IN0(\r60/CARRYB[17][12] ), 
        .IN1(\r60/SUMB[17][13] ), .COUT(\r60/CARRYB[18][12] ), .SUM(
        \r60/SUMB[18][12] ) );
  FADDER \r60/S2_18_11  ( .CIN(\r60/ab[18][11] ), .IN0(\r60/CARRYB[17][11] ), 
        .IN1(\r60/SUMB[17][12] ), .COUT(\r60/CARRYB[18][11] ), .SUM(
        \r60/SUMB[18][11] ) );
  FADDER \r60/S2_18_10  ( .CIN(\r60/ab[18][10] ), .IN0(\r60/CARRYB[17][10] ), 
        .IN1(\r60/SUMB[17][11] ), .COUT(\r60/CARRYB[18][10] ), .SUM(
        \r60/SUMB[18][10] ) );
  FADDER \r60/S2_18_9  ( .CIN(\r60/ab[18][9] ), .IN0(\r60/CARRYB[17][9] ), 
        .IN1(\r60/SUMB[17][10] ), .COUT(\r60/CARRYB[18][9] ), .SUM(
        \r60/SUMB[18][9] ) );
  FADDER \r60/S2_18_8  ( .CIN(\r60/ab[18][8] ), .IN0(\r60/CARRYB[17][8] ), 
        .IN1(\r60/SUMB[17][9] ), .COUT(\r60/CARRYB[18][8] ), .SUM(
        \r60/SUMB[18][8] ) );
  FADDER \r60/S2_18_7  ( .CIN(\r60/ab[18][7] ), .IN0(\r60/CARRYB[17][7] ), 
        .IN1(\r60/SUMB[17][8] ), .COUT(\r60/CARRYB[18][7] ), .SUM(
        \r60/SUMB[18][7] ) );
  FADDER \r60/S2_18_6  ( .CIN(\r60/ab[18][6] ), .IN0(\r60/CARRYB[17][6] ), 
        .IN1(\r60/SUMB[17][7] ), .COUT(\r60/CARRYB[18][6] ), .SUM(
        \r60/SUMB[18][6] ) );
  FADDER \r60/S2_18_5  ( .CIN(\r60/ab[18][5] ), .IN0(\r60/CARRYB[17][5] ), 
        .IN1(\r60/SUMB[17][6] ), .COUT(\r60/CARRYB[18][5] ), .SUM(
        \r60/SUMB[18][5] ) );
  FADDER \r60/S2_18_4  ( .CIN(\r60/ab[18][4] ), .IN0(\r60/CARRYB[17][4] ), 
        .IN1(\r60/SUMB[17][5] ), .COUT(\r60/CARRYB[18][4] ), .SUM(
        \r60/SUMB[18][4] ) );
  FADDER \r60/S2_18_3  ( .CIN(\r60/ab[18][3] ), .IN0(\r60/CARRYB[17][3] ), 
        .IN1(\r60/SUMB[17][4] ), .COUT(\r60/CARRYB[18][3] ), .SUM(
        \r60/SUMB[18][3] ) );
  FADDER \r60/S2_18_2  ( .CIN(\r60/ab[18][2] ), .IN0(\r60/CARRYB[17][2] ), 
        .IN1(\r60/SUMB[17][3] ), .COUT(\r60/CARRYB[18][2] ), .SUM(
        \r60/SUMB[18][2] ) );
  FADDER \r60/S2_18_1  ( .CIN(\r60/ab[18][1] ), .IN0(\r60/CARRYB[17][1] ), 
        .IN1(\r60/SUMB[17][2] ), .COUT(\r60/CARRYB[18][1] ), .SUM(
        \r60/SUMB[18][1] ) );
  FADDER \r60/S1_18_0  ( .CIN(\r60/ab[18][0] ), .IN0(\r60/CARRYB[17][0] ), 
        .IN1(\r60/SUMB[17][1] ), .COUT(\r60/CARRYB[18][0] ), .SUM(N135) );
  FADDER \r60/S3_19_30  ( .CIN(\r60/ab[19][30] ), .IN0(\r60/CARRYB[18][30] ), 
        .IN1(\r60/ab[18][31] ), .COUT(\r60/CARRYB[19][30] ), .SUM(
        \r60/SUMB[19][30] ) );
  FADDER \r60/S2_19_29  ( .CIN(\r60/ab[19][29] ), .IN0(\r60/CARRYB[18][29] ), 
        .IN1(\r60/SUMB[18][30] ), .COUT(\r60/CARRYB[19][29] ), .SUM(
        \r60/SUMB[19][29] ) );
  FADDER \r60/S2_19_28  ( .CIN(\r60/ab[19][28] ), .IN0(\r60/CARRYB[18][28] ), 
        .IN1(\r60/SUMB[18][29] ), .COUT(\r60/CARRYB[19][28] ), .SUM(
        \r60/SUMB[19][28] ) );
  FADDER \r60/S2_19_27  ( .CIN(\r60/ab[19][27] ), .IN0(\r60/CARRYB[18][27] ), 
        .IN1(\r60/SUMB[18][28] ), .COUT(\r60/CARRYB[19][27] ), .SUM(
        \r60/SUMB[19][27] ) );
  FADDER \r60/S2_19_26  ( .CIN(\r60/ab[19][26] ), .IN0(\r60/CARRYB[18][26] ), 
        .IN1(\r60/SUMB[18][27] ), .COUT(\r60/CARRYB[19][26] ), .SUM(
        \r60/SUMB[19][26] ) );
  FADDER \r60/S2_19_25  ( .CIN(\r60/ab[19][25] ), .IN0(\r60/CARRYB[18][25] ), 
        .IN1(\r60/SUMB[18][26] ), .COUT(\r60/CARRYB[19][25] ), .SUM(
        \r60/SUMB[19][25] ) );
  FADDER \r60/S2_19_24  ( .CIN(\r60/ab[19][24] ), .IN0(\r60/CARRYB[18][24] ), 
        .IN1(\r60/SUMB[18][25] ), .COUT(\r60/CARRYB[19][24] ), .SUM(
        \r60/SUMB[19][24] ) );
  FADDER \r60/S2_19_23  ( .CIN(\r60/ab[19][23] ), .IN0(\r60/CARRYB[18][23] ), 
        .IN1(\r60/SUMB[18][24] ), .COUT(\r60/CARRYB[19][23] ), .SUM(
        \r60/SUMB[19][23] ) );
  FADDER \r60/S2_19_22  ( .CIN(\r60/ab[19][22] ), .IN0(\r60/CARRYB[18][22] ), 
        .IN1(\r60/SUMB[18][23] ), .COUT(\r60/CARRYB[19][22] ), .SUM(
        \r60/SUMB[19][22] ) );
  FADDER \r60/S2_19_21  ( .CIN(\r60/ab[19][21] ), .IN0(\r60/CARRYB[18][21] ), 
        .IN1(\r60/SUMB[18][22] ), .COUT(\r60/CARRYB[19][21] ), .SUM(
        \r60/SUMB[19][21] ) );
  FADDER \r60/S2_19_20  ( .CIN(\r60/ab[19][20] ), .IN0(\r60/CARRYB[18][20] ), 
        .IN1(\r60/SUMB[18][21] ), .COUT(\r60/CARRYB[19][20] ), .SUM(
        \r60/SUMB[19][20] ) );
  FADDER \r60/S2_19_19  ( .CIN(\r60/ab[19][19] ), .IN0(\r60/CARRYB[18][19] ), 
        .IN1(\r60/SUMB[18][20] ), .COUT(\r60/CARRYB[19][19] ), .SUM(
        \r60/SUMB[19][19] ) );
  FADDER \r60/S2_19_18  ( .CIN(\r60/ab[19][18] ), .IN0(\r60/CARRYB[18][18] ), 
        .IN1(\r60/SUMB[18][19] ), .COUT(\r60/CARRYB[19][18] ), .SUM(
        \r60/SUMB[19][18] ) );
  FADDER \r60/S2_19_17  ( .CIN(\r60/ab[19][17] ), .IN0(\r60/CARRYB[18][17] ), 
        .IN1(\r60/SUMB[18][18] ), .COUT(\r60/CARRYB[19][17] ), .SUM(
        \r60/SUMB[19][17] ) );
  FADDER \r60/S2_19_16  ( .CIN(\r60/ab[19][16] ), .IN0(\r60/CARRYB[18][16] ), 
        .IN1(\r60/SUMB[18][17] ), .COUT(\r60/CARRYB[19][16] ), .SUM(
        \r60/SUMB[19][16] ) );
  FADDER \r60/S2_19_15  ( .CIN(\r60/ab[19][15] ), .IN0(\r60/CARRYB[18][15] ), 
        .IN1(\r60/SUMB[18][16] ), .COUT(\r60/CARRYB[19][15] ), .SUM(
        \r60/SUMB[19][15] ) );
  FADDER \r60/S2_19_14  ( .CIN(\r60/ab[19][14] ), .IN0(\r60/CARRYB[18][14] ), 
        .IN1(\r60/SUMB[18][15] ), .COUT(\r60/CARRYB[19][14] ), .SUM(
        \r60/SUMB[19][14] ) );
  FADDER \r60/S2_19_13  ( .CIN(\r60/ab[19][13] ), .IN0(\r60/CARRYB[18][13] ), 
        .IN1(\r60/SUMB[18][14] ), .COUT(\r60/CARRYB[19][13] ), .SUM(
        \r60/SUMB[19][13] ) );
  FADDER \r60/S2_19_12  ( .CIN(\r60/ab[19][12] ), .IN0(\r60/CARRYB[18][12] ), 
        .IN1(\r60/SUMB[18][13] ), .COUT(\r60/CARRYB[19][12] ), .SUM(
        \r60/SUMB[19][12] ) );
  FADDER \r60/S2_19_11  ( .CIN(\r60/ab[19][11] ), .IN0(\r60/CARRYB[18][11] ), 
        .IN1(\r60/SUMB[18][12] ), .COUT(\r60/CARRYB[19][11] ), .SUM(
        \r60/SUMB[19][11] ) );
  FADDER \r60/S2_19_10  ( .CIN(\r60/ab[19][10] ), .IN0(\r60/CARRYB[18][10] ), 
        .IN1(\r60/SUMB[18][11] ), .COUT(\r60/CARRYB[19][10] ), .SUM(
        \r60/SUMB[19][10] ) );
  FADDER \r60/S2_19_9  ( .CIN(\r60/ab[19][9] ), .IN0(\r60/CARRYB[18][9] ), 
        .IN1(\r60/SUMB[18][10] ), .COUT(\r60/CARRYB[19][9] ), .SUM(
        \r60/SUMB[19][9] ) );
  FADDER \r60/S2_19_8  ( .CIN(\r60/ab[19][8] ), .IN0(\r60/CARRYB[18][8] ), 
        .IN1(\r60/SUMB[18][9] ), .COUT(\r60/CARRYB[19][8] ), .SUM(
        \r60/SUMB[19][8] ) );
  FADDER \r60/S2_19_7  ( .CIN(\r60/ab[19][7] ), .IN0(\r60/CARRYB[18][7] ), 
        .IN1(\r60/SUMB[18][8] ), .COUT(\r60/CARRYB[19][7] ), .SUM(
        \r60/SUMB[19][7] ) );
  FADDER \r60/S2_19_6  ( .CIN(\r60/ab[19][6] ), .IN0(\r60/CARRYB[18][6] ), 
        .IN1(\r60/SUMB[18][7] ), .COUT(\r60/CARRYB[19][6] ), .SUM(
        \r60/SUMB[19][6] ) );
  FADDER \r60/S2_19_5  ( .CIN(\r60/ab[19][5] ), .IN0(\r60/CARRYB[18][5] ), 
        .IN1(\r60/SUMB[18][6] ), .COUT(\r60/CARRYB[19][5] ), .SUM(
        \r60/SUMB[19][5] ) );
  FADDER \r60/S2_19_4  ( .CIN(\r60/ab[19][4] ), .IN0(\r60/CARRYB[18][4] ), 
        .IN1(\r60/SUMB[18][5] ), .COUT(\r60/CARRYB[19][4] ), .SUM(
        \r60/SUMB[19][4] ) );
  FADDER \r60/S2_19_3  ( .CIN(\r60/ab[19][3] ), .IN0(\r60/CARRYB[18][3] ), 
        .IN1(\r60/SUMB[18][4] ), .COUT(\r60/CARRYB[19][3] ), .SUM(
        \r60/SUMB[19][3] ) );
  FADDER \r60/S2_19_2  ( .CIN(\r60/ab[19][2] ), .IN0(\r60/CARRYB[18][2] ), 
        .IN1(\r60/SUMB[18][3] ), .COUT(\r60/CARRYB[19][2] ), .SUM(
        \r60/SUMB[19][2] ) );
  FADDER \r60/S2_19_1  ( .CIN(\r60/ab[19][1] ), .IN0(\r60/CARRYB[18][1] ), 
        .IN1(\r60/SUMB[18][2] ), .COUT(\r60/CARRYB[19][1] ), .SUM(
        \r60/SUMB[19][1] ) );
  FADDER \r60/S1_19_0  ( .CIN(\r60/ab[19][0] ), .IN0(\r60/CARRYB[18][0] ), 
        .IN1(\r60/SUMB[18][1] ), .COUT(\r60/CARRYB[19][0] ), .SUM(N136) );
  FADDER \r60/S3_20_30  ( .CIN(\r60/ab[20][30] ), .IN0(\r60/CARRYB[19][30] ), 
        .IN1(\r60/ab[19][31] ), .COUT(\r60/CARRYB[20][30] ), .SUM(
        \r60/SUMB[20][30] ) );
  FADDER \r60/S2_20_29  ( .CIN(\r60/ab[20][29] ), .IN0(\r60/CARRYB[19][29] ), 
        .IN1(\r60/SUMB[19][30] ), .COUT(\r60/CARRYB[20][29] ), .SUM(
        \r60/SUMB[20][29] ) );
  FADDER \r60/S2_20_28  ( .CIN(\r60/ab[20][28] ), .IN0(\r60/CARRYB[19][28] ), 
        .IN1(\r60/SUMB[19][29] ), .COUT(\r60/CARRYB[20][28] ), .SUM(
        \r60/SUMB[20][28] ) );
  FADDER \r60/S2_20_27  ( .CIN(\r60/ab[20][27] ), .IN0(\r60/CARRYB[19][27] ), 
        .IN1(\r60/SUMB[19][28] ), .COUT(\r60/CARRYB[20][27] ), .SUM(
        \r60/SUMB[20][27] ) );
  FADDER \r60/S2_20_26  ( .CIN(\r60/ab[20][26] ), .IN0(\r60/CARRYB[19][26] ), 
        .IN1(\r60/SUMB[19][27] ), .COUT(\r60/CARRYB[20][26] ), .SUM(
        \r60/SUMB[20][26] ) );
  FADDER \r60/S2_20_25  ( .CIN(\r60/ab[20][25] ), .IN0(\r60/CARRYB[19][25] ), 
        .IN1(\r60/SUMB[19][26] ), .COUT(\r60/CARRYB[20][25] ), .SUM(
        \r60/SUMB[20][25] ) );
  FADDER \r60/S2_20_24  ( .CIN(\r60/ab[20][24] ), .IN0(\r60/CARRYB[19][24] ), 
        .IN1(\r60/SUMB[19][25] ), .COUT(\r60/CARRYB[20][24] ), .SUM(
        \r60/SUMB[20][24] ) );
  FADDER \r60/S2_20_23  ( .CIN(\r60/ab[20][23] ), .IN0(\r60/CARRYB[19][23] ), 
        .IN1(\r60/SUMB[19][24] ), .COUT(\r60/CARRYB[20][23] ), .SUM(
        \r60/SUMB[20][23] ) );
  FADDER \r60/S2_20_22  ( .CIN(\r60/ab[20][22] ), .IN0(\r60/CARRYB[19][22] ), 
        .IN1(\r60/SUMB[19][23] ), .COUT(\r60/CARRYB[20][22] ), .SUM(
        \r60/SUMB[20][22] ) );
  FADDER \r60/S2_20_21  ( .CIN(\r60/ab[20][21] ), .IN0(\r60/CARRYB[19][21] ), 
        .IN1(\r60/SUMB[19][22] ), .COUT(\r60/CARRYB[20][21] ), .SUM(
        \r60/SUMB[20][21] ) );
  FADDER \r60/S2_20_20  ( .CIN(\r60/ab[20][20] ), .IN0(\r60/CARRYB[19][20] ), 
        .IN1(\r60/SUMB[19][21] ), .COUT(\r60/CARRYB[20][20] ), .SUM(
        \r60/SUMB[20][20] ) );
  FADDER \r60/S2_20_19  ( .CIN(\r60/ab[20][19] ), .IN0(\r60/CARRYB[19][19] ), 
        .IN1(\r60/SUMB[19][20] ), .COUT(\r60/CARRYB[20][19] ), .SUM(
        \r60/SUMB[20][19] ) );
  FADDER \r60/S2_20_18  ( .CIN(\r60/ab[20][18] ), .IN0(\r60/CARRYB[19][18] ), 
        .IN1(\r60/SUMB[19][19] ), .COUT(\r60/CARRYB[20][18] ), .SUM(
        \r60/SUMB[20][18] ) );
  FADDER \r60/S2_20_17  ( .CIN(\r60/ab[20][17] ), .IN0(\r60/CARRYB[19][17] ), 
        .IN1(\r60/SUMB[19][18] ), .COUT(\r60/CARRYB[20][17] ), .SUM(
        \r60/SUMB[20][17] ) );
  FADDER \r60/S2_20_16  ( .CIN(\r60/ab[20][16] ), .IN0(\r60/CARRYB[19][16] ), 
        .IN1(\r60/SUMB[19][17] ), .COUT(\r60/CARRYB[20][16] ), .SUM(
        \r60/SUMB[20][16] ) );
  FADDER \r60/S2_20_15  ( .CIN(\r60/ab[20][15] ), .IN0(\r60/CARRYB[19][15] ), 
        .IN1(\r60/SUMB[19][16] ), .COUT(\r60/CARRYB[20][15] ), .SUM(
        \r60/SUMB[20][15] ) );
  FADDER \r60/S2_20_14  ( .CIN(\r60/ab[20][14] ), .IN0(\r60/CARRYB[19][14] ), 
        .IN1(\r60/SUMB[19][15] ), .COUT(\r60/CARRYB[20][14] ), .SUM(
        \r60/SUMB[20][14] ) );
  FADDER \r60/S2_20_13  ( .CIN(\r60/ab[20][13] ), .IN0(\r60/CARRYB[19][13] ), 
        .IN1(\r60/SUMB[19][14] ), .COUT(\r60/CARRYB[20][13] ), .SUM(
        \r60/SUMB[20][13] ) );
  FADDER \r60/S2_20_12  ( .CIN(\r60/ab[20][12] ), .IN0(\r60/CARRYB[19][12] ), 
        .IN1(\r60/SUMB[19][13] ), .COUT(\r60/CARRYB[20][12] ), .SUM(
        \r60/SUMB[20][12] ) );
  FADDER \r60/S2_20_11  ( .CIN(\r60/ab[20][11] ), .IN0(\r60/CARRYB[19][11] ), 
        .IN1(\r60/SUMB[19][12] ), .COUT(\r60/CARRYB[20][11] ), .SUM(
        \r60/SUMB[20][11] ) );
  FADDER \r60/S2_20_10  ( .CIN(\r60/ab[20][10] ), .IN0(\r60/CARRYB[19][10] ), 
        .IN1(\r60/SUMB[19][11] ), .COUT(\r60/CARRYB[20][10] ), .SUM(
        \r60/SUMB[20][10] ) );
  FADDER \r60/S2_20_9  ( .CIN(\r60/ab[20][9] ), .IN0(\r60/CARRYB[19][9] ), 
        .IN1(\r60/SUMB[19][10] ), .COUT(\r60/CARRYB[20][9] ), .SUM(
        \r60/SUMB[20][9] ) );
  FADDER \r60/S2_20_8  ( .CIN(\r60/ab[20][8] ), .IN0(\r60/CARRYB[19][8] ), 
        .IN1(\r60/SUMB[19][9] ), .COUT(\r60/CARRYB[20][8] ), .SUM(
        \r60/SUMB[20][8] ) );
  FADDER \r60/S2_20_7  ( .CIN(\r60/ab[20][7] ), .IN0(\r60/CARRYB[19][7] ), 
        .IN1(\r60/SUMB[19][8] ), .COUT(\r60/CARRYB[20][7] ), .SUM(
        \r60/SUMB[20][7] ) );
  FADDER \r60/S2_20_6  ( .CIN(\r60/ab[20][6] ), .IN0(\r60/CARRYB[19][6] ), 
        .IN1(\r60/SUMB[19][7] ), .COUT(\r60/CARRYB[20][6] ), .SUM(
        \r60/SUMB[20][6] ) );
  FADDER \r60/S2_20_5  ( .CIN(\r60/ab[20][5] ), .IN0(\r60/CARRYB[19][5] ), 
        .IN1(\r60/SUMB[19][6] ), .COUT(\r60/CARRYB[20][5] ), .SUM(
        \r60/SUMB[20][5] ) );
  FADDER \r60/S2_20_4  ( .CIN(\r60/ab[20][4] ), .IN0(\r60/CARRYB[19][4] ), 
        .IN1(\r60/SUMB[19][5] ), .COUT(\r60/CARRYB[20][4] ), .SUM(
        \r60/SUMB[20][4] ) );
  FADDER \r60/S2_20_3  ( .CIN(\r60/ab[20][3] ), .IN0(\r60/CARRYB[19][3] ), 
        .IN1(\r60/SUMB[19][4] ), .COUT(\r60/CARRYB[20][3] ), .SUM(
        \r60/SUMB[20][3] ) );
  FADDER \r60/S2_20_2  ( .CIN(\r60/ab[20][2] ), .IN0(\r60/CARRYB[19][2] ), 
        .IN1(\r60/SUMB[19][3] ), .COUT(\r60/CARRYB[20][2] ), .SUM(
        \r60/SUMB[20][2] ) );
  FADDER \r60/S2_20_1  ( .CIN(\r60/ab[20][1] ), .IN0(\r60/CARRYB[19][1] ), 
        .IN1(\r60/SUMB[19][2] ), .COUT(\r60/CARRYB[20][1] ), .SUM(
        \r60/SUMB[20][1] ) );
  FADDER \r60/S1_20_0  ( .CIN(\r60/ab[20][0] ), .IN0(\r60/CARRYB[19][0] ), 
        .IN1(\r60/SUMB[19][1] ), .COUT(\r60/CARRYB[20][0] ), .SUM(N137) );
  FADDER \r60/S3_21_30  ( .CIN(\r60/ab[21][30] ), .IN0(\r60/CARRYB[20][30] ), 
        .IN1(\r60/ab[20][31] ), .COUT(\r60/CARRYB[21][30] ), .SUM(
        \r60/SUMB[21][30] ) );
  FADDER \r60/S2_21_29  ( .CIN(\r60/ab[21][29] ), .IN0(\r60/CARRYB[20][29] ), 
        .IN1(\r60/SUMB[20][30] ), .COUT(\r60/CARRYB[21][29] ), .SUM(
        \r60/SUMB[21][29] ) );
  FADDER \r60/S2_21_28  ( .CIN(\r60/ab[21][28] ), .IN0(\r60/CARRYB[20][28] ), 
        .IN1(\r60/SUMB[20][29] ), .COUT(\r60/CARRYB[21][28] ), .SUM(
        \r60/SUMB[21][28] ) );
  FADDER \r60/S2_21_27  ( .CIN(\r60/ab[21][27] ), .IN0(\r60/CARRYB[20][27] ), 
        .IN1(\r60/SUMB[20][28] ), .COUT(\r60/CARRYB[21][27] ), .SUM(
        \r60/SUMB[21][27] ) );
  FADDER \r60/S2_21_26  ( .CIN(\r60/ab[21][26] ), .IN0(\r60/CARRYB[20][26] ), 
        .IN1(\r60/SUMB[20][27] ), .COUT(\r60/CARRYB[21][26] ), .SUM(
        \r60/SUMB[21][26] ) );
  FADDER \r60/S2_21_25  ( .CIN(\r60/ab[21][25] ), .IN0(\r60/CARRYB[20][25] ), 
        .IN1(\r60/SUMB[20][26] ), .COUT(\r60/CARRYB[21][25] ), .SUM(
        \r60/SUMB[21][25] ) );
  FADDER \r60/S2_21_24  ( .CIN(\r60/ab[21][24] ), .IN0(\r60/CARRYB[20][24] ), 
        .IN1(\r60/SUMB[20][25] ), .COUT(\r60/CARRYB[21][24] ), .SUM(
        \r60/SUMB[21][24] ) );
  FADDER \r60/S2_21_23  ( .CIN(\r60/ab[21][23] ), .IN0(\r60/CARRYB[20][23] ), 
        .IN1(\r60/SUMB[20][24] ), .COUT(\r60/CARRYB[21][23] ), .SUM(
        \r60/SUMB[21][23] ) );
  FADDER \r60/S2_21_22  ( .CIN(\r60/ab[21][22] ), .IN0(\r60/CARRYB[20][22] ), 
        .IN1(\r60/SUMB[20][23] ), .COUT(\r60/CARRYB[21][22] ), .SUM(
        \r60/SUMB[21][22] ) );
  FADDER \r60/S2_21_21  ( .CIN(\r60/ab[21][21] ), .IN0(\r60/CARRYB[20][21] ), 
        .IN1(\r60/SUMB[20][22] ), .COUT(\r60/CARRYB[21][21] ), .SUM(
        \r60/SUMB[21][21] ) );
  FADDER \r60/S2_21_20  ( .CIN(\r60/ab[21][20] ), .IN0(\r60/CARRYB[20][20] ), 
        .IN1(\r60/SUMB[20][21] ), .COUT(\r60/CARRYB[21][20] ), .SUM(
        \r60/SUMB[21][20] ) );
  FADDER \r60/S2_21_19  ( .CIN(\r60/ab[21][19] ), .IN0(\r60/CARRYB[20][19] ), 
        .IN1(\r60/SUMB[20][20] ), .COUT(\r60/CARRYB[21][19] ), .SUM(
        \r60/SUMB[21][19] ) );
  FADDER \r60/S2_21_18  ( .CIN(\r60/ab[21][18] ), .IN0(\r60/CARRYB[20][18] ), 
        .IN1(\r60/SUMB[20][19] ), .COUT(\r60/CARRYB[21][18] ), .SUM(
        \r60/SUMB[21][18] ) );
  FADDER \r60/S2_21_17  ( .CIN(\r60/ab[21][17] ), .IN0(\r60/CARRYB[20][17] ), 
        .IN1(\r60/SUMB[20][18] ), .COUT(\r60/CARRYB[21][17] ), .SUM(
        \r60/SUMB[21][17] ) );
  FADDER \r60/S2_21_16  ( .CIN(\r60/ab[21][16] ), .IN0(\r60/CARRYB[20][16] ), 
        .IN1(\r60/SUMB[20][17] ), .COUT(\r60/CARRYB[21][16] ), .SUM(
        \r60/SUMB[21][16] ) );
  FADDER \r60/S2_21_15  ( .CIN(\r60/ab[21][15] ), .IN0(\r60/CARRYB[20][15] ), 
        .IN1(\r60/SUMB[20][16] ), .COUT(\r60/CARRYB[21][15] ), .SUM(
        \r60/SUMB[21][15] ) );
  FADDER \r60/S2_21_14  ( .CIN(\r60/ab[21][14] ), .IN0(\r60/CARRYB[20][14] ), 
        .IN1(\r60/SUMB[20][15] ), .COUT(\r60/CARRYB[21][14] ), .SUM(
        \r60/SUMB[21][14] ) );
  FADDER \r60/S2_21_13  ( .CIN(\r60/ab[21][13] ), .IN0(\r60/CARRYB[20][13] ), 
        .IN1(\r60/SUMB[20][14] ), .COUT(\r60/CARRYB[21][13] ), .SUM(
        \r60/SUMB[21][13] ) );
  FADDER \r60/S2_21_12  ( .CIN(\r60/ab[21][12] ), .IN0(\r60/CARRYB[20][12] ), 
        .IN1(\r60/SUMB[20][13] ), .COUT(\r60/CARRYB[21][12] ), .SUM(
        \r60/SUMB[21][12] ) );
  FADDER \r60/S2_21_11  ( .CIN(\r60/ab[21][11] ), .IN0(\r60/CARRYB[20][11] ), 
        .IN1(\r60/SUMB[20][12] ), .COUT(\r60/CARRYB[21][11] ), .SUM(
        \r60/SUMB[21][11] ) );
  FADDER \r60/S2_21_10  ( .CIN(\r60/ab[21][10] ), .IN0(\r60/CARRYB[20][10] ), 
        .IN1(\r60/SUMB[20][11] ), .COUT(\r60/CARRYB[21][10] ), .SUM(
        \r60/SUMB[21][10] ) );
  FADDER \r60/S2_21_9  ( .CIN(\r60/ab[21][9] ), .IN0(\r60/CARRYB[20][9] ), 
        .IN1(\r60/SUMB[20][10] ), .COUT(\r60/CARRYB[21][9] ), .SUM(
        \r60/SUMB[21][9] ) );
  FADDER \r60/S2_21_8  ( .CIN(\r60/ab[21][8] ), .IN0(\r60/CARRYB[20][8] ), 
        .IN1(\r60/SUMB[20][9] ), .COUT(\r60/CARRYB[21][8] ), .SUM(
        \r60/SUMB[21][8] ) );
  FADDER \r60/S2_21_7  ( .CIN(\r60/ab[21][7] ), .IN0(\r60/CARRYB[20][7] ), 
        .IN1(\r60/SUMB[20][8] ), .COUT(\r60/CARRYB[21][7] ), .SUM(
        \r60/SUMB[21][7] ) );
  FADDER \r60/S2_21_6  ( .CIN(\r60/ab[21][6] ), .IN0(\r60/CARRYB[20][6] ), 
        .IN1(\r60/SUMB[20][7] ), .COUT(\r60/CARRYB[21][6] ), .SUM(
        \r60/SUMB[21][6] ) );
  FADDER \r60/S2_21_5  ( .CIN(\r60/ab[21][5] ), .IN0(\r60/CARRYB[20][5] ), 
        .IN1(\r60/SUMB[20][6] ), .COUT(\r60/CARRYB[21][5] ), .SUM(
        \r60/SUMB[21][5] ) );
  FADDER \r60/S2_21_4  ( .CIN(\r60/ab[21][4] ), .IN0(\r60/CARRYB[20][4] ), 
        .IN1(\r60/SUMB[20][5] ), .COUT(\r60/CARRYB[21][4] ), .SUM(
        \r60/SUMB[21][4] ) );
  FADDER \r60/S2_21_3  ( .CIN(\r60/ab[21][3] ), .IN0(\r60/CARRYB[20][3] ), 
        .IN1(\r60/SUMB[20][4] ), .COUT(\r60/CARRYB[21][3] ), .SUM(
        \r60/SUMB[21][3] ) );
  FADDER \r60/S2_21_2  ( .CIN(\r60/ab[21][2] ), .IN0(\r60/CARRYB[20][2] ), 
        .IN1(\r60/SUMB[20][3] ), .COUT(\r60/CARRYB[21][2] ), .SUM(
        \r60/SUMB[21][2] ) );
  FADDER \r60/S2_21_1  ( .CIN(\r60/ab[21][1] ), .IN0(\r60/CARRYB[20][1] ), 
        .IN1(\r60/SUMB[20][2] ), .COUT(\r60/CARRYB[21][1] ), .SUM(
        \r60/SUMB[21][1] ) );
  FADDER \r60/S1_21_0  ( .CIN(\r60/ab[21][0] ), .IN0(\r60/CARRYB[20][0] ), 
        .IN1(\r60/SUMB[20][1] ), .COUT(\r60/CARRYB[21][0] ), .SUM(N138) );
  FADDER \r60/S3_22_30  ( .CIN(\r60/ab[22][30] ), .IN0(\r60/CARRYB[21][30] ), 
        .IN1(\r60/ab[21][31] ), .COUT(\r60/CARRYB[22][30] ), .SUM(
        \r60/SUMB[22][30] ) );
  FADDER \r60/S2_22_29  ( .CIN(\r60/ab[22][29] ), .IN0(\r60/CARRYB[21][29] ), 
        .IN1(\r60/SUMB[21][30] ), .COUT(\r60/CARRYB[22][29] ), .SUM(
        \r60/SUMB[22][29] ) );
  FADDER \r60/S2_22_28  ( .CIN(\r60/ab[22][28] ), .IN0(\r60/CARRYB[21][28] ), 
        .IN1(\r60/SUMB[21][29] ), .COUT(\r60/CARRYB[22][28] ), .SUM(
        \r60/SUMB[22][28] ) );
  FADDER \r60/S2_22_27  ( .CIN(\r60/ab[22][27] ), .IN0(\r60/CARRYB[21][27] ), 
        .IN1(\r60/SUMB[21][28] ), .COUT(\r60/CARRYB[22][27] ), .SUM(
        \r60/SUMB[22][27] ) );
  FADDER \r60/S2_22_26  ( .CIN(\r60/ab[22][26] ), .IN0(\r60/CARRYB[21][26] ), 
        .IN1(\r60/SUMB[21][27] ), .COUT(\r60/CARRYB[22][26] ), .SUM(
        \r60/SUMB[22][26] ) );
  FADDER \r60/S2_22_25  ( .CIN(\r60/ab[22][25] ), .IN0(\r60/CARRYB[21][25] ), 
        .IN1(\r60/SUMB[21][26] ), .COUT(\r60/CARRYB[22][25] ), .SUM(
        \r60/SUMB[22][25] ) );
  FADDER \r60/S2_22_24  ( .CIN(\r60/ab[22][24] ), .IN0(\r60/CARRYB[21][24] ), 
        .IN1(\r60/SUMB[21][25] ), .COUT(\r60/CARRYB[22][24] ), .SUM(
        \r60/SUMB[22][24] ) );
  FADDER \r60/S2_22_23  ( .CIN(\r60/ab[22][23] ), .IN0(\r60/CARRYB[21][23] ), 
        .IN1(\r60/SUMB[21][24] ), .COUT(\r60/CARRYB[22][23] ), .SUM(
        \r60/SUMB[22][23] ) );
  FADDER \r60/S2_22_22  ( .CIN(\r60/ab[22][22] ), .IN0(\r60/CARRYB[21][22] ), 
        .IN1(\r60/SUMB[21][23] ), .COUT(\r60/CARRYB[22][22] ), .SUM(
        \r60/SUMB[22][22] ) );
  FADDER \r60/S2_22_21  ( .CIN(\r60/ab[22][21] ), .IN0(\r60/CARRYB[21][21] ), 
        .IN1(\r60/SUMB[21][22] ), .COUT(\r60/CARRYB[22][21] ), .SUM(
        \r60/SUMB[22][21] ) );
  FADDER \r60/S2_22_20  ( .CIN(\r60/ab[22][20] ), .IN0(\r60/CARRYB[21][20] ), 
        .IN1(\r60/SUMB[21][21] ), .COUT(\r60/CARRYB[22][20] ), .SUM(
        \r60/SUMB[22][20] ) );
  FADDER \r60/S2_22_19  ( .CIN(\r60/ab[22][19] ), .IN0(\r60/CARRYB[21][19] ), 
        .IN1(\r60/SUMB[21][20] ), .COUT(\r60/CARRYB[22][19] ), .SUM(
        \r60/SUMB[22][19] ) );
  FADDER \r60/S2_22_18  ( .CIN(\r60/ab[22][18] ), .IN0(\r60/CARRYB[21][18] ), 
        .IN1(\r60/SUMB[21][19] ), .COUT(\r60/CARRYB[22][18] ), .SUM(
        \r60/SUMB[22][18] ) );
  FADDER \r60/S2_22_17  ( .CIN(\r60/ab[22][17] ), .IN0(\r60/CARRYB[21][17] ), 
        .IN1(\r60/SUMB[21][18] ), .COUT(\r60/CARRYB[22][17] ), .SUM(
        \r60/SUMB[22][17] ) );
  FADDER \r60/S2_22_16  ( .CIN(\r60/ab[22][16] ), .IN0(\r60/CARRYB[21][16] ), 
        .IN1(\r60/SUMB[21][17] ), .COUT(\r60/CARRYB[22][16] ), .SUM(
        \r60/SUMB[22][16] ) );
  FADDER \r60/S2_22_15  ( .CIN(\r60/ab[22][15] ), .IN0(\r60/CARRYB[21][15] ), 
        .IN1(\r60/SUMB[21][16] ), .COUT(\r60/CARRYB[22][15] ), .SUM(
        \r60/SUMB[22][15] ) );
  FADDER \r60/S2_22_14  ( .CIN(\r60/ab[22][14] ), .IN0(\r60/CARRYB[21][14] ), 
        .IN1(\r60/SUMB[21][15] ), .COUT(\r60/CARRYB[22][14] ), .SUM(
        \r60/SUMB[22][14] ) );
  FADDER \r60/S2_22_13  ( .CIN(\r60/ab[22][13] ), .IN0(\r60/CARRYB[21][13] ), 
        .IN1(\r60/SUMB[21][14] ), .COUT(\r60/CARRYB[22][13] ), .SUM(
        \r60/SUMB[22][13] ) );
  FADDER \r60/S2_22_12  ( .CIN(\r60/ab[22][12] ), .IN0(\r60/CARRYB[21][12] ), 
        .IN1(\r60/SUMB[21][13] ), .COUT(\r60/CARRYB[22][12] ), .SUM(
        \r60/SUMB[22][12] ) );
  FADDER \r60/S2_22_11  ( .CIN(\r60/ab[22][11] ), .IN0(\r60/CARRYB[21][11] ), 
        .IN1(\r60/SUMB[21][12] ), .COUT(\r60/CARRYB[22][11] ), .SUM(
        \r60/SUMB[22][11] ) );
  FADDER \r60/S2_22_10  ( .CIN(\r60/ab[22][10] ), .IN0(\r60/CARRYB[21][10] ), 
        .IN1(\r60/SUMB[21][11] ), .COUT(\r60/CARRYB[22][10] ), .SUM(
        \r60/SUMB[22][10] ) );
  FADDER \r60/S2_22_9  ( .CIN(\r60/ab[22][9] ), .IN0(\r60/CARRYB[21][9] ), 
        .IN1(\r60/SUMB[21][10] ), .COUT(\r60/CARRYB[22][9] ), .SUM(
        \r60/SUMB[22][9] ) );
  FADDER \r60/S2_22_8  ( .CIN(\r60/ab[22][8] ), .IN0(\r60/CARRYB[21][8] ), 
        .IN1(\r60/SUMB[21][9] ), .COUT(\r60/CARRYB[22][8] ), .SUM(
        \r60/SUMB[22][8] ) );
  FADDER \r60/S2_22_7  ( .CIN(\r60/ab[22][7] ), .IN0(\r60/CARRYB[21][7] ), 
        .IN1(\r60/SUMB[21][8] ), .COUT(\r60/CARRYB[22][7] ), .SUM(
        \r60/SUMB[22][7] ) );
  FADDER \r60/S2_22_6  ( .CIN(\r60/ab[22][6] ), .IN0(\r60/CARRYB[21][6] ), 
        .IN1(\r60/SUMB[21][7] ), .COUT(\r60/CARRYB[22][6] ), .SUM(
        \r60/SUMB[22][6] ) );
  FADDER \r60/S2_22_5  ( .CIN(\r60/ab[22][5] ), .IN0(\r60/CARRYB[21][5] ), 
        .IN1(\r60/SUMB[21][6] ), .COUT(\r60/CARRYB[22][5] ), .SUM(
        \r60/SUMB[22][5] ) );
  FADDER \r60/S2_22_4  ( .CIN(\r60/ab[22][4] ), .IN0(\r60/CARRYB[21][4] ), 
        .IN1(\r60/SUMB[21][5] ), .COUT(\r60/CARRYB[22][4] ), .SUM(
        \r60/SUMB[22][4] ) );
  FADDER \r60/S2_22_3  ( .CIN(\r60/ab[22][3] ), .IN0(\r60/CARRYB[21][3] ), 
        .IN1(\r60/SUMB[21][4] ), .COUT(\r60/CARRYB[22][3] ), .SUM(
        \r60/SUMB[22][3] ) );
  FADDER \r60/S2_22_2  ( .CIN(\r60/ab[22][2] ), .IN0(\r60/CARRYB[21][2] ), 
        .IN1(\r60/SUMB[21][3] ), .COUT(\r60/CARRYB[22][2] ), .SUM(
        \r60/SUMB[22][2] ) );
  FADDER \r60/S2_22_1  ( .CIN(\r60/ab[22][1] ), .IN0(\r60/CARRYB[21][1] ), 
        .IN1(\r60/SUMB[21][2] ), .COUT(\r60/CARRYB[22][1] ), .SUM(
        \r60/SUMB[22][1] ) );
  FADDER \r60/S1_22_0  ( .CIN(\r60/ab[22][0] ), .IN0(\r60/CARRYB[21][0] ), 
        .IN1(\r60/SUMB[21][1] ), .COUT(\r60/CARRYB[22][0] ), .SUM(N139) );
  FADDER \r60/S3_23_30  ( .CIN(\r60/ab[23][30] ), .IN0(\r60/CARRYB[22][30] ), 
        .IN1(\r60/ab[22][31] ), .COUT(\r60/CARRYB[23][30] ), .SUM(
        \r60/SUMB[23][30] ) );
  FADDER \r60/S2_23_29  ( .CIN(\r60/ab[23][29] ), .IN0(\r60/CARRYB[22][29] ), 
        .IN1(\r60/SUMB[22][30] ), .COUT(\r60/CARRYB[23][29] ), .SUM(
        \r60/SUMB[23][29] ) );
  FADDER \r60/S2_23_28  ( .CIN(\r60/ab[23][28] ), .IN0(\r60/CARRYB[22][28] ), 
        .IN1(\r60/SUMB[22][29] ), .COUT(\r60/CARRYB[23][28] ), .SUM(
        \r60/SUMB[23][28] ) );
  FADDER \r60/S2_23_27  ( .CIN(\r60/ab[23][27] ), .IN0(\r60/CARRYB[22][27] ), 
        .IN1(\r60/SUMB[22][28] ), .COUT(\r60/CARRYB[23][27] ), .SUM(
        \r60/SUMB[23][27] ) );
  FADDER \r60/S2_23_26  ( .CIN(\r60/ab[23][26] ), .IN0(\r60/CARRYB[22][26] ), 
        .IN1(\r60/SUMB[22][27] ), .COUT(\r60/CARRYB[23][26] ), .SUM(
        \r60/SUMB[23][26] ) );
  FADDER \r60/S2_23_25  ( .CIN(\r60/ab[23][25] ), .IN0(\r60/CARRYB[22][25] ), 
        .IN1(\r60/SUMB[22][26] ), .COUT(\r60/CARRYB[23][25] ), .SUM(
        \r60/SUMB[23][25] ) );
  FADDER \r60/S2_23_24  ( .CIN(\r60/ab[23][24] ), .IN0(\r60/CARRYB[22][24] ), 
        .IN1(\r60/SUMB[22][25] ), .COUT(\r60/CARRYB[23][24] ), .SUM(
        \r60/SUMB[23][24] ) );
  FADDER \r60/S2_23_23  ( .CIN(\r60/ab[23][23] ), .IN0(\r60/CARRYB[22][23] ), 
        .IN1(\r60/SUMB[22][24] ), .COUT(\r60/CARRYB[23][23] ), .SUM(
        \r60/SUMB[23][23] ) );
  FADDER \r60/S2_23_22  ( .CIN(\r60/ab[23][22] ), .IN0(\r60/CARRYB[22][22] ), 
        .IN1(\r60/SUMB[22][23] ), .COUT(\r60/CARRYB[23][22] ), .SUM(
        \r60/SUMB[23][22] ) );
  FADDER \r60/S2_23_21  ( .CIN(\r60/ab[23][21] ), .IN0(\r60/CARRYB[22][21] ), 
        .IN1(\r60/SUMB[22][22] ), .COUT(\r60/CARRYB[23][21] ), .SUM(
        \r60/SUMB[23][21] ) );
  FADDER \r60/S2_23_20  ( .CIN(\r60/ab[23][20] ), .IN0(\r60/CARRYB[22][20] ), 
        .IN1(\r60/SUMB[22][21] ), .COUT(\r60/CARRYB[23][20] ), .SUM(
        \r60/SUMB[23][20] ) );
  FADDER \r60/S2_23_19  ( .CIN(\r60/ab[23][19] ), .IN0(\r60/CARRYB[22][19] ), 
        .IN1(\r60/SUMB[22][20] ), .COUT(\r60/CARRYB[23][19] ), .SUM(
        \r60/SUMB[23][19] ) );
  FADDER \r60/S2_23_18  ( .CIN(\r60/ab[23][18] ), .IN0(\r60/CARRYB[22][18] ), 
        .IN1(\r60/SUMB[22][19] ), .COUT(\r60/CARRYB[23][18] ), .SUM(
        \r60/SUMB[23][18] ) );
  FADDER \r60/S2_23_17  ( .CIN(\r60/ab[23][17] ), .IN0(\r60/CARRYB[22][17] ), 
        .IN1(\r60/SUMB[22][18] ), .COUT(\r60/CARRYB[23][17] ), .SUM(
        \r60/SUMB[23][17] ) );
  FADDER \r60/S2_23_16  ( .CIN(\r60/ab[23][16] ), .IN0(\r60/CARRYB[22][16] ), 
        .IN1(\r60/SUMB[22][17] ), .COUT(\r60/CARRYB[23][16] ), .SUM(
        \r60/SUMB[23][16] ) );
  FADDER \r60/S2_23_15  ( .CIN(\r60/ab[23][15] ), .IN0(\r60/CARRYB[22][15] ), 
        .IN1(\r60/SUMB[22][16] ), .COUT(\r60/CARRYB[23][15] ), .SUM(
        \r60/SUMB[23][15] ) );
  FADDER \r60/S2_23_14  ( .CIN(\r60/ab[23][14] ), .IN0(\r60/CARRYB[22][14] ), 
        .IN1(\r60/SUMB[22][15] ), .COUT(\r60/CARRYB[23][14] ), .SUM(
        \r60/SUMB[23][14] ) );
  FADDER \r60/S2_23_13  ( .CIN(\r60/ab[23][13] ), .IN0(\r60/CARRYB[22][13] ), 
        .IN1(\r60/SUMB[22][14] ), .COUT(\r60/CARRYB[23][13] ), .SUM(
        \r60/SUMB[23][13] ) );
  FADDER \r60/S2_23_12  ( .CIN(\r60/ab[23][12] ), .IN0(\r60/CARRYB[22][12] ), 
        .IN1(\r60/SUMB[22][13] ), .COUT(\r60/CARRYB[23][12] ), .SUM(
        \r60/SUMB[23][12] ) );
  FADDER \r60/S2_23_11  ( .CIN(\r60/ab[23][11] ), .IN0(\r60/CARRYB[22][11] ), 
        .IN1(\r60/SUMB[22][12] ), .COUT(\r60/CARRYB[23][11] ), .SUM(
        \r60/SUMB[23][11] ) );
  FADDER \r60/S2_23_10  ( .CIN(\r60/ab[23][10] ), .IN0(\r60/CARRYB[22][10] ), 
        .IN1(\r60/SUMB[22][11] ), .COUT(\r60/CARRYB[23][10] ), .SUM(
        \r60/SUMB[23][10] ) );
  FADDER \r60/S2_23_9  ( .CIN(\r60/ab[23][9] ), .IN0(\r60/CARRYB[22][9] ), 
        .IN1(\r60/SUMB[22][10] ), .COUT(\r60/CARRYB[23][9] ), .SUM(
        \r60/SUMB[23][9] ) );
  FADDER \r60/S2_23_8  ( .CIN(\r60/ab[23][8] ), .IN0(\r60/CARRYB[22][8] ), 
        .IN1(\r60/SUMB[22][9] ), .COUT(\r60/CARRYB[23][8] ), .SUM(
        \r60/SUMB[23][8] ) );
  FADDER \r60/S2_23_7  ( .CIN(\r60/ab[23][7] ), .IN0(\r60/CARRYB[22][7] ), 
        .IN1(\r60/SUMB[22][8] ), .COUT(\r60/CARRYB[23][7] ), .SUM(
        \r60/SUMB[23][7] ) );
  FADDER \r60/S2_23_6  ( .CIN(\r60/ab[23][6] ), .IN0(\r60/CARRYB[22][6] ), 
        .IN1(\r60/SUMB[22][7] ), .COUT(\r60/CARRYB[23][6] ), .SUM(
        \r60/SUMB[23][6] ) );
  FADDER \r60/S2_23_5  ( .CIN(\r60/ab[23][5] ), .IN0(\r60/CARRYB[22][5] ), 
        .IN1(\r60/SUMB[22][6] ), .COUT(\r60/CARRYB[23][5] ), .SUM(
        \r60/SUMB[23][5] ) );
  FADDER \r60/S2_23_4  ( .CIN(\r60/ab[23][4] ), .IN0(\r60/CARRYB[22][4] ), 
        .IN1(\r60/SUMB[22][5] ), .COUT(\r60/CARRYB[23][4] ), .SUM(
        \r60/SUMB[23][4] ) );
  FADDER \r60/S2_23_3  ( .CIN(\r60/ab[23][3] ), .IN0(\r60/CARRYB[22][3] ), 
        .IN1(\r60/SUMB[22][4] ), .COUT(\r60/CARRYB[23][3] ), .SUM(
        \r60/SUMB[23][3] ) );
  FADDER \r60/S2_23_2  ( .CIN(\r60/ab[23][2] ), .IN0(\r60/CARRYB[22][2] ), 
        .IN1(\r60/SUMB[22][3] ), .COUT(\r60/CARRYB[23][2] ), .SUM(
        \r60/SUMB[23][2] ) );
  FADDER \r60/S2_23_1  ( .CIN(\r60/ab[23][1] ), .IN0(\r60/CARRYB[22][1] ), 
        .IN1(\r60/SUMB[22][2] ), .COUT(\r60/CARRYB[23][1] ), .SUM(
        \r60/SUMB[23][1] ) );
  FADDER \r60/S1_23_0  ( .CIN(\r60/ab[23][0] ), .IN0(\r60/CARRYB[22][0] ), 
        .IN1(\r60/SUMB[22][1] ), .COUT(\r60/CARRYB[23][0] ), .SUM(N140) );
  FADDER \r60/S3_24_30  ( .CIN(\r60/ab[24][30] ), .IN0(\r60/CARRYB[23][30] ), 
        .IN1(\r60/ab[23][31] ), .COUT(\r60/CARRYB[24][30] ), .SUM(
        \r60/SUMB[24][30] ) );
  FADDER \r60/S2_24_29  ( .CIN(\r60/ab[24][29] ), .IN0(\r60/CARRYB[23][29] ), 
        .IN1(\r60/SUMB[23][30] ), .COUT(\r60/CARRYB[24][29] ), .SUM(
        \r60/SUMB[24][29] ) );
  FADDER \r60/S2_24_28  ( .CIN(\r60/ab[24][28] ), .IN0(\r60/CARRYB[23][28] ), 
        .IN1(\r60/SUMB[23][29] ), .COUT(\r60/CARRYB[24][28] ), .SUM(
        \r60/SUMB[24][28] ) );
  FADDER \r60/S2_24_27  ( .CIN(\r60/ab[24][27] ), .IN0(\r60/CARRYB[23][27] ), 
        .IN1(\r60/SUMB[23][28] ), .COUT(\r60/CARRYB[24][27] ), .SUM(
        \r60/SUMB[24][27] ) );
  FADDER \r60/S2_24_26  ( .CIN(\r60/ab[24][26] ), .IN0(\r60/CARRYB[23][26] ), 
        .IN1(\r60/SUMB[23][27] ), .COUT(\r60/CARRYB[24][26] ), .SUM(
        \r60/SUMB[24][26] ) );
  FADDER \r60/S2_24_25  ( .CIN(\r60/ab[24][25] ), .IN0(\r60/CARRYB[23][25] ), 
        .IN1(\r60/SUMB[23][26] ), .COUT(\r60/CARRYB[24][25] ), .SUM(
        \r60/SUMB[24][25] ) );
  FADDER \r60/S2_24_24  ( .CIN(\r60/ab[24][24] ), .IN0(\r60/CARRYB[23][24] ), 
        .IN1(\r60/SUMB[23][25] ), .COUT(\r60/CARRYB[24][24] ), .SUM(
        \r60/SUMB[24][24] ) );
  FADDER \r60/S2_24_23  ( .CIN(\r60/ab[24][23] ), .IN0(\r60/CARRYB[23][23] ), 
        .IN1(\r60/SUMB[23][24] ), .COUT(\r60/CARRYB[24][23] ), .SUM(
        \r60/SUMB[24][23] ) );
  FADDER \r60/S2_24_22  ( .CIN(\r60/ab[24][22] ), .IN0(\r60/CARRYB[23][22] ), 
        .IN1(\r60/SUMB[23][23] ), .COUT(\r60/CARRYB[24][22] ), .SUM(
        \r60/SUMB[24][22] ) );
  FADDER \r60/S2_24_21  ( .CIN(\r60/ab[24][21] ), .IN0(\r60/CARRYB[23][21] ), 
        .IN1(\r60/SUMB[23][22] ), .COUT(\r60/CARRYB[24][21] ), .SUM(
        \r60/SUMB[24][21] ) );
  FADDER \r60/S2_24_20  ( .CIN(\r60/ab[24][20] ), .IN0(\r60/CARRYB[23][20] ), 
        .IN1(\r60/SUMB[23][21] ), .COUT(\r60/CARRYB[24][20] ), .SUM(
        \r60/SUMB[24][20] ) );
  FADDER \r60/S2_24_19  ( .CIN(\r60/ab[24][19] ), .IN0(\r60/CARRYB[23][19] ), 
        .IN1(\r60/SUMB[23][20] ), .COUT(\r60/CARRYB[24][19] ), .SUM(
        \r60/SUMB[24][19] ) );
  FADDER \r60/S2_24_18  ( .CIN(\r60/ab[24][18] ), .IN0(\r60/CARRYB[23][18] ), 
        .IN1(\r60/SUMB[23][19] ), .COUT(\r60/CARRYB[24][18] ), .SUM(
        \r60/SUMB[24][18] ) );
  FADDER \r60/S2_24_17  ( .CIN(\r60/ab[24][17] ), .IN0(\r60/CARRYB[23][17] ), 
        .IN1(\r60/SUMB[23][18] ), .COUT(\r60/CARRYB[24][17] ), .SUM(
        \r60/SUMB[24][17] ) );
  FADDER \r60/S2_24_16  ( .CIN(\r60/ab[24][16] ), .IN0(\r60/CARRYB[23][16] ), 
        .IN1(\r60/SUMB[23][17] ), .COUT(\r60/CARRYB[24][16] ), .SUM(
        \r60/SUMB[24][16] ) );
  FADDER \r60/S2_24_15  ( .CIN(\r60/ab[24][15] ), .IN0(\r60/CARRYB[23][15] ), 
        .IN1(\r60/SUMB[23][16] ), .COUT(\r60/CARRYB[24][15] ), .SUM(
        \r60/SUMB[24][15] ) );
  FADDER \r60/S2_24_14  ( .CIN(\r60/ab[24][14] ), .IN0(\r60/CARRYB[23][14] ), 
        .IN1(\r60/SUMB[23][15] ), .COUT(\r60/CARRYB[24][14] ), .SUM(
        \r60/SUMB[24][14] ) );
  FADDER \r60/S2_24_13  ( .CIN(\r60/ab[24][13] ), .IN0(\r60/CARRYB[23][13] ), 
        .IN1(\r60/SUMB[23][14] ), .COUT(\r60/CARRYB[24][13] ), .SUM(
        \r60/SUMB[24][13] ) );
  FADDER \r60/S2_24_12  ( .CIN(\r60/ab[24][12] ), .IN0(\r60/CARRYB[23][12] ), 
        .IN1(\r60/SUMB[23][13] ), .COUT(\r60/CARRYB[24][12] ), .SUM(
        \r60/SUMB[24][12] ) );
  FADDER \r60/S2_24_11  ( .CIN(\r60/ab[24][11] ), .IN0(\r60/CARRYB[23][11] ), 
        .IN1(\r60/SUMB[23][12] ), .COUT(\r60/CARRYB[24][11] ), .SUM(
        \r60/SUMB[24][11] ) );
  FADDER \r60/S2_24_10  ( .CIN(\r60/ab[24][10] ), .IN0(\r60/CARRYB[23][10] ), 
        .IN1(\r60/SUMB[23][11] ), .COUT(\r60/CARRYB[24][10] ), .SUM(
        \r60/SUMB[24][10] ) );
  FADDER \r60/S2_24_9  ( .CIN(\r60/ab[24][9] ), .IN0(\r60/CARRYB[23][9] ), 
        .IN1(\r60/SUMB[23][10] ), .COUT(\r60/CARRYB[24][9] ), .SUM(
        \r60/SUMB[24][9] ) );
  FADDER \r60/S2_24_8  ( .CIN(\r60/ab[24][8] ), .IN0(\r60/CARRYB[23][8] ), 
        .IN1(\r60/SUMB[23][9] ), .COUT(\r60/CARRYB[24][8] ), .SUM(
        \r60/SUMB[24][8] ) );
  FADDER \r60/S2_24_7  ( .CIN(\r60/ab[24][7] ), .IN0(\r60/CARRYB[23][7] ), 
        .IN1(\r60/SUMB[23][8] ), .COUT(\r60/CARRYB[24][7] ), .SUM(
        \r60/SUMB[24][7] ) );
  FADDER \r60/S2_24_6  ( .CIN(\r60/ab[24][6] ), .IN0(\r60/CARRYB[23][6] ), 
        .IN1(\r60/SUMB[23][7] ), .COUT(\r60/CARRYB[24][6] ), .SUM(
        \r60/SUMB[24][6] ) );
  FADDER \r60/S2_24_5  ( .CIN(\r60/ab[24][5] ), .IN0(\r60/CARRYB[23][5] ), 
        .IN1(\r60/SUMB[23][6] ), .COUT(\r60/CARRYB[24][5] ), .SUM(
        \r60/SUMB[24][5] ) );
  FADDER \r60/S2_24_4  ( .CIN(\r60/ab[24][4] ), .IN0(\r60/CARRYB[23][4] ), 
        .IN1(\r60/SUMB[23][5] ), .COUT(\r60/CARRYB[24][4] ), .SUM(
        \r60/SUMB[24][4] ) );
  FADDER \r60/S2_24_3  ( .CIN(\r60/ab[24][3] ), .IN0(\r60/CARRYB[23][3] ), 
        .IN1(\r60/SUMB[23][4] ), .COUT(\r60/CARRYB[24][3] ), .SUM(
        \r60/SUMB[24][3] ) );
  FADDER \r60/S2_24_2  ( .CIN(\r60/ab[24][2] ), .IN0(\r60/CARRYB[23][2] ), 
        .IN1(\r60/SUMB[23][3] ), .COUT(\r60/CARRYB[24][2] ), .SUM(
        \r60/SUMB[24][2] ) );
  FADDER \r60/S2_24_1  ( .CIN(\r60/ab[24][1] ), .IN0(\r60/CARRYB[23][1] ), 
        .IN1(\r60/SUMB[23][2] ), .COUT(\r60/CARRYB[24][1] ), .SUM(
        \r60/SUMB[24][1] ) );
  FADDER \r60/S1_24_0  ( .CIN(\r60/ab[24][0] ), .IN0(\r60/CARRYB[23][0] ), 
        .IN1(\r60/SUMB[23][1] ), .COUT(\r60/CARRYB[24][0] ), .SUM(N141) );
  FADDER \r60/S3_25_30  ( .CIN(\r60/ab[25][30] ), .IN0(\r60/CARRYB[24][30] ), 
        .IN1(\r60/ab[24][31] ), .COUT(\r60/CARRYB[25][30] ), .SUM(
        \r60/SUMB[25][30] ) );
  FADDER \r60/S2_25_29  ( .CIN(\r60/ab[25][29] ), .IN0(\r60/CARRYB[24][29] ), 
        .IN1(\r60/SUMB[24][30] ), .COUT(\r60/CARRYB[25][29] ), .SUM(
        \r60/SUMB[25][29] ) );
  FADDER \r60/S2_25_28  ( .CIN(\r60/ab[25][28] ), .IN0(\r60/CARRYB[24][28] ), 
        .IN1(\r60/SUMB[24][29] ), .COUT(\r60/CARRYB[25][28] ), .SUM(
        \r60/SUMB[25][28] ) );
  FADDER \r60/S2_25_27  ( .CIN(\r60/ab[25][27] ), .IN0(\r60/CARRYB[24][27] ), 
        .IN1(\r60/SUMB[24][28] ), .COUT(\r60/CARRYB[25][27] ), .SUM(
        \r60/SUMB[25][27] ) );
  FADDER \r60/S2_25_26  ( .CIN(\r60/ab[25][26] ), .IN0(\r60/CARRYB[24][26] ), 
        .IN1(\r60/SUMB[24][27] ), .COUT(\r60/CARRYB[25][26] ), .SUM(
        \r60/SUMB[25][26] ) );
  FADDER \r60/S2_25_25  ( .CIN(\r60/ab[25][25] ), .IN0(\r60/CARRYB[24][25] ), 
        .IN1(\r60/SUMB[24][26] ), .COUT(\r60/CARRYB[25][25] ), .SUM(
        \r60/SUMB[25][25] ) );
  FADDER \r60/S2_25_24  ( .CIN(\r60/ab[25][24] ), .IN0(\r60/CARRYB[24][24] ), 
        .IN1(\r60/SUMB[24][25] ), .COUT(\r60/CARRYB[25][24] ), .SUM(
        \r60/SUMB[25][24] ) );
  FADDER \r60/S2_25_23  ( .CIN(\r60/ab[25][23] ), .IN0(\r60/CARRYB[24][23] ), 
        .IN1(\r60/SUMB[24][24] ), .COUT(\r60/CARRYB[25][23] ), .SUM(
        \r60/SUMB[25][23] ) );
  FADDER \r60/S2_25_22  ( .CIN(\r60/ab[25][22] ), .IN0(\r60/CARRYB[24][22] ), 
        .IN1(\r60/SUMB[24][23] ), .COUT(\r60/CARRYB[25][22] ), .SUM(
        \r60/SUMB[25][22] ) );
  FADDER \r60/S2_25_21  ( .CIN(\r60/ab[25][21] ), .IN0(\r60/CARRYB[24][21] ), 
        .IN1(\r60/SUMB[24][22] ), .COUT(\r60/CARRYB[25][21] ), .SUM(
        \r60/SUMB[25][21] ) );
  FADDER \r60/S2_25_20  ( .CIN(\r60/ab[25][20] ), .IN0(\r60/CARRYB[24][20] ), 
        .IN1(\r60/SUMB[24][21] ), .COUT(\r60/CARRYB[25][20] ), .SUM(
        \r60/SUMB[25][20] ) );
  FADDER \r60/S2_25_19  ( .CIN(\r60/ab[25][19] ), .IN0(\r60/CARRYB[24][19] ), 
        .IN1(\r60/SUMB[24][20] ), .COUT(\r60/CARRYB[25][19] ), .SUM(
        \r60/SUMB[25][19] ) );
  FADDER \r60/S2_25_18  ( .CIN(\r60/ab[25][18] ), .IN0(\r60/CARRYB[24][18] ), 
        .IN1(\r60/SUMB[24][19] ), .COUT(\r60/CARRYB[25][18] ), .SUM(
        \r60/SUMB[25][18] ) );
  FADDER \r60/S2_25_17  ( .CIN(\r60/ab[25][17] ), .IN0(\r60/CARRYB[24][17] ), 
        .IN1(\r60/SUMB[24][18] ), .COUT(\r60/CARRYB[25][17] ), .SUM(
        \r60/SUMB[25][17] ) );
  FADDER \r60/S2_25_16  ( .CIN(\r60/ab[25][16] ), .IN0(\r60/CARRYB[24][16] ), 
        .IN1(\r60/SUMB[24][17] ), .COUT(\r60/CARRYB[25][16] ), .SUM(
        \r60/SUMB[25][16] ) );
  FADDER \r60/S2_25_15  ( .CIN(\r60/ab[25][15] ), .IN0(\r60/CARRYB[24][15] ), 
        .IN1(\r60/SUMB[24][16] ), .COUT(\r60/CARRYB[25][15] ), .SUM(
        \r60/SUMB[25][15] ) );
  FADDER \r60/S2_25_14  ( .CIN(\r60/ab[25][14] ), .IN0(\r60/CARRYB[24][14] ), 
        .IN1(\r60/SUMB[24][15] ), .COUT(\r60/CARRYB[25][14] ), .SUM(
        \r60/SUMB[25][14] ) );
  FADDER \r60/S2_25_13  ( .CIN(\r60/ab[25][13] ), .IN0(\r60/CARRYB[24][13] ), 
        .IN1(\r60/SUMB[24][14] ), .COUT(\r60/CARRYB[25][13] ), .SUM(
        \r60/SUMB[25][13] ) );
  FADDER \r60/S2_25_12  ( .CIN(\r60/ab[25][12] ), .IN0(\r60/CARRYB[24][12] ), 
        .IN1(\r60/SUMB[24][13] ), .COUT(\r60/CARRYB[25][12] ), .SUM(
        \r60/SUMB[25][12] ) );
  FADDER \r60/S2_25_11  ( .CIN(\r60/ab[25][11] ), .IN0(\r60/CARRYB[24][11] ), 
        .IN1(\r60/SUMB[24][12] ), .COUT(\r60/CARRYB[25][11] ), .SUM(
        \r60/SUMB[25][11] ) );
  FADDER \r60/S2_25_10  ( .CIN(\r60/ab[25][10] ), .IN0(\r60/CARRYB[24][10] ), 
        .IN1(\r60/SUMB[24][11] ), .COUT(\r60/CARRYB[25][10] ), .SUM(
        \r60/SUMB[25][10] ) );
  FADDER \r60/S2_25_9  ( .CIN(\r60/ab[25][9] ), .IN0(\r60/CARRYB[24][9] ), 
        .IN1(\r60/SUMB[24][10] ), .COUT(\r60/CARRYB[25][9] ), .SUM(
        \r60/SUMB[25][9] ) );
  FADDER \r60/S2_25_8  ( .CIN(\r60/ab[25][8] ), .IN0(\r60/CARRYB[24][8] ), 
        .IN1(\r60/SUMB[24][9] ), .COUT(\r60/CARRYB[25][8] ), .SUM(
        \r60/SUMB[25][8] ) );
  FADDER \r60/S2_25_7  ( .CIN(\r60/ab[25][7] ), .IN0(\r60/CARRYB[24][7] ), 
        .IN1(\r60/SUMB[24][8] ), .COUT(\r60/CARRYB[25][7] ), .SUM(
        \r60/SUMB[25][7] ) );
  FADDER \r60/S2_25_6  ( .CIN(\r60/ab[25][6] ), .IN0(\r60/CARRYB[24][6] ), 
        .IN1(\r60/SUMB[24][7] ), .COUT(\r60/CARRYB[25][6] ), .SUM(
        \r60/SUMB[25][6] ) );
  FADDER \r60/S2_25_5  ( .CIN(\r60/ab[25][5] ), .IN0(\r60/CARRYB[24][5] ), 
        .IN1(\r60/SUMB[24][6] ), .COUT(\r60/CARRYB[25][5] ), .SUM(
        \r60/SUMB[25][5] ) );
  FADDER \r60/S2_25_4  ( .CIN(\r60/ab[25][4] ), .IN0(\r60/CARRYB[24][4] ), 
        .IN1(\r60/SUMB[24][5] ), .COUT(\r60/CARRYB[25][4] ), .SUM(
        \r60/SUMB[25][4] ) );
  FADDER \r60/S2_25_3  ( .CIN(\r60/ab[25][3] ), .IN0(\r60/CARRYB[24][3] ), 
        .IN1(\r60/SUMB[24][4] ), .COUT(\r60/CARRYB[25][3] ), .SUM(
        \r60/SUMB[25][3] ) );
  FADDER \r60/S2_25_2  ( .CIN(\r60/ab[25][2] ), .IN0(\r60/CARRYB[24][2] ), 
        .IN1(\r60/SUMB[24][3] ), .COUT(\r60/CARRYB[25][2] ), .SUM(
        \r60/SUMB[25][2] ) );
  FADDER \r60/S2_25_1  ( .CIN(\r60/ab[25][1] ), .IN0(\r60/CARRYB[24][1] ), 
        .IN1(\r60/SUMB[24][2] ), .COUT(\r60/CARRYB[25][1] ), .SUM(
        \r60/SUMB[25][1] ) );
  FADDER \r60/S1_25_0  ( .CIN(\r60/ab[25][0] ), .IN0(\r60/CARRYB[24][0] ), 
        .IN1(\r60/SUMB[24][1] ), .COUT(\r60/CARRYB[25][0] ), .SUM(N142) );
  FADDER \r60/S3_26_30  ( .CIN(\r60/ab[26][30] ), .IN0(\r60/CARRYB[25][30] ), 
        .IN1(\r60/ab[25][31] ), .COUT(\r60/CARRYB[26][30] ), .SUM(
        \r60/SUMB[26][30] ) );
  FADDER \r60/S2_26_29  ( .CIN(\r60/ab[26][29] ), .IN0(\r60/CARRYB[25][29] ), 
        .IN1(\r60/SUMB[25][30] ), .COUT(\r60/CARRYB[26][29] ), .SUM(
        \r60/SUMB[26][29] ) );
  FADDER \r60/S2_26_28  ( .CIN(\r60/ab[26][28] ), .IN0(\r60/CARRYB[25][28] ), 
        .IN1(\r60/SUMB[25][29] ), .COUT(\r60/CARRYB[26][28] ), .SUM(
        \r60/SUMB[26][28] ) );
  FADDER \r60/S2_26_27  ( .CIN(\r60/ab[26][27] ), .IN0(\r60/CARRYB[25][27] ), 
        .IN1(\r60/SUMB[25][28] ), .COUT(\r60/CARRYB[26][27] ), .SUM(
        \r60/SUMB[26][27] ) );
  FADDER \r60/S2_26_26  ( .CIN(\r60/ab[26][26] ), .IN0(\r60/CARRYB[25][26] ), 
        .IN1(\r60/SUMB[25][27] ), .COUT(\r60/CARRYB[26][26] ), .SUM(
        \r60/SUMB[26][26] ) );
  FADDER \r60/S2_26_25  ( .CIN(\r60/ab[26][25] ), .IN0(\r60/CARRYB[25][25] ), 
        .IN1(\r60/SUMB[25][26] ), .COUT(\r60/CARRYB[26][25] ), .SUM(
        \r60/SUMB[26][25] ) );
  FADDER \r60/S2_26_24  ( .CIN(\r60/ab[26][24] ), .IN0(\r60/CARRYB[25][24] ), 
        .IN1(\r60/SUMB[25][25] ), .COUT(\r60/CARRYB[26][24] ), .SUM(
        \r60/SUMB[26][24] ) );
  FADDER \r60/S2_26_23  ( .CIN(\r60/ab[26][23] ), .IN0(\r60/CARRYB[25][23] ), 
        .IN1(\r60/SUMB[25][24] ), .COUT(\r60/CARRYB[26][23] ), .SUM(
        \r60/SUMB[26][23] ) );
  FADDER \r60/S2_26_22  ( .CIN(\r60/ab[26][22] ), .IN0(\r60/CARRYB[25][22] ), 
        .IN1(\r60/SUMB[25][23] ), .COUT(\r60/CARRYB[26][22] ), .SUM(
        \r60/SUMB[26][22] ) );
  FADDER \r60/S2_26_21  ( .CIN(\r60/ab[26][21] ), .IN0(\r60/CARRYB[25][21] ), 
        .IN1(\r60/SUMB[25][22] ), .COUT(\r60/CARRYB[26][21] ), .SUM(
        \r60/SUMB[26][21] ) );
  FADDER \r60/S2_26_20  ( .CIN(\r60/ab[26][20] ), .IN0(\r60/CARRYB[25][20] ), 
        .IN1(\r60/SUMB[25][21] ), .COUT(\r60/CARRYB[26][20] ), .SUM(
        \r60/SUMB[26][20] ) );
  FADDER \r60/S2_26_19  ( .CIN(\r60/ab[26][19] ), .IN0(\r60/CARRYB[25][19] ), 
        .IN1(\r60/SUMB[25][20] ), .COUT(\r60/CARRYB[26][19] ), .SUM(
        \r60/SUMB[26][19] ) );
  FADDER \r60/S2_26_18  ( .CIN(\r60/ab[26][18] ), .IN0(\r60/CARRYB[25][18] ), 
        .IN1(\r60/SUMB[25][19] ), .COUT(\r60/CARRYB[26][18] ), .SUM(
        \r60/SUMB[26][18] ) );
  FADDER \r60/S2_26_17  ( .CIN(\r60/ab[26][17] ), .IN0(\r60/CARRYB[25][17] ), 
        .IN1(\r60/SUMB[25][18] ), .COUT(\r60/CARRYB[26][17] ), .SUM(
        \r60/SUMB[26][17] ) );
  FADDER \r60/S2_26_16  ( .CIN(\r60/ab[26][16] ), .IN0(\r60/CARRYB[25][16] ), 
        .IN1(\r60/SUMB[25][17] ), .COUT(\r60/CARRYB[26][16] ), .SUM(
        \r60/SUMB[26][16] ) );
  FADDER \r60/S2_26_15  ( .CIN(\r60/ab[26][15] ), .IN0(\r60/CARRYB[25][15] ), 
        .IN1(\r60/SUMB[25][16] ), .COUT(\r60/CARRYB[26][15] ), .SUM(
        \r60/SUMB[26][15] ) );
  FADDER \r60/S2_26_14  ( .CIN(\r60/ab[26][14] ), .IN0(\r60/CARRYB[25][14] ), 
        .IN1(\r60/SUMB[25][15] ), .COUT(\r60/CARRYB[26][14] ), .SUM(
        \r60/SUMB[26][14] ) );
  FADDER \r60/S2_26_13  ( .CIN(\r60/ab[26][13] ), .IN0(\r60/CARRYB[25][13] ), 
        .IN1(\r60/SUMB[25][14] ), .COUT(\r60/CARRYB[26][13] ), .SUM(
        \r60/SUMB[26][13] ) );
  FADDER \r60/S2_26_12  ( .CIN(\r60/ab[26][12] ), .IN0(\r60/CARRYB[25][12] ), 
        .IN1(\r60/SUMB[25][13] ), .COUT(\r60/CARRYB[26][12] ), .SUM(
        \r60/SUMB[26][12] ) );
  FADDER \r60/S2_26_11  ( .CIN(\r60/ab[26][11] ), .IN0(\r60/CARRYB[25][11] ), 
        .IN1(\r60/SUMB[25][12] ), .COUT(\r60/CARRYB[26][11] ), .SUM(
        \r60/SUMB[26][11] ) );
  FADDER \r60/S2_26_10  ( .CIN(\r60/ab[26][10] ), .IN0(\r60/CARRYB[25][10] ), 
        .IN1(\r60/SUMB[25][11] ), .COUT(\r60/CARRYB[26][10] ), .SUM(
        \r60/SUMB[26][10] ) );
  FADDER \r60/S2_26_9  ( .CIN(\r60/ab[26][9] ), .IN0(\r60/CARRYB[25][9] ), 
        .IN1(\r60/SUMB[25][10] ), .COUT(\r60/CARRYB[26][9] ), .SUM(
        \r60/SUMB[26][9] ) );
  FADDER \r60/S2_26_8  ( .CIN(\r60/ab[26][8] ), .IN0(\r60/CARRYB[25][8] ), 
        .IN1(\r60/SUMB[25][9] ), .COUT(\r60/CARRYB[26][8] ), .SUM(
        \r60/SUMB[26][8] ) );
  FADDER \r60/S2_26_7  ( .CIN(\r60/ab[26][7] ), .IN0(\r60/CARRYB[25][7] ), 
        .IN1(\r60/SUMB[25][8] ), .COUT(\r60/CARRYB[26][7] ), .SUM(
        \r60/SUMB[26][7] ) );
  FADDER \r60/S2_26_6  ( .CIN(\r60/ab[26][6] ), .IN0(\r60/CARRYB[25][6] ), 
        .IN1(\r60/SUMB[25][7] ), .COUT(\r60/CARRYB[26][6] ), .SUM(
        \r60/SUMB[26][6] ) );
  FADDER \r60/S2_26_5  ( .CIN(\r60/ab[26][5] ), .IN0(\r60/CARRYB[25][5] ), 
        .IN1(\r60/SUMB[25][6] ), .COUT(\r60/CARRYB[26][5] ), .SUM(
        \r60/SUMB[26][5] ) );
  FADDER \r60/S2_26_4  ( .CIN(\r60/ab[26][4] ), .IN0(\r60/CARRYB[25][4] ), 
        .IN1(\r60/SUMB[25][5] ), .COUT(\r60/CARRYB[26][4] ), .SUM(
        \r60/SUMB[26][4] ) );
  FADDER \r60/S2_26_3  ( .CIN(\r60/ab[26][3] ), .IN0(\r60/CARRYB[25][3] ), 
        .IN1(\r60/SUMB[25][4] ), .COUT(\r60/CARRYB[26][3] ), .SUM(
        \r60/SUMB[26][3] ) );
  FADDER \r60/S2_26_2  ( .CIN(\r60/ab[26][2] ), .IN0(\r60/CARRYB[25][2] ), 
        .IN1(\r60/SUMB[25][3] ), .COUT(\r60/CARRYB[26][2] ), .SUM(
        \r60/SUMB[26][2] ) );
  FADDER \r60/S2_26_1  ( .CIN(\r60/ab[26][1] ), .IN0(\r60/CARRYB[25][1] ), 
        .IN1(\r60/SUMB[25][2] ), .COUT(\r60/CARRYB[26][1] ), .SUM(
        \r60/SUMB[26][1] ) );
  FADDER \r60/S1_26_0  ( .CIN(\r60/ab[26][0] ), .IN0(\r60/CARRYB[25][0] ), 
        .IN1(\r60/SUMB[25][1] ), .COUT(\r60/CARRYB[26][0] ), .SUM(N143) );
  FADDER \r60/S3_27_30  ( .CIN(\r60/ab[27][30] ), .IN0(\r60/CARRYB[26][30] ), 
        .IN1(\r60/ab[26][31] ), .COUT(\r60/CARRYB[27][30] ), .SUM(
        \r60/SUMB[27][30] ) );
  FADDER \r60/S2_27_29  ( .CIN(\r60/ab[27][29] ), .IN0(\r60/CARRYB[26][29] ), 
        .IN1(\r60/SUMB[26][30] ), .COUT(\r60/CARRYB[27][29] ), .SUM(
        \r60/SUMB[27][29] ) );
  FADDER \r60/S2_27_28  ( .CIN(\r60/ab[27][28] ), .IN0(\r60/CARRYB[26][28] ), 
        .IN1(\r60/SUMB[26][29] ), .COUT(\r60/CARRYB[27][28] ), .SUM(
        \r60/SUMB[27][28] ) );
  FADDER \r60/S2_27_27  ( .CIN(\r60/ab[27][27] ), .IN0(\r60/CARRYB[26][27] ), 
        .IN1(\r60/SUMB[26][28] ), .COUT(\r60/CARRYB[27][27] ), .SUM(
        \r60/SUMB[27][27] ) );
  FADDER \r60/S2_27_26  ( .CIN(\r60/ab[27][26] ), .IN0(\r60/CARRYB[26][26] ), 
        .IN1(\r60/SUMB[26][27] ), .COUT(\r60/CARRYB[27][26] ), .SUM(
        \r60/SUMB[27][26] ) );
  FADDER \r60/S2_27_25  ( .CIN(\r60/ab[27][25] ), .IN0(\r60/CARRYB[26][25] ), 
        .IN1(\r60/SUMB[26][26] ), .COUT(\r60/CARRYB[27][25] ), .SUM(
        \r60/SUMB[27][25] ) );
  FADDER \r60/S2_27_24  ( .CIN(\r60/ab[27][24] ), .IN0(\r60/CARRYB[26][24] ), 
        .IN1(\r60/SUMB[26][25] ), .COUT(\r60/CARRYB[27][24] ), .SUM(
        \r60/SUMB[27][24] ) );
  FADDER \r60/S2_27_23  ( .CIN(\r60/ab[27][23] ), .IN0(\r60/CARRYB[26][23] ), 
        .IN1(\r60/SUMB[26][24] ), .COUT(\r60/CARRYB[27][23] ), .SUM(
        \r60/SUMB[27][23] ) );
  FADDER \r60/S2_27_22  ( .CIN(\r60/ab[27][22] ), .IN0(\r60/CARRYB[26][22] ), 
        .IN1(\r60/SUMB[26][23] ), .COUT(\r60/CARRYB[27][22] ), .SUM(
        \r60/SUMB[27][22] ) );
  FADDER \r60/S2_27_21  ( .CIN(\r60/ab[27][21] ), .IN0(\r60/CARRYB[26][21] ), 
        .IN1(\r60/SUMB[26][22] ), .COUT(\r60/CARRYB[27][21] ), .SUM(
        \r60/SUMB[27][21] ) );
  FADDER \r60/S2_27_20  ( .CIN(\r60/ab[27][20] ), .IN0(\r60/CARRYB[26][20] ), 
        .IN1(\r60/SUMB[26][21] ), .COUT(\r60/CARRYB[27][20] ), .SUM(
        \r60/SUMB[27][20] ) );
  FADDER \r60/S2_27_19  ( .CIN(\r60/ab[27][19] ), .IN0(\r60/CARRYB[26][19] ), 
        .IN1(\r60/SUMB[26][20] ), .COUT(\r60/CARRYB[27][19] ), .SUM(
        \r60/SUMB[27][19] ) );
  FADDER \r60/S2_27_18  ( .CIN(\r60/ab[27][18] ), .IN0(\r60/CARRYB[26][18] ), 
        .IN1(\r60/SUMB[26][19] ), .COUT(\r60/CARRYB[27][18] ), .SUM(
        \r60/SUMB[27][18] ) );
  FADDER \r60/S2_27_17  ( .CIN(\r60/ab[27][17] ), .IN0(\r60/CARRYB[26][17] ), 
        .IN1(\r60/SUMB[26][18] ), .COUT(\r60/CARRYB[27][17] ), .SUM(
        \r60/SUMB[27][17] ) );
  FADDER \r60/S2_27_16  ( .CIN(\r60/ab[27][16] ), .IN0(\r60/CARRYB[26][16] ), 
        .IN1(\r60/SUMB[26][17] ), .COUT(\r60/CARRYB[27][16] ), .SUM(
        \r60/SUMB[27][16] ) );
  FADDER \r60/S2_27_15  ( .CIN(\r60/ab[27][15] ), .IN0(\r60/CARRYB[26][15] ), 
        .IN1(\r60/SUMB[26][16] ), .COUT(\r60/CARRYB[27][15] ), .SUM(
        \r60/SUMB[27][15] ) );
  FADDER \r60/S2_27_14  ( .CIN(\r60/ab[27][14] ), .IN0(\r60/CARRYB[26][14] ), 
        .IN1(\r60/SUMB[26][15] ), .COUT(\r60/CARRYB[27][14] ), .SUM(
        \r60/SUMB[27][14] ) );
  FADDER \r60/S2_27_13  ( .CIN(\r60/ab[27][13] ), .IN0(\r60/CARRYB[26][13] ), 
        .IN1(\r60/SUMB[26][14] ), .COUT(\r60/CARRYB[27][13] ), .SUM(
        \r60/SUMB[27][13] ) );
  FADDER \r60/S2_27_12  ( .CIN(\r60/ab[27][12] ), .IN0(\r60/CARRYB[26][12] ), 
        .IN1(\r60/SUMB[26][13] ), .COUT(\r60/CARRYB[27][12] ), .SUM(
        \r60/SUMB[27][12] ) );
  FADDER \r60/S2_27_11  ( .CIN(\r60/ab[27][11] ), .IN0(\r60/CARRYB[26][11] ), 
        .IN1(\r60/SUMB[26][12] ), .COUT(\r60/CARRYB[27][11] ), .SUM(
        \r60/SUMB[27][11] ) );
  FADDER \r60/S2_27_10  ( .CIN(\r60/ab[27][10] ), .IN0(\r60/CARRYB[26][10] ), 
        .IN1(\r60/SUMB[26][11] ), .COUT(\r60/CARRYB[27][10] ), .SUM(
        \r60/SUMB[27][10] ) );
  FADDER \r60/S2_27_9  ( .CIN(\r60/ab[27][9] ), .IN0(\r60/CARRYB[26][9] ), 
        .IN1(\r60/SUMB[26][10] ), .COUT(\r60/CARRYB[27][9] ), .SUM(
        \r60/SUMB[27][9] ) );
  FADDER \r60/S2_27_8  ( .CIN(\r60/ab[27][8] ), .IN0(\r60/CARRYB[26][8] ), 
        .IN1(\r60/SUMB[26][9] ), .COUT(\r60/CARRYB[27][8] ), .SUM(
        \r60/SUMB[27][8] ) );
  FADDER \r60/S2_27_7  ( .CIN(\r60/ab[27][7] ), .IN0(\r60/CARRYB[26][7] ), 
        .IN1(\r60/SUMB[26][8] ), .COUT(\r60/CARRYB[27][7] ), .SUM(
        \r60/SUMB[27][7] ) );
  FADDER \r60/S2_27_6  ( .CIN(\r60/ab[27][6] ), .IN0(\r60/CARRYB[26][6] ), 
        .IN1(\r60/SUMB[26][7] ), .COUT(\r60/CARRYB[27][6] ), .SUM(
        \r60/SUMB[27][6] ) );
  FADDER \r60/S2_27_5  ( .CIN(\r60/ab[27][5] ), .IN0(\r60/CARRYB[26][5] ), 
        .IN1(\r60/SUMB[26][6] ), .COUT(\r60/CARRYB[27][5] ), .SUM(
        \r60/SUMB[27][5] ) );
  FADDER \r60/S2_27_4  ( .CIN(\r60/ab[27][4] ), .IN0(\r60/CARRYB[26][4] ), 
        .IN1(\r60/SUMB[26][5] ), .COUT(\r60/CARRYB[27][4] ), .SUM(
        \r60/SUMB[27][4] ) );
  FADDER \r60/S2_27_3  ( .CIN(\r60/ab[27][3] ), .IN0(\r60/CARRYB[26][3] ), 
        .IN1(\r60/SUMB[26][4] ), .COUT(\r60/CARRYB[27][3] ), .SUM(
        \r60/SUMB[27][3] ) );
  FADDER \r60/S2_27_2  ( .CIN(\r60/ab[27][2] ), .IN0(\r60/CARRYB[26][2] ), 
        .IN1(\r60/SUMB[26][3] ), .COUT(\r60/CARRYB[27][2] ), .SUM(
        \r60/SUMB[27][2] ) );
  FADDER \r60/S2_27_1  ( .CIN(\r60/ab[27][1] ), .IN0(\r60/CARRYB[26][1] ), 
        .IN1(\r60/SUMB[26][2] ), .COUT(\r60/CARRYB[27][1] ), .SUM(
        \r60/SUMB[27][1] ) );
  FADDER \r60/S1_27_0  ( .CIN(\r60/ab[27][0] ), .IN0(\r60/CARRYB[26][0] ), 
        .IN1(\r60/SUMB[26][1] ), .COUT(\r60/CARRYB[27][0] ), .SUM(N144) );
  FADDER \r60/S3_28_30  ( .CIN(\r60/ab[28][30] ), .IN0(\r60/CARRYB[27][30] ), 
        .IN1(\r60/ab[27][31] ), .COUT(\r60/CARRYB[28][30] ), .SUM(
        \r60/SUMB[28][30] ) );
  FADDER \r60/S2_28_29  ( .CIN(\r60/ab[28][29] ), .IN0(\r60/CARRYB[27][29] ), 
        .IN1(\r60/SUMB[27][30] ), .COUT(\r60/CARRYB[28][29] ), .SUM(
        \r60/SUMB[28][29] ) );
  FADDER \r60/S2_28_28  ( .CIN(\r60/ab[28][28] ), .IN0(\r60/CARRYB[27][28] ), 
        .IN1(\r60/SUMB[27][29] ), .COUT(\r60/CARRYB[28][28] ), .SUM(
        \r60/SUMB[28][28] ) );
  FADDER \r60/S2_28_27  ( .CIN(\r60/ab[28][27] ), .IN0(\r60/CARRYB[27][27] ), 
        .IN1(\r60/SUMB[27][28] ), .COUT(\r60/CARRYB[28][27] ), .SUM(
        \r60/SUMB[28][27] ) );
  FADDER \r60/S2_28_26  ( .CIN(\r60/ab[28][26] ), .IN0(\r60/CARRYB[27][26] ), 
        .IN1(\r60/SUMB[27][27] ), .COUT(\r60/CARRYB[28][26] ), .SUM(
        \r60/SUMB[28][26] ) );
  FADDER \r60/S2_28_25  ( .CIN(\r60/ab[28][25] ), .IN0(\r60/CARRYB[27][25] ), 
        .IN1(\r60/SUMB[27][26] ), .COUT(\r60/CARRYB[28][25] ), .SUM(
        \r60/SUMB[28][25] ) );
  FADDER \r60/S2_28_24  ( .CIN(\r60/ab[28][24] ), .IN0(\r60/CARRYB[27][24] ), 
        .IN1(\r60/SUMB[27][25] ), .COUT(\r60/CARRYB[28][24] ), .SUM(
        \r60/SUMB[28][24] ) );
  FADDER \r60/S2_28_23  ( .CIN(\r60/ab[28][23] ), .IN0(\r60/CARRYB[27][23] ), 
        .IN1(\r60/SUMB[27][24] ), .COUT(\r60/CARRYB[28][23] ), .SUM(
        \r60/SUMB[28][23] ) );
  FADDER \r60/S2_28_22  ( .CIN(\r60/ab[28][22] ), .IN0(\r60/CARRYB[27][22] ), 
        .IN1(\r60/SUMB[27][23] ), .COUT(\r60/CARRYB[28][22] ), .SUM(
        \r60/SUMB[28][22] ) );
  FADDER \r60/S2_28_21  ( .CIN(\r60/ab[28][21] ), .IN0(\r60/CARRYB[27][21] ), 
        .IN1(\r60/SUMB[27][22] ), .COUT(\r60/CARRYB[28][21] ), .SUM(
        \r60/SUMB[28][21] ) );
  FADDER \r60/S2_28_20  ( .CIN(\r60/ab[28][20] ), .IN0(\r60/CARRYB[27][20] ), 
        .IN1(\r60/SUMB[27][21] ), .COUT(\r60/CARRYB[28][20] ), .SUM(
        \r60/SUMB[28][20] ) );
  FADDER \r60/S2_28_19  ( .CIN(\r60/ab[28][19] ), .IN0(\r60/CARRYB[27][19] ), 
        .IN1(\r60/SUMB[27][20] ), .COUT(\r60/CARRYB[28][19] ), .SUM(
        \r60/SUMB[28][19] ) );
  FADDER \r60/S2_28_18  ( .CIN(\r60/ab[28][18] ), .IN0(\r60/CARRYB[27][18] ), 
        .IN1(\r60/SUMB[27][19] ), .COUT(\r60/CARRYB[28][18] ), .SUM(
        \r60/SUMB[28][18] ) );
  FADDER \r60/S2_28_17  ( .CIN(\r60/ab[28][17] ), .IN0(\r60/CARRYB[27][17] ), 
        .IN1(\r60/SUMB[27][18] ), .COUT(\r60/CARRYB[28][17] ), .SUM(
        \r60/SUMB[28][17] ) );
  FADDER \r60/S2_28_16  ( .CIN(\r60/ab[28][16] ), .IN0(\r60/CARRYB[27][16] ), 
        .IN1(\r60/SUMB[27][17] ), .COUT(\r60/CARRYB[28][16] ), .SUM(
        \r60/SUMB[28][16] ) );
  FADDER \r60/S2_28_15  ( .CIN(\r60/ab[28][15] ), .IN0(\r60/CARRYB[27][15] ), 
        .IN1(\r60/SUMB[27][16] ), .COUT(\r60/CARRYB[28][15] ), .SUM(
        \r60/SUMB[28][15] ) );
  FADDER \r60/S2_28_14  ( .CIN(\r60/ab[28][14] ), .IN0(\r60/CARRYB[27][14] ), 
        .IN1(\r60/SUMB[27][15] ), .COUT(\r60/CARRYB[28][14] ), .SUM(
        \r60/SUMB[28][14] ) );
  FADDER \r60/S2_28_13  ( .CIN(\r60/ab[28][13] ), .IN0(\r60/CARRYB[27][13] ), 
        .IN1(\r60/SUMB[27][14] ), .COUT(\r60/CARRYB[28][13] ), .SUM(
        \r60/SUMB[28][13] ) );
  FADDER \r60/S2_28_12  ( .CIN(\r60/ab[28][12] ), .IN0(\r60/CARRYB[27][12] ), 
        .IN1(\r60/SUMB[27][13] ), .COUT(\r60/CARRYB[28][12] ), .SUM(
        \r60/SUMB[28][12] ) );
  FADDER \r60/S2_28_11  ( .CIN(\r60/ab[28][11] ), .IN0(\r60/CARRYB[27][11] ), 
        .IN1(\r60/SUMB[27][12] ), .COUT(\r60/CARRYB[28][11] ), .SUM(
        \r60/SUMB[28][11] ) );
  FADDER \r60/S2_28_10  ( .CIN(\r60/ab[28][10] ), .IN0(\r60/CARRYB[27][10] ), 
        .IN1(\r60/SUMB[27][11] ), .COUT(\r60/CARRYB[28][10] ), .SUM(
        \r60/SUMB[28][10] ) );
  FADDER \r60/S2_28_9  ( .CIN(\r60/ab[28][9] ), .IN0(\r60/CARRYB[27][9] ), 
        .IN1(\r60/SUMB[27][10] ), .COUT(\r60/CARRYB[28][9] ), .SUM(
        \r60/SUMB[28][9] ) );
  FADDER \r60/S2_28_8  ( .CIN(\r60/ab[28][8] ), .IN0(\r60/CARRYB[27][8] ), 
        .IN1(\r60/SUMB[27][9] ), .COUT(\r60/CARRYB[28][8] ), .SUM(
        \r60/SUMB[28][8] ) );
  FADDER \r60/S2_28_7  ( .CIN(\r60/ab[28][7] ), .IN0(\r60/CARRYB[27][7] ), 
        .IN1(\r60/SUMB[27][8] ), .COUT(\r60/CARRYB[28][7] ), .SUM(
        \r60/SUMB[28][7] ) );
  FADDER \r60/S2_28_6  ( .CIN(\r60/ab[28][6] ), .IN0(\r60/CARRYB[27][6] ), 
        .IN1(\r60/SUMB[27][7] ), .COUT(\r60/CARRYB[28][6] ), .SUM(
        \r60/SUMB[28][6] ) );
  FADDER \r60/S2_28_5  ( .CIN(\r60/ab[28][5] ), .IN0(\r60/CARRYB[27][5] ), 
        .IN1(\r60/SUMB[27][6] ), .COUT(\r60/CARRYB[28][5] ), .SUM(
        \r60/SUMB[28][5] ) );
  FADDER \r60/S2_28_4  ( .CIN(\r60/ab[28][4] ), .IN0(\r60/CARRYB[27][4] ), 
        .IN1(\r60/SUMB[27][5] ), .COUT(\r60/CARRYB[28][4] ), .SUM(
        \r60/SUMB[28][4] ) );
  FADDER \r60/S2_28_3  ( .CIN(\r60/ab[28][3] ), .IN0(\r60/CARRYB[27][3] ), 
        .IN1(\r60/SUMB[27][4] ), .COUT(\r60/CARRYB[28][3] ), .SUM(
        \r60/SUMB[28][3] ) );
  FADDER \r60/S2_28_2  ( .CIN(\r60/ab[28][2] ), .IN0(\r60/CARRYB[27][2] ), 
        .IN1(\r60/SUMB[27][3] ), .COUT(\r60/CARRYB[28][2] ), .SUM(
        \r60/SUMB[28][2] ) );
  FADDER \r60/S2_28_1  ( .CIN(\r60/ab[28][1] ), .IN0(\r60/CARRYB[27][1] ), 
        .IN1(\r60/SUMB[27][2] ), .COUT(\r60/CARRYB[28][1] ), .SUM(
        \r60/SUMB[28][1] ) );
  FADDER \r60/S1_28_0  ( .CIN(\r60/ab[28][0] ), .IN0(\r60/CARRYB[27][0] ), 
        .IN1(\r60/SUMB[27][1] ), .COUT(\r60/CARRYB[28][0] ), .SUM(N145) );
  FADDER \r60/S3_29_30  ( .CIN(\r60/ab[29][30] ), .IN0(\r60/CARRYB[28][30] ), 
        .IN1(\r60/ab[28][31] ), .COUT(\r60/CARRYB[29][30] ), .SUM(
        \r60/SUMB[29][30] ) );
  FADDER \r60/S2_29_29  ( .CIN(\r60/ab[29][29] ), .IN0(\r60/CARRYB[28][29] ), 
        .IN1(\r60/SUMB[28][30] ), .COUT(\r60/CARRYB[29][29] ), .SUM(
        \r60/SUMB[29][29] ) );
  FADDER \r60/S2_29_28  ( .CIN(\r60/ab[29][28] ), .IN0(\r60/CARRYB[28][28] ), 
        .IN1(\r60/SUMB[28][29] ), .COUT(\r60/CARRYB[29][28] ), .SUM(
        \r60/SUMB[29][28] ) );
  FADDER \r60/S2_29_27  ( .CIN(\r60/ab[29][27] ), .IN0(\r60/CARRYB[28][27] ), 
        .IN1(\r60/SUMB[28][28] ), .COUT(\r60/CARRYB[29][27] ), .SUM(
        \r60/SUMB[29][27] ) );
  FADDER \r60/S2_29_26  ( .CIN(\r60/ab[29][26] ), .IN0(\r60/CARRYB[28][26] ), 
        .IN1(\r60/SUMB[28][27] ), .COUT(\r60/CARRYB[29][26] ), .SUM(
        \r60/SUMB[29][26] ) );
  FADDER \r60/S2_29_25  ( .CIN(\r60/ab[29][25] ), .IN0(\r60/CARRYB[28][25] ), 
        .IN1(\r60/SUMB[28][26] ), .COUT(\r60/CARRYB[29][25] ), .SUM(
        \r60/SUMB[29][25] ) );
  FADDER \r60/S2_29_24  ( .CIN(\r60/ab[29][24] ), .IN0(\r60/CARRYB[28][24] ), 
        .IN1(\r60/SUMB[28][25] ), .COUT(\r60/CARRYB[29][24] ), .SUM(
        \r60/SUMB[29][24] ) );
  FADDER \r60/S2_29_23  ( .CIN(\r60/ab[29][23] ), .IN0(\r60/CARRYB[28][23] ), 
        .IN1(\r60/SUMB[28][24] ), .COUT(\r60/CARRYB[29][23] ), .SUM(
        \r60/SUMB[29][23] ) );
  FADDER \r60/S2_29_22  ( .CIN(\r60/ab[29][22] ), .IN0(\r60/CARRYB[28][22] ), 
        .IN1(\r60/SUMB[28][23] ), .COUT(\r60/CARRYB[29][22] ), .SUM(
        \r60/SUMB[29][22] ) );
  FADDER \r60/S2_29_21  ( .CIN(\r60/ab[29][21] ), .IN0(\r60/CARRYB[28][21] ), 
        .IN1(\r60/SUMB[28][22] ), .COUT(\r60/CARRYB[29][21] ), .SUM(
        \r60/SUMB[29][21] ) );
  FADDER \r60/S2_29_20  ( .CIN(\r60/ab[29][20] ), .IN0(\r60/CARRYB[28][20] ), 
        .IN1(\r60/SUMB[28][21] ), .COUT(\r60/CARRYB[29][20] ), .SUM(
        \r60/SUMB[29][20] ) );
  FADDER \r60/S2_29_19  ( .CIN(\r60/ab[29][19] ), .IN0(\r60/CARRYB[28][19] ), 
        .IN1(\r60/SUMB[28][20] ), .COUT(\r60/CARRYB[29][19] ), .SUM(
        \r60/SUMB[29][19] ) );
  FADDER \r60/S2_29_18  ( .CIN(\r60/ab[29][18] ), .IN0(\r60/CARRYB[28][18] ), 
        .IN1(\r60/SUMB[28][19] ), .COUT(\r60/CARRYB[29][18] ), .SUM(
        \r60/SUMB[29][18] ) );
  FADDER \r60/S2_29_17  ( .CIN(\r60/ab[29][17] ), .IN0(\r60/CARRYB[28][17] ), 
        .IN1(\r60/SUMB[28][18] ), .COUT(\r60/CARRYB[29][17] ), .SUM(
        \r60/SUMB[29][17] ) );
  FADDER \r60/S2_29_16  ( .CIN(\r60/ab[29][16] ), .IN0(\r60/CARRYB[28][16] ), 
        .IN1(\r60/SUMB[28][17] ), .COUT(\r60/CARRYB[29][16] ), .SUM(
        \r60/SUMB[29][16] ) );
  FADDER \r60/S2_29_15  ( .CIN(\r60/ab[29][15] ), .IN0(\r60/CARRYB[28][15] ), 
        .IN1(\r60/SUMB[28][16] ), .COUT(\r60/CARRYB[29][15] ), .SUM(
        \r60/SUMB[29][15] ) );
  FADDER \r60/S2_29_14  ( .CIN(\r60/ab[29][14] ), .IN0(\r60/CARRYB[28][14] ), 
        .IN1(\r60/SUMB[28][15] ), .COUT(\r60/CARRYB[29][14] ), .SUM(
        \r60/SUMB[29][14] ) );
  FADDER \r60/S2_29_13  ( .CIN(\r60/ab[29][13] ), .IN0(\r60/CARRYB[28][13] ), 
        .IN1(\r60/SUMB[28][14] ), .COUT(\r60/CARRYB[29][13] ), .SUM(
        \r60/SUMB[29][13] ) );
  FADDER \r60/S2_29_12  ( .CIN(\r60/ab[29][12] ), .IN0(\r60/CARRYB[28][12] ), 
        .IN1(\r60/SUMB[28][13] ), .COUT(\r60/CARRYB[29][12] ), .SUM(
        \r60/SUMB[29][12] ) );
  FADDER \r60/S2_29_11  ( .CIN(\r60/ab[29][11] ), .IN0(\r60/CARRYB[28][11] ), 
        .IN1(\r60/SUMB[28][12] ), .COUT(\r60/CARRYB[29][11] ), .SUM(
        \r60/SUMB[29][11] ) );
  FADDER \r60/S2_29_10  ( .CIN(\r60/ab[29][10] ), .IN0(\r60/CARRYB[28][10] ), 
        .IN1(\r60/SUMB[28][11] ), .COUT(\r60/CARRYB[29][10] ), .SUM(
        \r60/SUMB[29][10] ) );
  FADDER \r60/S2_29_9  ( .CIN(\r60/ab[29][9] ), .IN0(\r60/CARRYB[28][9] ), 
        .IN1(\r60/SUMB[28][10] ), .COUT(\r60/CARRYB[29][9] ), .SUM(
        \r60/SUMB[29][9] ) );
  FADDER \r60/S2_29_8  ( .CIN(\r60/ab[29][8] ), .IN0(\r60/CARRYB[28][8] ), 
        .IN1(\r60/SUMB[28][9] ), .COUT(\r60/CARRYB[29][8] ), .SUM(
        \r60/SUMB[29][8] ) );
  FADDER \r60/S2_29_7  ( .CIN(\r60/ab[29][7] ), .IN0(\r60/CARRYB[28][7] ), 
        .IN1(\r60/SUMB[28][8] ), .COUT(\r60/CARRYB[29][7] ), .SUM(
        \r60/SUMB[29][7] ) );
  FADDER \r60/S2_29_6  ( .CIN(\r60/ab[29][6] ), .IN0(\r60/CARRYB[28][6] ), 
        .IN1(\r60/SUMB[28][7] ), .COUT(\r60/CARRYB[29][6] ), .SUM(
        \r60/SUMB[29][6] ) );
  FADDER \r60/S2_29_5  ( .CIN(\r60/ab[29][5] ), .IN0(\r60/CARRYB[28][5] ), 
        .IN1(\r60/SUMB[28][6] ), .COUT(\r60/CARRYB[29][5] ), .SUM(
        \r60/SUMB[29][5] ) );
  FADDER \r60/S2_29_4  ( .CIN(\r60/ab[29][4] ), .IN0(\r60/CARRYB[28][4] ), 
        .IN1(\r60/SUMB[28][5] ), .COUT(\r60/CARRYB[29][4] ), .SUM(
        \r60/SUMB[29][4] ) );
  FADDER \r60/S2_29_3  ( .CIN(\r60/ab[29][3] ), .IN0(\r60/CARRYB[28][3] ), 
        .IN1(\r60/SUMB[28][4] ), .COUT(\r60/CARRYB[29][3] ), .SUM(
        \r60/SUMB[29][3] ) );
  FADDER \r60/S2_29_2  ( .CIN(\r60/ab[29][2] ), .IN0(\r60/CARRYB[28][2] ), 
        .IN1(\r60/SUMB[28][3] ), .COUT(\r60/CARRYB[29][2] ), .SUM(
        \r60/SUMB[29][2] ) );
  FADDER \r60/S2_29_1  ( .CIN(\r60/ab[29][1] ), .IN0(\r60/CARRYB[28][1] ), 
        .IN1(\r60/SUMB[28][2] ), .COUT(\r60/CARRYB[29][1] ), .SUM(
        \r60/SUMB[29][1] ) );
  FADDER \r60/S1_29_0  ( .CIN(\r60/ab[29][0] ), .IN0(\r60/CARRYB[28][0] ), 
        .IN1(\r60/SUMB[28][1] ), .COUT(\r60/CARRYB[29][0] ), .SUM(N146) );
  FADDER \r60/S3_30_30  ( .CIN(\r60/ab[30][30] ), .IN0(\r60/CARRYB[29][30] ), 
        .IN1(\r60/ab[29][31] ), .COUT(\r60/CARRYB[30][30] ), .SUM(
        \r60/SUMB[30][30] ) );
  FADDER \r60/S2_30_29  ( .CIN(\r60/ab[30][29] ), .IN0(\r60/CARRYB[29][29] ), 
        .IN1(\r60/SUMB[29][30] ), .COUT(\r60/CARRYB[30][29] ), .SUM(
        \r60/SUMB[30][29] ) );
  FADDER \r60/S2_30_28  ( .CIN(\r60/ab[30][28] ), .IN0(\r60/CARRYB[29][28] ), 
        .IN1(\r60/SUMB[29][29] ), .COUT(\r60/CARRYB[30][28] ), .SUM(
        \r60/SUMB[30][28] ) );
  FADDER \r60/S2_30_27  ( .CIN(\r60/ab[30][27] ), .IN0(\r60/CARRYB[29][27] ), 
        .IN1(\r60/SUMB[29][28] ), .COUT(\r60/CARRYB[30][27] ), .SUM(
        \r60/SUMB[30][27] ) );
  FADDER \r60/S2_30_26  ( .CIN(\r60/ab[30][26] ), .IN0(\r60/CARRYB[29][26] ), 
        .IN1(\r60/SUMB[29][27] ), .COUT(\r60/CARRYB[30][26] ), .SUM(
        \r60/SUMB[30][26] ) );
  FADDER \r60/S2_30_25  ( .CIN(\r60/ab[30][25] ), .IN0(\r60/CARRYB[29][25] ), 
        .IN1(\r60/SUMB[29][26] ), .COUT(\r60/CARRYB[30][25] ), .SUM(
        \r60/SUMB[30][25] ) );
  FADDER \r60/S2_30_24  ( .CIN(\r60/ab[30][24] ), .IN0(\r60/CARRYB[29][24] ), 
        .IN1(\r60/SUMB[29][25] ), .COUT(\r60/CARRYB[30][24] ), .SUM(
        \r60/SUMB[30][24] ) );
  FADDER \r60/S2_30_23  ( .CIN(\r60/ab[30][23] ), .IN0(\r60/CARRYB[29][23] ), 
        .IN1(\r60/SUMB[29][24] ), .COUT(\r60/CARRYB[30][23] ), .SUM(
        \r60/SUMB[30][23] ) );
  FADDER \r60/S2_30_22  ( .CIN(\r60/ab[30][22] ), .IN0(\r60/CARRYB[29][22] ), 
        .IN1(\r60/SUMB[29][23] ), .COUT(\r60/CARRYB[30][22] ), .SUM(
        \r60/SUMB[30][22] ) );
  FADDER \r60/S2_30_21  ( .CIN(\r60/ab[30][21] ), .IN0(\r60/CARRYB[29][21] ), 
        .IN1(\r60/SUMB[29][22] ), .COUT(\r60/CARRYB[30][21] ), .SUM(
        \r60/SUMB[30][21] ) );
  FADDER \r60/S2_30_20  ( .CIN(\r60/ab[30][20] ), .IN0(\r60/CARRYB[29][20] ), 
        .IN1(\r60/SUMB[29][21] ), .COUT(\r60/CARRYB[30][20] ), .SUM(
        \r60/SUMB[30][20] ) );
  FADDER \r60/S2_30_19  ( .CIN(\r60/ab[30][19] ), .IN0(\r60/CARRYB[29][19] ), 
        .IN1(\r60/SUMB[29][20] ), .COUT(\r60/CARRYB[30][19] ), .SUM(
        \r60/SUMB[30][19] ) );
  FADDER \r60/S2_30_18  ( .CIN(\r60/ab[30][18] ), .IN0(\r60/CARRYB[29][18] ), 
        .IN1(\r60/SUMB[29][19] ), .COUT(\r60/CARRYB[30][18] ), .SUM(
        \r60/SUMB[30][18] ) );
  FADDER \r60/S2_30_17  ( .CIN(\r60/ab[30][17] ), .IN0(\r60/CARRYB[29][17] ), 
        .IN1(\r60/SUMB[29][18] ), .COUT(\r60/CARRYB[30][17] ), .SUM(
        \r60/SUMB[30][17] ) );
  FADDER \r60/S2_30_16  ( .CIN(\r60/ab[30][16] ), .IN0(\r60/CARRYB[29][16] ), 
        .IN1(\r60/SUMB[29][17] ), .COUT(\r60/CARRYB[30][16] ), .SUM(
        \r60/SUMB[30][16] ) );
  FADDER \r60/S2_30_15  ( .CIN(\r60/ab[30][15] ), .IN0(\r60/CARRYB[29][15] ), 
        .IN1(\r60/SUMB[29][16] ), .COUT(\r60/CARRYB[30][15] ), .SUM(
        \r60/SUMB[30][15] ) );
  FADDER \r60/S2_30_14  ( .CIN(\r60/ab[30][14] ), .IN0(\r60/CARRYB[29][14] ), 
        .IN1(\r60/SUMB[29][15] ), .COUT(\r60/CARRYB[30][14] ), .SUM(
        \r60/SUMB[30][14] ) );
  FADDER \r60/S2_30_13  ( .CIN(\r60/ab[30][13] ), .IN0(\r60/CARRYB[29][13] ), 
        .IN1(\r60/SUMB[29][14] ), .COUT(\r60/CARRYB[30][13] ), .SUM(
        \r60/SUMB[30][13] ) );
  FADDER \r60/S2_30_12  ( .CIN(\r60/ab[30][12] ), .IN0(\r60/CARRYB[29][12] ), 
        .IN1(\r60/SUMB[29][13] ), .COUT(\r60/CARRYB[30][12] ), .SUM(
        \r60/SUMB[30][12] ) );
  FADDER \r60/S2_30_11  ( .CIN(\r60/ab[30][11] ), .IN0(\r60/CARRYB[29][11] ), 
        .IN1(\r60/SUMB[29][12] ), .COUT(\r60/CARRYB[30][11] ), .SUM(
        \r60/SUMB[30][11] ) );
  FADDER \r60/S2_30_10  ( .CIN(\r60/ab[30][10] ), .IN0(\r60/CARRYB[29][10] ), 
        .IN1(\r60/SUMB[29][11] ), .COUT(\r60/CARRYB[30][10] ), .SUM(
        \r60/SUMB[30][10] ) );
  FADDER \r60/S2_30_9  ( .CIN(\r60/ab[30][9] ), .IN0(\r60/CARRYB[29][9] ), 
        .IN1(\r60/SUMB[29][10] ), .COUT(\r60/CARRYB[30][9] ), .SUM(
        \r60/SUMB[30][9] ) );
  FADDER \r60/S2_30_8  ( .CIN(\r60/ab[30][8] ), .IN0(\r60/CARRYB[29][8] ), 
        .IN1(\r60/SUMB[29][9] ), .COUT(\r60/CARRYB[30][8] ), .SUM(
        \r60/SUMB[30][8] ) );
  FADDER \r60/S2_30_7  ( .CIN(\r60/ab[30][7] ), .IN0(\r60/CARRYB[29][7] ), 
        .IN1(\r60/SUMB[29][8] ), .COUT(\r60/CARRYB[30][7] ), .SUM(
        \r60/SUMB[30][7] ) );
  FADDER \r60/S2_30_6  ( .CIN(\r60/ab[30][6] ), .IN0(\r60/CARRYB[29][6] ), 
        .IN1(\r60/SUMB[29][7] ), .COUT(\r60/CARRYB[30][6] ), .SUM(
        \r60/SUMB[30][6] ) );
  FADDER \r60/S2_30_5  ( .CIN(\r60/ab[30][5] ), .IN0(\r60/CARRYB[29][5] ), 
        .IN1(\r60/SUMB[29][6] ), .COUT(\r60/CARRYB[30][5] ), .SUM(
        \r60/SUMB[30][5] ) );
  FADDER \r60/S2_30_4  ( .CIN(\r60/ab[30][4] ), .IN0(\r60/CARRYB[29][4] ), 
        .IN1(\r60/SUMB[29][5] ), .COUT(\r60/CARRYB[30][4] ), .SUM(
        \r60/SUMB[30][4] ) );
  FADDER \r60/S2_30_3  ( .CIN(\r60/ab[30][3] ), .IN0(\r60/CARRYB[29][3] ), 
        .IN1(\r60/SUMB[29][4] ), .COUT(\r60/CARRYB[30][3] ), .SUM(
        \r60/SUMB[30][3] ) );
  FADDER \r60/S2_30_2  ( .CIN(\r60/ab[30][2] ), .IN0(\r60/CARRYB[29][2] ), 
        .IN1(\r60/SUMB[29][3] ), .COUT(\r60/CARRYB[30][2] ), .SUM(
        \r60/SUMB[30][2] ) );
  FADDER \r60/S2_30_1  ( .CIN(\r60/ab[30][1] ), .IN0(\r60/CARRYB[29][1] ), 
        .IN1(\r60/SUMB[29][2] ), .COUT(\r60/CARRYB[30][1] ), .SUM(
        \r60/SUMB[30][1] ) );
  FADDER \r60/S1_30_0  ( .CIN(\r60/ab[30][0] ), .IN0(\r60/CARRYB[29][0] ), 
        .IN1(\r60/SUMB[29][1] ), .COUT(\r60/CARRYB[30][0] ), .SUM(N147) );
  FADDER \r60/S14_31  ( .CIN(\r60/QA ), .IN0(\r60/QB ), .IN1(\r60/ab[31][31] ), 
        .COUT(\r60/CARRYB[31][31] ), .SUM(\r60/SUMB[31][31] ) );
  FADDER \r60/S5_30  ( .CIN(\r60/ab[31][30] ), .IN0(\r60/CARRYB[30][30] ), 
        .IN1(\r60/ab[30][31] ), .COUT(\r60/CARRYB[31][30] ), .SUM(
        \r60/SUMB[31][30] ) );
  FADDER \r60/S4_29  ( .CIN(\r60/ab[31][29] ), .IN0(\r60/CARRYB[30][29] ), 
        .IN1(\r60/SUMB[30][30] ), .COUT(\r60/CARRYB[31][29] ), .SUM(
        \r60/SUMB[31][29] ) );
  FADDER \r60/S4_28  ( .CIN(\r60/ab[31][28] ), .IN0(\r60/CARRYB[30][28] ), 
        .IN1(\r60/SUMB[30][29] ), .COUT(\r60/CARRYB[31][28] ), .SUM(
        \r60/SUMB[31][28] ) );
  FADDER \r60/S4_27  ( .CIN(\r60/ab[31][27] ), .IN0(\r60/CARRYB[30][27] ), 
        .IN1(\r60/SUMB[30][28] ), .COUT(\r60/CARRYB[31][27] ), .SUM(
        \r60/SUMB[31][27] ) );
  FADDER \r60/S4_26  ( .CIN(\r60/ab[31][26] ), .IN0(\r60/CARRYB[30][26] ), 
        .IN1(\r60/SUMB[30][27] ), .COUT(\r60/CARRYB[31][26] ), .SUM(
        \r60/SUMB[31][26] ) );
  FADDER \r60/S4_25  ( .CIN(\r60/ab[31][25] ), .IN0(\r60/CARRYB[30][25] ), 
        .IN1(\r60/SUMB[30][26] ), .COUT(\r60/CARRYB[31][25] ), .SUM(
        \r60/SUMB[31][25] ) );
  FADDER \r60/S4_24  ( .CIN(\r60/ab[31][24] ), .IN0(\r60/CARRYB[30][24] ), 
        .IN1(\r60/SUMB[30][25] ), .COUT(\r60/CARRYB[31][24] ), .SUM(
        \r60/SUMB[31][24] ) );
  FADDER \r60/S4_23  ( .CIN(\r60/ab[31][23] ), .IN0(\r60/CARRYB[30][23] ), 
        .IN1(\r60/SUMB[30][24] ), .COUT(\r60/CARRYB[31][23] ), .SUM(
        \r60/SUMB[31][23] ) );
  FADDER \r60/S4_22  ( .CIN(\r60/ab[31][22] ), .IN0(\r60/CARRYB[30][22] ), 
        .IN1(\r60/SUMB[30][23] ), .COUT(\r60/CARRYB[31][22] ), .SUM(
        \r60/SUMB[31][22] ) );
  FADDER \r60/S4_21  ( .CIN(\r60/ab[31][21] ), .IN0(\r60/CARRYB[30][21] ), 
        .IN1(\r60/SUMB[30][22] ), .COUT(\r60/CARRYB[31][21] ), .SUM(
        \r60/SUMB[31][21] ) );
  FADDER \r60/S4_20  ( .CIN(\r60/ab[31][20] ), .IN0(\r60/CARRYB[30][20] ), 
        .IN1(\r60/SUMB[30][21] ), .COUT(\r60/CARRYB[31][20] ), .SUM(
        \r60/SUMB[31][20] ) );
  FADDER \r60/S4_19  ( .CIN(\r60/ab[31][19] ), .IN0(\r60/CARRYB[30][19] ), 
        .IN1(\r60/SUMB[30][20] ), .COUT(\r60/CARRYB[31][19] ), .SUM(
        \r60/SUMB[31][19] ) );
  FADDER \r60/S4_18  ( .CIN(\r60/ab[31][18] ), .IN0(\r60/CARRYB[30][18] ), 
        .IN1(\r60/SUMB[30][19] ), .COUT(\r60/CARRYB[31][18] ), .SUM(
        \r60/SUMB[31][18] ) );
  FADDER \r60/S4_17  ( .CIN(\r60/ab[31][17] ), .IN0(\r60/CARRYB[30][17] ), 
        .IN1(\r60/SUMB[30][18] ), .COUT(\r60/CARRYB[31][17] ), .SUM(
        \r60/SUMB[31][17] ) );
  FADDER \r60/S4_16  ( .CIN(\r60/ab[31][16] ), .IN0(\r60/CARRYB[30][16] ), 
        .IN1(\r60/SUMB[30][17] ), .COUT(\r60/CARRYB[31][16] ), .SUM(
        \r60/SUMB[31][16] ) );
  FADDER \r60/S4_15  ( .CIN(\r60/ab[31][15] ), .IN0(\r60/CARRYB[30][15] ), 
        .IN1(\r60/SUMB[30][16] ), .COUT(\r60/CARRYB[31][15] ), .SUM(
        \r60/SUMB[31][15] ) );
  FADDER \r60/S4_14  ( .CIN(\r60/ab[31][14] ), .IN0(\r60/CARRYB[30][14] ), 
        .IN1(\r60/SUMB[30][15] ), .COUT(\r60/CARRYB[31][14] ), .SUM(
        \r60/SUMB[31][14] ) );
  FADDER \r60/S4_13  ( .CIN(\r60/ab[31][13] ), .IN0(\r60/CARRYB[30][13] ), 
        .IN1(\r60/SUMB[30][14] ), .COUT(\r60/CARRYB[31][13] ), .SUM(
        \r60/SUMB[31][13] ) );
  FADDER \r60/S4_12  ( .CIN(\r60/ab[31][12] ), .IN0(\r60/CARRYB[30][12] ), 
        .IN1(\r60/SUMB[30][13] ), .COUT(\r60/CARRYB[31][12] ), .SUM(
        \r60/SUMB[31][12] ) );
  FADDER \r60/S4_11  ( .CIN(\r60/ab[31][11] ), .IN0(\r60/CARRYB[30][11] ), 
        .IN1(\r60/SUMB[30][12] ), .COUT(\r60/CARRYB[31][11] ), .SUM(
        \r60/SUMB[31][11] ) );
  FADDER \r60/S4_10  ( .CIN(\r60/ab[31][10] ), .IN0(\r60/CARRYB[30][10] ), 
        .IN1(\r60/SUMB[30][11] ), .COUT(\r60/CARRYB[31][10] ), .SUM(
        \r60/SUMB[31][10] ) );
  FADDER \r60/S4_9  ( .CIN(\r60/ab[31][9] ), .IN0(\r60/CARRYB[30][9] ), .IN1(
        \r60/SUMB[30][10] ), .COUT(\r60/CARRYB[31][9] ), .SUM(
        \r60/SUMB[31][9] ) );
  FADDER \r60/S4_8  ( .CIN(\r60/ab[31][8] ), .IN0(\r60/CARRYB[30][8] ), .IN1(
        \r60/SUMB[30][9] ), .COUT(\r60/CARRYB[31][8] ), .SUM(\r60/SUMB[31][8] ) );
  FADDER \r60/S4_7  ( .CIN(\r60/ab[31][7] ), .IN0(\r60/CARRYB[30][7] ), .IN1(
        \r60/SUMB[30][8] ), .COUT(\r60/CARRYB[31][7] ), .SUM(\r60/SUMB[31][7] ) );
  FADDER \r60/S4_6  ( .CIN(\r60/ab[31][6] ), .IN0(\r60/CARRYB[30][6] ), .IN1(
        \r60/SUMB[30][7] ), .COUT(\r60/CARRYB[31][6] ), .SUM(\r60/SUMB[31][6] ) );
  FADDER \r60/S4_5  ( .CIN(\r60/ab[31][5] ), .IN0(\r60/CARRYB[30][5] ), .IN1(
        \r60/SUMB[30][6] ), .COUT(\r60/CARRYB[31][5] ), .SUM(\r60/SUMB[31][5] ) );
  FADDER \r60/S4_4  ( .CIN(\r60/ab[31][4] ), .IN0(\r60/CARRYB[30][4] ), .IN1(
        \r60/SUMB[30][5] ), .COUT(\r60/CARRYB[31][4] ), .SUM(\r60/SUMB[31][4] ) );
  FADDER \r60/S4_3  ( .CIN(\r60/ab[31][3] ), .IN0(\r60/CARRYB[30][3] ), .IN1(
        \r60/SUMB[30][4] ), .COUT(\r60/CARRYB[31][3] ), .SUM(\r60/SUMB[31][3] ) );
  FADDER \r60/S4_2  ( .CIN(\r60/ab[31][2] ), .IN0(\r60/CARRYB[30][2] ), .IN1(
        \r60/SUMB[30][3] ), .COUT(\r60/CARRYB[31][2] ), .SUM(\r60/SUMB[31][2] ) );
  FADDER \r60/S4_1  ( .CIN(\r60/ab[31][1] ), .IN0(\r60/CARRYB[30][1] ), .IN1(
        \r60/SUMB[30][2] ), .COUT(\r60/CARRYB[31][1] ), .SUM(\r60/SUMB[31][1] ) );
  FADDER \r60/S4_0  ( .CIN(\r60/ab[31][0] ), .IN0(\r60/CARRYB[30][0] ), .IN1(
        \r60/SUMB[30][1] ), .COUT(\r60/CARRYB[31][0] ), .SUM(\r60/SUMB[31][0] ) );
  FADDER \r60/S14_31_0  ( .CIN(\r60/ZA ), .IN0(\r60/ZB ), .IN1(
        \r60/SUMB[31][0] ), .COUT(\r60/A2[30] ), .SUM(N148) );
  AND U710 ( .A(\r60/SUMB[31][1] ), .B(\r60/CARRYB[31][0] ), .Z(\r60/A2[31] )
         );
  XOR U711 ( .A(\r60/SUMB[31][1] ), .B(\r60/CARRYB[31][0] ), .Z(\r60/A1[30] )
         );
  AND U712 ( .A(\r60/SUMB[31][2] ), .B(\r60/CARRYB[31][1] ), .Z(\r60/A2[32] )
         );
  XOR U713 ( .A(\r60/SUMB[31][2] ), .B(\r60/CARRYB[31][1] ), .Z(\r60/A1[31] )
         );
  AND U714 ( .A(\r60/SUMB[31][3] ), .B(\r60/CARRYB[31][2] ), .Z(\r60/A2[33] )
         );
  XOR U715 ( .A(\r60/SUMB[31][3] ), .B(\r60/CARRYB[31][2] ), .Z(\r60/A1[32] )
         );
  AND U716 ( .A(\r60/SUMB[31][4] ), .B(\r60/CARRYB[31][3] ), .Z(\r60/A2[34] )
         );
  XOR U717 ( .A(\r60/SUMB[31][4] ), .B(\r60/CARRYB[31][3] ), .Z(\r60/A1[33] )
         );
  AND U718 ( .A(\r60/SUMB[31][5] ), .B(\r60/CARRYB[31][4] ), .Z(\r60/A2[35] )
         );
  XOR U719 ( .A(\r60/SUMB[31][5] ), .B(\r60/CARRYB[31][4] ), .Z(\r60/A1[34] )
         );
  AND U720 ( .A(\r60/SUMB[31][6] ), .B(\r60/CARRYB[31][5] ), .Z(\r60/A2[36] )
         );
  XOR U721 ( .A(\r60/SUMB[31][6] ), .B(\r60/CARRYB[31][5] ), .Z(\r60/A1[35] )
         );
  AND U722 ( .A(\r60/SUMB[31][7] ), .B(\r60/CARRYB[31][6] ), .Z(\r60/A2[37] )
         );
  XOR U723 ( .A(\r60/SUMB[31][7] ), .B(\r60/CARRYB[31][6] ), .Z(\r60/A1[36] )
         );
  AND U724 ( .A(\r60/SUMB[31][8] ), .B(\r60/CARRYB[31][7] ), .Z(\r60/A2[38] )
         );
  XOR U725 ( .A(\r60/SUMB[31][8] ), .B(\r60/CARRYB[31][7] ), .Z(\r60/A1[37] )
         );
  AND U726 ( .A(\r60/SUMB[31][9] ), .B(\r60/CARRYB[31][8] ), .Z(\r60/A2[39] )
         );
  XOR U727 ( .A(\r60/SUMB[31][9] ), .B(\r60/CARRYB[31][8] ), .Z(\r60/A1[38] )
         );
  AND U728 ( .A(\r60/SUMB[31][10] ), .B(\r60/CARRYB[31][9] ), .Z(\r60/A2[40] )
         );
  XOR U729 ( .A(\r60/SUMB[31][10] ), .B(\r60/CARRYB[31][9] ), .Z(\r60/A1[39] )
         );
  AND U730 ( .A(\r60/SUMB[31][11] ), .B(\r60/CARRYB[31][10] ), .Z(\r60/A2[41] ) );
  XOR U731 ( .A(\r60/SUMB[31][11] ), .B(\r60/CARRYB[31][10] ), .Z(\r60/A1[40] ) );
  AND U732 ( .A(\r60/SUMB[31][12] ), .B(\r60/CARRYB[31][11] ), .Z(\r60/A2[42] ) );
  XOR U733 ( .A(\r60/SUMB[31][12] ), .B(\r60/CARRYB[31][11] ), .Z(\r60/A1[41] ) );
  AND U734 ( .A(\r60/SUMB[31][13] ), .B(\r60/CARRYB[31][12] ), .Z(\r60/A2[43] ) );
  XOR U735 ( .A(\r60/SUMB[31][13] ), .B(\r60/CARRYB[31][12] ), .Z(\r60/A1[42] ) );
  AND U736 ( .A(\r60/SUMB[31][14] ), .B(\r60/CARRYB[31][13] ), .Z(\r60/A2[44] ) );
  XOR U737 ( .A(\r60/SUMB[31][14] ), .B(\r60/CARRYB[31][13] ), .Z(\r60/A1[43] ) );
  AND U738 ( .A(\r60/SUMB[31][15] ), .B(\r60/CARRYB[31][14] ), .Z(\r60/A2[45] ) );
  XOR U739 ( .A(\r60/SUMB[31][15] ), .B(\r60/CARRYB[31][14] ), .Z(\r60/A1[44] ) );
  AND U740 ( .A(\r60/SUMB[31][16] ), .B(\r60/CARRYB[31][15] ), .Z(\r60/A2[46] ) );
  XOR U741 ( .A(\r60/SUMB[31][16] ), .B(\r60/CARRYB[31][15] ), .Z(\r60/A1[45] ) );
  AND U742 ( .A(\r60/SUMB[31][17] ), .B(\r60/CARRYB[31][16] ), .Z(\r60/A2[47] ) );
  XOR U743 ( .A(\r60/SUMB[31][17] ), .B(\r60/CARRYB[31][16] ), .Z(\r60/A1[46] ) );
  AND U744 ( .A(\r60/SUMB[31][18] ), .B(\r60/CARRYB[31][17] ), .Z(\r60/A2[48] ) );
  XOR U745 ( .A(\r60/SUMB[31][18] ), .B(\r60/CARRYB[31][17] ), .Z(\r60/A1[47] ) );
  AND U746 ( .A(\r60/SUMB[31][19] ), .B(\r60/CARRYB[31][18] ), .Z(\r60/A2[49] ) );
  XOR U747 ( .A(\r60/SUMB[31][19] ), .B(\r60/CARRYB[31][18] ), .Z(\r60/A1[48] ) );
  AND U748 ( .A(\r60/SUMB[31][20] ), .B(\r60/CARRYB[31][19] ), .Z(\r60/A2[50] ) );
  XOR U749 ( .A(\r60/SUMB[31][20] ), .B(\r60/CARRYB[31][19] ), .Z(\r60/A1[49] ) );
  AND U750 ( .A(\r60/SUMB[31][21] ), .B(\r60/CARRYB[31][20] ), .Z(\r60/A2[51] ) );
  XOR U751 ( .A(\r60/SUMB[31][21] ), .B(\r60/CARRYB[31][20] ), .Z(\r60/A1[50] ) );
  AND U752 ( .A(\r60/SUMB[31][22] ), .B(\r60/CARRYB[31][21] ), .Z(\r60/A2[52] ) );
  XOR U753 ( .A(\r60/SUMB[31][22] ), .B(\r60/CARRYB[31][21] ), .Z(\r60/A1[51] ) );
  AND U754 ( .A(\r60/SUMB[31][23] ), .B(\r60/CARRYB[31][22] ), .Z(\r60/A2[53] ) );
  XOR U755 ( .A(\r60/SUMB[31][23] ), .B(\r60/CARRYB[31][22] ), .Z(\r60/A1[52] ) );
  AND U756 ( .A(\r60/SUMB[31][24] ), .B(\r60/CARRYB[31][23] ), .Z(\r60/A2[54] ) );
  XOR U757 ( .A(\r60/SUMB[31][24] ), .B(\r60/CARRYB[31][23] ), .Z(\r60/A1[53] ) );
  AND U758 ( .A(\r60/SUMB[31][25] ), .B(\r60/CARRYB[31][24] ), .Z(\r60/A2[55] ) );
  XOR U759 ( .A(\r60/SUMB[31][25] ), .B(\r60/CARRYB[31][24] ), .Z(\r60/A1[54] ) );
  AND U760 ( .A(\r60/SUMB[31][26] ), .B(\r60/CARRYB[31][25] ), .Z(\r60/A2[56] ) );
  XOR U761 ( .A(\r60/SUMB[31][26] ), .B(\r60/CARRYB[31][25] ), .Z(\r60/A1[55] ) );
  AND U762 ( .A(\r60/SUMB[31][27] ), .B(\r60/CARRYB[31][26] ), .Z(\r60/A2[57] ) );
  XOR U763 ( .A(\r60/SUMB[31][27] ), .B(\r60/CARRYB[31][26] ), .Z(\r60/A1[56] ) );
  AND U764 ( .A(\r60/SUMB[31][28] ), .B(\r60/CARRYB[31][27] ), .Z(\r60/A2[58] ) );
  XOR U765 ( .A(\r60/SUMB[31][28] ), .B(\r60/CARRYB[31][27] ), .Z(\r60/A1[57] ) );
  AND U766 ( .A(\r60/SUMB[31][29] ), .B(\r60/CARRYB[31][28] ), .Z(\r60/A2[59] ) );
  XOR U767 ( .A(\r60/SUMB[31][29] ), .B(\r60/CARRYB[31][28] ), .Z(\r60/A1[58] ) );
  AND U768 ( .A(\r60/SUMB[31][30] ), .B(\r60/CARRYB[31][29] ), .Z(\r60/A2[60] ) );
  XOR U769 ( .A(\r60/SUMB[31][30] ), .B(\r60/CARRYB[31][29] ), .Z(\r60/A1[59] ) );
  AND U770 ( .A(\r60/SUMB[31][31] ), .B(\r60/CARRYB[31][30] ), .Z(\r60/A2[61] ) );
  XOR U771 ( .A(\r60/SUMB[31][31] ), .B(\r60/CARRYB[31][30] ), .Z(\r60/A1[60] ) );
  XOR U772 ( .A(\r60/CARRYB[31][31] ), .B(\U3/U1/Z_0 ), .Z(\r60/A1[61] ) );
  AND U773 ( .A(\r60/ab[0][1] ), .B(\r60/ab[1][0] ), .Z(\r60/CARRYB[1][0] ) );
  XOR U774 ( .A(\r60/ab[0][1] ), .B(\r60/ab[1][0] ), .Z(N118) );
  AND U775 ( .A(\r60/ab[1][1] ), .B(\r60/ab[0][2] ), .Z(\r60/CARRYB[1][1] ) );
  XOR U776 ( .A(\r60/ab[0][2] ), .B(\r60/ab[1][1] ), .Z(\r60/SUMB[1][1] ) );
  AND U777 ( .A(\r60/ab[1][2] ), .B(\r60/ab[0][3] ), .Z(\r60/CARRYB[1][2] ) );
  XOR U778 ( .A(\r60/ab[0][3] ), .B(\r60/ab[1][2] ), .Z(\r60/SUMB[1][2] ) );
  AND U779 ( .A(\r60/ab[1][3] ), .B(\r60/ab[0][4] ), .Z(\r60/CARRYB[1][3] ) );
  XOR U780 ( .A(\r60/ab[0][4] ), .B(\r60/ab[1][3] ), .Z(\r60/SUMB[1][3] ) );
  AND U781 ( .A(\r60/ab[1][4] ), .B(\r60/ab[0][5] ), .Z(\r60/CARRYB[1][4] ) );
  XOR U782 ( .A(\r60/ab[0][5] ), .B(\r60/ab[1][4] ), .Z(\r60/SUMB[1][4] ) );
  AND U783 ( .A(\r60/ab[1][5] ), .B(\r60/ab[0][6] ), .Z(\r60/CARRYB[1][5] ) );
  XOR U784 ( .A(\r60/ab[0][6] ), .B(\r60/ab[1][5] ), .Z(\r60/SUMB[1][5] ) );
  AND U785 ( .A(\r60/ab[1][6] ), .B(\r60/ab[0][7] ), .Z(\r60/CARRYB[1][6] ) );
  XOR U786 ( .A(\r60/ab[0][7] ), .B(\r60/ab[1][6] ), .Z(\r60/SUMB[1][6] ) );
  AND U787 ( .A(\r60/ab[1][7] ), .B(\r60/ab[0][8] ), .Z(\r60/CARRYB[1][7] ) );
  XOR U788 ( .A(\r60/ab[0][8] ), .B(\r60/ab[1][7] ), .Z(\r60/SUMB[1][7] ) );
  AND U789 ( .A(\r60/ab[1][8] ), .B(\r60/ab[0][9] ), .Z(\r60/CARRYB[1][8] ) );
  XOR U790 ( .A(\r60/ab[0][9] ), .B(\r60/ab[1][8] ), .Z(\r60/SUMB[1][8] ) );
  AND U791 ( .A(\r60/ab[1][9] ), .B(\r60/ab[0][10] ), .Z(\r60/CARRYB[1][9] )
         );
  XOR U792 ( .A(\r60/ab[0][10] ), .B(\r60/ab[1][9] ), .Z(\r60/SUMB[1][9] ) );
  AND U793 ( .A(\r60/ab[1][10] ), .B(\r60/ab[0][11] ), .Z(\r60/CARRYB[1][10] )
         );
  XOR U794 ( .A(\r60/ab[0][11] ), .B(\r60/ab[1][10] ), .Z(\r60/SUMB[1][10] )
         );
  AND U795 ( .A(\r60/ab[1][11] ), .B(\r60/ab[0][12] ), .Z(\r60/CARRYB[1][11] )
         );
  XOR U796 ( .A(\r60/ab[0][12] ), .B(\r60/ab[1][11] ), .Z(\r60/SUMB[1][11] )
         );
  AND U797 ( .A(\r60/ab[1][12] ), .B(\r60/ab[0][13] ), .Z(\r60/CARRYB[1][12] )
         );
  XOR U798 ( .A(\r60/ab[0][13] ), .B(\r60/ab[1][12] ), .Z(\r60/SUMB[1][12] )
         );
  AND U799 ( .A(\r60/ab[1][13] ), .B(\r60/ab[0][14] ), .Z(\r60/CARRYB[1][13] )
         );
  XOR U800 ( .A(\r60/ab[0][14] ), .B(\r60/ab[1][13] ), .Z(\r60/SUMB[1][13] )
         );
  AND U801 ( .A(\r60/ab[1][14] ), .B(\r60/ab[0][15] ), .Z(\r60/CARRYB[1][14] )
         );
  XOR U802 ( .A(\r60/ab[0][15] ), .B(\r60/ab[1][14] ), .Z(\r60/SUMB[1][14] )
         );
  AND U803 ( .A(\r60/ab[1][15] ), .B(\r60/ab[0][16] ), .Z(\r60/CARRYB[1][15] )
         );
  XOR U804 ( .A(\r60/ab[0][16] ), .B(\r60/ab[1][15] ), .Z(\r60/SUMB[1][15] )
         );
  AND U805 ( .A(\r60/ab[1][16] ), .B(\r60/ab[0][17] ), .Z(\r60/CARRYB[1][16] )
         );
  XOR U806 ( .A(\r60/ab[0][17] ), .B(\r60/ab[1][16] ), .Z(\r60/SUMB[1][16] )
         );
  AND U807 ( .A(\r60/ab[1][17] ), .B(\r60/ab[0][18] ), .Z(\r60/CARRYB[1][17] )
         );
  XOR U808 ( .A(\r60/ab[0][18] ), .B(\r60/ab[1][17] ), .Z(\r60/SUMB[1][17] )
         );
  AND U809 ( .A(\r60/ab[1][18] ), .B(\r60/ab[0][19] ), .Z(\r60/CARRYB[1][18] )
         );
  XOR U810 ( .A(\r60/ab[0][19] ), .B(\r60/ab[1][18] ), .Z(\r60/SUMB[1][18] )
         );
  AND U811 ( .A(\r60/ab[1][19] ), .B(\r60/ab[0][20] ), .Z(\r60/CARRYB[1][19] )
         );
  XOR U812 ( .A(\r60/ab[0][20] ), .B(\r60/ab[1][19] ), .Z(\r60/SUMB[1][19] )
         );
  AND U813 ( .A(\r60/ab[1][20] ), .B(\r60/ab[0][21] ), .Z(\r60/CARRYB[1][20] )
         );
  XOR U814 ( .A(\r60/ab[0][21] ), .B(\r60/ab[1][20] ), .Z(\r60/SUMB[1][20] )
         );
  AND U815 ( .A(\r60/ab[1][21] ), .B(\r60/ab[0][22] ), .Z(\r60/CARRYB[1][21] )
         );
  XOR U816 ( .A(\r60/ab[0][22] ), .B(\r60/ab[1][21] ), .Z(\r60/SUMB[1][21] )
         );
  AND U817 ( .A(\r60/ab[1][22] ), .B(\r60/ab[0][23] ), .Z(\r60/CARRYB[1][22] )
         );
  XOR U818 ( .A(\r60/ab[0][23] ), .B(\r60/ab[1][22] ), .Z(\r60/SUMB[1][22] )
         );
  AND U819 ( .A(\r60/ab[1][23] ), .B(\r60/ab[0][24] ), .Z(\r60/CARRYB[1][23] )
         );
  XOR U820 ( .A(\r60/ab[0][24] ), .B(\r60/ab[1][23] ), .Z(\r60/SUMB[1][23] )
         );
  AND U821 ( .A(\r60/ab[1][24] ), .B(\r60/ab[0][25] ), .Z(\r60/CARRYB[1][24] )
         );
  XOR U822 ( .A(\r60/ab[0][25] ), .B(\r60/ab[1][24] ), .Z(\r60/SUMB[1][24] )
         );
  AND U823 ( .A(\r60/ab[1][25] ), .B(\r60/ab[0][26] ), .Z(\r60/CARRYB[1][25] )
         );
  XOR U824 ( .A(\r60/ab[0][26] ), .B(\r60/ab[1][25] ), .Z(\r60/SUMB[1][25] )
         );
  AND U825 ( .A(\r60/ab[1][26] ), .B(\r60/ab[0][27] ), .Z(\r60/CARRYB[1][26] )
         );
  XOR U826 ( .A(\r60/ab[0][27] ), .B(\r60/ab[1][26] ), .Z(\r60/SUMB[1][26] )
         );
  AND U827 ( .A(\r60/ab[1][27] ), .B(\r60/ab[0][28] ), .Z(\r60/CARRYB[1][27] )
         );
  XOR U828 ( .A(\r60/ab[0][28] ), .B(\r60/ab[1][27] ), .Z(\r60/SUMB[1][27] )
         );
  AND U829 ( .A(\r60/ab[1][28] ), .B(\r60/ab[0][29] ), .Z(\r60/CARRYB[1][28] )
         );
  XOR U830 ( .A(\r60/ab[0][29] ), .B(\r60/ab[1][28] ), .Z(\r60/SUMB[1][28] )
         );
  AND U831 ( .A(\r60/ab[1][29] ), .B(\r60/ab[0][30] ), .Z(\r60/CARRYB[1][29] )
         );
  XOR U832 ( .A(\r60/ab[0][30] ), .B(\r60/ab[1][29] ), .Z(\r60/SUMB[1][29] )
         );
  AND U833 ( .A(\r60/ab[1][30] ), .B(\r60/ab[0][31] ), .Z(\r60/CARRYB[1][30] )
         );
  XOR U834 ( .A(\r60/ab[0][31] ), .B(\r60/ab[1][30] ), .Z(\r60/SUMB[1][30] )
         );
  AND U835 ( .A(a[9]), .B(b[9]), .Z(\r60/ab[9][9] ) );
  AND U836 ( .A(a[9]), .B(b[8]), .Z(\r60/ab[9][8] ) );
  AND U837 ( .A(a[9]), .B(b[7]), .Z(\r60/ab[9][7] ) );
  AND U838 ( .A(a[9]), .B(b[6]), .Z(\r60/ab[9][6] ) );
  AND U839 ( .A(a[9]), .B(b[5]), .Z(\r60/ab[9][5] ) );
  AND U840 ( .A(a[9]), .B(b[4]), .Z(\r60/ab[9][4] ) );
  AND U841 ( .A(a[9]), .B(b[3]), .Z(\r60/ab[9][3] ) );
  MUX U842 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[9]), .F(\r60/ab[9][31] ) );
  AND U843 ( .A(a[9]), .B(b[30]), .Z(\r60/ab[9][30] ) );
  AND U844 ( .A(a[9]), .B(b[2]), .Z(\r60/ab[9][2] ) );
  AND U845 ( .A(a[9]), .B(b[29]), .Z(\r60/ab[9][29] ) );
  AND U846 ( .A(a[9]), .B(b[28]), .Z(\r60/ab[9][28] ) );
  AND U847 ( .A(a[9]), .B(b[27]), .Z(\r60/ab[9][27] ) );
  AND U848 ( .A(a[9]), .B(b[26]), .Z(\r60/ab[9][26] ) );
  AND U849 ( .A(a[9]), .B(b[25]), .Z(\r60/ab[9][25] ) );
  AND U850 ( .A(a[9]), .B(b[24]), .Z(\r60/ab[9][24] ) );
  AND U851 ( .A(a[9]), .B(b[23]), .Z(\r60/ab[9][23] ) );
  AND U852 ( .A(a[9]), .B(b[22]), .Z(\r60/ab[9][22] ) );
  AND U853 ( .A(a[9]), .B(b[21]), .Z(\r60/ab[9][21] ) );
  AND U854 ( .A(a[9]), .B(b[20]), .Z(\r60/ab[9][20] ) );
  AND U855 ( .A(a[9]), .B(b[1]), .Z(\r60/ab[9][1] ) );
  AND U856 ( .A(a[9]), .B(b[19]), .Z(\r60/ab[9][19] ) );
  AND U857 ( .A(a[9]), .B(b[18]), .Z(\r60/ab[9][18] ) );
  AND U858 ( .A(a[9]), .B(b[17]), .Z(\r60/ab[9][17] ) );
  AND U859 ( .A(a[9]), .B(b[16]), .Z(\r60/ab[9][16] ) );
  AND U860 ( .A(a[9]), .B(b[15]), .Z(\r60/ab[9][15] ) );
  AND U861 ( .A(a[9]), .B(b[14]), .Z(\r60/ab[9][14] ) );
  AND U862 ( .A(a[9]), .B(b[13]), .Z(\r60/ab[9][13] ) );
  AND U863 ( .A(a[9]), .B(b[12]), .Z(\r60/ab[9][12] ) );
  AND U864 ( .A(a[9]), .B(b[11]), .Z(\r60/ab[9][11] ) );
  AND U865 ( .A(a[9]), .B(b[10]), .Z(\r60/ab[9][10] ) );
  AND U866 ( .A(a[9]), .B(b[0]), .Z(\r60/ab[9][0] ) );
  AND U867 ( .A(b[9]), .B(a[8]), .Z(\r60/ab[8][9] ) );
  AND U868 ( .A(b[8]), .B(a[8]), .Z(\r60/ab[8][8] ) );
  AND U869 ( .A(b[7]), .B(a[8]), .Z(\r60/ab[8][7] ) );
  AND U870 ( .A(b[6]), .B(a[8]), .Z(\r60/ab[8][6] ) );
  AND U871 ( .A(b[5]), .B(a[8]), .Z(\r60/ab[8][5] ) );
  AND U872 ( .A(b[4]), .B(a[8]), .Z(\r60/ab[8][4] ) );
  AND U873 ( .A(b[3]), .B(a[8]), .Z(\r60/ab[8][3] ) );
  MUX U874 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[8]), .F(\r60/ab[8][31] ) );
  AND U875 ( .A(b[30]), .B(a[8]), .Z(\r60/ab[8][30] ) );
  AND U876 ( .A(b[2]), .B(a[8]), .Z(\r60/ab[8][2] ) );
  AND U877 ( .A(b[29]), .B(a[8]), .Z(\r60/ab[8][29] ) );
  AND U878 ( .A(b[28]), .B(a[8]), .Z(\r60/ab[8][28] ) );
  AND U879 ( .A(b[27]), .B(a[8]), .Z(\r60/ab[8][27] ) );
  AND U880 ( .A(b[26]), .B(a[8]), .Z(\r60/ab[8][26] ) );
  AND U881 ( .A(b[25]), .B(a[8]), .Z(\r60/ab[8][25] ) );
  AND U882 ( .A(b[24]), .B(a[8]), .Z(\r60/ab[8][24] ) );
  AND U883 ( .A(b[23]), .B(a[8]), .Z(\r60/ab[8][23] ) );
  AND U884 ( .A(b[22]), .B(a[8]), .Z(\r60/ab[8][22] ) );
  AND U885 ( .A(b[21]), .B(a[8]), .Z(\r60/ab[8][21] ) );
  AND U886 ( .A(b[20]), .B(a[8]), .Z(\r60/ab[8][20] ) );
  AND U887 ( .A(b[1]), .B(a[8]), .Z(\r60/ab[8][1] ) );
  AND U888 ( .A(b[19]), .B(a[8]), .Z(\r60/ab[8][19] ) );
  AND U889 ( .A(b[18]), .B(a[8]), .Z(\r60/ab[8][18] ) );
  AND U890 ( .A(b[17]), .B(a[8]), .Z(\r60/ab[8][17] ) );
  AND U891 ( .A(b[16]), .B(a[8]), .Z(\r60/ab[8][16] ) );
  AND U892 ( .A(b[15]), .B(a[8]), .Z(\r60/ab[8][15] ) );
  AND U893 ( .A(b[14]), .B(a[8]), .Z(\r60/ab[8][14] ) );
  AND U894 ( .A(b[13]), .B(a[8]), .Z(\r60/ab[8][13] ) );
  AND U895 ( .A(b[12]), .B(a[8]), .Z(\r60/ab[8][12] ) );
  AND U896 ( .A(b[11]), .B(a[8]), .Z(\r60/ab[8][11] ) );
  AND U897 ( .A(b[10]), .B(a[8]), .Z(\r60/ab[8][10] ) );
  AND U898 ( .A(b[0]), .B(a[8]), .Z(\r60/ab[8][0] ) );
  AND U899 ( .A(b[9]), .B(a[7]), .Z(\r60/ab[7][9] ) );
  AND U900 ( .A(b[8]), .B(a[7]), .Z(\r60/ab[7][8] ) );
  AND U901 ( .A(b[7]), .B(a[7]), .Z(\r60/ab[7][7] ) );
  AND U902 ( .A(b[6]), .B(a[7]), .Z(\r60/ab[7][6] ) );
  AND U903 ( .A(b[5]), .B(a[7]), .Z(\r60/ab[7][5] ) );
  AND U904 ( .A(b[4]), .B(a[7]), .Z(\r60/ab[7][4] ) );
  AND U905 ( .A(b[3]), .B(a[7]), .Z(\r60/ab[7][3] ) );
  MUX U906 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[7]), .F(\r60/ab[7][31] ) );
  AND U907 ( .A(b[30]), .B(a[7]), .Z(\r60/ab[7][30] ) );
  AND U908 ( .A(b[2]), .B(a[7]), .Z(\r60/ab[7][2] ) );
  AND U909 ( .A(b[29]), .B(a[7]), .Z(\r60/ab[7][29] ) );
  AND U910 ( .A(b[28]), .B(a[7]), .Z(\r60/ab[7][28] ) );
  AND U911 ( .A(b[27]), .B(a[7]), .Z(\r60/ab[7][27] ) );
  AND U912 ( .A(b[26]), .B(a[7]), .Z(\r60/ab[7][26] ) );
  AND U913 ( .A(b[25]), .B(a[7]), .Z(\r60/ab[7][25] ) );
  AND U914 ( .A(b[24]), .B(a[7]), .Z(\r60/ab[7][24] ) );
  AND U915 ( .A(b[23]), .B(a[7]), .Z(\r60/ab[7][23] ) );
  AND U916 ( .A(b[22]), .B(a[7]), .Z(\r60/ab[7][22] ) );
  AND U917 ( .A(b[21]), .B(a[7]), .Z(\r60/ab[7][21] ) );
  AND U918 ( .A(b[20]), .B(a[7]), .Z(\r60/ab[7][20] ) );
  AND U919 ( .A(b[1]), .B(a[7]), .Z(\r60/ab[7][1] ) );
  AND U920 ( .A(b[19]), .B(a[7]), .Z(\r60/ab[7][19] ) );
  AND U921 ( .A(b[18]), .B(a[7]), .Z(\r60/ab[7][18] ) );
  AND U922 ( .A(b[17]), .B(a[7]), .Z(\r60/ab[7][17] ) );
  AND U923 ( .A(b[16]), .B(a[7]), .Z(\r60/ab[7][16] ) );
  AND U924 ( .A(b[15]), .B(a[7]), .Z(\r60/ab[7][15] ) );
  AND U925 ( .A(b[14]), .B(a[7]), .Z(\r60/ab[7][14] ) );
  AND U926 ( .A(b[13]), .B(a[7]), .Z(\r60/ab[7][13] ) );
  AND U927 ( .A(b[12]), .B(a[7]), .Z(\r60/ab[7][12] ) );
  AND U928 ( .A(b[11]), .B(a[7]), .Z(\r60/ab[7][11] ) );
  AND U929 ( .A(b[10]), .B(a[7]), .Z(\r60/ab[7][10] ) );
  AND U930 ( .A(b[0]), .B(a[7]), .Z(\r60/ab[7][0] ) );
  AND U931 ( .A(b[9]), .B(a[6]), .Z(\r60/ab[6][9] ) );
  AND U932 ( .A(b[8]), .B(a[6]), .Z(\r60/ab[6][8] ) );
  AND U933 ( .A(b[7]), .B(a[6]), .Z(\r60/ab[6][7] ) );
  AND U934 ( .A(b[6]), .B(a[6]), .Z(\r60/ab[6][6] ) );
  AND U935 ( .A(b[5]), .B(a[6]), .Z(\r60/ab[6][5] ) );
  AND U936 ( .A(b[4]), .B(a[6]), .Z(\r60/ab[6][4] ) );
  AND U937 ( .A(b[3]), .B(a[6]), .Z(\r60/ab[6][3] ) );
  MUX U938 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[6]), .F(\r60/ab[6][31] ) );
  AND U939 ( .A(b[30]), .B(a[6]), .Z(\r60/ab[6][30] ) );
  AND U940 ( .A(b[2]), .B(a[6]), .Z(\r60/ab[6][2] ) );
  AND U941 ( .A(b[29]), .B(a[6]), .Z(\r60/ab[6][29] ) );
  AND U942 ( .A(b[28]), .B(a[6]), .Z(\r60/ab[6][28] ) );
  AND U943 ( .A(b[27]), .B(a[6]), .Z(\r60/ab[6][27] ) );
  AND U944 ( .A(b[26]), .B(a[6]), .Z(\r60/ab[6][26] ) );
  AND U945 ( .A(b[25]), .B(a[6]), .Z(\r60/ab[6][25] ) );
  AND U946 ( .A(b[24]), .B(a[6]), .Z(\r60/ab[6][24] ) );
  AND U947 ( .A(b[23]), .B(a[6]), .Z(\r60/ab[6][23] ) );
  AND U948 ( .A(b[22]), .B(a[6]), .Z(\r60/ab[6][22] ) );
  AND U949 ( .A(b[21]), .B(a[6]), .Z(\r60/ab[6][21] ) );
  AND U950 ( .A(b[20]), .B(a[6]), .Z(\r60/ab[6][20] ) );
  AND U951 ( .A(b[1]), .B(a[6]), .Z(\r60/ab[6][1] ) );
  AND U952 ( .A(b[19]), .B(a[6]), .Z(\r60/ab[6][19] ) );
  AND U953 ( .A(b[18]), .B(a[6]), .Z(\r60/ab[6][18] ) );
  AND U954 ( .A(b[17]), .B(a[6]), .Z(\r60/ab[6][17] ) );
  AND U955 ( .A(b[16]), .B(a[6]), .Z(\r60/ab[6][16] ) );
  AND U956 ( .A(b[15]), .B(a[6]), .Z(\r60/ab[6][15] ) );
  AND U957 ( .A(b[14]), .B(a[6]), .Z(\r60/ab[6][14] ) );
  AND U958 ( .A(b[13]), .B(a[6]), .Z(\r60/ab[6][13] ) );
  AND U959 ( .A(b[12]), .B(a[6]), .Z(\r60/ab[6][12] ) );
  AND U960 ( .A(b[11]), .B(a[6]), .Z(\r60/ab[6][11] ) );
  AND U961 ( .A(b[10]), .B(a[6]), .Z(\r60/ab[6][10] ) );
  AND U962 ( .A(b[0]), .B(a[6]), .Z(\r60/ab[6][0] ) );
  AND U963 ( .A(b[9]), .B(a[5]), .Z(\r60/ab[5][9] ) );
  AND U964 ( .A(b[8]), .B(a[5]), .Z(\r60/ab[5][8] ) );
  AND U965 ( .A(b[7]), .B(a[5]), .Z(\r60/ab[5][7] ) );
  AND U966 ( .A(b[6]), .B(a[5]), .Z(\r60/ab[5][6] ) );
  AND U967 ( .A(b[5]), .B(a[5]), .Z(\r60/ab[5][5] ) );
  AND U968 ( .A(b[4]), .B(a[5]), .Z(\r60/ab[5][4] ) );
  AND U969 ( .A(b[3]), .B(a[5]), .Z(\r60/ab[5][3] ) );
  MUX U970 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[5]), .F(\r60/ab[5][31] ) );
  AND U971 ( .A(b[30]), .B(a[5]), .Z(\r60/ab[5][30] ) );
  AND U972 ( .A(b[2]), .B(a[5]), .Z(\r60/ab[5][2] ) );
  AND U973 ( .A(b[29]), .B(a[5]), .Z(\r60/ab[5][29] ) );
  AND U974 ( .A(b[28]), .B(a[5]), .Z(\r60/ab[5][28] ) );
  AND U975 ( .A(b[27]), .B(a[5]), .Z(\r60/ab[5][27] ) );
  AND U976 ( .A(b[26]), .B(a[5]), .Z(\r60/ab[5][26] ) );
  AND U977 ( .A(b[25]), .B(a[5]), .Z(\r60/ab[5][25] ) );
  AND U978 ( .A(b[24]), .B(a[5]), .Z(\r60/ab[5][24] ) );
  AND U979 ( .A(b[23]), .B(a[5]), .Z(\r60/ab[5][23] ) );
  AND U980 ( .A(b[22]), .B(a[5]), .Z(\r60/ab[5][22] ) );
  AND U981 ( .A(b[21]), .B(a[5]), .Z(\r60/ab[5][21] ) );
  AND U982 ( .A(b[20]), .B(a[5]), .Z(\r60/ab[5][20] ) );
  AND U983 ( .A(b[1]), .B(a[5]), .Z(\r60/ab[5][1] ) );
  AND U984 ( .A(b[19]), .B(a[5]), .Z(\r60/ab[5][19] ) );
  AND U985 ( .A(b[18]), .B(a[5]), .Z(\r60/ab[5][18] ) );
  AND U986 ( .A(b[17]), .B(a[5]), .Z(\r60/ab[5][17] ) );
  AND U987 ( .A(b[16]), .B(a[5]), .Z(\r60/ab[5][16] ) );
  AND U988 ( .A(b[15]), .B(a[5]), .Z(\r60/ab[5][15] ) );
  AND U989 ( .A(b[14]), .B(a[5]), .Z(\r60/ab[5][14] ) );
  AND U990 ( .A(b[13]), .B(a[5]), .Z(\r60/ab[5][13] ) );
  AND U991 ( .A(b[12]), .B(a[5]), .Z(\r60/ab[5][12] ) );
  AND U992 ( .A(b[11]), .B(a[5]), .Z(\r60/ab[5][11] ) );
  AND U993 ( .A(b[10]), .B(a[5]), .Z(\r60/ab[5][10] ) );
  AND U994 ( .A(b[0]), .B(a[5]), .Z(\r60/ab[5][0] ) );
  AND U995 ( .A(b[9]), .B(a[4]), .Z(\r60/ab[4][9] ) );
  AND U996 ( .A(b[8]), .B(a[4]), .Z(\r60/ab[4][8] ) );
  AND U997 ( .A(b[7]), .B(a[4]), .Z(\r60/ab[4][7] ) );
  AND U998 ( .A(b[6]), .B(a[4]), .Z(\r60/ab[4][6] ) );
  AND U999 ( .A(b[5]), .B(a[4]), .Z(\r60/ab[4][5] ) );
  AND U1000 ( .A(b[4]), .B(a[4]), .Z(\r60/ab[4][4] ) );
  AND U1001 ( .A(b[3]), .B(a[4]), .Z(\r60/ab[4][3] ) );
  MUX U1002 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[4]), .F(\r60/ab[4][31] ) );
  AND U1003 ( .A(b[30]), .B(a[4]), .Z(\r60/ab[4][30] ) );
  AND U1004 ( .A(b[2]), .B(a[4]), .Z(\r60/ab[4][2] ) );
  AND U1005 ( .A(b[29]), .B(a[4]), .Z(\r60/ab[4][29] ) );
  AND U1006 ( .A(b[28]), .B(a[4]), .Z(\r60/ab[4][28] ) );
  AND U1007 ( .A(b[27]), .B(a[4]), .Z(\r60/ab[4][27] ) );
  AND U1008 ( .A(b[26]), .B(a[4]), .Z(\r60/ab[4][26] ) );
  AND U1009 ( .A(b[25]), .B(a[4]), .Z(\r60/ab[4][25] ) );
  AND U1010 ( .A(b[24]), .B(a[4]), .Z(\r60/ab[4][24] ) );
  AND U1011 ( .A(b[23]), .B(a[4]), .Z(\r60/ab[4][23] ) );
  AND U1012 ( .A(b[22]), .B(a[4]), .Z(\r60/ab[4][22] ) );
  AND U1013 ( .A(b[21]), .B(a[4]), .Z(\r60/ab[4][21] ) );
  AND U1014 ( .A(b[20]), .B(a[4]), .Z(\r60/ab[4][20] ) );
  AND U1015 ( .A(b[1]), .B(a[4]), .Z(\r60/ab[4][1] ) );
  AND U1016 ( .A(b[19]), .B(a[4]), .Z(\r60/ab[4][19] ) );
  AND U1017 ( .A(b[18]), .B(a[4]), .Z(\r60/ab[4][18] ) );
  AND U1018 ( .A(b[17]), .B(a[4]), .Z(\r60/ab[4][17] ) );
  AND U1019 ( .A(b[16]), .B(a[4]), .Z(\r60/ab[4][16] ) );
  AND U1020 ( .A(b[15]), .B(a[4]), .Z(\r60/ab[4][15] ) );
  AND U1021 ( .A(b[14]), .B(a[4]), .Z(\r60/ab[4][14] ) );
  AND U1022 ( .A(b[13]), .B(a[4]), .Z(\r60/ab[4][13] ) );
  AND U1023 ( .A(b[12]), .B(a[4]), .Z(\r60/ab[4][12] ) );
  AND U1024 ( .A(b[11]), .B(a[4]), .Z(\r60/ab[4][11] ) );
  AND U1025 ( .A(b[10]), .B(a[4]), .Z(\r60/ab[4][10] ) );
  AND U1026 ( .A(b[0]), .B(a[4]), .Z(\r60/ab[4][0] ) );
  AND U1027 ( .A(b[9]), .B(a[3]), .Z(\r60/ab[3][9] ) );
  AND U1028 ( .A(b[8]), .B(a[3]), .Z(\r60/ab[3][8] ) );
  AND U1029 ( .A(b[7]), .B(a[3]), .Z(\r60/ab[3][7] ) );
  AND U1030 ( .A(b[6]), .B(a[3]), .Z(\r60/ab[3][6] ) );
  AND U1031 ( .A(b[5]), .B(a[3]), .Z(\r60/ab[3][5] ) );
  AND U1032 ( .A(b[4]), .B(a[3]), .Z(\r60/ab[3][4] ) );
  AND U1033 ( .A(b[3]), .B(a[3]), .Z(\r60/ab[3][3] ) );
  MUX U1034 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[3]), .F(\r60/ab[3][31] ) );
  AND U1035 ( .A(b[30]), .B(a[3]), .Z(\r60/ab[3][30] ) );
  AND U1036 ( .A(b[2]), .B(a[3]), .Z(\r60/ab[3][2] ) );
  AND U1037 ( .A(b[29]), .B(a[3]), .Z(\r60/ab[3][29] ) );
  AND U1038 ( .A(b[28]), .B(a[3]), .Z(\r60/ab[3][28] ) );
  AND U1039 ( .A(b[27]), .B(a[3]), .Z(\r60/ab[3][27] ) );
  AND U1040 ( .A(b[26]), .B(a[3]), .Z(\r60/ab[3][26] ) );
  AND U1041 ( .A(b[25]), .B(a[3]), .Z(\r60/ab[3][25] ) );
  AND U1042 ( .A(b[24]), .B(a[3]), .Z(\r60/ab[3][24] ) );
  AND U1043 ( .A(b[23]), .B(a[3]), .Z(\r60/ab[3][23] ) );
  AND U1044 ( .A(b[22]), .B(a[3]), .Z(\r60/ab[3][22] ) );
  AND U1045 ( .A(b[21]), .B(a[3]), .Z(\r60/ab[3][21] ) );
  AND U1046 ( .A(b[20]), .B(a[3]), .Z(\r60/ab[3][20] ) );
  AND U1047 ( .A(b[1]), .B(a[3]), .Z(\r60/ab[3][1] ) );
  AND U1048 ( .A(b[19]), .B(a[3]), .Z(\r60/ab[3][19] ) );
  AND U1049 ( .A(b[18]), .B(a[3]), .Z(\r60/ab[3][18] ) );
  AND U1050 ( .A(b[17]), .B(a[3]), .Z(\r60/ab[3][17] ) );
  AND U1051 ( .A(b[16]), .B(a[3]), .Z(\r60/ab[3][16] ) );
  AND U1052 ( .A(b[15]), .B(a[3]), .Z(\r60/ab[3][15] ) );
  AND U1053 ( .A(b[14]), .B(a[3]), .Z(\r60/ab[3][14] ) );
  AND U1054 ( .A(b[13]), .B(a[3]), .Z(\r60/ab[3][13] ) );
  AND U1055 ( .A(b[12]), .B(a[3]), .Z(\r60/ab[3][12] ) );
  AND U1056 ( .A(b[11]), .B(a[3]), .Z(\r60/ab[3][11] ) );
  AND U1057 ( .A(b[10]), .B(a[3]), .Z(\r60/ab[3][10] ) );
  AND U1058 ( .A(b[0]), .B(a[3]), .Z(\r60/ab[3][0] ) );
  MUX U1059 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[9]), .F(\r60/ab[31][9] ) );
  MUX U1060 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[8]), .F(\r60/ab[31][8] ) );
  MUX U1061 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[7]), .F(\r60/ab[31][7] ) );
  MUX U1062 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[6]), .F(\r60/ab[31][6] ) );
  MUX U1063 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[5]), .F(\r60/ab[31][5] ) );
  MUX U1064 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[4]), .F(\r60/ab[31][4] ) );
  MUX U1065 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[3]), .F(\r60/ab[31][3] ) );
  ANDN U1066 ( .B(b[31]), .A(n682), .Z(\r60/ab[31][31] ) );
  MUX U1067 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[30]), .F(\r60/ab[31][30] ) );
  MUX U1068 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[2]), .F(\r60/ab[31][2] ) );
  MUX U1069 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[29]), .F(\r60/ab[31][29] ) );
  MUX U1070 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[28]), .F(\r60/ab[31][28] ) );
  MUX U1071 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[27]), .F(\r60/ab[31][27] ) );
  MUX U1072 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[26]), .F(\r60/ab[31][26] ) );
  MUX U1073 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[25]), .F(\r60/ab[31][25] ) );
  MUX U1074 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[24]), .F(\r60/ab[31][24] ) );
  MUX U1075 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[23]), .F(\r60/ab[31][23] ) );
  MUX U1076 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[22]), .F(\r60/ab[31][22] ) );
  MUX U1077 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[21]), .F(\r60/ab[31][21] ) );
  MUX U1078 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[20]), .F(\r60/ab[31][20] ) );
  MUX U1079 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[1]), .F(\r60/ab[31][1] ) );
  MUX U1080 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[19]), .F(\r60/ab[31][19] ) );
  MUX U1081 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[18]), .F(\r60/ab[31][18] ) );
  MUX U1082 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[17]), .F(\r60/ab[31][17] ) );
  MUX U1083 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[16]), .F(\r60/ab[31][16] ) );
  MUX U1084 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[15]), .F(\r60/ab[31][15] ) );
  MUX U1085 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[14]), .F(\r60/ab[31][14] ) );
  MUX U1086 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[13]), .F(\r60/ab[31][13] ) );
  MUX U1087 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[12]), .F(\r60/ab[31][12] ) );
  MUX U1088 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[11]), .F(\r60/ab[31][11] ) );
  MUX U1089 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[10]), .F(\r60/ab[31][10] ) );
  MUX U1090 ( .IN0(\r60/ZA ), .IN1(n681), .SEL(b[0]), .F(\r60/ab[31][0] ) );
  NOR U1091 ( .A(n682), .B(\U3/U1/Z_0 ), .Z(n681) );
  AND U1092 ( .A(b[9]), .B(a[30]), .Z(\r60/ab[30][9] ) );
  AND U1093 ( .A(b[8]), .B(a[30]), .Z(\r60/ab[30][8] ) );
  AND U1094 ( .A(b[7]), .B(a[30]), .Z(\r60/ab[30][7] ) );
  AND U1095 ( .A(b[6]), .B(a[30]), .Z(\r60/ab[30][6] ) );
  AND U1096 ( .A(b[5]), .B(a[30]), .Z(\r60/ab[30][5] ) );
  AND U1097 ( .A(b[4]), .B(a[30]), .Z(\r60/ab[30][4] ) );
  AND U1098 ( .A(b[3]), .B(a[30]), .Z(\r60/ab[30][3] ) );
  MUX U1099 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[30]), .F(\r60/ab[30][31] ) );
  AND U1100 ( .A(b[30]), .B(a[30]), .Z(\r60/ab[30][30] ) );
  AND U1101 ( .A(b[2]), .B(a[30]), .Z(\r60/ab[30][2] ) );
  AND U1102 ( .A(b[29]), .B(a[30]), .Z(\r60/ab[30][29] ) );
  AND U1103 ( .A(b[28]), .B(a[30]), .Z(\r60/ab[30][28] ) );
  AND U1104 ( .A(b[27]), .B(a[30]), .Z(\r60/ab[30][27] ) );
  AND U1105 ( .A(b[26]), .B(a[30]), .Z(\r60/ab[30][26] ) );
  AND U1106 ( .A(b[25]), .B(a[30]), .Z(\r60/ab[30][25] ) );
  AND U1107 ( .A(b[24]), .B(a[30]), .Z(\r60/ab[30][24] ) );
  AND U1108 ( .A(b[23]), .B(a[30]), .Z(\r60/ab[30][23] ) );
  AND U1109 ( .A(b[22]), .B(a[30]), .Z(\r60/ab[30][22] ) );
  AND U1110 ( .A(b[21]), .B(a[30]), .Z(\r60/ab[30][21] ) );
  AND U1111 ( .A(b[20]), .B(a[30]), .Z(\r60/ab[30][20] ) );
  AND U1112 ( .A(b[1]), .B(a[30]), .Z(\r60/ab[30][1] ) );
  AND U1113 ( .A(b[19]), .B(a[30]), .Z(\r60/ab[30][19] ) );
  AND U1114 ( .A(b[18]), .B(a[30]), .Z(\r60/ab[30][18] ) );
  AND U1115 ( .A(b[17]), .B(a[30]), .Z(\r60/ab[30][17] ) );
  AND U1116 ( .A(b[16]), .B(a[30]), .Z(\r60/ab[30][16] ) );
  AND U1117 ( .A(b[15]), .B(a[30]), .Z(\r60/ab[30][15] ) );
  AND U1118 ( .A(b[14]), .B(a[30]), .Z(\r60/ab[30][14] ) );
  AND U1119 ( .A(b[13]), .B(a[30]), .Z(\r60/ab[30][13] ) );
  AND U1120 ( .A(b[12]), .B(a[30]), .Z(\r60/ab[30][12] ) );
  AND U1121 ( .A(b[11]), .B(a[30]), .Z(\r60/ab[30][11] ) );
  AND U1122 ( .A(b[10]), .B(a[30]), .Z(\r60/ab[30][10] ) );
  AND U1123 ( .A(b[0]), .B(a[30]), .Z(\r60/ab[30][0] ) );
  AND U1124 ( .A(b[9]), .B(a[2]), .Z(\r60/ab[2][9] ) );
  AND U1125 ( .A(b[8]), .B(a[2]), .Z(\r60/ab[2][8] ) );
  AND U1126 ( .A(b[7]), .B(a[2]), .Z(\r60/ab[2][7] ) );
  AND U1127 ( .A(b[6]), .B(a[2]), .Z(\r60/ab[2][6] ) );
  AND U1128 ( .A(b[5]), .B(a[2]), .Z(\r60/ab[2][5] ) );
  AND U1129 ( .A(b[4]), .B(a[2]), .Z(\r60/ab[2][4] ) );
  AND U1130 ( .A(b[3]), .B(a[2]), .Z(\r60/ab[2][3] ) );
  MUX U1131 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[2]), .F(\r60/ab[2][31] ) );
  AND U1132 ( .A(b[30]), .B(a[2]), .Z(\r60/ab[2][30] ) );
  AND U1133 ( .A(b[2]), .B(a[2]), .Z(\r60/ab[2][2] ) );
  AND U1134 ( .A(b[29]), .B(a[2]), .Z(\r60/ab[2][29] ) );
  AND U1135 ( .A(b[28]), .B(a[2]), .Z(\r60/ab[2][28] ) );
  AND U1136 ( .A(b[27]), .B(a[2]), .Z(\r60/ab[2][27] ) );
  AND U1137 ( .A(b[26]), .B(a[2]), .Z(\r60/ab[2][26] ) );
  AND U1138 ( .A(b[25]), .B(a[2]), .Z(\r60/ab[2][25] ) );
  AND U1139 ( .A(b[24]), .B(a[2]), .Z(\r60/ab[2][24] ) );
  AND U1140 ( .A(b[23]), .B(a[2]), .Z(\r60/ab[2][23] ) );
  AND U1141 ( .A(b[22]), .B(a[2]), .Z(\r60/ab[2][22] ) );
  AND U1142 ( .A(b[21]), .B(a[2]), .Z(\r60/ab[2][21] ) );
  AND U1143 ( .A(b[20]), .B(a[2]), .Z(\r60/ab[2][20] ) );
  AND U1144 ( .A(b[1]), .B(a[2]), .Z(\r60/ab[2][1] ) );
  AND U1145 ( .A(b[19]), .B(a[2]), .Z(\r60/ab[2][19] ) );
  AND U1146 ( .A(b[18]), .B(a[2]), .Z(\r60/ab[2][18] ) );
  AND U1147 ( .A(b[17]), .B(a[2]), .Z(\r60/ab[2][17] ) );
  AND U1148 ( .A(b[16]), .B(a[2]), .Z(\r60/ab[2][16] ) );
  AND U1149 ( .A(b[15]), .B(a[2]), .Z(\r60/ab[2][15] ) );
  AND U1150 ( .A(b[14]), .B(a[2]), .Z(\r60/ab[2][14] ) );
  AND U1151 ( .A(b[13]), .B(a[2]), .Z(\r60/ab[2][13] ) );
  AND U1152 ( .A(b[12]), .B(a[2]), .Z(\r60/ab[2][12] ) );
  AND U1153 ( .A(b[11]), .B(a[2]), .Z(\r60/ab[2][11] ) );
  AND U1154 ( .A(b[10]), .B(a[2]), .Z(\r60/ab[2][10] ) );
  AND U1155 ( .A(b[0]), .B(a[2]), .Z(\r60/ab[2][0] ) );
  AND U1156 ( .A(b[9]), .B(a[29]), .Z(\r60/ab[29][9] ) );
  AND U1157 ( .A(b[8]), .B(a[29]), .Z(\r60/ab[29][8] ) );
  AND U1158 ( .A(b[7]), .B(a[29]), .Z(\r60/ab[29][7] ) );
  AND U1159 ( .A(b[6]), .B(a[29]), .Z(\r60/ab[29][6] ) );
  AND U1160 ( .A(b[5]), .B(a[29]), .Z(\r60/ab[29][5] ) );
  AND U1161 ( .A(b[4]), .B(a[29]), .Z(\r60/ab[29][4] ) );
  AND U1162 ( .A(b[3]), .B(a[29]), .Z(\r60/ab[29][3] ) );
  MUX U1163 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[29]), .F(\r60/ab[29][31] ) );
  AND U1164 ( .A(b[30]), .B(a[29]), .Z(\r60/ab[29][30] ) );
  AND U1165 ( .A(b[2]), .B(a[29]), .Z(\r60/ab[29][2] ) );
  AND U1166 ( .A(b[29]), .B(a[29]), .Z(\r60/ab[29][29] ) );
  AND U1167 ( .A(b[28]), .B(a[29]), .Z(\r60/ab[29][28] ) );
  AND U1168 ( .A(b[27]), .B(a[29]), .Z(\r60/ab[29][27] ) );
  AND U1169 ( .A(b[26]), .B(a[29]), .Z(\r60/ab[29][26] ) );
  AND U1170 ( .A(b[25]), .B(a[29]), .Z(\r60/ab[29][25] ) );
  AND U1171 ( .A(b[24]), .B(a[29]), .Z(\r60/ab[29][24] ) );
  AND U1172 ( .A(b[23]), .B(a[29]), .Z(\r60/ab[29][23] ) );
  AND U1173 ( .A(b[22]), .B(a[29]), .Z(\r60/ab[29][22] ) );
  AND U1174 ( .A(b[21]), .B(a[29]), .Z(\r60/ab[29][21] ) );
  AND U1175 ( .A(b[20]), .B(a[29]), .Z(\r60/ab[29][20] ) );
  AND U1176 ( .A(b[1]), .B(a[29]), .Z(\r60/ab[29][1] ) );
  AND U1177 ( .A(b[19]), .B(a[29]), .Z(\r60/ab[29][19] ) );
  AND U1178 ( .A(b[18]), .B(a[29]), .Z(\r60/ab[29][18] ) );
  AND U1179 ( .A(b[17]), .B(a[29]), .Z(\r60/ab[29][17] ) );
  AND U1180 ( .A(b[16]), .B(a[29]), .Z(\r60/ab[29][16] ) );
  AND U1181 ( .A(b[15]), .B(a[29]), .Z(\r60/ab[29][15] ) );
  AND U1182 ( .A(b[14]), .B(a[29]), .Z(\r60/ab[29][14] ) );
  AND U1183 ( .A(b[13]), .B(a[29]), .Z(\r60/ab[29][13] ) );
  AND U1184 ( .A(b[12]), .B(a[29]), .Z(\r60/ab[29][12] ) );
  AND U1185 ( .A(b[11]), .B(a[29]), .Z(\r60/ab[29][11] ) );
  AND U1186 ( .A(b[10]), .B(a[29]), .Z(\r60/ab[29][10] ) );
  AND U1187 ( .A(b[0]), .B(a[29]), .Z(\r60/ab[29][0] ) );
  AND U1188 ( .A(b[9]), .B(a[28]), .Z(\r60/ab[28][9] ) );
  AND U1189 ( .A(b[8]), .B(a[28]), .Z(\r60/ab[28][8] ) );
  AND U1190 ( .A(b[7]), .B(a[28]), .Z(\r60/ab[28][7] ) );
  AND U1191 ( .A(b[6]), .B(a[28]), .Z(\r60/ab[28][6] ) );
  AND U1192 ( .A(b[5]), .B(a[28]), .Z(\r60/ab[28][5] ) );
  AND U1193 ( .A(b[4]), .B(a[28]), .Z(\r60/ab[28][4] ) );
  AND U1194 ( .A(b[3]), .B(a[28]), .Z(\r60/ab[28][3] ) );
  MUX U1195 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[28]), .F(\r60/ab[28][31] ) );
  AND U1196 ( .A(b[30]), .B(a[28]), .Z(\r60/ab[28][30] ) );
  AND U1197 ( .A(b[2]), .B(a[28]), .Z(\r60/ab[28][2] ) );
  AND U1198 ( .A(b[29]), .B(a[28]), .Z(\r60/ab[28][29] ) );
  AND U1199 ( .A(b[28]), .B(a[28]), .Z(\r60/ab[28][28] ) );
  AND U1200 ( .A(b[27]), .B(a[28]), .Z(\r60/ab[28][27] ) );
  AND U1201 ( .A(b[26]), .B(a[28]), .Z(\r60/ab[28][26] ) );
  AND U1202 ( .A(b[25]), .B(a[28]), .Z(\r60/ab[28][25] ) );
  AND U1203 ( .A(b[24]), .B(a[28]), .Z(\r60/ab[28][24] ) );
  AND U1204 ( .A(b[23]), .B(a[28]), .Z(\r60/ab[28][23] ) );
  AND U1205 ( .A(b[22]), .B(a[28]), .Z(\r60/ab[28][22] ) );
  AND U1206 ( .A(b[21]), .B(a[28]), .Z(\r60/ab[28][21] ) );
  AND U1207 ( .A(b[20]), .B(a[28]), .Z(\r60/ab[28][20] ) );
  AND U1208 ( .A(b[1]), .B(a[28]), .Z(\r60/ab[28][1] ) );
  AND U1209 ( .A(b[19]), .B(a[28]), .Z(\r60/ab[28][19] ) );
  AND U1210 ( .A(b[18]), .B(a[28]), .Z(\r60/ab[28][18] ) );
  AND U1211 ( .A(b[17]), .B(a[28]), .Z(\r60/ab[28][17] ) );
  AND U1212 ( .A(b[16]), .B(a[28]), .Z(\r60/ab[28][16] ) );
  AND U1213 ( .A(b[15]), .B(a[28]), .Z(\r60/ab[28][15] ) );
  AND U1214 ( .A(b[14]), .B(a[28]), .Z(\r60/ab[28][14] ) );
  AND U1215 ( .A(b[13]), .B(a[28]), .Z(\r60/ab[28][13] ) );
  AND U1216 ( .A(b[12]), .B(a[28]), .Z(\r60/ab[28][12] ) );
  AND U1217 ( .A(b[11]), .B(a[28]), .Z(\r60/ab[28][11] ) );
  AND U1218 ( .A(b[10]), .B(a[28]), .Z(\r60/ab[28][10] ) );
  AND U1219 ( .A(b[0]), .B(a[28]), .Z(\r60/ab[28][0] ) );
  AND U1220 ( .A(b[9]), .B(a[27]), .Z(\r60/ab[27][9] ) );
  AND U1221 ( .A(b[8]), .B(a[27]), .Z(\r60/ab[27][8] ) );
  AND U1222 ( .A(b[7]), .B(a[27]), .Z(\r60/ab[27][7] ) );
  AND U1223 ( .A(b[6]), .B(a[27]), .Z(\r60/ab[27][6] ) );
  AND U1224 ( .A(b[5]), .B(a[27]), .Z(\r60/ab[27][5] ) );
  AND U1225 ( .A(b[4]), .B(a[27]), .Z(\r60/ab[27][4] ) );
  AND U1226 ( .A(b[3]), .B(a[27]), .Z(\r60/ab[27][3] ) );
  MUX U1227 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[27]), .F(\r60/ab[27][31] ) );
  AND U1228 ( .A(b[30]), .B(a[27]), .Z(\r60/ab[27][30] ) );
  AND U1229 ( .A(b[2]), .B(a[27]), .Z(\r60/ab[27][2] ) );
  AND U1230 ( .A(b[29]), .B(a[27]), .Z(\r60/ab[27][29] ) );
  AND U1231 ( .A(b[28]), .B(a[27]), .Z(\r60/ab[27][28] ) );
  AND U1232 ( .A(b[27]), .B(a[27]), .Z(\r60/ab[27][27] ) );
  AND U1233 ( .A(b[26]), .B(a[27]), .Z(\r60/ab[27][26] ) );
  AND U1234 ( .A(b[25]), .B(a[27]), .Z(\r60/ab[27][25] ) );
  AND U1235 ( .A(b[24]), .B(a[27]), .Z(\r60/ab[27][24] ) );
  AND U1236 ( .A(b[23]), .B(a[27]), .Z(\r60/ab[27][23] ) );
  AND U1237 ( .A(b[22]), .B(a[27]), .Z(\r60/ab[27][22] ) );
  AND U1238 ( .A(b[21]), .B(a[27]), .Z(\r60/ab[27][21] ) );
  AND U1239 ( .A(b[20]), .B(a[27]), .Z(\r60/ab[27][20] ) );
  AND U1240 ( .A(b[1]), .B(a[27]), .Z(\r60/ab[27][1] ) );
  AND U1241 ( .A(b[19]), .B(a[27]), .Z(\r60/ab[27][19] ) );
  AND U1242 ( .A(b[18]), .B(a[27]), .Z(\r60/ab[27][18] ) );
  AND U1243 ( .A(b[17]), .B(a[27]), .Z(\r60/ab[27][17] ) );
  AND U1244 ( .A(b[16]), .B(a[27]), .Z(\r60/ab[27][16] ) );
  AND U1245 ( .A(b[15]), .B(a[27]), .Z(\r60/ab[27][15] ) );
  AND U1246 ( .A(b[14]), .B(a[27]), .Z(\r60/ab[27][14] ) );
  AND U1247 ( .A(b[13]), .B(a[27]), .Z(\r60/ab[27][13] ) );
  AND U1248 ( .A(b[12]), .B(a[27]), .Z(\r60/ab[27][12] ) );
  AND U1249 ( .A(b[11]), .B(a[27]), .Z(\r60/ab[27][11] ) );
  AND U1250 ( .A(b[10]), .B(a[27]), .Z(\r60/ab[27][10] ) );
  AND U1251 ( .A(b[0]), .B(a[27]), .Z(\r60/ab[27][0] ) );
  AND U1252 ( .A(b[9]), .B(a[26]), .Z(\r60/ab[26][9] ) );
  AND U1253 ( .A(b[8]), .B(a[26]), .Z(\r60/ab[26][8] ) );
  AND U1254 ( .A(b[7]), .B(a[26]), .Z(\r60/ab[26][7] ) );
  AND U1255 ( .A(b[6]), .B(a[26]), .Z(\r60/ab[26][6] ) );
  AND U1256 ( .A(b[5]), .B(a[26]), .Z(\r60/ab[26][5] ) );
  AND U1257 ( .A(b[4]), .B(a[26]), .Z(\r60/ab[26][4] ) );
  AND U1258 ( .A(b[3]), .B(a[26]), .Z(\r60/ab[26][3] ) );
  MUX U1259 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[26]), .F(\r60/ab[26][31] ) );
  AND U1260 ( .A(b[30]), .B(a[26]), .Z(\r60/ab[26][30] ) );
  AND U1261 ( .A(b[2]), .B(a[26]), .Z(\r60/ab[26][2] ) );
  AND U1262 ( .A(b[29]), .B(a[26]), .Z(\r60/ab[26][29] ) );
  AND U1263 ( .A(b[28]), .B(a[26]), .Z(\r60/ab[26][28] ) );
  AND U1264 ( .A(b[27]), .B(a[26]), .Z(\r60/ab[26][27] ) );
  AND U1265 ( .A(b[26]), .B(a[26]), .Z(\r60/ab[26][26] ) );
  AND U1266 ( .A(b[25]), .B(a[26]), .Z(\r60/ab[26][25] ) );
  AND U1267 ( .A(b[24]), .B(a[26]), .Z(\r60/ab[26][24] ) );
  AND U1268 ( .A(b[23]), .B(a[26]), .Z(\r60/ab[26][23] ) );
  AND U1269 ( .A(b[22]), .B(a[26]), .Z(\r60/ab[26][22] ) );
  AND U1270 ( .A(b[21]), .B(a[26]), .Z(\r60/ab[26][21] ) );
  AND U1271 ( .A(b[20]), .B(a[26]), .Z(\r60/ab[26][20] ) );
  AND U1272 ( .A(b[1]), .B(a[26]), .Z(\r60/ab[26][1] ) );
  AND U1273 ( .A(b[19]), .B(a[26]), .Z(\r60/ab[26][19] ) );
  AND U1274 ( .A(b[18]), .B(a[26]), .Z(\r60/ab[26][18] ) );
  AND U1275 ( .A(b[17]), .B(a[26]), .Z(\r60/ab[26][17] ) );
  AND U1276 ( .A(b[16]), .B(a[26]), .Z(\r60/ab[26][16] ) );
  AND U1277 ( .A(b[15]), .B(a[26]), .Z(\r60/ab[26][15] ) );
  AND U1278 ( .A(b[14]), .B(a[26]), .Z(\r60/ab[26][14] ) );
  AND U1279 ( .A(b[13]), .B(a[26]), .Z(\r60/ab[26][13] ) );
  AND U1280 ( .A(b[12]), .B(a[26]), .Z(\r60/ab[26][12] ) );
  AND U1281 ( .A(b[11]), .B(a[26]), .Z(\r60/ab[26][11] ) );
  AND U1282 ( .A(b[10]), .B(a[26]), .Z(\r60/ab[26][10] ) );
  AND U1283 ( .A(b[0]), .B(a[26]), .Z(\r60/ab[26][0] ) );
  AND U1284 ( .A(b[9]), .B(a[25]), .Z(\r60/ab[25][9] ) );
  AND U1285 ( .A(b[8]), .B(a[25]), .Z(\r60/ab[25][8] ) );
  AND U1286 ( .A(b[7]), .B(a[25]), .Z(\r60/ab[25][7] ) );
  AND U1287 ( .A(b[6]), .B(a[25]), .Z(\r60/ab[25][6] ) );
  AND U1288 ( .A(b[5]), .B(a[25]), .Z(\r60/ab[25][5] ) );
  AND U1289 ( .A(b[4]), .B(a[25]), .Z(\r60/ab[25][4] ) );
  AND U1290 ( .A(b[3]), .B(a[25]), .Z(\r60/ab[25][3] ) );
  MUX U1291 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[25]), .F(\r60/ab[25][31] ) );
  AND U1292 ( .A(b[30]), .B(a[25]), .Z(\r60/ab[25][30] ) );
  AND U1293 ( .A(b[2]), .B(a[25]), .Z(\r60/ab[25][2] ) );
  AND U1294 ( .A(b[29]), .B(a[25]), .Z(\r60/ab[25][29] ) );
  AND U1295 ( .A(b[28]), .B(a[25]), .Z(\r60/ab[25][28] ) );
  AND U1296 ( .A(b[27]), .B(a[25]), .Z(\r60/ab[25][27] ) );
  AND U1297 ( .A(b[26]), .B(a[25]), .Z(\r60/ab[25][26] ) );
  AND U1298 ( .A(b[25]), .B(a[25]), .Z(\r60/ab[25][25] ) );
  AND U1299 ( .A(b[24]), .B(a[25]), .Z(\r60/ab[25][24] ) );
  AND U1300 ( .A(b[23]), .B(a[25]), .Z(\r60/ab[25][23] ) );
  AND U1301 ( .A(b[22]), .B(a[25]), .Z(\r60/ab[25][22] ) );
  AND U1302 ( .A(b[21]), .B(a[25]), .Z(\r60/ab[25][21] ) );
  AND U1303 ( .A(b[20]), .B(a[25]), .Z(\r60/ab[25][20] ) );
  AND U1304 ( .A(b[1]), .B(a[25]), .Z(\r60/ab[25][1] ) );
  AND U1305 ( .A(b[19]), .B(a[25]), .Z(\r60/ab[25][19] ) );
  AND U1306 ( .A(b[18]), .B(a[25]), .Z(\r60/ab[25][18] ) );
  AND U1307 ( .A(b[17]), .B(a[25]), .Z(\r60/ab[25][17] ) );
  AND U1308 ( .A(b[16]), .B(a[25]), .Z(\r60/ab[25][16] ) );
  AND U1309 ( .A(b[15]), .B(a[25]), .Z(\r60/ab[25][15] ) );
  AND U1310 ( .A(b[14]), .B(a[25]), .Z(\r60/ab[25][14] ) );
  AND U1311 ( .A(b[13]), .B(a[25]), .Z(\r60/ab[25][13] ) );
  AND U1312 ( .A(b[12]), .B(a[25]), .Z(\r60/ab[25][12] ) );
  AND U1313 ( .A(b[11]), .B(a[25]), .Z(\r60/ab[25][11] ) );
  AND U1314 ( .A(b[10]), .B(a[25]), .Z(\r60/ab[25][10] ) );
  AND U1315 ( .A(b[0]), .B(a[25]), .Z(\r60/ab[25][0] ) );
  AND U1316 ( .A(b[9]), .B(a[24]), .Z(\r60/ab[24][9] ) );
  AND U1317 ( .A(b[8]), .B(a[24]), .Z(\r60/ab[24][8] ) );
  AND U1318 ( .A(b[7]), .B(a[24]), .Z(\r60/ab[24][7] ) );
  AND U1319 ( .A(b[6]), .B(a[24]), .Z(\r60/ab[24][6] ) );
  AND U1320 ( .A(b[5]), .B(a[24]), .Z(\r60/ab[24][5] ) );
  AND U1321 ( .A(b[4]), .B(a[24]), .Z(\r60/ab[24][4] ) );
  AND U1322 ( .A(b[3]), .B(a[24]), .Z(\r60/ab[24][3] ) );
  MUX U1323 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[24]), .F(\r60/ab[24][31] ) );
  AND U1324 ( .A(b[30]), .B(a[24]), .Z(\r60/ab[24][30] ) );
  AND U1325 ( .A(b[2]), .B(a[24]), .Z(\r60/ab[24][2] ) );
  AND U1326 ( .A(b[29]), .B(a[24]), .Z(\r60/ab[24][29] ) );
  AND U1327 ( .A(b[28]), .B(a[24]), .Z(\r60/ab[24][28] ) );
  AND U1328 ( .A(b[27]), .B(a[24]), .Z(\r60/ab[24][27] ) );
  AND U1329 ( .A(b[26]), .B(a[24]), .Z(\r60/ab[24][26] ) );
  AND U1330 ( .A(b[25]), .B(a[24]), .Z(\r60/ab[24][25] ) );
  AND U1331 ( .A(b[24]), .B(a[24]), .Z(\r60/ab[24][24] ) );
  AND U1332 ( .A(b[23]), .B(a[24]), .Z(\r60/ab[24][23] ) );
  AND U1333 ( .A(b[22]), .B(a[24]), .Z(\r60/ab[24][22] ) );
  AND U1334 ( .A(b[21]), .B(a[24]), .Z(\r60/ab[24][21] ) );
  AND U1335 ( .A(b[20]), .B(a[24]), .Z(\r60/ab[24][20] ) );
  AND U1336 ( .A(b[1]), .B(a[24]), .Z(\r60/ab[24][1] ) );
  AND U1337 ( .A(b[19]), .B(a[24]), .Z(\r60/ab[24][19] ) );
  AND U1338 ( .A(b[18]), .B(a[24]), .Z(\r60/ab[24][18] ) );
  AND U1339 ( .A(b[17]), .B(a[24]), .Z(\r60/ab[24][17] ) );
  AND U1340 ( .A(b[16]), .B(a[24]), .Z(\r60/ab[24][16] ) );
  AND U1341 ( .A(b[15]), .B(a[24]), .Z(\r60/ab[24][15] ) );
  AND U1342 ( .A(b[14]), .B(a[24]), .Z(\r60/ab[24][14] ) );
  AND U1343 ( .A(b[13]), .B(a[24]), .Z(\r60/ab[24][13] ) );
  AND U1344 ( .A(b[12]), .B(a[24]), .Z(\r60/ab[24][12] ) );
  AND U1345 ( .A(b[11]), .B(a[24]), .Z(\r60/ab[24][11] ) );
  AND U1346 ( .A(b[10]), .B(a[24]), .Z(\r60/ab[24][10] ) );
  AND U1347 ( .A(b[0]), .B(a[24]), .Z(\r60/ab[24][0] ) );
  AND U1348 ( .A(b[9]), .B(a[23]), .Z(\r60/ab[23][9] ) );
  AND U1349 ( .A(b[8]), .B(a[23]), .Z(\r60/ab[23][8] ) );
  AND U1350 ( .A(b[7]), .B(a[23]), .Z(\r60/ab[23][7] ) );
  AND U1351 ( .A(b[6]), .B(a[23]), .Z(\r60/ab[23][6] ) );
  AND U1352 ( .A(b[5]), .B(a[23]), .Z(\r60/ab[23][5] ) );
  AND U1353 ( .A(b[4]), .B(a[23]), .Z(\r60/ab[23][4] ) );
  AND U1354 ( .A(b[3]), .B(a[23]), .Z(\r60/ab[23][3] ) );
  MUX U1355 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[23]), .F(\r60/ab[23][31] ) );
  AND U1356 ( .A(b[30]), .B(a[23]), .Z(\r60/ab[23][30] ) );
  AND U1357 ( .A(b[2]), .B(a[23]), .Z(\r60/ab[23][2] ) );
  AND U1358 ( .A(b[29]), .B(a[23]), .Z(\r60/ab[23][29] ) );
  AND U1359 ( .A(b[28]), .B(a[23]), .Z(\r60/ab[23][28] ) );
  AND U1360 ( .A(b[27]), .B(a[23]), .Z(\r60/ab[23][27] ) );
  AND U1361 ( .A(b[26]), .B(a[23]), .Z(\r60/ab[23][26] ) );
  AND U1362 ( .A(b[25]), .B(a[23]), .Z(\r60/ab[23][25] ) );
  AND U1363 ( .A(b[24]), .B(a[23]), .Z(\r60/ab[23][24] ) );
  AND U1364 ( .A(b[23]), .B(a[23]), .Z(\r60/ab[23][23] ) );
  AND U1365 ( .A(b[22]), .B(a[23]), .Z(\r60/ab[23][22] ) );
  AND U1366 ( .A(b[21]), .B(a[23]), .Z(\r60/ab[23][21] ) );
  AND U1367 ( .A(b[20]), .B(a[23]), .Z(\r60/ab[23][20] ) );
  AND U1368 ( .A(b[1]), .B(a[23]), .Z(\r60/ab[23][1] ) );
  AND U1369 ( .A(b[19]), .B(a[23]), .Z(\r60/ab[23][19] ) );
  AND U1370 ( .A(b[18]), .B(a[23]), .Z(\r60/ab[23][18] ) );
  AND U1371 ( .A(b[17]), .B(a[23]), .Z(\r60/ab[23][17] ) );
  AND U1372 ( .A(b[16]), .B(a[23]), .Z(\r60/ab[23][16] ) );
  AND U1373 ( .A(b[15]), .B(a[23]), .Z(\r60/ab[23][15] ) );
  AND U1374 ( .A(b[14]), .B(a[23]), .Z(\r60/ab[23][14] ) );
  AND U1375 ( .A(b[13]), .B(a[23]), .Z(\r60/ab[23][13] ) );
  AND U1376 ( .A(b[12]), .B(a[23]), .Z(\r60/ab[23][12] ) );
  AND U1377 ( .A(b[11]), .B(a[23]), .Z(\r60/ab[23][11] ) );
  AND U1378 ( .A(b[10]), .B(a[23]), .Z(\r60/ab[23][10] ) );
  AND U1379 ( .A(b[0]), .B(a[23]), .Z(\r60/ab[23][0] ) );
  AND U1380 ( .A(b[9]), .B(a[22]), .Z(\r60/ab[22][9] ) );
  AND U1381 ( .A(b[8]), .B(a[22]), .Z(\r60/ab[22][8] ) );
  AND U1382 ( .A(b[7]), .B(a[22]), .Z(\r60/ab[22][7] ) );
  AND U1383 ( .A(b[6]), .B(a[22]), .Z(\r60/ab[22][6] ) );
  AND U1384 ( .A(b[5]), .B(a[22]), .Z(\r60/ab[22][5] ) );
  AND U1385 ( .A(b[4]), .B(a[22]), .Z(\r60/ab[22][4] ) );
  AND U1386 ( .A(b[3]), .B(a[22]), .Z(\r60/ab[22][3] ) );
  MUX U1387 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[22]), .F(\r60/ab[22][31] ) );
  AND U1388 ( .A(b[30]), .B(a[22]), .Z(\r60/ab[22][30] ) );
  AND U1389 ( .A(b[2]), .B(a[22]), .Z(\r60/ab[22][2] ) );
  AND U1390 ( .A(b[29]), .B(a[22]), .Z(\r60/ab[22][29] ) );
  AND U1391 ( .A(b[28]), .B(a[22]), .Z(\r60/ab[22][28] ) );
  AND U1392 ( .A(b[27]), .B(a[22]), .Z(\r60/ab[22][27] ) );
  AND U1393 ( .A(b[26]), .B(a[22]), .Z(\r60/ab[22][26] ) );
  AND U1394 ( .A(b[25]), .B(a[22]), .Z(\r60/ab[22][25] ) );
  AND U1395 ( .A(b[24]), .B(a[22]), .Z(\r60/ab[22][24] ) );
  AND U1396 ( .A(b[23]), .B(a[22]), .Z(\r60/ab[22][23] ) );
  AND U1397 ( .A(b[22]), .B(a[22]), .Z(\r60/ab[22][22] ) );
  AND U1398 ( .A(b[21]), .B(a[22]), .Z(\r60/ab[22][21] ) );
  AND U1399 ( .A(b[20]), .B(a[22]), .Z(\r60/ab[22][20] ) );
  AND U1400 ( .A(b[1]), .B(a[22]), .Z(\r60/ab[22][1] ) );
  AND U1401 ( .A(b[19]), .B(a[22]), .Z(\r60/ab[22][19] ) );
  AND U1402 ( .A(b[18]), .B(a[22]), .Z(\r60/ab[22][18] ) );
  AND U1403 ( .A(b[17]), .B(a[22]), .Z(\r60/ab[22][17] ) );
  AND U1404 ( .A(b[16]), .B(a[22]), .Z(\r60/ab[22][16] ) );
  AND U1405 ( .A(b[15]), .B(a[22]), .Z(\r60/ab[22][15] ) );
  AND U1406 ( .A(b[14]), .B(a[22]), .Z(\r60/ab[22][14] ) );
  AND U1407 ( .A(b[13]), .B(a[22]), .Z(\r60/ab[22][13] ) );
  AND U1408 ( .A(b[12]), .B(a[22]), .Z(\r60/ab[22][12] ) );
  AND U1409 ( .A(b[11]), .B(a[22]), .Z(\r60/ab[22][11] ) );
  AND U1410 ( .A(b[10]), .B(a[22]), .Z(\r60/ab[22][10] ) );
  AND U1411 ( .A(b[0]), .B(a[22]), .Z(\r60/ab[22][0] ) );
  AND U1412 ( .A(b[9]), .B(a[21]), .Z(\r60/ab[21][9] ) );
  AND U1413 ( .A(b[8]), .B(a[21]), .Z(\r60/ab[21][8] ) );
  AND U1414 ( .A(b[7]), .B(a[21]), .Z(\r60/ab[21][7] ) );
  AND U1415 ( .A(b[6]), .B(a[21]), .Z(\r60/ab[21][6] ) );
  AND U1416 ( .A(b[5]), .B(a[21]), .Z(\r60/ab[21][5] ) );
  AND U1417 ( .A(b[4]), .B(a[21]), .Z(\r60/ab[21][4] ) );
  AND U1418 ( .A(b[3]), .B(a[21]), .Z(\r60/ab[21][3] ) );
  MUX U1419 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[21]), .F(\r60/ab[21][31] ) );
  AND U1420 ( .A(b[30]), .B(a[21]), .Z(\r60/ab[21][30] ) );
  AND U1421 ( .A(b[2]), .B(a[21]), .Z(\r60/ab[21][2] ) );
  AND U1422 ( .A(b[29]), .B(a[21]), .Z(\r60/ab[21][29] ) );
  AND U1423 ( .A(b[28]), .B(a[21]), .Z(\r60/ab[21][28] ) );
  AND U1424 ( .A(b[27]), .B(a[21]), .Z(\r60/ab[21][27] ) );
  AND U1425 ( .A(b[26]), .B(a[21]), .Z(\r60/ab[21][26] ) );
  AND U1426 ( .A(b[25]), .B(a[21]), .Z(\r60/ab[21][25] ) );
  AND U1427 ( .A(b[24]), .B(a[21]), .Z(\r60/ab[21][24] ) );
  AND U1428 ( .A(b[23]), .B(a[21]), .Z(\r60/ab[21][23] ) );
  AND U1429 ( .A(b[22]), .B(a[21]), .Z(\r60/ab[21][22] ) );
  AND U1430 ( .A(b[21]), .B(a[21]), .Z(\r60/ab[21][21] ) );
  AND U1431 ( .A(b[20]), .B(a[21]), .Z(\r60/ab[21][20] ) );
  AND U1432 ( .A(b[1]), .B(a[21]), .Z(\r60/ab[21][1] ) );
  AND U1433 ( .A(b[19]), .B(a[21]), .Z(\r60/ab[21][19] ) );
  AND U1434 ( .A(b[18]), .B(a[21]), .Z(\r60/ab[21][18] ) );
  AND U1435 ( .A(b[17]), .B(a[21]), .Z(\r60/ab[21][17] ) );
  AND U1436 ( .A(b[16]), .B(a[21]), .Z(\r60/ab[21][16] ) );
  AND U1437 ( .A(b[15]), .B(a[21]), .Z(\r60/ab[21][15] ) );
  AND U1438 ( .A(b[14]), .B(a[21]), .Z(\r60/ab[21][14] ) );
  AND U1439 ( .A(b[13]), .B(a[21]), .Z(\r60/ab[21][13] ) );
  AND U1440 ( .A(b[12]), .B(a[21]), .Z(\r60/ab[21][12] ) );
  AND U1441 ( .A(b[11]), .B(a[21]), .Z(\r60/ab[21][11] ) );
  AND U1442 ( .A(b[10]), .B(a[21]), .Z(\r60/ab[21][10] ) );
  AND U1443 ( .A(b[0]), .B(a[21]), .Z(\r60/ab[21][0] ) );
  AND U1444 ( .A(b[9]), .B(a[20]), .Z(\r60/ab[20][9] ) );
  AND U1445 ( .A(b[8]), .B(a[20]), .Z(\r60/ab[20][8] ) );
  AND U1446 ( .A(b[7]), .B(a[20]), .Z(\r60/ab[20][7] ) );
  AND U1447 ( .A(b[6]), .B(a[20]), .Z(\r60/ab[20][6] ) );
  AND U1448 ( .A(b[5]), .B(a[20]), .Z(\r60/ab[20][5] ) );
  AND U1449 ( .A(b[4]), .B(a[20]), .Z(\r60/ab[20][4] ) );
  AND U1450 ( .A(b[3]), .B(a[20]), .Z(\r60/ab[20][3] ) );
  MUX U1451 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[20]), .F(\r60/ab[20][31] ) );
  AND U1452 ( .A(b[30]), .B(a[20]), .Z(\r60/ab[20][30] ) );
  AND U1453 ( .A(b[2]), .B(a[20]), .Z(\r60/ab[20][2] ) );
  AND U1454 ( .A(b[29]), .B(a[20]), .Z(\r60/ab[20][29] ) );
  AND U1455 ( .A(b[28]), .B(a[20]), .Z(\r60/ab[20][28] ) );
  AND U1456 ( .A(b[27]), .B(a[20]), .Z(\r60/ab[20][27] ) );
  AND U1457 ( .A(b[26]), .B(a[20]), .Z(\r60/ab[20][26] ) );
  AND U1458 ( .A(b[25]), .B(a[20]), .Z(\r60/ab[20][25] ) );
  AND U1459 ( .A(b[24]), .B(a[20]), .Z(\r60/ab[20][24] ) );
  AND U1460 ( .A(b[23]), .B(a[20]), .Z(\r60/ab[20][23] ) );
  AND U1461 ( .A(b[22]), .B(a[20]), .Z(\r60/ab[20][22] ) );
  AND U1462 ( .A(b[21]), .B(a[20]), .Z(\r60/ab[20][21] ) );
  AND U1463 ( .A(b[20]), .B(a[20]), .Z(\r60/ab[20][20] ) );
  AND U1464 ( .A(b[1]), .B(a[20]), .Z(\r60/ab[20][1] ) );
  AND U1465 ( .A(b[19]), .B(a[20]), .Z(\r60/ab[20][19] ) );
  AND U1466 ( .A(b[18]), .B(a[20]), .Z(\r60/ab[20][18] ) );
  AND U1467 ( .A(b[17]), .B(a[20]), .Z(\r60/ab[20][17] ) );
  AND U1468 ( .A(b[16]), .B(a[20]), .Z(\r60/ab[20][16] ) );
  AND U1469 ( .A(b[15]), .B(a[20]), .Z(\r60/ab[20][15] ) );
  AND U1470 ( .A(b[14]), .B(a[20]), .Z(\r60/ab[20][14] ) );
  AND U1471 ( .A(b[13]), .B(a[20]), .Z(\r60/ab[20][13] ) );
  AND U1472 ( .A(b[12]), .B(a[20]), .Z(\r60/ab[20][12] ) );
  AND U1473 ( .A(b[11]), .B(a[20]), .Z(\r60/ab[20][11] ) );
  AND U1474 ( .A(b[10]), .B(a[20]), .Z(\r60/ab[20][10] ) );
  AND U1475 ( .A(b[0]), .B(a[20]), .Z(\r60/ab[20][0] ) );
  AND U1476 ( .A(b[9]), .B(a[1]), .Z(\r60/ab[1][9] ) );
  AND U1477 ( .A(b[8]), .B(a[1]), .Z(\r60/ab[1][8] ) );
  AND U1478 ( .A(b[7]), .B(a[1]), .Z(\r60/ab[1][7] ) );
  AND U1479 ( .A(b[6]), .B(a[1]), .Z(\r60/ab[1][6] ) );
  AND U1480 ( .A(b[5]), .B(a[1]), .Z(\r60/ab[1][5] ) );
  AND U1481 ( .A(b[4]), .B(a[1]), .Z(\r60/ab[1][4] ) );
  AND U1482 ( .A(b[3]), .B(a[1]), .Z(\r60/ab[1][3] ) );
  MUX U1483 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[1]), .F(\r60/ab[1][31] ) );
  AND U1484 ( .A(b[30]), .B(a[1]), .Z(\r60/ab[1][30] ) );
  AND U1485 ( .A(b[2]), .B(a[1]), .Z(\r60/ab[1][2] ) );
  AND U1486 ( .A(b[29]), .B(a[1]), .Z(\r60/ab[1][29] ) );
  AND U1487 ( .A(b[28]), .B(a[1]), .Z(\r60/ab[1][28] ) );
  AND U1488 ( .A(b[27]), .B(a[1]), .Z(\r60/ab[1][27] ) );
  AND U1489 ( .A(b[26]), .B(a[1]), .Z(\r60/ab[1][26] ) );
  AND U1490 ( .A(b[25]), .B(a[1]), .Z(\r60/ab[1][25] ) );
  AND U1491 ( .A(b[24]), .B(a[1]), .Z(\r60/ab[1][24] ) );
  AND U1492 ( .A(b[23]), .B(a[1]), .Z(\r60/ab[1][23] ) );
  AND U1493 ( .A(b[22]), .B(a[1]), .Z(\r60/ab[1][22] ) );
  AND U1494 ( .A(b[21]), .B(a[1]), .Z(\r60/ab[1][21] ) );
  AND U1495 ( .A(b[20]), .B(a[1]), .Z(\r60/ab[1][20] ) );
  AND U1496 ( .A(b[1]), .B(a[1]), .Z(\r60/ab[1][1] ) );
  AND U1497 ( .A(b[19]), .B(a[1]), .Z(\r60/ab[1][19] ) );
  AND U1498 ( .A(b[18]), .B(a[1]), .Z(\r60/ab[1][18] ) );
  AND U1499 ( .A(b[17]), .B(a[1]), .Z(\r60/ab[1][17] ) );
  AND U1500 ( .A(b[16]), .B(a[1]), .Z(\r60/ab[1][16] ) );
  AND U1501 ( .A(b[15]), .B(a[1]), .Z(\r60/ab[1][15] ) );
  AND U1502 ( .A(b[14]), .B(a[1]), .Z(\r60/ab[1][14] ) );
  AND U1503 ( .A(b[13]), .B(a[1]), .Z(\r60/ab[1][13] ) );
  AND U1504 ( .A(b[12]), .B(a[1]), .Z(\r60/ab[1][12] ) );
  AND U1505 ( .A(b[11]), .B(a[1]), .Z(\r60/ab[1][11] ) );
  AND U1506 ( .A(b[10]), .B(a[1]), .Z(\r60/ab[1][10] ) );
  AND U1507 ( .A(b[0]), .B(a[1]), .Z(\r60/ab[1][0] ) );
  AND U1508 ( .A(b[9]), .B(a[19]), .Z(\r60/ab[19][9] ) );
  AND U1509 ( .A(b[8]), .B(a[19]), .Z(\r60/ab[19][8] ) );
  AND U1510 ( .A(b[7]), .B(a[19]), .Z(\r60/ab[19][7] ) );
  AND U1511 ( .A(b[6]), .B(a[19]), .Z(\r60/ab[19][6] ) );
  AND U1512 ( .A(b[5]), .B(a[19]), .Z(\r60/ab[19][5] ) );
  AND U1513 ( .A(b[4]), .B(a[19]), .Z(\r60/ab[19][4] ) );
  AND U1514 ( .A(b[3]), .B(a[19]), .Z(\r60/ab[19][3] ) );
  MUX U1515 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[19]), .F(\r60/ab[19][31] ) );
  AND U1516 ( .A(b[30]), .B(a[19]), .Z(\r60/ab[19][30] ) );
  AND U1517 ( .A(b[2]), .B(a[19]), .Z(\r60/ab[19][2] ) );
  AND U1518 ( .A(b[29]), .B(a[19]), .Z(\r60/ab[19][29] ) );
  AND U1519 ( .A(b[28]), .B(a[19]), .Z(\r60/ab[19][28] ) );
  AND U1520 ( .A(b[27]), .B(a[19]), .Z(\r60/ab[19][27] ) );
  AND U1521 ( .A(b[26]), .B(a[19]), .Z(\r60/ab[19][26] ) );
  AND U1522 ( .A(b[25]), .B(a[19]), .Z(\r60/ab[19][25] ) );
  AND U1523 ( .A(b[24]), .B(a[19]), .Z(\r60/ab[19][24] ) );
  AND U1524 ( .A(b[23]), .B(a[19]), .Z(\r60/ab[19][23] ) );
  AND U1525 ( .A(b[22]), .B(a[19]), .Z(\r60/ab[19][22] ) );
  AND U1526 ( .A(b[21]), .B(a[19]), .Z(\r60/ab[19][21] ) );
  AND U1527 ( .A(b[20]), .B(a[19]), .Z(\r60/ab[19][20] ) );
  AND U1528 ( .A(b[1]), .B(a[19]), .Z(\r60/ab[19][1] ) );
  AND U1529 ( .A(b[19]), .B(a[19]), .Z(\r60/ab[19][19] ) );
  AND U1530 ( .A(b[18]), .B(a[19]), .Z(\r60/ab[19][18] ) );
  AND U1531 ( .A(b[17]), .B(a[19]), .Z(\r60/ab[19][17] ) );
  AND U1532 ( .A(b[16]), .B(a[19]), .Z(\r60/ab[19][16] ) );
  AND U1533 ( .A(b[15]), .B(a[19]), .Z(\r60/ab[19][15] ) );
  AND U1534 ( .A(b[14]), .B(a[19]), .Z(\r60/ab[19][14] ) );
  AND U1535 ( .A(b[13]), .B(a[19]), .Z(\r60/ab[19][13] ) );
  AND U1536 ( .A(b[12]), .B(a[19]), .Z(\r60/ab[19][12] ) );
  AND U1537 ( .A(b[11]), .B(a[19]), .Z(\r60/ab[19][11] ) );
  AND U1538 ( .A(b[10]), .B(a[19]), .Z(\r60/ab[19][10] ) );
  AND U1539 ( .A(b[0]), .B(a[19]), .Z(\r60/ab[19][0] ) );
  AND U1540 ( .A(b[9]), .B(a[18]), .Z(\r60/ab[18][9] ) );
  AND U1541 ( .A(b[8]), .B(a[18]), .Z(\r60/ab[18][8] ) );
  AND U1542 ( .A(b[7]), .B(a[18]), .Z(\r60/ab[18][7] ) );
  AND U1543 ( .A(b[6]), .B(a[18]), .Z(\r60/ab[18][6] ) );
  AND U1544 ( .A(b[5]), .B(a[18]), .Z(\r60/ab[18][5] ) );
  AND U1545 ( .A(b[4]), .B(a[18]), .Z(\r60/ab[18][4] ) );
  AND U1546 ( .A(b[3]), .B(a[18]), .Z(\r60/ab[18][3] ) );
  MUX U1547 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[18]), .F(\r60/ab[18][31] ) );
  AND U1548 ( .A(b[30]), .B(a[18]), .Z(\r60/ab[18][30] ) );
  AND U1549 ( .A(b[2]), .B(a[18]), .Z(\r60/ab[18][2] ) );
  AND U1550 ( .A(b[29]), .B(a[18]), .Z(\r60/ab[18][29] ) );
  AND U1551 ( .A(b[28]), .B(a[18]), .Z(\r60/ab[18][28] ) );
  AND U1552 ( .A(b[27]), .B(a[18]), .Z(\r60/ab[18][27] ) );
  AND U1553 ( .A(b[26]), .B(a[18]), .Z(\r60/ab[18][26] ) );
  AND U1554 ( .A(b[25]), .B(a[18]), .Z(\r60/ab[18][25] ) );
  AND U1555 ( .A(b[24]), .B(a[18]), .Z(\r60/ab[18][24] ) );
  AND U1556 ( .A(b[23]), .B(a[18]), .Z(\r60/ab[18][23] ) );
  AND U1557 ( .A(b[22]), .B(a[18]), .Z(\r60/ab[18][22] ) );
  AND U1558 ( .A(b[21]), .B(a[18]), .Z(\r60/ab[18][21] ) );
  AND U1559 ( .A(b[20]), .B(a[18]), .Z(\r60/ab[18][20] ) );
  AND U1560 ( .A(b[1]), .B(a[18]), .Z(\r60/ab[18][1] ) );
  AND U1561 ( .A(b[19]), .B(a[18]), .Z(\r60/ab[18][19] ) );
  AND U1562 ( .A(b[18]), .B(a[18]), .Z(\r60/ab[18][18] ) );
  AND U1563 ( .A(b[17]), .B(a[18]), .Z(\r60/ab[18][17] ) );
  AND U1564 ( .A(b[16]), .B(a[18]), .Z(\r60/ab[18][16] ) );
  AND U1565 ( .A(b[15]), .B(a[18]), .Z(\r60/ab[18][15] ) );
  AND U1566 ( .A(b[14]), .B(a[18]), .Z(\r60/ab[18][14] ) );
  AND U1567 ( .A(b[13]), .B(a[18]), .Z(\r60/ab[18][13] ) );
  AND U1568 ( .A(b[12]), .B(a[18]), .Z(\r60/ab[18][12] ) );
  AND U1569 ( .A(b[11]), .B(a[18]), .Z(\r60/ab[18][11] ) );
  AND U1570 ( .A(b[10]), .B(a[18]), .Z(\r60/ab[18][10] ) );
  AND U1571 ( .A(b[0]), .B(a[18]), .Z(\r60/ab[18][0] ) );
  AND U1572 ( .A(b[9]), .B(a[17]), .Z(\r60/ab[17][9] ) );
  AND U1573 ( .A(b[8]), .B(a[17]), .Z(\r60/ab[17][8] ) );
  AND U1574 ( .A(b[7]), .B(a[17]), .Z(\r60/ab[17][7] ) );
  AND U1575 ( .A(b[6]), .B(a[17]), .Z(\r60/ab[17][6] ) );
  AND U1576 ( .A(b[5]), .B(a[17]), .Z(\r60/ab[17][5] ) );
  AND U1577 ( .A(b[4]), .B(a[17]), .Z(\r60/ab[17][4] ) );
  AND U1578 ( .A(b[3]), .B(a[17]), .Z(\r60/ab[17][3] ) );
  MUX U1579 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[17]), .F(\r60/ab[17][31] ) );
  AND U1580 ( .A(b[30]), .B(a[17]), .Z(\r60/ab[17][30] ) );
  AND U1581 ( .A(b[2]), .B(a[17]), .Z(\r60/ab[17][2] ) );
  AND U1582 ( .A(b[29]), .B(a[17]), .Z(\r60/ab[17][29] ) );
  AND U1583 ( .A(b[28]), .B(a[17]), .Z(\r60/ab[17][28] ) );
  AND U1584 ( .A(b[27]), .B(a[17]), .Z(\r60/ab[17][27] ) );
  AND U1585 ( .A(b[26]), .B(a[17]), .Z(\r60/ab[17][26] ) );
  AND U1586 ( .A(b[25]), .B(a[17]), .Z(\r60/ab[17][25] ) );
  AND U1587 ( .A(b[24]), .B(a[17]), .Z(\r60/ab[17][24] ) );
  AND U1588 ( .A(b[23]), .B(a[17]), .Z(\r60/ab[17][23] ) );
  AND U1589 ( .A(b[22]), .B(a[17]), .Z(\r60/ab[17][22] ) );
  AND U1590 ( .A(b[21]), .B(a[17]), .Z(\r60/ab[17][21] ) );
  AND U1591 ( .A(b[20]), .B(a[17]), .Z(\r60/ab[17][20] ) );
  AND U1592 ( .A(b[1]), .B(a[17]), .Z(\r60/ab[17][1] ) );
  AND U1593 ( .A(b[19]), .B(a[17]), .Z(\r60/ab[17][19] ) );
  AND U1594 ( .A(b[18]), .B(a[17]), .Z(\r60/ab[17][18] ) );
  AND U1595 ( .A(b[17]), .B(a[17]), .Z(\r60/ab[17][17] ) );
  AND U1596 ( .A(b[16]), .B(a[17]), .Z(\r60/ab[17][16] ) );
  AND U1597 ( .A(b[15]), .B(a[17]), .Z(\r60/ab[17][15] ) );
  AND U1598 ( .A(b[14]), .B(a[17]), .Z(\r60/ab[17][14] ) );
  AND U1599 ( .A(b[13]), .B(a[17]), .Z(\r60/ab[17][13] ) );
  AND U1600 ( .A(b[12]), .B(a[17]), .Z(\r60/ab[17][12] ) );
  AND U1601 ( .A(b[11]), .B(a[17]), .Z(\r60/ab[17][11] ) );
  AND U1602 ( .A(b[10]), .B(a[17]), .Z(\r60/ab[17][10] ) );
  AND U1603 ( .A(b[0]), .B(a[17]), .Z(\r60/ab[17][0] ) );
  AND U1604 ( .A(b[9]), .B(a[16]), .Z(\r60/ab[16][9] ) );
  AND U1605 ( .A(b[8]), .B(a[16]), .Z(\r60/ab[16][8] ) );
  AND U1606 ( .A(b[7]), .B(a[16]), .Z(\r60/ab[16][7] ) );
  AND U1607 ( .A(b[6]), .B(a[16]), .Z(\r60/ab[16][6] ) );
  AND U1608 ( .A(b[5]), .B(a[16]), .Z(\r60/ab[16][5] ) );
  AND U1609 ( .A(b[4]), .B(a[16]), .Z(\r60/ab[16][4] ) );
  AND U1610 ( .A(b[3]), .B(a[16]), .Z(\r60/ab[16][3] ) );
  MUX U1611 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[16]), .F(\r60/ab[16][31] ) );
  AND U1612 ( .A(b[30]), .B(a[16]), .Z(\r60/ab[16][30] ) );
  AND U1613 ( .A(b[2]), .B(a[16]), .Z(\r60/ab[16][2] ) );
  AND U1614 ( .A(b[29]), .B(a[16]), .Z(\r60/ab[16][29] ) );
  AND U1615 ( .A(b[28]), .B(a[16]), .Z(\r60/ab[16][28] ) );
  AND U1616 ( .A(b[27]), .B(a[16]), .Z(\r60/ab[16][27] ) );
  AND U1617 ( .A(b[26]), .B(a[16]), .Z(\r60/ab[16][26] ) );
  AND U1618 ( .A(b[25]), .B(a[16]), .Z(\r60/ab[16][25] ) );
  AND U1619 ( .A(b[24]), .B(a[16]), .Z(\r60/ab[16][24] ) );
  AND U1620 ( .A(b[23]), .B(a[16]), .Z(\r60/ab[16][23] ) );
  AND U1621 ( .A(b[22]), .B(a[16]), .Z(\r60/ab[16][22] ) );
  AND U1622 ( .A(b[21]), .B(a[16]), .Z(\r60/ab[16][21] ) );
  AND U1623 ( .A(b[20]), .B(a[16]), .Z(\r60/ab[16][20] ) );
  AND U1624 ( .A(b[1]), .B(a[16]), .Z(\r60/ab[16][1] ) );
  AND U1625 ( .A(b[19]), .B(a[16]), .Z(\r60/ab[16][19] ) );
  AND U1626 ( .A(b[18]), .B(a[16]), .Z(\r60/ab[16][18] ) );
  AND U1627 ( .A(b[17]), .B(a[16]), .Z(\r60/ab[16][17] ) );
  AND U1628 ( .A(b[16]), .B(a[16]), .Z(\r60/ab[16][16] ) );
  AND U1629 ( .A(b[15]), .B(a[16]), .Z(\r60/ab[16][15] ) );
  AND U1630 ( .A(b[14]), .B(a[16]), .Z(\r60/ab[16][14] ) );
  AND U1631 ( .A(b[13]), .B(a[16]), .Z(\r60/ab[16][13] ) );
  AND U1632 ( .A(b[12]), .B(a[16]), .Z(\r60/ab[16][12] ) );
  AND U1633 ( .A(b[11]), .B(a[16]), .Z(\r60/ab[16][11] ) );
  AND U1634 ( .A(b[10]), .B(a[16]), .Z(\r60/ab[16][10] ) );
  AND U1635 ( .A(b[0]), .B(a[16]), .Z(\r60/ab[16][0] ) );
  AND U1636 ( .A(b[9]), .B(a[15]), .Z(\r60/ab[15][9] ) );
  AND U1637 ( .A(b[8]), .B(a[15]), .Z(\r60/ab[15][8] ) );
  AND U1638 ( .A(b[7]), .B(a[15]), .Z(\r60/ab[15][7] ) );
  AND U1639 ( .A(b[6]), .B(a[15]), .Z(\r60/ab[15][6] ) );
  AND U1640 ( .A(b[5]), .B(a[15]), .Z(\r60/ab[15][5] ) );
  AND U1641 ( .A(b[4]), .B(a[15]), .Z(\r60/ab[15][4] ) );
  AND U1642 ( .A(b[3]), .B(a[15]), .Z(\r60/ab[15][3] ) );
  MUX U1643 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[15]), .F(\r60/ab[15][31] ) );
  AND U1644 ( .A(b[30]), .B(a[15]), .Z(\r60/ab[15][30] ) );
  AND U1645 ( .A(b[2]), .B(a[15]), .Z(\r60/ab[15][2] ) );
  AND U1646 ( .A(b[29]), .B(a[15]), .Z(\r60/ab[15][29] ) );
  AND U1647 ( .A(b[28]), .B(a[15]), .Z(\r60/ab[15][28] ) );
  AND U1648 ( .A(b[27]), .B(a[15]), .Z(\r60/ab[15][27] ) );
  AND U1649 ( .A(b[26]), .B(a[15]), .Z(\r60/ab[15][26] ) );
  AND U1650 ( .A(b[25]), .B(a[15]), .Z(\r60/ab[15][25] ) );
  AND U1651 ( .A(b[24]), .B(a[15]), .Z(\r60/ab[15][24] ) );
  AND U1652 ( .A(b[23]), .B(a[15]), .Z(\r60/ab[15][23] ) );
  AND U1653 ( .A(b[22]), .B(a[15]), .Z(\r60/ab[15][22] ) );
  AND U1654 ( .A(b[21]), .B(a[15]), .Z(\r60/ab[15][21] ) );
  AND U1655 ( .A(b[20]), .B(a[15]), .Z(\r60/ab[15][20] ) );
  AND U1656 ( .A(b[1]), .B(a[15]), .Z(\r60/ab[15][1] ) );
  AND U1657 ( .A(b[19]), .B(a[15]), .Z(\r60/ab[15][19] ) );
  AND U1658 ( .A(b[18]), .B(a[15]), .Z(\r60/ab[15][18] ) );
  AND U1659 ( .A(b[17]), .B(a[15]), .Z(\r60/ab[15][17] ) );
  AND U1660 ( .A(b[16]), .B(a[15]), .Z(\r60/ab[15][16] ) );
  AND U1661 ( .A(b[15]), .B(a[15]), .Z(\r60/ab[15][15] ) );
  AND U1662 ( .A(b[14]), .B(a[15]), .Z(\r60/ab[15][14] ) );
  AND U1663 ( .A(b[13]), .B(a[15]), .Z(\r60/ab[15][13] ) );
  AND U1664 ( .A(b[12]), .B(a[15]), .Z(\r60/ab[15][12] ) );
  AND U1665 ( .A(b[11]), .B(a[15]), .Z(\r60/ab[15][11] ) );
  AND U1666 ( .A(b[10]), .B(a[15]), .Z(\r60/ab[15][10] ) );
  AND U1667 ( .A(b[0]), .B(a[15]), .Z(\r60/ab[15][0] ) );
  AND U1668 ( .A(b[9]), .B(a[14]), .Z(\r60/ab[14][9] ) );
  AND U1669 ( .A(b[8]), .B(a[14]), .Z(\r60/ab[14][8] ) );
  AND U1670 ( .A(b[7]), .B(a[14]), .Z(\r60/ab[14][7] ) );
  AND U1671 ( .A(b[6]), .B(a[14]), .Z(\r60/ab[14][6] ) );
  AND U1672 ( .A(b[5]), .B(a[14]), .Z(\r60/ab[14][5] ) );
  AND U1673 ( .A(b[4]), .B(a[14]), .Z(\r60/ab[14][4] ) );
  AND U1674 ( .A(b[3]), .B(a[14]), .Z(\r60/ab[14][3] ) );
  MUX U1675 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[14]), .F(\r60/ab[14][31] ) );
  AND U1676 ( .A(b[30]), .B(a[14]), .Z(\r60/ab[14][30] ) );
  AND U1677 ( .A(b[2]), .B(a[14]), .Z(\r60/ab[14][2] ) );
  AND U1678 ( .A(b[29]), .B(a[14]), .Z(\r60/ab[14][29] ) );
  AND U1679 ( .A(b[28]), .B(a[14]), .Z(\r60/ab[14][28] ) );
  AND U1680 ( .A(b[27]), .B(a[14]), .Z(\r60/ab[14][27] ) );
  AND U1681 ( .A(b[26]), .B(a[14]), .Z(\r60/ab[14][26] ) );
  AND U1682 ( .A(b[25]), .B(a[14]), .Z(\r60/ab[14][25] ) );
  AND U1683 ( .A(b[24]), .B(a[14]), .Z(\r60/ab[14][24] ) );
  AND U1684 ( .A(b[23]), .B(a[14]), .Z(\r60/ab[14][23] ) );
  AND U1685 ( .A(b[22]), .B(a[14]), .Z(\r60/ab[14][22] ) );
  AND U1686 ( .A(b[21]), .B(a[14]), .Z(\r60/ab[14][21] ) );
  AND U1687 ( .A(b[20]), .B(a[14]), .Z(\r60/ab[14][20] ) );
  AND U1688 ( .A(b[1]), .B(a[14]), .Z(\r60/ab[14][1] ) );
  AND U1689 ( .A(b[19]), .B(a[14]), .Z(\r60/ab[14][19] ) );
  AND U1690 ( .A(b[18]), .B(a[14]), .Z(\r60/ab[14][18] ) );
  AND U1691 ( .A(b[17]), .B(a[14]), .Z(\r60/ab[14][17] ) );
  AND U1692 ( .A(b[16]), .B(a[14]), .Z(\r60/ab[14][16] ) );
  AND U1693 ( .A(b[15]), .B(a[14]), .Z(\r60/ab[14][15] ) );
  AND U1694 ( .A(b[14]), .B(a[14]), .Z(\r60/ab[14][14] ) );
  AND U1695 ( .A(b[13]), .B(a[14]), .Z(\r60/ab[14][13] ) );
  AND U1696 ( .A(b[12]), .B(a[14]), .Z(\r60/ab[14][12] ) );
  AND U1697 ( .A(b[11]), .B(a[14]), .Z(\r60/ab[14][11] ) );
  AND U1698 ( .A(b[10]), .B(a[14]), .Z(\r60/ab[14][10] ) );
  AND U1699 ( .A(b[0]), .B(a[14]), .Z(\r60/ab[14][0] ) );
  AND U1700 ( .A(b[9]), .B(a[13]), .Z(\r60/ab[13][9] ) );
  AND U1701 ( .A(b[8]), .B(a[13]), .Z(\r60/ab[13][8] ) );
  AND U1702 ( .A(b[7]), .B(a[13]), .Z(\r60/ab[13][7] ) );
  AND U1703 ( .A(b[6]), .B(a[13]), .Z(\r60/ab[13][6] ) );
  AND U1704 ( .A(b[5]), .B(a[13]), .Z(\r60/ab[13][5] ) );
  AND U1705 ( .A(b[4]), .B(a[13]), .Z(\r60/ab[13][4] ) );
  AND U1706 ( .A(b[3]), .B(a[13]), .Z(\r60/ab[13][3] ) );
  MUX U1707 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[13]), .F(\r60/ab[13][31] ) );
  AND U1708 ( .A(b[30]), .B(a[13]), .Z(\r60/ab[13][30] ) );
  AND U1709 ( .A(b[2]), .B(a[13]), .Z(\r60/ab[13][2] ) );
  AND U1710 ( .A(b[29]), .B(a[13]), .Z(\r60/ab[13][29] ) );
  AND U1711 ( .A(b[28]), .B(a[13]), .Z(\r60/ab[13][28] ) );
  AND U1712 ( .A(b[27]), .B(a[13]), .Z(\r60/ab[13][27] ) );
  AND U1713 ( .A(b[26]), .B(a[13]), .Z(\r60/ab[13][26] ) );
  AND U1714 ( .A(b[25]), .B(a[13]), .Z(\r60/ab[13][25] ) );
  AND U1715 ( .A(b[24]), .B(a[13]), .Z(\r60/ab[13][24] ) );
  AND U1716 ( .A(b[23]), .B(a[13]), .Z(\r60/ab[13][23] ) );
  AND U1717 ( .A(b[22]), .B(a[13]), .Z(\r60/ab[13][22] ) );
  AND U1718 ( .A(b[21]), .B(a[13]), .Z(\r60/ab[13][21] ) );
  AND U1719 ( .A(b[20]), .B(a[13]), .Z(\r60/ab[13][20] ) );
  AND U1720 ( .A(b[1]), .B(a[13]), .Z(\r60/ab[13][1] ) );
  AND U1721 ( .A(b[19]), .B(a[13]), .Z(\r60/ab[13][19] ) );
  AND U1722 ( .A(b[18]), .B(a[13]), .Z(\r60/ab[13][18] ) );
  AND U1723 ( .A(b[17]), .B(a[13]), .Z(\r60/ab[13][17] ) );
  AND U1724 ( .A(b[16]), .B(a[13]), .Z(\r60/ab[13][16] ) );
  AND U1725 ( .A(b[15]), .B(a[13]), .Z(\r60/ab[13][15] ) );
  AND U1726 ( .A(b[14]), .B(a[13]), .Z(\r60/ab[13][14] ) );
  AND U1727 ( .A(b[13]), .B(a[13]), .Z(\r60/ab[13][13] ) );
  AND U1728 ( .A(b[12]), .B(a[13]), .Z(\r60/ab[13][12] ) );
  AND U1729 ( .A(b[11]), .B(a[13]), .Z(\r60/ab[13][11] ) );
  AND U1730 ( .A(b[10]), .B(a[13]), .Z(\r60/ab[13][10] ) );
  AND U1731 ( .A(b[0]), .B(a[13]), .Z(\r60/ab[13][0] ) );
  AND U1732 ( .A(b[9]), .B(a[12]), .Z(\r60/ab[12][9] ) );
  AND U1733 ( .A(b[8]), .B(a[12]), .Z(\r60/ab[12][8] ) );
  AND U1734 ( .A(b[7]), .B(a[12]), .Z(\r60/ab[12][7] ) );
  AND U1735 ( .A(b[6]), .B(a[12]), .Z(\r60/ab[12][6] ) );
  AND U1736 ( .A(b[5]), .B(a[12]), .Z(\r60/ab[12][5] ) );
  AND U1737 ( .A(b[4]), .B(a[12]), .Z(\r60/ab[12][4] ) );
  AND U1738 ( .A(b[3]), .B(a[12]), .Z(\r60/ab[12][3] ) );
  MUX U1739 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[12]), .F(\r60/ab[12][31] ) );
  AND U1740 ( .A(b[30]), .B(a[12]), .Z(\r60/ab[12][30] ) );
  AND U1741 ( .A(b[2]), .B(a[12]), .Z(\r60/ab[12][2] ) );
  AND U1742 ( .A(b[29]), .B(a[12]), .Z(\r60/ab[12][29] ) );
  AND U1743 ( .A(b[28]), .B(a[12]), .Z(\r60/ab[12][28] ) );
  AND U1744 ( .A(b[27]), .B(a[12]), .Z(\r60/ab[12][27] ) );
  AND U1745 ( .A(b[26]), .B(a[12]), .Z(\r60/ab[12][26] ) );
  AND U1746 ( .A(b[25]), .B(a[12]), .Z(\r60/ab[12][25] ) );
  AND U1747 ( .A(b[24]), .B(a[12]), .Z(\r60/ab[12][24] ) );
  AND U1748 ( .A(b[23]), .B(a[12]), .Z(\r60/ab[12][23] ) );
  AND U1749 ( .A(b[22]), .B(a[12]), .Z(\r60/ab[12][22] ) );
  AND U1750 ( .A(b[21]), .B(a[12]), .Z(\r60/ab[12][21] ) );
  AND U1751 ( .A(b[20]), .B(a[12]), .Z(\r60/ab[12][20] ) );
  AND U1752 ( .A(b[1]), .B(a[12]), .Z(\r60/ab[12][1] ) );
  AND U1753 ( .A(b[19]), .B(a[12]), .Z(\r60/ab[12][19] ) );
  AND U1754 ( .A(b[18]), .B(a[12]), .Z(\r60/ab[12][18] ) );
  AND U1755 ( .A(b[17]), .B(a[12]), .Z(\r60/ab[12][17] ) );
  AND U1756 ( .A(b[16]), .B(a[12]), .Z(\r60/ab[12][16] ) );
  AND U1757 ( .A(b[15]), .B(a[12]), .Z(\r60/ab[12][15] ) );
  AND U1758 ( .A(b[14]), .B(a[12]), .Z(\r60/ab[12][14] ) );
  AND U1759 ( .A(b[13]), .B(a[12]), .Z(\r60/ab[12][13] ) );
  AND U1760 ( .A(b[12]), .B(a[12]), .Z(\r60/ab[12][12] ) );
  AND U1761 ( .A(b[11]), .B(a[12]), .Z(\r60/ab[12][11] ) );
  AND U1762 ( .A(b[10]), .B(a[12]), .Z(\r60/ab[12][10] ) );
  AND U1763 ( .A(b[0]), .B(a[12]), .Z(\r60/ab[12][0] ) );
  AND U1764 ( .A(b[9]), .B(a[11]), .Z(\r60/ab[11][9] ) );
  AND U1765 ( .A(b[8]), .B(a[11]), .Z(\r60/ab[11][8] ) );
  AND U1766 ( .A(b[7]), .B(a[11]), .Z(\r60/ab[11][7] ) );
  AND U1767 ( .A(b[6]), .B(a[11]), .Z(\r60/ab[11][6] ) );
  AND U1768 ( .A(b[5]), .B(a[11]), .Z(\r60/ab[11][5] ) );
  AND U1769 ( .A(b[4]), .B(a[11]), .Z(\r60/ab[11][4] ) );
  AND U1770 ( .A(b[3]), .B(a[11]), .Z(\r60/ab[11][3] ) );
  MUX U1771 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[11]), .F(\r60/ab[11][31] ) );
  AND U1772 ( .A(b[30]), .B(a[11]), .Z(\r60/ab[11][30] ) );
  AND U1773 ( .A(b[2]), .B(a[11]), .Z(\r60/ab[11][2] ) );
  AND U1774 ( .A(b[29]), .B(a[11]), .Z(\r60/ab[11][29] ) );
  AND U1775 ( .A(b[28]), .B(a[11]), .Z(\r60/ab[11][28] ) );
  AND U1776 ( .A(b[27]), .B(a[11]), .Z(\r60/ab[11][27] ) );
  AND U1777 ( .A(b[26]), .B(a[11]), .Z(\r60/ab[11][26] ) );
  AND U1778 ( .A(b[25]), .B(a[11]), .Z(\r60/ab[11][25] ) );
  AND U1779 ( .A(b[24]), .B(a[11]), .Z(\r60/ab[11][24] ) );
  AND U1780 ( .A(b[23]), .B(a[11]), .Z(\r60/ab[11][23] ) );
  AND U1781 ( .A(b[22]), .B(a[11]), .Z(\r60/ab[11][22] ) );
  AND U1782 ( .A(b[21]), .B(a[11]), .Z(\r60/ab[11][21] ) );
  AND U1783 ( .A(b[20]), .B(a[11]), .Z(\r60/ab[11][20] ) );
  AND U1784 ( .A(b[1]), .B(a[11]), .Z(\r60/ab[11][1] ) );
  AND U1785 ( .A(b[19]), .B(a[11]), .Z(\r60/ab[11][19] ) );
  AND U1786 ( .A(b[18]), .B(a[11]), .Z(\r60/ab[11][18] ) );
  AND U1787 ( .A(b[17]), .B(a[11]), .Z(\r60/ab[11][17] ) );
  AND U1788 ( .A(b[16]), .B(a[11]), .Z(\r60/ab[11][16] ) );
  AND U1789 ( .A(b[15]), .B(a[11]), .Z(\r60/ab[11][15] ) );
  AND U1790 ( .A(b[14]), .B(a[11]), .Z(\r60/ab[11][14] ) );
  AND U1791 ( .A(b[13]), .B(a[11]), .Z(\r60/ab[11][13] ) );
  AND U1792 ( .A(b[12]), .B(a[11]), .Z(\r60/ab[11][12] ) );
  AND U1793 ( .A(b[11]), .B(a[11]), .Z(\r60/ab[11][11] ) );
  AND U1794 ( .A(b[10]), .B(a[11]), .Z(\r60/ab[11][10] ) );
  AND U1795 ( .A(b[0]), .B(a[11]), .Z(\r60/ab[11][0] ) );
  AND U1796 ( .A(b[9]), .B(a[10]), .Z(\r60/ab[10][9] ) );
  AND U1797 ( .A(b[8]), .B(a[10]), .Z(\r60/ab[10][8] ) );
  AND U1798 ( .A(b[7]), .B(a[10]), .Z(\r60/ab[10][7] ) );
  AND U1799 ( .A(b[6]), .B(a[10]), .Z(\r60/ab[10][6] ) );
  AND U1800 ( .A(b[5]), .B(a[10]), .Z(\r60/ab[10][5] ) );
  AND U1801 ( .A(b[4]), .B(a[10]), .Z(\r60/ab[10][4] ) );
  AND U1802 ( .A(b[3]), .B(a[10]), .Z(\r60/ab[10][3] ) );
  MUX U1803 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[10]), .F(\r60/ab[10][31] ) );
  AND U1804 ( .A(b[30]), .B(a[10]), .Z(\r60/ab[10][30] ) );
  AND U1805 ( .A(b[2]), .B(a[10]), .Z(\r60/ab[10][2] ) );
  AND U1806 ( .A(b[29]), .B(a[10]), .Z(\r60/ab[10][29] ) );
  AND U1807 ( .A(b[28]), .B(a[10]), .Z(\r60/ab[10][28] ) );
  AND U1808 ( .A(b[27]), .B(a[10]), .Z(\r60/ab[10][27] ) );
  AND U1809 ( .A(b[26]), .B(a[10]), .Z(\r60/ab[10][26] ) );
  AND U1810 ( .A(b[25]), .B(a[10]), .Z(\r60/ab[10][25] ) );
  AND U1811 ( .A(b[24]), .B(a[10]), .Z(\r60/ab[10][24] ) );
  AND U1812 ( .A(b[23]), .B(a[10]), .Z(\r60/ab[10][23] ) );
  AND U1813 ( .A(b[22]), .B(a[10]), .Z(\r60/ab[10][22] ) );
  AND U1814 ( .A(b[21]), .B(a[10]), .Z(\r60/ab[10][21] ) );
  AND U1815 ( .A(b[20]), .B(a[10]), .Z(\r60/ab[10][20] ) );
  AND U1816 ( .A(b[1]), .B(a[10]), .Z(\r60/ab[10][1] ) );
  AND U1817 ( .A(b[19]), .B(a[10]), .Z(\r60/ab[10][19] ) );
  AND U1818 ( .A(b[18]), .B(a[10]), .Z(\r60/ab[10][18] ) );
  AND U1819 ( .A(b[17]), .B(a[10]), .Z(\r60/ab[10][17] ) );
  AND U1820 ( .A(b[16]), .B(a[10]), .Z(\r60/ab[10][16] ) );
  AND U1821 ( .A(b[15]), .B(a[10]), .Z(\r60/ab[10][15] ) );
  AND U1822 ( .A(b[14]), .B(a[10]), .Z(\r60/ab[10][14] ) );
  AND U1823 ( .A(b[13]), .B(a[10]), .Z(\r60/ab[10][13] ) );
  AND U1824 ( .A(b[12]), .B(a[10]), .Z(\r60/ab[10][12] ) );
  AND U1825 ( .A(b[11]), .B(a[10]), .Z(\r60/ab[10][11] ) );
  AND U1826 ( .A(b[10]), .B(a[10]), .Z(\r60/ab[10][10] ) );
  AND U1827 ( .A(b[0]), .B(a[10]), .Z(\r60/ab[10][0] ) );
  ANDN U1828 ( .B(b[9]), .A(n683), .Z(\r60/ab[0][9] ) );
  ANDN U1829 ( .B(b[8]), .A(n683), .Z(\r60/ab[0][8] ) );
  ANDN U1830 ( .B(b[7]), .A(n683), .Z(\r60/ab[0][7] ) );
  ANDN U1831 ( .B(b[6]), .A(n683), .Z(\r60/ab[0][6] ) );
  ANDN U1832 ( .B(b[5]), .A(n683), .Z(\r60/ab[0][5] ) );
  ANDN U1833 ( .B(b[4]), .A(n683), .Z(\r60/ab[0][4] ) );
  ANDN U1834 ( .B(b[3]), .A(n683), .Z(\r60/ab[0][3] ) );
  MUX U1835 ( .IN0(\r60/ZB ), .IN1(n680), .SEL(a[0]), .F(\r60/ab[0][31] ) );
  ANDN U1836 ( .B(b[31]), .A(\U3/U1/Z_0 ), .Z(n680) );
  ANDN U1837 ( .B(b[30]), .A(n683), .Z(\r60/ab[0][30] ) );
  ANDN U1838 ( .B(b[2]), .A(n683), .Z(\r60/ab[0][2] ) );
  ANDN U1839 ( .B(b[29]), .A(n683), .Z(\r60/ab[0][29] ) );
  ANDN U1840 ( .B(b[28]), .A(n683), .Z(\r60/ab[0][28] ) );
  ANDN U1841 ( .B(b[27]), .A(n683), .Z(\r60/ab[0][27] ) );
  ANDN U1842 ( .B(b[26]), .A(n683), .Z(\r60/ab[0][26] ) );
  ANDN U1843 ( .B(b[25]), .A(n683), .Z(\r60/ab[0][25] ) );
  ANDN U1844 ( .B(b[24]), .A(n683), .Z(\r60/ab[0][24] ) );
  ANDN U1845 ( .B(b[23]), .A(n683), .Z(\r60/ab[0][23] ) );
  ANDN U1846 ( .B(b[22]), .A(n683), .Z(\r60/ab[0][22] ) );
  ANDN U1847 ( .B(b[21]), .A(n683), .Z(\r60/ab[0][21] ) );
  ANDN U1848 ( .B(b[20]), .A(n683), .Z(\r60/ab[0][20] ) );
  ANDN U1849 ( .B(b[1]), .A(n683), .Z(\r60/ab[0][1] ) );
  ANDN U1850 ( .B(b[19]), .A(n683), .Z(\r60/ab[0][19] ) );
  ANDN U1851 ( .B(b[18]), .A(n683), .Z(\r60/ab[0][18] ) );
  ANDN U1852 ( .B(b[17]), .A(n683), .Z(\r60/ab[0][17] ) );
  ANDN U1853 ( .B(b[16]), .A(n683), .Z(\r60/ab[0][16] ) );
  ANDN U1854 ( .B(b[15]), .A(n683), .Z(\r60/ab[0][15] ) );
  ANDN U1855 ( .B(b[14]), .A(n683), .Z(\r60/ab[0][14] ) );
  ANDN U1856 ( .B(b[13]), .A(n683), .Z(\r60/ab[0][13] ) );
  ANDN U1857 ( .B(b[12]), .A(n683), .Z(\r60/ab[0][12] ) );
  ANDN U1858 ( .B(b[11]), .A(n683), .Z(\r60/ab[0][11] ) );
  ANDN U1859 ( .B(b[10]), .A(n683), .Z(\r60/ab[0][10] ) );
  AND U1860 ( .A(\U3/U1/Z_0 ), .B(b[31]), .Z(\r60/ZB ) );
  ANDN U1861 ( .B(\U3/U1/Z_0 ), .A(n682), .Z(\r60/ZA ) );
  ANDN U1862 ( .B(\U3/U1/Z_0 ), .A(b[31]), .Z(\r60/QB ) );
  ANDN U1863 ( .B(\U3/U1/Z_0 ), .A(a[31]), .Z(\r60/QA ) );
  MUX U1864 ( .IN0(n684), .IN1(Hi[31]), .SEL(n685), .F(n679) );
  NANDN U1865 ( .A(n686), .B(n687), .Z(n684) );
  AND U1866 ( .A(n688), .B(n689), .Z(n687) );
  NANDN U1867 ( .A(n690), .B(n691), .Z(n689) );
  NANDN U1868 ( .A(n690), .B(\U3/U1/Z_0 ), .Z(n688) );
  XNOR U1869 ( .A(n692), .B(n693), .Z(n690) );
  ANDN U1870 ( .B(n694), .A(n695), .Z(n693) );
  NANDN U1871 ( .A(n696), .B(n697), .Z(n694) );
  XNOR U1872 ( .A(\r60/A2[61] ), .B(\r60/A1[61] ), .Z(n692) );
  MUX U1873 ( .IN0(n698), .IN1(Hi[30]), .SEL(n685), .F(n678) );
  NANDN U1874 ( .A(n699), .B(n700), .Z(n698) );
  AND U1875 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U1876 ( .A(n703), .B(n691), .Z(n702) );
  NANDN U1877 ( .A(n703), .B(\U3/U1/Z_0 ), .Z(n701) );
  XOR U1878 ( .A(n704), .B(n697), .Z(n703) );
  NANDN U1879 ( .A(n705), .B(n706), .Z(n697) );
  NANDN U1880 ( .A(n707), .B(n708), .Z(n706) );
  OR U1881 ( .A(n696), .B(n695), .Z(n704) );
  AND U1882 ( .A(\r60/A1[60] ), .B(\r60/A2[60] ), .Z(n695) );
  NOR U1883 ( .A(\r60/A2[60] ), .B(\r60/A1[60] ), .Z(n696) );
  MUX U1884 ( .IN0(n709), .IN1(Hi[29]), .SEL(n685), .F(n677) );
  NANDN U1885 ( .A(n710), .B(n711), .Z(n709) );
  AND U1886 ( .A(n712), .B(n713), .Z(n711) );
  NANDN U1887 ( .A(n714), .B(n691), .Z(n713) );
  NANDN U1888 ( .A(n714), .B(\U3/U1/Z_0 ), .Z(n712) );
  XOR U1889 ( .A(n715), .B(n708), .Z(n714) );
  NANDN U1890 ( .A(n716), .B(n717), .Z(n708) );
  NANDN U1891 ( .A(n718), .B(n719), .Z(n717) );
  OR U1892 ( .A(n707), .B(n705), .Z(n715) );
  AND U1893 ( .A(\r60/A1[59] ), .B(\r60/A2[59] ), .Z(n705) );
  NOR U1894 ( .A(\r60/A2[59] ), .B(\r60/A1[59] ), .Z(n707) );
  MUX U1895 ( .IN0(n720), .IN1(Hi[28]), .SEL(n685), .F(n676) );
  NANDN U1896 ( .A(n721), .B(n722), .Z(n720) );
  AND U1897 ( .A(n723), .B(n724), .Z(n722) );
  NANDN U1898 ( .A(n725), .B(n691), .Z(n724) );
  NANDN U1899 ( .A(n725), .B(\U3/U1/Z_0 ), .Z(n723) );
  XOR U1900 ( .A(n726), .B(n719), .Z(n725) );
  NANDN U1901 ( .A(n727), .B(n728), .Z(n719) );
  NANDN U1902 ( .A(n729), .B(n730), .Z(n728) );
  OR U1903 ( .A(n718), .B(n716), .Z(n726) );
  AND U1904 ( .A(\r60/A1[58] ), .B(\r60/A2[58] ), .Z(n716) );
  NOR U1905 ( .A(\r60/A2[58] ), .B(\r60/A1[58] ), .Z(n718) );
  MUX U1906 ( .IN0(n731), .IN1(Hi[27]), .SEL(n685), .F(n675) );
  NANDN U1907 ( .A(n732), .B(n733), .Z(n731) );
  AND U1908 ( .A(n734), .B(n735), .Z(n733) );
  NANDN U1909 ( .A(n736), .B(n691), .Z(n735) );
  NANDN U1910 ( .A(n736), .B(\U3/U1/Z_0 ), .Z(n734) );
  XOR U1911 ( .A(n737), .B(n730), .Z(n736) );
  NANDN U1912 ( .A(n738), .B(n739), .Z(n730) );
  NANDN U1913 ( .A(n740), .B(n741), .Z(n739) );
  OR U1914 ( .A(n729), .B(n727), .Z(n737) );
  AND U1915 ( .A(\r60/A1[57] ), .B(\r60/A2[57] ), .Z(n727) );
  NOR U1916 ( .A(\r60/A2[57] ), .B(\r60/A1[57] ), .Z(n729) );
  MUX U1917 ( .IN0(n742), .IN1(Hi[26]), .SEL(n685), .F(n674) );
  NANDN U1918 ( .A(n743), .B(n744), .Z(n742) );
  AND U1919 ( .A(n745), .B(n746), .Z(n744) );
  NANDN U1920 ( .A(n747), .B(n691), .Z(n746) );
  NANDN U1921 ( .A(n747), .B(\U3/U1/Z_0 ), .Z(n745) );
  XOR U1922 ( .A(n748), .B(n741), .Z(n747) );
  NANDN U1923 ( .A(n749), .B(n750), .Z(n741) );
  NANDN U1924 ( .A(n751), .B(n752), .Z(n750) );
  OR U1925 ( .A(n740), .B(n738), .Z(n748) );
  AND U1926 ( .A(\r60/A1[56] ), .B(\r60/A2[56] ), .Z(n738) );
  NOR U1927 ( .A(\r60/A2[56] ), .B(\r60/A1[56] ), .Z(n740) );
  MUX U1928 ( .IN0(n753), .IN1(Hi[25]), .SEL(n685), .F(n673) );
  NANDN U1929 ( .A(n754), .B(n755), .Z(n753) );
  AND U1930 ( .A(n756), .B(n757), .Z(n755) );
  NANDN U1931 ( .A(n758), .B(n691), .Z(n757) );
  NANDN U1932 ( .A(n758), .B(\U3/U1/Z_0 ), .Z(n756) );
  XOR U1933 ( .A(n759), .B(n752), .Z(n758) );
  NANDN U1934 ( .A(n760), .B(n761), .Z(n752) );
  NANDN U1935 ( .A(n762), .B(n763), .Z(n761) );
  OR U1936 ( .A(n751), .B(n749), .Z(n759) );
  AND U1937 ( .A(\r60/A1[55] ), .B(\r60/A2[55] ), .Z(n749) );
  NOR U1938 ( .A(\r60/A2[55] ), .B(\r60/A1[55] ), .Z(n751) );
  MUX U1939 ( .IN0(n764), .IN1(Hi[24]), .SEL(n685), .F(n672) );
  NANDN U1940 ( .A(n765), .B(n766), .Z(n764) );
  AND U1941 ( .A(n767), .B(n768), .Z(n766) );
  NANDN U1942 ( .A(n769), .B(n691), .Z(n768) );
  NANDN U1943 ( .A(n769), .B(\U3/U1/Z_0 ), .Z(n767) );
  XOR U1944 ( .A(n770), .B(n763), .Z(n769) );
  NANDN U1945 ( .A(n771), .B(n772), .Z(n763) );
  NANDN U1946 ( .A(n773), .B(n774), .Z(n772) );
  OR U1947 ( .A(n762), .B(n760), .Z(n770) );
  AND U1948 ( .A(\r60/A1[54] ), .B(\r60/A2[54] ), .Z(n760) );
  NOR U1949 ( .A(\r60/A2[54] ), .B(\r60/A1[54] ), .Z(n762) );
  MUX U1950 ( .IN0(n775), .IN1(Hi[23]), .SEL(n685), .F(n671) );
  NANDN U1951 ( .A(n776), .B(n777), .Z(n775) );
  AND U1952 ( .A(n778), .B(n779), .Z(n777) );
  NANDN U1953 ( .A(n780), .B(n691), .Z(n779) );
  NANDN U1954 ( .A(n780), .B(\U3/U1/Z_0 ), .Z(n778) );
  XOR U1955 ( .A(n781), .B(n774), .Z(n780) );
  NANDN U1956 ( .A(n782), .B(n783), .Z(n774) );
  NANDN U1957 ( .A(n784), .B(n785), .Z(n783) );
  OR U1958 ( .A(n773), .B(n771), .Z(n781) );
  AND U1959 ( .A(\r60/A1[53] ), .B(\r60/A2[53] ), .Z(n771) );
  NOR U1960 ( .A(\r60/A2[53] ), .B(\r60/A1[53] ), .Z(n773) );
  MUX U1961 ( .IN0(n786), .IN1(Hi[22]), .SEL(n685), .F(n670) );
  NANDN U1962 ( .A(n787), .B(n788), .Z(n786) );
  AND U1963 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U1964 ( .A(n791), .B(n691), .Z(n790) );
  NANDN U1965 ( .A(n791), .B(\U3/U1/Z_0 ), .Z(n789) );
  XOR U1966 ( .A(n792), .B(n785), .Z(n791) );
  NANDN U1967 ( .A(n793), .B(n794), .Z(n785) );
  NANDN U1968 ( .A(n795), .B(n796), .Z(n794) );
  OR U1969 ( .A(n784), .B(n782), .Z(n792) );
  AND U1970 ( .A(\r60/A1[52] ), .B(\r60/A2[52] ), .Z(n782) );
  NOR U1971 ( .A(\r60/A2[52] ), .B(\r60/A1[52] ), .Z(n784) );
  MUX U1972 ( .IN0(n797), .IN1(Hi[21]), .SEL(n685), .F(n669) );
  NANDN U1973 ( .A(n798), .B(n799), .Z(n797) );
  AND U1974 ( .A(n800), .B(n801), .Z(n799) );
  NANDN U1975 ( .A(n802), .B(n691), .Z(n801) );
  NANDN U1976 ( .A(n802), .B(\U3/U1/Z_0 ), .Z(n800) );
  XOR U1977 ( .A(n803), .B(n796), .Z(n802) );
  NANDN U1978 ( .A(n804), .B(n805), .Z(n796) );
  NANDN U1979 ( .A(n806), .B(n807), .Z(n805) );
  OR U1980 ( .A(n795), .B(n793), .Z(n803) );
  AND U1981 ( .A(\r60/A1[51] ), .B(\r60/A2[51] ), .Z(n793) );
  NOR U1982 ( .A(\r60/A2[51] ), .B(\r60/A1[51] ), .Z(n795) );
  MUX U1983 ( .IN0(n808), .IN1(Hi[20]), .SEL(n685), .F(n668) );
  NANDN U1984 ( .A(n809), .B(n810), .Z(n808) );
  AND U1985 ( .A(n811), .B(n812), .Z(n810) );
  NANDN U1986 ( .A(n813), .B(n691), .Z(n812) );
  NANDN U1987 ( .A(n813), .B(\U3/U1/Z_0 ), .Z(n811) );
  XOR U1988 ( .A(n814), .B(n807), .Z(n813) );
  NANDN U1989 ( .A(n815), .B(n816), .Z(n807) );
  NANDN U1990 ( .A(n817), .B(n818), .Z(n816) );
  OR U1991 ( .A(n806), .B(n804), .Z(n814) );
  AND U1992 ( .A(\r60/A1[50] ), .B(\r60/A2[50] ), .Z(n804) );
  NOR U1993 ( .A(\r60/A2[50] ), .B(\r60/A1[50] ), .Z(n806) );
  MUX U1994 ( .IN0(n819), .IN1(Hi[19]), .SEL(n685), .F(n667) );
  NANDN U1995 ( .A(n820), .B(n821), .Z(n819) );
  AND U1996 ( .A(n822), .B(n823), .Z(n821) );
  NANDN U1997 ( .A(n824), .B(n691), .Z(n823) );
  NANDN U1998 ( .A(n824), .B(\U3/U1/Z_0 ), .Z(n822) );
  XOR U1999 ( .A(n825), .B(n818), .Z(n824) );
  NANDN U2000 ( .A(n826), .B(n827), .Z(n818) );
  NANDN U2001 ( .A(n828), .B(n829), .Z(n827) );
  OR U2002 ( .A(n817), .B(n815), .Z(n825) );
  AND U2003 ( .A(\r60/A1[49] ), .B(\r60/A2[49] ), .Z(n815) );
  NOR U2004 ( .A(\r60/A2[49] ), .B(\r60/A1[49] ), .Z(n817) );
  MUX U2005 ( .IN0(n830), .IN1(Hi[18]), .SEL(n685), .F(n666) );
  NANDN U2006 ( .A(n831), .B(n832), .Z(n830) );
  AND U2007 ( .A(n833), .B(n834), .Z(n832) );
  NANDN U2008 ( .A(n835), .B(n691), .Z(n834) );
  NANDN U2009 ( .A(n835), .B(\U3/U1/Z_0 ), .Z(n833) );
  XOR U2010 ( .A(n836), .B(n829), .Z(n835) );
  NANDN U2011 ( .A(n837), .B(n838), .Z(n829) );
  NAND U2012 ( .A(n839), .B(n840), .Z(n838) );
  NAND U2013 ( .A(n841), .B(n842), .Z(n839) );
  NAND U2014 ( .A(n843), .B(n844), .Z(n841) );
  NAND U2015 ( .A(n845), .B(n846), .Z(n843) );
  NAND U2016 ( .A(n847), .B(n848), .Z(n845) );
  NAND U2017 ( .A(n849), .B(n850), .Z(n847) );
  NAND U2018 ( .A(n851), .B(n852), .Z(n849) );
  NAND U2019 ( .A(n853), .B(n854), .Z(n851) );
  NANDN U2020 ( .A(n855), .B(n856), .Z(n853) );
  NAND U2021 ( .A(n857), .B(n858), .Z(n856) );
  AND U2022 ( .A(n859), .B(n860), .Z(n857) );
  NANDN U2023 ( .A(n861), .B(n862), .Z(n860) );
  NAND U2024 ( .A(n862), .B(n863), .Z(n859) );
  OR U2025 ( .A(n828), .B(n826), .Z(n836) );
  AND U2026 ( .A(\r60/A1[48] ), .B(\r60/A2[48] ), .Z(n826) );
  NOR U2027 ( .A(\r60/A2[48] ), .B(\r60/A1[48] ), .Z(n828) );
  MUX U2028 ( .IN0(n864), .IN1(Hi[17]), .SEL(n685), .F(n665) );
  NANDN U2029 ( .A(n865), .B(n866), .Z(n864) );
  AND U2030 ( .A(n867), .B(n868), .Z(n866) );
  NANDN U2031 ( .A(n869), .B(n691), .Z(n868) );
  NANDN U2032 ( .A(n869), .B(\U3/U1/Z_0 ), .Z(n867) );
  XNOR U2033 ( .A(n870), .B(n871), .Z(n869) );
  AND U2034 ( .A(n842), .B(n872), .Z(n871) );
  NAND U2035 ( .A(n844), .B(n873), .Z(n872) );
  NANDN U2036 ( .A(n837), .B(n840), .Z(n870) );
  OR U2037 ( .A(\r60/A1[47] ), .B(\r60/A2[47] ), .Z(n840) );
  AND U2038 ( .A(\r60/A1[47] ), .B(\r60/A2[47] ), .Z(n837) );
  MUX U2039 ( .IN0(n874), .IN1(Hi[16]), .SEL(n685), .F(n664) );
  NANDN U2040 ( .A(n875), .B(n876), .Z(n874) );
  AND U2041 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U2042 ( .A(n879), .B(n691), .Z(n878) );
  NANDN U2043 ( .A(n879), .B(\U3/U1/Z_0 ), .Z(n877) );
  XOR U2044 ( .A(n880), .B(n873), .Z(n879) );
  NAND U2045 ( .A(n881), .B(n846), .Z(n873) );
  NAND U2046 ( .A(n848), .B(n882), .Z(n881) );
  NAND U2047 ( .A(n842), .B(n844), .Z(n880) );
  OR U2048 ( .A(\r60/A2[46] ), .B(\r60/A1[46] ), .Z(n844) );
  NAND U2049 ( .A(\r60/A2[46] ), .B(\r60/A1[46] ), .Z(n842) );
  MUX U2050 ( .IN0(n883), .IN1(Hi[15]), .SEL(n685), .F(n663) );
  NANDN U2051 ( .A(n884), .B(n885), .Z(n883) );
  AND U2052 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U2053 ( .A(n888), .B(n691), .Z(n887) );
  NANDN U2054 ( .A(n888), .B(\U3/U1/Z_0 ), .Z(n886) );
  XOR U2055 ( .A(n889), .B(n882), .Z(n888) );
  NAND U2056 ( .A(n890), .B(n850), .Z(n882) );
  NANDN U2057 ( .A(n891), .B(n852), .Z(n890) );
  NAND U2058 ( .A(n846), .B(n848), .Z(n889) );
  OR U2059 ( .A(\r60/A2[45] ), .B(\r60/A1[45] ), .Z(n848) );
  NAND U2060 ( .A(\r60/A2[45] ), .B(\r60/A1[45] ), .Z(n846) );
  MUX U2061 ( .IN0(n892), .IN1(Hi[14]), .SEL(n685), .F(n662) );
  NANDN U2062 ( .A(n893), .B(n894), .Z(n892) );
  AND U2063 ( .A(n895), .B(n896), .Z(n894) );
  NANDN U2064 ( .A(n897), .B(n691), .Z(n896) );
  NANDN U2065 ( .A(n897), .B(\U3/U1/Z_0 ), .Z(n895) );
  XNOR U2066 ( .A(n898), .B(n891), .Z(n897) );
  AND U2067 ( .A(n854), .B(n899), .Z(n891) );
  OR U2068 ( .A(n900), .B(n855), .Z(n899) );
  NAND U2069 ( .A(n901), .B(n902), .Z(n855) );
  AND U2070 ( .A(n903), .B(n904), .Z(n902) );
  AND U2071 ( .A(n905), .B(n906), .Z(n901) );
  ANDN U2072 ( .B(n907), .A(n908), .Z(n854) );
  NAND U2073 ( .A(n909), .B(n905), .Z(n907) );
  NAND U2074 ( .A(n910), .B(n911), .Z(n909) );
  NAND U2075 ( .A(n912), .B(n904), .Z(n910) );
  NANDN U2076 ( .A(n913), .B(n914), .Z(n912) );
  NANDN U2077 ( .A(n915), .B(n903), .Z(n914) );
  IV U2078 ( .A(n916), .Z(n915) );
  NAND U2079 ( .A(n850), .B(n852), .Z(n898) );
  OR U2080 ( .A(\r60/A2[44] ), .B(\r60/A1[44] ), .Z(n852) );
  NAND U2081 ( .A(\r60/A2[44] ), .B(\r60/A1[44] ), .Z(n850) );
  MUX U2082 ( .IN0(n917), .IN1(Hi[13]), .SEL(n685), .F(n661) );
  NANDN U2083 ( .A(n918), .B(n919), .Z(n917) );
  AND U2084 ( .A(n920), .B(n921), .Z(n919) );
  NANDN U2085 ( .A(n922), .B(n691), .Z(n921) );
  NANDN U2086 ( .A(n922), .B(\U3/U1/Z_0 ), .Z(n920) );
  XNOR U2087 ( .A(n923), .B(n924), .Z(n922) );
  AND U2088 ( .A(n911), .B(n925), .Z(n924) );
  NAND U2089 ( .A(n904), .B(n926), .Z(n925) );
  NANDN U2090 ( .A(n908), .B(n905), .Z(n923) );
  OR U2091 ( .A(\r60/A2[43] ), .B(\r60/A1[43] ), .Z(n905) );
  AND U2092 ( .A(\r60/A2[43] ), .B(\r60/A1[43] ), .Z(n908) );
  MUX U2093 ( .IN0(n927), .IN1(Hi[12]), .SEL(n685), .F(n660) );
  NANDN U2094 ( .A(n928), .B(n929), .Z(n927) );
  AND U2095 ( .A(n930), .B(n931), .Z(n929) );
  NANDN U2096 ( .A(n932), .B(n691), .Z(n931) );
  NANDN U2097 ( .A(n932), .B(\U3/U1/Z_0 ), .Z(n930) );
  XOR U2098 ( .A(n933), .B(n926), .Z(n932) );
  NAND U2099 ( .A(n934), .B(n935), .Z(n926) );
  NANDN U2100 ( .A(n936), .B(n903), .Z(n935) );
  IV U2101 ( .A(n913), .Z(n934) );
  NAND U2102 ( .A(n904), .B(n911), .Z(n933) );
  NAND U2103 ( .A(\r60/A2[42] ), .B(\r60/A1[42] ), .Z(n911) );
  OR U2104 ( .A(\r60/A2[42] ), .B(\r60/A1[42] ), .Z(n904) );
  MUX U2105 ( .IN0(n937), .IN1(Hi[11]), .SEL(n685), .F(n659) );
  NANDN U2106 ( .A(n938), .B(n939), .Z(n937) );
  AND U2107 ( .A(n940), .B(n941), .Z(n939) );
  NANDN U2108 ( .A(n942), .B(n691), .Z(n941) );
  NANDN U2109 ( .A(n942), .B(\U3/U1/Z_0 ), .Z(n940) );
  XNOR U2110 ( .A(n943), .B(n936), .Z(n942) );
  ANDN U2111 ( .B(n944), .A(n916), .Z(n936) );
  NANDN U2112 ( .A(n900), .B(n906), .Z(n944) );
  NANDN U2113 ( .A(n913), .B(n903), .Z(n943) );
  OR U2114 ( .A(\r60/A1[41] ), .B(\r60/A2[41] ), .Z(n903) );
  AND U2115 ( .A(\r60/A1[41] ), .B(\r60/A2[41] ), .Z(n913) );
  MUX U2116 ( .IN0(n945), .IN1(Hi[10]), .SEL(n685), .F(n658) );
  NANDN U2117 ( .A(n946), .B(n947), .Z(n945) );
  AND U2118 ( .A(n948), .B(n949), .Z(n947) );
  NANDN U2119 ( .A(n950), .B(n691), .Z(n949) );
  NANDN U2120 ( .A(n950), .B(\U3/U1/Z_0 ), .Z(n948) );
  XNOR U2121 ( .A(n951), .B(n900), .Z(n950) );
  AND U2122 ( .A(n858), .B(n952), .Z(n900) );
  NAND U2123 ( .A(n953), .B(n862), .Z(n952) );
  AND U2124 ( .A(n954), .B(n955), .Z(n862) );
  AND U2125 ( .A(n956), .B(n957), .Z(n955) );
  AND U2126 ( .A(n958), .B(n959), .Z(n954) );
  ANDN U2127 ( .B(n960), .A(n961), .Z(n858) );
  NAND U2128 ( .A(n962), .B(n958), .Z(n960) );
  NAND U2129 ( .A(n963), .B(n964), .Z(n962) );
  NAND U2130 ( .A(n965), .B(n957), .Z(n963) );
  NANDN U2131 ( .A(n966), .B(n967), .Z(n965) );
  NANDN U2132 ( .A(n968), .B(n956), .Z(n967) );
  NANDN U2133 ( .A(n916), .B(n906), .Z(n951) );
  OR U2134 ( .A(\r60/A2[40] ), .B(\r60/A1[40] ), .Z(n906) );
  AND U2135 ( .A(\r60/A2[40] ), .B(\r60/A1[40] ), .Z(n916) );
  MUX U2136 ( .IN0(n969), .IN1(Hi[9]), .SEL(n685), .F(n657) );
  NANDN U2137 ( .A(n970), .B(n971), .Z(n969) );
  AND U2138 ( .A(n972), .B(n973), .Z(n971) );
  NANDN U2139 ( .A(n974), .B(n691), .Z(n973) );
  NANDN U2140 ( .A(n974), .B(\U3/U1/Z_0 ), .Z(n972) );
  XNOR U2141 ( .A(n975), .B(n976), .Z(n974) );
  AND U2142 ( .A(n964), .B(n977), .Z(n976) );
  NAND U2143 ( .A(n957), .B(n978), .Z(n977) );
  NANDN U2144 ( .A(n961), .B(n958), .Z(n975) );
  OR U2145 ( .A(\r60/A2[39] ), .B(\r60/A1[39] ), .Z(n958) );
  AND U2146 ( .A(\r60/A1[39] ), .B(\r60/A2[39] ), .Z(n961) );
  MUX U2147 ( .IN0(n979), .IN1(Hi[8]), .SEL(n685), .F(n656) );
  NANDN U2148 ( .A(n980), .B(n981), .Z(n979) );
  AND U2149 ( .A(n982), .B(n983), .Z(n981) );
  NANDN U2150 ( .A(n984), .B(n691), .Z(n983) );
  NANDN U2151 ( .A(n984), .B(\U3/U1/Z_0 ), .Z(n982) );
  XOR U2152 ( .A(n985), .B(n978), .Z(n984) );
  NAND U2153 ( .A(n986), .B(n987), .Z(n978) );
  NANDN U2154 ( .A(n988), .B(n956), .Z(n987) );
  NAND U2155 ( .A(n957), .B(n964), .Z(n985) );
  NAND U2156 ( .A(\r60/A2[38] ), .B(\r60/A1[38] ), .Z(n964) );
  OR U2157 ( .A(\r60/A1[38] ), .B(\r60/A2[38] ), .Z(n957) );
  MUX U2158 ( .IN0(n989), .IN1(Hi[7]), .SEL(n685), .F(n655) );
  NANDN U2159 ( .A(n990), .B(n991), .Z(n989) );
  AND U2160 ( .A(n992), .B(n993), .Z(n991) );
  NANDN U2161 ( .A(n994), .B(n691), .Z(n993) );
  NANDN U2162 ( .A(n994), .B(\U3/U1/Z_0 ), .Z(n992) );
  XNOR U2163 ( .A(n995), .B(n988), .Z(n994) );
  AND U2164 ( .A(n996), .B(n968), .Z(n988) );
  NAND U2165 ( .A(n959), .B(n953), .Z(n996) );
  NANDN U2166 ( .A(n966), .B(n956), .Z(n995) );
  OR U2167 ( .A(\r60/A1[37] ), .B(\r60/A2[37] ), .Z(n956) );
  IV U2168 ( .A(n986), .Z(n966) );
  NAND U2169 ( .A(\r60/A2[37] ), .B(\r60/A1[37] ), .Z(n986) );
  MUX U2170 ( .IN0(n997), .IN1(Hi[6]), .SEL(n685), .F(n654) );
  NANDN U2171 ( .A(n998), .B(n999), .Z(n997) );
  AND U2172 ( .A(n1000), .B(n1001), .Z(n999) );
  NANDN U2173 ( .A(n1002), .B(n691), .Z(n1001) );
  NANDN U2174 ( .A(n1002), .B(\U3/U1/Z_0 ), .Z(n1000) );
  XOR U2175 ( .A(n1003), .B(n953), .Z(n1002) );
  NANDN U2176 ( .A(n863), .B(n861), .Z(n953) );
  NAND U2177 ( .A(n1004), .B(n1005), .Z(n861) );
  AND U2178 ( .A(n1006), .B(n1007), .Z(n1005) );
  AND U2179 ( .A(n1008), .B(n1009), .Z(n1007) );
  AND U2180 ( .A(n1010), .B(n1011), .Z(n1004) );
  NANDN U2181 ( .A(n1012), .B(n1013), .Z(n863) );
  NAND U2182 ( .A(n1014), .B(n1010), .Z(n1013) );
  NAND U2183 ( .A(n1015), .B(n1016), .Z(n1014) );
  NAND U2184 ( .A(n1017), .B(n1006), .Z(n1015) );
  NANDN U2185 ( .A(n1018), .B(n1019), .Z(n1017) );
  NANDN U2186 ( .A(n1020), .B(n1011), .Z(n1019) );
  NAND U2187 ( .A(n968), .B(n959), .Z(n1003) );
  OR U2188 ( .A(\r60/A1[36] ), .B(\r60/A2[36] ), .Z(n959) );
  NAND U2189 ( .A(\r60/A2[36] ), .B(\r60/A1[36] ), .Z(n968) );
  MUX U2190 ( .IN0(n1021), .IN1(Hi[5]), .SEL(n685), .F(n653) );
  NANDN U2191 ( .A(n1022), .B(n1023), .Z(n1021) );
  AND U2192 ( .A(n1024), .B(n1025), .Z(n1023) );
  NANDN U2193 ( .A(n1026), .B(n691), .Z(n1025) );
  NANDN U2194 ( .A(n1026), .B(\U3/U1/Z_0 ), .Z(n1024) );
  XNOR U2195 ( .A(n1027), .B(n1028), .Z(n1026) );
  AND U2196 ( .A(n1016), .B(n1029), .Z(n1028) );
  NAND U2197 ( .A(n1006), .B(n1030), .Z(n1029) );
  NANDN U2198 ( .A(n1012), .B(n1010), .Z(n1027) );
  OR U2199 ( .A(\r60/A2[35] ), .B(\r60/A1[35] ), .Z(n1010) );
  AND U2200 ( .A(\r60/A2[35] ), .B(\r60/A1[35] ), .Z(n1012) );
  MUX U2201 ( .IN0(n1031), .IN1(Hi[4]), .SEL(n685), .F(n652) );
  NANDN U2202 ( .A(n1032), .B(n1033), .Z(n1031) );
  AND U2203 ( .A(n1034), .B(n1035), .Z(n1033) );
  NANDN U2204 ( .A(n1036), .B(n691), .Z(n1035) );
  NANDN U2205 ( .A(n1036), .B(\U3/U1/Z_0 ), .Z(n1034) );
  XOR U2206 ( .A(n1037), .B(n1030), .Z(n1036) );
  NAND U2207 ( .A(n1038), .B(n1039), .Z(n1030) );
  NAND U2208 ( .A(n1011), .B(n1040), .Z(n1039) );
  IV U2209 ( .A(n1018), .Z(n1038) );
  NAND U2210 ( .A(n1006), .B(n1016), .Z(n1037) );
  NAND U2211 ( .A(\r60/A1[34] ), .B(\r60/A2[34] ), .Z(n1016) );
  OR U2212 ( .A(\r60/A1[34] ), .B(\r60/A2[34] ), .Z(n1006) );
  MUX U2213 ( .IN0(n1041), .IN1(Hi[3]), .SEL(n685), .F(n651) );
  NANDN U2214 ( .A(n1042), .B(n1043), .Z(n1041) );
  AND U2215 ( .A(n1044), .B(n1045), .Z(n1043) );
  NANDN U2216 ( .A(n1046), .B(n691), .Z(n1045) );
  NANDN U2217 ( .A(n1046), .B(\U3/U1/Z_0 ), .Z(n1044) );
  XOR U2218 ( .A(n1047), .B(n1040), .Z(n1046) );
  NAND U2219 ( .A(n1048), .B(n1020), .Z(n1040) );
  NAND U2220 ( .A(n1009), .B(n1008), .Z(n1048) );
  NANDN U2221 ( .A(n1018), .B(n1011), .Z(n1047) );
  OR U2222 ( .A(\r60/A1[33] ), .B(\r60/A2[33] ), .Z(n1011) );
  AND U2223 ( .A(\r60/A1[33] ), .B(\r60/A2[33] ), .Z(n1018) );
  MUX U2224 ( .IN0(n1049), .IN1(Hi[2]), .SEL(n685), .F(n650) );
  NANDN U2225 ( .A(n1050), .B(n1051), .Z(n1049) );
  AND U2226 ( .A(n1052), .B(n1053), .Z(n1051) );
  NANDN U2227 ( .A(n1054), .B(n691), .Z(n1053) );
  NANDN U2228 ( .A(n1054), .B(\U3/U1/Z_0 ), .Z(n1052) );
  XOR U2229 ( .A(n1055), .B(n1008), .Z(n1054) );
  NANDN U2230 ( .A(n1056), .B(n1057), .Z(n1008) );
  NANDN U2231 ( .A(n1058), .B(n1059), .Z(n1057) );
  NAND U2232 ( .A(n1020), .B(n1009), .Z(n1055) );
  OR U2233 ( .A(\r60/A1[32] ), .B(\r60/A2[32] ), .Z(n1009) );
  NAND U2234 ( .A(\r60/A2[32] ), .B(\r60/A1[32] ), .Z(n1020) );
  MUX U2235 ( .IN0(n1060), .IN1(Hi[1]), .SEL(n685), .F(n649) );
  NANDN U2236 ( .A(n1061), .B(n1062), .Z(n1060) );
  AND U2237 ( .A(n1063), .B(n1064), .Z(n1062) );
  NANDN U2238 ( .A(n1065), .B(n691), .Z(n1064) );
  NANDN U2239 ( .A(n1065), .B(\U3/U1/Z_0 ), .Z(n1063) );
  XNOR U2240 ( .A(n1066), .B(n1058), .Z(n1065) );
  NANDN U2241 ( .A(n1056), .B(n1059), .Z(n1066) );
  OR U2242 ( .A(\r60/A2[31] ), .B(\r60/A1[31] ), .Z(n1059) );
  AND U2243 ( .A(\r60/A2[31] ), .B(\r60/A1[31] ), .Z(n1056) );
  MUX U2244 ( .IN0(n1067), .IN1(Hi[0]), .SEL(n685), .F(n648) );
  ANDN U2245 ( .B(n1068), .A(n1069), .Z(n685) );
  AND U2246 ( .A(n1070), .B(n1071), .Z(n1068) );
  NANDN U2247 ( .A(n1072), .B(n1073), .Z(n1071) );
  NANDN U2248 ( .A(n1074), .B(n1075), .Z(n1067) );
  AND U2249 ( .A(n1076), .B(n1077), .Z(n1075) );
  NAND U2250 ( .A(n1078), .B(n691), .Z(n1077) );
  NAND U2251 ( .A(\U3/U1/Z_0 ), .B(n1078), .Z(n1076) );
  AND U2252 ( .A(n1079), .B(n1058), .Z(n1078) );
  NAND U2253 ( .A(\r60/A2[30] ), .B(\r60/A1[30] ), .Z(n1058) );
  OR U2254 ( .A(\r60/A1[30] ), .B(\r60/A2[30] ), .Z(n1079) );
  MUX U2255 ( .IN0(n1080), .IN1(Lo[31]), .SEL(n1081), .F(n647) );
  NAND U2256 ( .A(n1082), .B(n1083), .Z(n1080) );
  NAND U2257 ( .A(\U3/U1/Z_0 ), .B(N148), .Z(n1083) );
  ANDN U2258 ( .B(n1084), .A(n686), .Z(n1082) );
  NOR U2259 ( .A(n682), .B(n1085), .Z(n686) );
  IV U2260 ( .A(a[31]), .Z(n682) );
  NAND U2261 ( .A(n691), .B(N148), .Z(n1084) );
  MUX U2262 ( .IN0(n1086), .IN1(Lo[30]), .SEL(n1081), .F(n646) );
  NAND U2263 ( .A(n1087), .B(n1088), .Z(n1086) );
  NAND U2264 ( .A(\U3/U1/Z_0 ), .B(N147), .Z(n1088) );
  ANDN U2265 ( .B(n1089), .A(n699), .Z(n1087) );
  ANDN U2266 ( .B(a[30]), .A(n1085), .Z(n699) );
  NAND U2267 ( .A(n691), .B(N147), .Z(n1089) );
  MUX U2268 ( .IN0(n1090), .IN1(Lo[29]), .SEL(n1081), .F(n645) );
  NAND U2269 ( .A(n1091), .B(n1092), .Z(n1090) );
  NAND U2270 ( .A(\U3/U1/Z_0 ), .B(N146), .Z(n1092) );
  ANDN U2271 ( .B(n1093), .A(n710), .Z(n1091) );
  ANDN U2272 ( .B(a[29]), .A(n1085), .Z(n710) );
  NAND U2273 ( .A(n691), .B(N146), .Z(n1093) );
  MUX U2274 ( .IN0(n1094), .IN1(Lo[28]), .SEL(n1081), .F(n644) );
  NAND U2275 ( .A(n1095), .B(n1096), .Z(n1094) );
  NAND U2276 ( .A(\U3/U1/Z_0 ), .B(N145), .Z(n1096) );
  ANDN U2277 ( .B(n1097), .A(n721), .Z(n1095) );
  ANDN U2278 ( .B(a[28]), .A(n1085), .Z(n721) );
  NAND U2279 ( .A(n691), .B(N145), .Z(n1097) );
  MUX U2280 ( .IN0(n1098), .IN1(Lo[27]), .SEL(n1081), .F(n643) );
  NAND U2281 ( .A(n1099), .B(n1100), .Z(n1098) );
  NAND U2282 ( .A(\U3/U1/Z_0 ), .B(N144), .Z(n1100) );
  ANDN U2283 ( .B(n1101), .A(n732), .Z(n1099) );
  ANDN U2284 ( .B(a[27]), .A(n1085), .Z(n732) );
  NAND U2285 ( .A(n691), .B(N144), .Z(n1101) );
  MUX U2286 ( .IN0(n1102), .IN1(Lo[26]), .SEL(n1081), .F(n642) );
  NAND U2287 ( .A(n1103), .B(n1104), .Z(n1102) );
  NAND U2288 ( .A(\U3/U1/Z_0 ), .B(N143), .Z(n1104) );
  ANDN U2289 ( .B(n1105), .A(n743), .Z(n1103) );
  ANDN U2290 ( .B(a[26]), .A(n1085), .Z(n743) );
  NAND U2291 ( .A(n691), .B(N143), .Z(n1105) );
  MUX U2292 ( .IN0(n1106), .IN1(Lo[25]), .SEL(n1081), .F(n641) );
  NAND U2293 ( .A(n1107), .B(n1108), .Z(n1106) );
  NAND U2294 ( .A(\U3/U1/Z_0 ), .B(N142), .Z(n1108) );
  ANDN U2295 ( .B(n1109), .A(n754), .Z(n1107) );
  ANDN U2296 ( .B(a[25]), .A(n1085), .Z(n754) );
  NAND U2297 ( .A(n691), .B(N142), .Z(n1109) );
  MUX U2298 ( .IN0(n1110), .IN1(Lo[24]), .SEL(n1081), .F(n640) );
  NAND U2299 ( .A(n1111), .B(n1112), .Z(n1110) );
  NAND U2300 ( .A(\U3/U1/Z_0 ), .B(N141), .Z(n1112) );
  ANDN U2301 ( .B(n1113), .A(n765), .Z(n1111) );
  ANDN U2302 ( .B(a[24]), .A(n1085), .Z(n765) );
  NAND U2303 ( .A(n691), .B(N141), .Z(n1113) );
  MUX U2304 ( .IN0(n1114), .IN1(Lo[23]), .SEL(n1081), .F(n639) );
  NAND U2305 ( .A(n1115), .B(n1116), .Z(n1114) );
  NAND U2306 ( .A(\U3/U1/Z_0 ), .B(N140), .Z(n1116) );
  ANDN U2307 ( .B(n1117), .A(n776), .Z(n1115) );
  ANDN U2308 ( .B(a[23]), .A(n1085), .Z(n776) );
  NAND U2309 ( .A(n691), .B(N140), .Z(n1117) );
  MUX U2310 ( .IN0(n1118), .IN1(Lo[22]), .SEL(n1081), .F(n638) );
  NAND U2311 ( .A(n1119), .B(n1120), .Z(n1118) );
  NAND U2312 ( .A(\U3/U1/Z_0 ), .B(N139), .Z(n1120) );
  ANDN U2313 ( .B(n1121), .A(n787), .Z(n1119) );
  ANDN U2314 ( .B(a[22]), .A(n1085), .Z(n787) );
  NAND U2315 ( .A(n691), .B(N139), .Z(n1121) );
  MUX U2316 ( .IN0(n1122), .IN1(Lo[21]), .SEL(n1081), .F(n637) );
  NAND U2317 ( .A(n1123), .B(n1124), .Z(n1122) );
  NAND U2318 ( .A(\U3/U1/Z_0 ), .B(N138), .Z(n1124) );
  ANDN U2319 ( .B(n1125), .A(n798), .Z(n1123) );
  ANDN U2320 ( .B(a[21]), .A(n1085), .Z(n798) );
  NAND U2321 ( .A(n691), .B(N138), .Z(n1125) );
  MUX U2322 ( .IN0(n1126), .IN1(Lo[20]), .SEL(n1081), .F(n636) );
  NAND U2323 ( .A(n1127), .B(n1128), .Z(n1126) );
  NAND U2324 ( .A(\U3/U1/Z_0 ), .B(N137), .Z(n1128) );
  ANDN U2325 ( .B(n1129), .A(n809), .Z(n1127) );
  ANDN U2326 ( .B(a[20]), .A(n1085), .Z(n809) );
  NAND U2327 ( .A(n691), .B(N137), .Z(n1129) );
  MUX U2328 ( .IN0(n1130), .IN1(Lo[19]), .SEL(n1081), .F(n635) );
  NAND U2329 ( .A(n1131), .B(n1132), .Z(n1130) );
  NAND U2330 ( .A(\U3/U1/Z_0 ), .B(N136), .Z(n1132) );
  ANDN U2331 ( .B(n1133), .A(n820), .Z(n1131) );
  ANDN U2332 ( .B(a[19]), .A(n1085), .Z(n820) );
  NAND U2333 ( .A(n691), .B(N136), .Z(n1133) );
  MUX U2334 ( .IN0(n1134), .IN1(Lo[18]), .SEL(n1081), .F(n634) );
  NAND U2335 ( .A(n1135), .B(n1136), .Z(n1134) );
  NAND U2336 ( .A(\U3/U1/Z_0 ), .B(N135), .Z(n1136) );
  ANDN U2337 ( .B(n1137), .A(n831), .Z(n1135) );
  ANDN U2338 ( .B(a[18]), .A(n1085), .Z(n831) );
  NAND U2339 ( .A(n691), .B(N135), .Z(n1137) );
  MUX U2340 ( .IN0(n1138), .IN1(Lo[17]), .SEL(n1081), .F(n633) );
  NAND U2341 ( .A(n1139), .B(n1140), .Z(n1138) );
  NAND U2342 ( .A(\U3/U1/Z_0 ), .B(N134), .Z(n1140) );
  ANDN U2343 ( .B(n1141), .A(n865), .Z(n1139) );
  ANDN U2344 ( .B(a[17]), .A(n1085), .Z(n865) );
  NAND U2345 ( .A(n691), .B(N134), .Z(n1141) );
  MUX U2346 ( .IN0(n1142), .IN1(Lo[16]), .SEL(n1081), .F(n632) );
  NAND U2347 ( .A(n1143), .B(n1144), .Z(n1142) );
  NAND U2348 ( .A(\U3/U1/Z_0 ), .B(N133), .Z(n1144) );
  ANDN U2349 ( .B(n1145), .A(n875), .Z(n1143) );
  ANDN U2350 ( .B(a[16]), .A(n1085), .Z(n875) );
  NAND U2351 ( .A(n691), .B(N133), .Z(n1145) );
  MUX U2352 ( .IN0(n1146), .IN1(Lo[15]), .SEL(n1081), .F(n631) );
  NAND U2353 ( .A(n1147), .B(n1148), .Z(n1146) );
  NAND U2354 ( .A(\U3/U1/Z_0 ), .B(N132), .Z(n1148) );
  ANDN U2355 ( .B(n1149), .A(n884), .Z(n1147) );
  ANDN U2356 ( .B(a[15]), .A(n1085), .Z(n884) );
  NAND U2357 ( .A(n691), .B(N132), .Z(n1149) );
  MUX U2358 ( .IN0(n1150), .IN1(Lo[14]), .SEL(n1081), .F(n630) );
  NAND U2359 ( .A(n1151), .B(n1152), .Z(n1150) );
  NAND U2360 ( .A(\U3/U1/Z_0 ), .B(N131), .Z(n1152) );
  ANDN U2361 ( .B(n1153), .A(n893), .Z(n1151) );
  ANDN U2362 ( .B(a[14]), .A(n1085), .Z(n893) );
  NAND U2363 ( .A(n691), .B(N131), .Z(n1153) );
  MUX U2364 ( .IN0(n1154), .IN1(Lo[13]), .SEL(n1081), .F(n629) );
  NAND U2365 ( .A(n1155), .B(n1156), .Z(n1154) );
  NAND U2366 ( .A(\U3/U1/Z_0 ), .B(N130), .Z(n1156) );
  ANDN U2367 ( .B(n1157), .A(n918), .Z(n1155) );
  ANDN U2368 ( .B(a[13]), .A(n1085), .Z(n918) );
  NAND U2369 ( .A(n691), .B(N130), .Z(n1157) );
  MUX U2370 ( .IN0(n1158), .IN1(Lo[12]), .SEL(n1081), .F(n628) );
  NAND U2371 ( .A(n1159), .B(n1160), .Z(n1158) );
  NAND U2372 ( .A(\U3/U1/Z_0 ), .B(N129), .Z(n1160) );
  ANDN U2373 ( .B(n1161), .A(n928), .Z(n1159) );
  ANDN U2374 ( .B(a[12]), .A(n1085), .Z(n928) );
  NAND U2375 ( .A(n691), .B(N129), .Z(n1161) );
  MUX U2376 ( .IN0(n1162), .IN1(Lo[11]), .SEL(n1081), .F(n627) );
  NAND U2377 ( .A(n1163), .B(n1164), .Z(n1162) );
  NAND U2378 ( .A(\U3/U1/Z_0 ), .B(N128), .Z(n1164) );
  ANDN U2379 ( .B(n1165), .A(n938), .Z(n1163) );
  ANDN U2380 ( .B(a[11]), .A(n1085), .Z(n938) );
  NAND U2381 ( .A(n691), .B(N128), .Z(n1165) );
  MUX U2382 ( .IN0(n1166), .IN1(Lo[10]), .SEL(n1081), .F(n626) );
  NAND U2383 ( .A(n1167), .B(n1168), .Z(n1166) );
  NAND U2384 ( .A(\U3/U1/Z_0 ), .B(N127), .Z(n1168) );
  ANDN U2385 ( .B(n1169), .A(n946), .Z(n1167) );
  ANDN U2386 ( .B(a[10]), .A(n1085), .Z(n946) );
  NAND U2387 ( .A(n691), .B(N127), .Z(n1169) );
  MUX U2388 ( .IN0(n1170), .IN1(Lo[9]), .SEL(n1081), .F(n625) );
  NAND U2389 ( .A(n1171), .B(n1172), .Z(n1170) );
  NAND U2390 ( .A(\U3/U1/Z_0 ), .B(N126), .Z(n1172) );
  ANDN U2391 ( .B(n1173), .A(n970), .Z(n1171) );
  ANDN U2392 ( .B(a[9]), .A(n1085), .Z(n970) );
  NAND U2393 ( .A(n691), .B(N126), .Z(n1173) );
  MUX U2394 ( .IN0(n1174), .IN1(Lo[8]), .SEL(n1081), .F(n624) );
  NAND U2395 ( .A(n1175), .B(n1176), .Z(n1174) );
  NAND U2396 ( .A(\U3/U1/Z_0 ), .B(N125), .Z(n1176) );
  ANDN U2397 ( .B(n1177), .A(n980), .Z(n1175) );
  ANDN U2398 ( .B(a[8]), .A(n1085), .Z(n980) );
  NAND U2399 ( .A(n691), .B(N125), .Z(n1177) );
  MUX U2400 ( .IN0(n1178), .IN1(Lo[7]), .SEL(n1081), .F(n623) );
  NAND U2401 ( .A(n1179), .B(n1180), .Z(n1178) );
  NAND U2402 ( .A(\U3/U1/Z_0 ), .B(N124), .Z(n1180) );
  ANDN U2403 ( .B(n1181), .A(n990), .Z(n1179) );
  ANDN U2404 ( .B(a[7]), .A(n1085), .Z(n990) );
  NAND U2405 ( .A(n691), .B(N124), .Z(n1181) );
  MUX U2406 ( .IN0(n1182), .IN1(Lo[6]), .SEL(n1081), .F(n622) );
  NAND U2407 ( .A(n1183), .B(n1184), .Z(n1182) );
  NAND U2408 ( .A(\U3/U1/Z_0 ), .B(N123), .Z(n1184) );
  ANDN U2409 ( .B(n1185), .A(n998), .Z(n1183) );
  ANDN U2410 ( .B(a[6]), .A(n1085), .Z(n998) );
  NAND U2411 ( .A(n691), .B(N123), .Z(n1185) );
  MUX U2412 ( .IN0(n1186), .IN1(Lo[5]), .SEL(n1081), .F(n621) );
  NAND U2413 ( .A(n1187), .B(n1188), .Z(n1186) );
  NAND U2414 ( .A(\U3/U1/Z_0 ), .B(N122), .Z(n1188) );
  ANDN U2415 ( .B(n1189), .A(n1022), .Z(n1187) );
  ANDN U2416 ( .B(a[5]), .A(n1085), .Z(n1022) );
  NAND U2417 ( .A(n691), .B(N122), .Z(n1189) );
  MUX U2418 ( .IN0(n1190), .IN1(Lo[4]), .SEL(n1081), .F(n620) );
  NAND U2419 ( .A(n1191), .B(n1192), .Z(n1190) );
  NAND U2420 ( .A(\U3/U1/Z_0 ), .B(N121), .Z(n1192) );
  ANDN U2421 ( .B(n1193), .A(n1032), .Z(n1191) );
  ANDN U2422 ( .B(a[4]), .A(n1085), .Z(n1032) );
  NAND U2423 ( .A(n691), .B(N121), .Z(n1193) );
  MUX U2424 ( .IN0(n1194), .IN1(Lo[3]), .SEL(n1081), .F(n619) );
  NAND U2425 ( .A(n1195), .B(n1196), .Z(n1194) );
  NAND U2426 ( .A(\U3/U1/Z_0 ), .B(N120), .Z(n1196) );
  ANDN U2427 ( .B(n1197), .A(n1042), .Z(n1195) );
  ANDN U2428 ( .B(a[3]), .A(n1085), .Z(n1042) );
  NAND U2429 ( .A(n691), .B(N120), .Z(n1197) );
  MUX U2430 ( .IN0(n1198), .IN1(Lo[2]), .SEL(n1081), .F(n618) );
  NAND U2431 ( .A(n1199), .B(n1200), .Z(n1198) );
  NAND U2432 ( .A(\U3/U1/Z_0 ), .B(N119), .Z(n1200) );
  ANDN U2433 ( .B(n1201), .A(n1050), .Z(n1199) );
  ANDN U2434 ( .B(a[2]), .A(n1085), .Z(n1050) );
  NAND U2435 ( .A(n691), .B(N119), .Z(n1201) );
  MUX U2436 ( .IN0(n1202), .IN1(Lo[1]), .SEL(n1081), .F(n617) );
  NAND U2437 ( .A(n1203), .B(n1204), .Z(n1202) );
  NAND U2438 ( .A(\U3/U1/Z_0 ), .B(N118), .Z(n1204) );
  ANDN U2439 ( .B(n1205), .A(n1061), .Z(n1203) );
  ANDN U2440 ( .B(a[1]), .A(n1085), .Z(n1061) );
  NAND U2441 ( .A(n691), .B(N118), .Z(n1205) );
  MUX U2442 ( .IN0(n1206), .IN1(Lo[0]), .SEL(n1081), .F(n616) );
  ANDN U2443 ( .B(n1207), .A(n1069), .Z(n1081) );
  NAND U2444 ( .A(n1208), .B(n1209), .Z(n1069) );
  OR U2445 ( .A(n1210), .B(n1211), .Z(n1209) );
  OR U2446 ( .A(n1210), .B(n1212), .Z(n1208) );
  AND U2447 ( .A(n1213), .B(n1214), .Z(n1210) );
  AND U2448 ( .A(n1215), .B(n1216), .Z(n1214) );
  AND U2449 ( .A(n1217), .B(n1218), .Z(n1216) );
  AND U2450 ( .A(n1219), .B(n1220), .Z(n1218) );
  NOR U2451 ( .A(b[8]), .B(b[9]), .Z(n1220) );
  NOR U2452 ( .A(b[6]), .B(b[7]), .Z(n1219) );
  AND U2453 ( .A(n1221), .B(n1222), .Z(n1217) );
  NOR U2454 ( .A(b[4]), .B(b[5]), .Z(n1222) );
  NOR U2455 ( .A(b[31]), .B(b[3]), .Z(n1221) );
  AND U2456 ( .A(n1223), .B(n1224), .Z(n1215) );
  AND U2457 ( .A(n1225), .B(n1226), .Z(n1224) );
  NOR U2458 ( .A(b[2]), .B(b[30]), .Z(n1226) );
  NOR U2459 ( .A(b[28]), .B(b[29]), .Z(n1225) );
  AND U2460 ( .A(n1227), .B(n1228), .Z(n1223) );
  NOR U2461 ( .A(b[26]), .B(b[27]), .Z(n1228) );
  NOR U2462 ( .A(b[24]), .B(b[25]), .Z(n1227) );
  AND U2463 ( .A(n1229), .B(n1230), .Z(n1213) );
  AND U2464 ( .A(n1231), .B(n1232), .Z(n1230) );
  AND U2465 ( .A(n1233), .B(n1234), .Z(n1232) );
  NOR U2466 ( .A(b[22]), .B(b[23]), .Z(n1234) );
  NOR U2467 ( .A(b[20]), .B(b[21]), .Z(n1233) );
  AND U2468 ( .A(n1235), .B(n1236), .Z(n1231) );
  NOR U2469 ( .A(b[19]), .B(b[1]), .Z(n1236) );
  NOR U2470 ( .A(b[17]), .B(b[18]), .Z(n1235) );
  AND U2471 ( .A(n1237), .B(n1238), .Z(n1229) );
  AND U2472 ( .A(n1239), .B(n1240), .Z(n1238) );
  NOR U2473 ( .A(b[15]), .B(b[16]), .Z(n1240) );
  NOR U2474 ( .A(b[13]), .B(b[14]), .Z(n1239) );
  AND U2475 ( .A(n1241), .B(n1242), .Z(n1237) );
  NOR U2476 ( .A(b[11]), .B(b[12]), .Z(n1242) );
  NOR U2477 ( .A(b[0]), .B(b[10]), .Z(n1241) );
  AND U2478 ( .A(n1070), .B(n1243), .Z(n1207) );
  NANDN U2479 ( .A(n1244), .B(n1245), .Z(n1243) );
  NOR U2480 ( .A(\U3/U1/Z_0 ), .B(n691), .Z(n1070) );
  NAND U2481 ( .A(n1246), .B(n1247), .Z(n1206) );
  NANDN U2482 ( .A(n1248), .B(\U3/U1/Z_0 ), .Z(n1247) );
  ANDN U2483 ( .B(n1249), .A(n1074), .Z(n1246) );
  ANDN U2484 ( .B(a[0]), .A(n1085), .Z(n1074) );
  NANDN U2485 ( .A(n1250), .B(n1251), .Z(n1085) );
  AND U2486 ( .A(n1212), .B(n1252), .Z(n1251) );
  NAND U2487 ( .A(n1253), .B(mult_func[3]), .Z(n1212) );
  NOR U2488 ( .A(mult_func[2]), .B(n1072), .Z(n1253) );
  OR U2489 ( .A(mult_func[0]), .B(mult_func[1]), .Z(n1072) );
  NANDN U2490 ( .A(n1248), .B(n691), .Z(n1249) );
  NOR U2491 ( .A(n1250), .B(n1252), .Z(n691) );
  NANDN U2492 ( .A(n683), .B(b[0]), .Z(n1248) );
  IV U2493 ( .A(a[0]), .Z(n683) );
  NAND U2494 ( .A(n1254), .B(n1255), .Z(c_mult[9]) );
  NANDN U2495 ( .A(n1256), .B(Hi[9]), .Z(n1255) );
  NANDN U2496 ( .A(n1257), .B(Lo[9]), .Z(n1254) );
  NAND U2497 ( .A(n1258), .B(n1259), .Z(c_mult[8]) );
  NANDN U2498 ( .A(n1256), .B(Hi[8]), .Z(n1259) );
  NANDN U2499 ( .A(n1257), .B(Lo[8]), .Z(n1258) );
  NAND U2500 ( .A(n1260), .B(n1261), .Z(c_mult[7]) );
  NANDN U2501 ( .A(n1256), .B(Hi[7]), .Z(n1261) );
  NANDN U2502 ( .A(n1257), .B(Lo[7]), .Z(n1260) );
  NAND U2503 ( .A(n1262), .B(n1263), .Z(c_mult[6]) );
  NANDN U2504 ( .A(n1256), .B(Hi[6]), .Z(n1263) );
  NANDN U2505 ( .A(n1257), .B(Lo[6]), .Z(n1262) );
  NAND U2506 ( .A(n1264), .B(n1265), .Z(c_mult[5]) );
  NANDN U2507 ( .A(n1256), .B(Hi[5]), .Z(n1265) );
  NANDN U2508 ( .A(n1257), .B(Lo[5]), .Z(n1264) );
  NAND U2509 ( .A(n1266), .B(n1267), .Z(c_mult[4]) );
  NANDN U2510 ( .A(n1256), .B(Hi[4]), .Z(n1267) );
  NANDN U2511 ( .A(n1257), .B(Lo[4]), .Z(n1266) );
  NAND U2512 ( .A(n1268), .B(n1269), .Z(c_mult[3]) );
  NANDN U2513 ( .A(n1256), .B(Hi[3]), .Z(n1269) );
  NANDN U2514 ( .A(n1257), .B(Lo[3]), .Z(n1268) );
  NAND U2515 ( .A(n1270), .B(n1271), .Z(c_mult[31]) );
  NANDN U2516 ( .A(n1256), .B(Hi[31]), .Z(n1271) );
  NANDN U2517 ( .A(n1257), .B(Lo[31]), .Z(n1270) );
  NAND U2518 ( .A(n1272), .B(n1273), .Z(c_mult[30]) );
  NANDN U2519 ( .A(n1256), .B(Hi[30]), .Z(n1273) );
  NANDN U2520 ( .A(n1257), .B(Lo[30]), .Z(n1272) );
  NAND U2521 ( .A(n1274), .B(n1275), .Z(c_mult[2]) );
  NANDN U2522 ( .A(n1256), .B(Hi[2]), .Z(n1275) );
  NANDN U2523 ( .A(n1257), .B(Lo[2]), .Z(n1274) );
  NAND U2524 ( .A(n1276), .B(n1277), .Z(c_mult[29]) );
  NANDN U2525 ( .A(n1256), .B(Hi[29]), .Z(n1277) );
  NANDN U2526 ( .A(n1257), .B(Lo[29]), .Z(n1276) );
  NAND U2527 ( .A(n1278), .B(n1279), .Z(c_mult[28]) );
  NANDN U2528 ( .A(n1256), .B(Hi[28]), .Z(n1279) );
  NANDN U2529 ( .A(n1257), .B(Lo[28]), .Z(n1278) );
  NAND U2530 ( .A(n1280), .B(n1281), .Z(c_mult[27]) );
  NANDN U2531 ( .A(n1256), .B(Hi[27]), .Z(n1281) );
  NANDN U2532 ( .A(n1257), .B(Lo[27]), .Z(n1280) );
  NAND U2533 ( .A(n1282), .B(n1283), .Z(c_mult[26]) );
  NANDN U2534 ( .A(n1256), .B(Hi[26]), .Z(n1283) );
  NANDN U2535 ( .A(n1257), .B(Lo[26]), .Z(n1282) );
  NAND U2536 ( .A(n1284), .B(n1285), .Z(c_mult[25]) );
  NANDN U2537 ( .A(n1256), .B(Hi[25]), .Z(n1285) );
  NANDN U2538 ( .A(n1257), .B(Lo[25]), .Z(n1284) );
  NAND U2539 ( .A(n1286), .B(n1287), .Z(c_mult[24]) );
  NANDN U2540 ( .A(n1256), .B(Hi[24]), .Z(n1287) );
  NANDN U2541 ( .A(n1257), .B(Lo[24]), .Z(n1286) );
  NAND U2542 ( .A(n1288), .B(n1289), .Z(c_mult[23]) );
  NANDN U2543 ( .A(n1256), .B(Hi[23]), .Z(n1289) );
  NANDN U2544 ( .A(n1257), .B(Lo[23]), .Z(n1288) );
  NAND U2545 ( .A(n1290), .B(n1291), .Z(c_mult[22]) );
  NANDN U2546 ( .A(n1256), .B(Hi[22]), .Z(n1291) );
  NANDN U2547 ( .A(n1257), .B(Lo[22]), .Z(n1290) );
  NAND U2548 ( .A(n1292), .B(n1293), .Z(c_mult[21]) );
  NANDN U2549 ( .A(n1256), .B(Hi[21]), .Z(n1293) );
  NANDN U2550 ( .A(n1257), .B(Lo[21]), .Z(n1292) );
  NAND U2551 ( .A(n1294), .B(n1295), .Z(c_mult[20]) );
  NANDN U2552 ( .A(n1256), .B(Hi[20]), .Z(n1295) );
  NANDN U2553 ( .A(n1257), .B(Lo[20]), .Z(n1294) );
  NAND U2554 ( .A(n1296), .B(n1297), .Z(c_mult[1]) );
  NANDN U2555 ( .A(n1256), .B(Hi[1]), .Z(n1297) );
  NANDN U2556 ( .A(n1257), .B(Lo[1]), .Z(n1296) );
  NAND U2557 ( .A(n1298), .B(n1299), .Z(c_mult[19]) );
  NANDN U2558 ( .A(n1256), .B(Hi[19]), .Z(n1299) );
  NANDN U2559 ( .A(n1257), .B(Lo[19]), .Z(n1298) );
  NAND U2560 ( .A(n1300), .B(n1301), .Z(c_mult[18]) );
  NANDN U2561 ( .A(n1256), .B(Hi[18]), .Z(n1301) );
  NANDN U2562 ( .A(n1257), .B(Lo[18]), .Z(n1300) );
  NAND U2563 ( .A(n1302), .B(n1303), .Z(c_mult[17]) );
  NANDN U2564 ( .A(n1256), .B(Hi[17]), .Z(n1303) );
  NANDN U2565 ( .A(n1257), .B(Lo[17]), .Z(n1302) );
  NAND U2566 ( .A(n1304), .B(n1305), .Z(c_mult[16]) );
  NANDN U2567 ( .A(n1256), .B(Hi[16]), .Z(n1305) );
  NANDN U2568 ( .A(n1257), .B(Lo[16]), .Z(n1304) );
  NAND U2569 ( .A(n1306), .B(n1307), .Z(c_mult[15]) );
  NANDN U2570 ( .A(n1256), .B(Hi[15]), .Z(n1307) );
  NANDN U2571 ( .A(n1257), .B(Lo[15]), .Z(n1306) );
  NAND U2572 ( .A(n1308), .B(n1309), .Z(c_mult[14]) );
  NANDN U2573 ( .A(n1256), .B(Hi[14]), .Z(n1309) );
  NANDN U2574 ( .A(n1257), .B(Lo[14]), .Z(n1308) );
  NAND U2575 ( .A(n1310), .B(n1311), .Z(c_mult[13]) );
  NANDN U2576 ( .A(n1256), .B(Hi[13]), .Z(n1311) );
  NANDN U2577 ( .A(n1257), .B(Lo[13]), .Z(n1310) );
  NAND U2578 ( .A(n1312), .B(n1313), .Z(c_mult[12]) );
  NANDN U2579 ( .A(n1256), .B(Hi[12]), .Z(n1313) );
  NANDN U2580 ( .A(n1257), .B(Lo[12]), .Z(n1312) );
  NAND U2581 ( .A(n1314), .B(n1315), .Z(c_mult[11]) );
  NANDN U2582 ( .A(n1256), .B(Hi[11]), .Z(n1315) );
  NANDN U2583 ( .A(n1257), .B(Lo[11]), .Z(n1314) );
  NAND U2584 ( .A(n1316), .B(n1317), .Z(c_mult[10]) );
  NANDN U2585 ( .A(n1256), .B(Hi[10]), .Z(n1317) );
  NANDN U2586 ( .A(n1257), .B(Lo[10]), .Z(n1316) );
  NAND U2587 ( .A(n1318), .B(n1319), .Z(c_mult[0]) );
  NANDN U2588 ( .A(n1256), .B(Hi[0]), .Z(n1319) );
  NAND U2589 ( .A(n1320), .B(n1245), .Z(n1256) );
  NANDN U2590 ( .A(n1257), .B(Lo[0]), .Z(n1318) );
  NAND U2591 ( .A(n1321), .B(n1245), .Z(n1257) );
  NOR U2592 ( .A(mult_func[2]), .B(mult_func[3]), .Z(n1245) );
  AND U2593 ( .A(n1252), .B(n1250), .Z(\U3/U1/Z_0 ) );
  IV U2594 ( .A(n1211), .Z(n1250) );
  AND U2595 ( .A(n1322), .B(n1323), .Z(n1211) );
  NAND U2596 ( .A(n1073), .B(n1320), .Z(n1322) );
  ANDN U2597 ( .B(mult_func[1]), .A(mult_func[0]), .Z(n1320) );
  AND U2598 ( .A(n1324), .B(n1323), .Z(n1252) );
  NANDN U2599 ( .A(n1244), .B(n1073), .Z(n1323) );
  NANDN U2600 ( .A(n1325), .B(mult_func[0]), .Z(n1244) );
  NAND U2601 ( .A(n1073), .B(n1321), .Z(n1324) );
  AND U2602 ( .A(mult_func[0]), .B(n1325), .Z(n1321) );
  IV U2603 ( .A(mult_func[1]), .Z(n1325) );
  ANDN U2604 ( .B(mult_func[2]), .A(mult_func[3]), .Z(n1073) );
endmodule

