
module mult_N64_CC16 ( clk, rst, a, b, c );
  input [63:0] a;
  input [3:0] b;
  output [63:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674;
  wire   [63:4] swire;
  wire   [127:64] sreg;

  DFF \sreg_reg[64]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[65]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[66]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[67]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[68]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[69]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[70]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[71]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[72]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[73]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[74]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[75]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[76]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[77]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[78]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[79]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[80]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[81]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[82]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[83]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[84]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[85]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[86]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[87]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[88]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[89]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[90]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[91]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[92]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[93]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[94]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[95]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[96]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[96]) );
  DFF \sreg_reg[97]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[97]) );
  DFF \sreg_reg[98]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[98]) );
  DFF \sreg_reg[99]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[99]) );
  DFF \sreg_reg[100]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[100]) );
  DFF \sreg_reg[101]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[101]) );
  DFF \sreg_reg[102]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[102]) );
  DFF \sreg_reg[103]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[103]) );
  DFF \sreg_reg[104]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[104]) );
  DFF \sreg_reg[105]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[105]) );
  DFF \sreg_reg[106]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[106]) );
  DFF \sreg_reg[107]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[107]) );
  DFF \sreg_reg[108]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[108]) );
  DFF \sreg_reg[109]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[109]) );
  DFF \sreg_reg[110]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[110]) );
  DFF \sreg_reg[111]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[111]) );
  DFF \sreg_reg[112]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[112]) );
  DFF \sreg_reg[113]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[113]) );
  DFF \sreg_reg[114]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[114]) );
  DFF \sreg_reg[115]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[115]) );
  DFF \sreg_reg[116]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[116]) );
  DFF \sreg_reg[117]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[117]) );
  DFF \sreg_reg[118]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[118]) );
  DFF \sreg_reg[119]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[119]) );
  DFF \sreg_reg[120]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[120]) );
  DFF \sreg_reg[121]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[121]) );
  DFF \sreg_reg[122]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[122]) );
  DFF \sreg_reg[123]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[123]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U7 ( .A(n664), .B(n655), .Z(n663) );
  NAND U8 ( .A(n31), .B(n30), .Z(n21) );
  XOR U9 ( .A(n1), .B(n2), .Z(swire[9]) );
  XOR U10 ( .A(n3), .B(n4), .Z(swire[8]) );
  XOR U11 ( .A(n5), .B(n6), .Z(swire[7]) );
  XOR U12 ( .A(n7), .B(n8), .Z(swire[6]) );
  XOR U13 ( .A(n9), .B(n10), .Z(swire[63]) );
  XOR U14 ( .A(n11), .B(n12), .Z(n10) );
  AND U15 ( .A(a[63]), .B(b[0]), .Z(n12) );
  AND U16 ( .A(b[1]), .B(a[62]), .Z(n11) );
  XOR U17 ( .A(n13), .B(n14), .Z(n9) );
  AND U18 ( .A(b[2]), .B(a[61]), .Z(n14) );
  AND U19 ( .A(b[3]), .B(a[60]), .Z(n13) );
  XOR U20 ( .A(n15), .B(n16), .Z(swire[62]) );
  XOR U21 ( .A(n17), .B(n18), .Z(n16) );
  AND U22 ( .A(a[62]), .B(b[0]), .Z(n18) );
  AND U23 ( .A(b[1]), .B(a[61]), .Z(n17) );
  XOR U24 ( .A(n19), .B(n20), .Z(n15) );
  AND U25 ( .A(b[2]), .B(a[60]), .Z(n20) );
  AND U26 ( .A(b[3]), .B(a[59]), .Z(n19) );
  XNOR U27 ( .A(n21), .B(n22), .Z(swire[61]) );
  XOR U28 ( .A(n23), .B(n24), .Z(n22) );
  XNOR U29 ( .A(n25), .B(n21), .Z(n24) );
  AND U30 ( .A(a[61]), .B(b[0]), .Z(n25) );
  XOR U31 ( .A(n26), .B(n27), .Z(n23) );
  XOR U32 ( .A(n28), .B(n29), .Z(n27) );
  AND U33 ( .A(a[59]), .B(b[2]), .Z(n29) );
  AND U34 ( .A(a[58]), .B(b[3]), .Z(n28) );
  AND U35 ( .A(a[60]), .B(b[1]), .Z(n26) );
  XNOR U36 ( .A(n30), .B(n31), .Z(swire[60]) );
  XOR U37 ( .A(n32), .B(n33), .Z(n31) );
  XNOR U38 ( .A(n34), .B(n30), .Z(n33) );
  AND U39 ( .A(b[0]), .B(a[60]), .Z(n34) );
  XOR U40 ( .A(n35), .B(n36), .Z(n32) );
  XOR U41 ( .A(n37), .B(n38), .Z(n36) );
  AND U42 ( .A(b[2]), .B(a[58]), .Z(n38) );
  AND U43 ( .A(a[57]), .B(b[3]), .Z(n37) );
  AND U44 ( .A(b[1]), .B(a[59]), .Z(n35) );
  XNOR U45 ( .A(n39), .B(n40), .Z(n30) );
  NOR U46 ( .A(n41), .B(n42), .Z(n39) );
  XOR U47 ( .A(n43), .B(n44), .Z(swire[5]) );
  XOR U48 ( .A(n42), .B(n41), .Z(swire[59]) );
  XOR U49 ( .A(sreg[123]), .B(n40), .Z(n41) );
  XOR U50 ( .A(n45), .B(n46), .Z(n42) );
  XOR U51 ( .A(n47), .B(n40), .Z(n46) );
  XOR U52 ( .A(n48), .B(n49), .Z(n40) );
  NOR U53 ( .A(n50), .B(n51), .Z(n48) );
  AND U54 ( .A(b[0]), .B(a[59]), .Z(n47) );
  XOR U55 ( .A(n52), .B(n53), .Z(n45) );
  XOR U56 ( .A(n54), .B(n55), .Z(n53) );
  AND U57 ( .A(b[2]), .B(a[57]), .Z(n55) );
  AND U58 ( .A(a[56]), .B(b[3]), .Z(n54) );
  AND U59 ( .A(b[1]), .B(a[58]), .Z(n52) );
  XOR U60 ( .A(n51), .B(n50), .Z(swire[58]) );
  XOR U61 ( .A(sreg[122]), .B(n49), .Z(n50) );
  XOR U62 ( .A(n56), .B(n57), .Z(n51) );
  XOR U63 ( .A(n58), .B(n49), .Z(n57) );
  XOR U64 ( .A(n59), .B(n60), .Z(n49) );
  NOR U65 ( .A(n61), .B(n62), .Z(n59) );
  AND U66 ( .A(b[0]), .B(a[58]), .Z(n58) );
  XOR U67 ( .A(n63), .B(n64), .Z(n56) );
  XOR U68 ( .A(n65), .B(n66), .Z(n64) );
  AND U69 ( .A(b[2]), .B(a[56]), .Z(n66) );
  AND U70 ( .A(a[55]), .B(b[3]), .Z(n65) );
  AND U71 ( .A(b[1]), .B(a[57]), .Z(n63) );
  XOR U72 ( .A(n62), .B(n61), .Z(swire[57]) );
  XOR U73 ( .A(sreg[121]), .B(n60), .Z(n61) );
  XOR U74 ( .A(n67), .B(n68), .Z(n62) );
  XOR U75 ( .A(n69), .B(n60), .Z(n68) );
  XOR U76 ( .A(n70), .B(n71), .Z(n60) );
  NOR U77 ( .A(n72), .B(n73), .Z(n70) );
  AND U78 ( .A(b[0]), .B(a[57]), .Z(n69) );
  XOR U79 ( .A(n74), .B(n75), .Z(n67) );
  XOR U80 ( .A(n76), .B(n77), .Z(n75) );
  AND U81 ( .A(b[2]), .B(a[55]), .Z(n77) );
  AND U82 ( .A(a[54]), .B(b[3]), .Z(n76) );
  AND U83 ( .A(b[1]), .B(a[56]), .Z(n74) );
  XOR U84 ( .A(n73), .B(n72), .Z(swire[56]) );
  XOR U85 ( .A(sreg[120]), .B(n71), .Z(n72) );
  XOR U86 ( .A(n78), .B(n79), .Z(n73) );
  XOR U87 ( .A(n80), .B(n71), .Z(n79) );
  XOR U88 ( .A(n81), .B(n82), .Z(n71) );
  NOR U89 ( .A(n83), .B(n84), .Z(n81) );
  AND U90 ( .A(b[0]), .B(a[56]), .Z(n80) );
  XOR U91 ( .A(n85), .B(n86), .Z(n78) );
  XOR U92 ( .A(n87), .B(n88), .Z(n86) );
  AND U93 ( .A(b[2]), .B(a[54]), .Z(n88) );
  AND U94 ( .A(a[53]), .B(b[3]), .Z(n87) );
  AND U95 ( .A(b[1]), .B(a[55]), .Z(n85) );
  XOR U96 ( .A(n84), .B(n83), .Z(swire[55]) );
  XOR U97 ( .A(sreg[119]), .B(n82), .Z(n83) );
  XOR U98 ( .A(n89), .B(n90), .Z(n84) );
  XOR U99 ( .A(n91), .B(n82), .Z(n90) );
  XOR U100 ( .A(n92), .B(n93), .Z(n82) );
  NOR U101 ( .A(n94), .B(n95), .Z(n92) );
  AND U102 ( .A(b[0]), .B(a[55]), .Z(n91) );
  XOR U103 ( .A(n96), .B(n97), .Z(n89) );
  XOR U104 ( .A(n98), .B(n99), .Z(n97) );
  AND U105 ( .A(b[2]), .B(a[53]), .Z(n99) );
  AND U106 ( .A(a[52]), .B(b[3]), .Z(n98) );
  AND U107 ( .A(b[1]), .B(a[54]), .Z(n96) );
  XOR U108 ( .A(n95), .B(n94), .Z(swire[54]) );
  XOR U109 ( .A(sreg[118]), .B(n93), .Z(n94) );
  XOR U110 ( .A(n100), .B(n101), .Z(n95) );
  XOR U111 ( .A(n102), .B(n93), .Z(n101) );
  XOR U112 ( .A(n103), .B(n104), .Z(n93) );
  NOR U113 ( .A(n105), .B(n106), .Z(n103) );
  AND U114 ( .A(b[0]), .B(a[54]), .Z(n102) );
  XOR U115 ( .A(n107), .B(n108), .Z(n100) );
  XOR U116 ( .A(n109), .B(n110), .Z(n108) );
  AND U117 ( .A(b[2]), .B(a[52]), .Z(n110) );
  AND U118 ( .A(a[51]), .B(b[3]), .Z(n109) );
  AND U119 ( .A(b[1]), .B(a[53]), .Z(n107) );
  XOR U120 ( .A(n106), .B(n105), .Z(swire[53]) );
  XOR U121 ( .A(sreg[117]), .B(n104), .Z(n105) );
  XOR U122 ( .A(n111), .B(n112), .Z(n106) );
  XOR U123 ( .A(n113), .B(n104), .Z(n112) );
  XOR U124 ( .A(n114), .B(n115), .Z(n104) );
  NOR U125 ( .A(n116), .B(n117), .Z(n114) );
  AND U126 ( .A(b[0]), .B(a[53]), .Z(n113) );
  XOR U127 ( .A(n118), .B(n119), .Z(n111) );
  XOR U128 ( .A(n120), .B(n121), .Z(n119) );
  AND U129 ( .A(b[2]), .B(a[51]), .Z(n121) );
  AND U130 ( .A(a[50]), .B(b[3]), .Z(n120) );
  AND U131 ( .A(b[1]), .B(a[52]), .Z(n118) );
  XOR U132 ( .A(n117), .B(n116), .Z(swire[52]) );
  XOR U133 ( .A(sreg[116]), .B(n115), .Z(n116) );
  XOR U134 ( .A(n122), .B(n123), .Z(n117) );
  XOR U135 ( .A(n124), .B(n115), .Z(n123) );
  XOR U136 ( .A(n125), .B(n126), .Z(n115) );
  NOR U137 ( .A(n127), .B(n128), .Z(n125) );
  AND U138 ( .A(b[0]), .B(a[52]), .Z(n124) );
  XOR U139 ( .A(n129), .B(n130), .Z(n122) );
  XOR U140 ( .A(n131), .B(n132), .Z(n130) );
  AND U141 ( .A(b[2]), .B(a[50]), .Z(n132) );
  AND U142 ( .A(a[49]), .B(b[3]), .Z(n131) );
  AND U143 ( .A(b[1]), .B(a[51]), .Z(n129) );
  XOR U144 ( .A(n128), .B(n127), .Z(swire[51]) );
  XOR U145 ( .A(sreg[115]), .B(n126), .Z(n127) );
  XOR U146 ( .A(n133), .B(n134), .Z(n128) );
  XOR U147 ( .A(n135), .B(n126), .Z(n134) );
  XOR U148 ( .A(n136), .B(n137), .Z(n126) );
  NOR U149 ( .A(n138), .B(n139), .Z(n136) );
  AND U150 ( .A(b[0]), .B(a[51]), .Z(n135) );
  XOR U151 ( .A(n140), .B(n141), .Z(n133) );
  XOR U152 ( .A(n142), .B(n143), .Z(n141) );
  AND U153 ( .A(b[2]), .B(a[49]), .Z(n143) );
  AND U154 ( .A(a[48]), .B(b[3]), .Z(n142) );
  AND U155 ( .A(b[1]), .B(a[50]), .Z(n140) );
  XOR U156 ( .A(n139), .B(n138), .Z(swire[50]) );
  XOR U157 ( .A(sreg[114]), .B(n137), .Z(n138) );
  XOR U158 ( .A(n144), .B(n145), .Z(n139) );
  XOR U159 ( .A(n146), .B(n137), .Z(n145) );
  XOR U160 ( .A(n147), .B(n148), .Z(n137) );
  NOR U161 ( .A(n149), .B(n150), .Z(n147) );
  AND U162 ( .A(b[0]), .B(a[50]), .Z(n146) );
  XOR U163 ( .A(n151), .B(n152), .Z(n144) );
  XOR U164 ( .A(n153), .B(n154), .Z(n152) );
  AND U165 ( .A(b[2]), .B(a[48]), .Z(n154) );
  AND U166 ( .A(a[47]), .B(b[3]), .Z(n153) );
  AND U167 ( .A(b[1]), .B(a[49]), .Z(n151) );
  XOR U168 ( .A(n155), .B(n156), .Z(swire[4]) );
  XOR U169 ( .A(n150), .B(n149), .Z(swire[49]) );
  XOR U170 ( .A(sreg[113]), .B(n148), .Z(n149) );
  XOR U171 ( .A(n157), .B(n158), .Z(n150) );
  XOR U172 ( .A(n159), .B(n148), .Z(n158) );
  XOR U173 ( .A(n160), .B(n161), .Z(n148) );
  NOR U174 ( .A(n162), .B(n163), .Z(n160) );
  AND U175 ( .A(b[0]), .B(a[49]), .Z(n159) );
  XOR U176 ( .A(n164), .B(n165), .Z(n157) );
  XOR U177 ( .A(n166), .B(n167), .Z(n165) );
  AND U178 ( .A(b[2]), .B(a[47]), .Z(n167) );
  AND U179 ( .A(a[46]), .B(b[3]), .Z(n166) );
  AND U180 ( .A(b[1]), .B(a[48]), .Z(n164) );
  XOR U181 ( .A(n163), .B(n162), .Z(swire[48]) );
  XOR U182 ( .A(sreg[112]), .B(n161), .Z(n162) );
  XOR U183 ( .A(n168), .B(n169), .Z(n163) );
  XOR U184 ( .A(n170), .B(n161), .Z(n169) );
  XOR U185 ( .A(n171), .B(n172), .Z(n161) );
  NOR U186 ( .A(n173), .B(n174), .Z(n171) );
  AND U187 ( .A(b[0]), .B(a[48]), .Z(n170) );
  XOR U188 ( .A(n175), .B(n176), .Z(n168) );
  XOR U189 ( .A(n177), .B(n178), .Z(n176) );
  AND U190 ( .A(b[2]), .B(a[46]), .Z(n178) );
  AND U191 ( .A(a[45]), .B(b[3]), .Z(n177) );
  AND U192 ( .A(b[1]), .B(a[47]), .Z(n175) );
  XOR U193 ( .A(n174), .B(n173), .Z(swire[47]) );
  XOR U194 ( .A(sreg[111]), .B(n172), .Z(n173) );
  XOR U195 ( .A(n179), .B(n180), .Z(n174) );
  XOR U196 ( .A(n181), .B(n172), .Z(n180) );
  XOR U197 ( .A(n182), .B(n183), .Z(n172) );
  NOR U198 ( .A(n184), .B(n185), .Z(n182) );
  AND U199 ( .A(b[0]), .B(a[47]), .Z(n181) );
  XOR U200 ( .A(n186), .B(n187), .Z(n179) );
  XOR U201 ( .A(n188), .B(n189), .Z(n187) );
  AND U202 ( .A(b[2]), .B(a[45]), .Z(n189) );
  AND U203 ( .A(a[44]), .B(b[3]), .Z(n188) );
  AND U204 ( .A(b[1]), .B(a[46]), .Z(n186) );
  XOR U205 ( .A(n185), .B(n184), .Z(swire[46]) );
  XOR U206 ( .A(sreg[110]), .B(n183), .Z(n184) );
  XOR U207 ( .A(n190), .B(n191), .Z(n185) );
  XOR U208 ( .A(n192), .B(n183), .Z(n191) );
  XOR U209 ( .A(n193), .B(n194), .Z(n183) );
  NOR U210 ( .A(n195), .B(n196), .Z(n193) );
  AND U211 ( .A(b[0]), .B(a[46]), .Z(n192) );
  XOR U212 ( .A(n197), .B(n198), .Z(n190) );
  XOR U213 ( .A(n199), .B(n200), .Z(n198) );
  AND U214 ( .A(b[2]), .B(a[44]), .Z(n200) );
  AND U215 ( .A(a[43]), .B(b[3]), .Z(n199) );
  AND U216 ( .A(b[1]), .B(a[45]), .Z(n197) );
  XOR U217 ( .A(n196), .B(n195), .Z(swire[45]) );
  XOR U218 ( .A(sreg[109]), .B(n194), .Z(n195) );
  XOR U219 ( .A(n201), .B(n202), .Z(n196) );
  XOR U220 ( .A(n203), .B(n194), .Z(n202) );
  XOR U221 ( .A(n204), .B(n205), .Z(n194) );
  NOR U222 ( .A(n206), .B(n207), .Z(n204) );
  AND U223 ( .A(b[0]), .B(a[45]), .Z(n203) );
  XOR U224 ( .A(n208), .B(n209), .Z(n201) );
  XOR U225 ( .A(n210), .B(n211), .Z(n209) );
  AND U226 ( .A(b[2]), .B(a[43]), .Z(n211) );
  AND U227 ( .A(a[42]), .B(b[3]), .Z(n210) );
  AND U228 ( .A(b[1]), .B(a[44]), .Z(n208) );
  XOR U229 ( .A(n207), .B(n206), .Z(swire[44]) );
  XOR U230 ( .A(sreg[108]), .B(n205), .Z(n206) );
  XOR U231 ( .A(n212), .B(n213), .Z(n207) );
  XOR U232 ( .A(n214), .B(n205), .Z(n213) );
  XOR U233 ( .A(n215), .B(n216), .Z(n205) );
  NOR U234 ( .A(n217), .B(n218), .Z(n215) );
  AND U235 ( .A(b[0]), .B(a[44]), .Z(n214) );
  XOR U236 ( .A(n219), .B(n220), .Z(n212) );
  XOR U237 ( .A(n221), .B(n222), .Z(n220) );
  AND U238 ( .A(b[2]), .B(a[42]), .Z(n222) );
  AND U239 ( .A(a[41]), .B(b[3]), .Z(n221) );
  AND U240 ( .A(b[1]), .B(a[43]), .Z(n219) );
  XOR U241 ( .A(n218), .B(n217), .Z(swire[43]) );
  XOR U242 ( .A(sreg[107]), .B(n216), .Z(n217) );
  XOR U243 ( .A(n223), .B(n224), .Z(n218) );
  XOR U244 ( .A(n225), .B(n216), .Z(n224) );
  XOR U245 ( .A(n226), .B(n227), .Z(n216) );
  NOR U246 ( .A(n228), .B(n229), .Z(n226) );
  AND U247 ( .A(b[0]), .B(a[43]), .Z(n225) );
  XOR U248 ( .A(n230), .B(n231), .Z(n223) );
  XOR U249 ( .A(n232), .B(n233), .Z(n231) );
  AND U250 ( .A(b[2]), .B(a[41]), .Z(n233) );
  AND U251 ( .A(a[40]), .B(b[3]), .Z(n232) );
  AND U252 ( .A(b[1]), .B(a[42]), .Z(n230) );
  XOR U253 ( .A(n229), .B(n228), .Z(swire[42]) );
  XOR U254 ( .A(sreg[106]), .B(n227), .Z(n228) );
  XOR U255 ( .A(n234), .B(n235), .Z(n229) );
  XOR U256 ( .A(n236), .B(n227), .Z(n235) );
  XOR U257 ( .A(n237), .B(n238), .Z(n227) );
  NOR U258 ( .A(n239), .B(n240), .Z(n237) );
  AND U259 ( .A(b[0]), .B(a[42]), .Z(n236) );
  XOR U260 ( .A(n241), .B(n242), .Z(n234) );
  XOR U261 ( .A(n243), .B(n244), .Z(n242) );
  AND U262 ( .A(b[2]), .B(a[40]), .Z(n244) );
  AND U263 ( .A(a[39]), .B(b[3]), .Z(n243) );
  AND U264 ( .A(b[1]), .B(a[41]), .Z(n241) );
  XOR U265 ( .A(n240), .B(n239), .Z(swire[41]) );
  XOR U266 ( .A(sreg[105]), .B(n238), .Z(n239) );
  XOR U267 ( .A(n245), .B(n246), .Z(n240) );
  XOR U268 ( .A(n247), .B(n238), .Z(n246) );
  XOR U269 ( .A(n248), .B(n249), .Z(n238) );
  NOR U270 ( .A(n250), .B(n251), .Z(n248) );
  AND U271 ( .A(b[0]), .B(a[41]), .Z(n247) );
  XOR U272 ( .A(n252), .B(n253), .Z(n245) );
  XOR U273 ( .A(n254), .B(n255), .Z(n253) );
  AND U274 ( .A(b[2]), .B(a[39]), .Z(n255) );
  AND U275 ( .A(a[38]), .B(b[3]), .Z(n254) );
  AND U276 ( .A(b[1]), .B(a[40]), .Z(n252) );
  XOR U277 ( .A(n251), .B(n250), .Z(swire[40]) );
  XOR U278 ( .A(sreg[104]), .B(n249), .Z(n250) );
  XOR U279 ( .A(n256), .B(n257), .Z(n251) );
  XOR U280 ( .A(n258), .B(n249), .Z(n257) );
  XOR U281 ( .A(n259), .B(n260), .Z(n249) );
  NOR U282 ( .A(n261), .B(n262), .Z(n259) );
  AND U283 ( .A(b[0]), .B(a[40]), .Z(n258) );
  XOR U284 ( .A(n263), .B(n264), .Z(n256) );
  XOR U285 ( .A(n265), .B(n266), .Z(n264) );
  AND U286 ( .A(b[2]), .B(a[38]), .Z(n266) );
  AND U287 ( .A(a[37]), .B(b[3]), .Z(n265) );
  AND U288 ( .A(b[1]), .B(a[39]), .Z(n263) );
  XOR U289 ( .A(n262), .B(n261), .Z(swire[39]) );
  XOR U290 ( .A(sreg[103]), .B(n260), .Z(n261) );
  XOR U291 ( .A(n267), .B(n268), .Z(n262) );
  XOR U292 ( .A(n269), .B(n260), .Z(n268) );
  XOR U293 ( .A(n270), .B(n271), .Z(n260) );
  NOR U294 ( .A(n272), .B(n273), .Z(n270) );
  AND U295 ( .A(b[0]), .B(a[39]), .Z(n269) );
  XOR U296 ( .A(n274), .B(n275), .Z(n267) );
  XOR U297 ( .A(n276), .B(n277), .Z(n275) );
  AND U298 ( .A(b[2]), .B(a[37]), .Z(n277) );
  AND U299 ( .A(a[36]), .B(b[3]), .Z(n276) );
  AND U300 ( .A(b[1]), .B(a[38]), .Z(n274) );
  XOR U301 ( .A(n273), .B(n272), .Z(swire[38]) );
  XOR U302 ( .A(sreg[102]), .B(n271), .Z(n272) );
  XOR U303 ( .A(n278), .B(n279), .Z(n273) );
  XOR U304 ( .A(n280), .B(n271), .Z(n279) );
  XOR U305 ( .A(n281), .B(n282), .Z(n271) );
  NOR U306 ( .A(n283), .B(n284), .Z(n281) );
  AND U307 ( .A(b[0]), .B(a[38]), .Z(n280) );
  XOR U308 ( .A(n285), .B(n286), .Z(n278) );
  XOR U309 ( .A(n287), .B(n288), .Z(n286) );
  AND U310 ( .A(b[2]), .B(a[36]), .Z(n288) );
  AND U311 ( .A(a[35]), .B(b[3]), .Z(n287) );
  AND U312 ( .A(b[1]), .B(a[37]), .Z(n285) );
  XOR U313 ( .A(n284), .B(n283), .Z(swire[37]) );
  XOR U314 ( .A(sreg[101]), .B(n282), .Z(n283) );
  XOR U315 ( .A(n289), .B(n290), .Z(n284) );
  XOR U316 ( .A(n291), .B(n282), .Z(n290) );
  XOR U317 ( .A(n292), .B(n293), .Z(n282) );
  NOR U318 ( .A(n294), .B(n295), .Z(n292) );
  AND U319 ( .A(b[0]), .B(a[37]), .Z(n291) );
  XOR U320 ( .A(n296), .B(n297), .Z(n289) );
  XOR U321 ( .A(n298), .B(n299), .Z(n297) );
  AND U322 ( .A(b[2]), .B(a[35]), .Z(n299) );
  AND U323 ( .A(a[34]), .B(b[3]), .Z(n298) );
  AND U324 ( .A(b[1]), .B(a[36]), .Z(n296) );
  XOR U325 ( .A(n295), .B(n294), .Z(swire[36]) );
  XOR U326 ( .A(sreg[100]), .B(n293), .Z(n294) );
  XOR U327 ( .A(n300), .B(n301), .Z(n295) );
  XOR U328 ( .A(n302), .B(n293), .Z(n301) );
  XOR U329 ( .A(n303), .B(n304), .Z(n293) );
  NOR U330 ( .A(n305), .B(n306), .Z(n303) );
  AND U331 ( .A(b[0]), .B(a[36]), .Z(n302) );
  XOR U332 ( .A(n307), .B(n308), .Z(n300) );
  XOR U333 ( .A(n309), .B(n310), .Z(n308) );
  AND U334 ( .A(b[2]), .B(a[34]), .Z(n310) );
  AND U335 ( .A(a[33]), .B(b[3]), .Z(n309) );
  AND U336 ( .A(b[1]), .B(a[35]), .Z(n307) );
  XOR U337 ( .A(n306), .B(n305), .Z(swire[35]) );
  XOR U338 ( .A(sreg[99]), .B(n304), .Z(n305) );
  XOR U339 ( .A(n311), .B(n312), .Z(n306) );
  XOR U340 ( .A(n313), .B(n304), .Z(n312) );
  XOR U341 ( .A(n314), .B(n315), .Z(n304) );
  NOR U342 ( .A(n316), .B(n317), .Z(n314) );
  AND U343 ( .A(b[0]), .B(a[35]), .Z(n313) );
  XOR U344 ( .A(n318), .B(n319), .Z(n311) );
  XOR U345 ( .A(n320), .B(n321), .Z(n319) );
  AND U346 ( .A(b[2]), .B(a[33]), .Z(n321) );
  AND U347 ( .A(a[32]), .B(b[3]), .Z(n320) );
  AND U348 ( .A(b[1]), .B(a[34]), .Z(n318) );
  XOR U349 ( .A(n317), .B(n316), .Z(swire[34]) );
  XOR U350 ( .A(sreg[98]), .B(n315), .Z(n316) );
  XOR U351 ( .A(n322), .B(n323), .Z(n317) );
  XOR U352 ( .A(n324), .B(n315), .Z(n323) );
  XOR U353 ( .A(n325), .B(n326), .Z(n315) );
  NOR U354 ( .A(n327), .B(n328), .Z(n325) );
  AND U355 ( .A(b[0]), .B(a[34]), .Z(n324) );
  XOR U356 ( .A(n329), .B(n330), .Z(n322) );
  XOR U357 ( .A(n331), .B(n332), .Z(n330) );
  AND U358 ( .A(b[2]), .B(a[32]), .Z(n332) );
  AND U359 ( .A(a[31]), .B(b[3]), .Z(n331) );
  AND U360 ( .A(b[1]), .B(a[33]), .Z(n329) );
  XOR U361 ( .A(n328), .B(n327), .Z(swire[33]) );
  XOR U362 ( .A(sreg[97]), .B(n326), .Z(n327) );
  XOR U363 ( .A(n333), .B(n334), .Z(n328) );
  XOR U364 ( .A(n335), .B(n326), .Z(n334) );
  XOR U365 ( .A(n336), .B(n337), .Z(n326) );
  NOR U366 ( .A(n338), .B(n339), .Z(n336) );
  AND U367 ( .A(b[0]), .B(a[33]), .Z(n335) );
  XOR U368 ( .A(n340), .B(n341), .Z(n333) );
  XOR U369 ( .A(n342), .B(n343), .Z(n341) );
  AND U370 ( .A(b[2]), .B(a[31]), .Z(n343) );
  AND U371 ( .A(a[30]), .B(b[3]), .Z(n342) );
  AND U372 ( .A(b[1]), .B(a[32]), .Z(n340) );
  XOR U373 ( .A(n339), .B(n338), .Z(swire[32]) );
  XOR U374 ( .A(sreg[96]), .B(n337), .Z(n338) );
  XOR U375 ( .A(n344), .B(n345), .Z(n339) );
  XOR U376 ( .A(n346), .B(n337), .Z(n345) );
  XOR U377 ( .A(n347), .B(n348), .Z(n337) );
  NOR U378 ( .A(n349), .B(n350), .Z(n347) );
  AND U379 ( .A(b[0]), .B(a[32]), .Z(n346) );
  XOR U380 ( .A(n351), .B(n352), .Z(n344) );
  XOR U381 ( .A(n353), .B(n354), .Z(n352) );
  AND U382 ( .A(b[2]), .B(a[30]), .Z(n354) );
  AND U383 ( .A(a[29]), .B(b[3]), .Z(n353) );
  AND U384 ( .A(b[1]), .B(a[31]), .Z(n351) );
  XOR U385 ( .A(n350), .B(n349), .Z(swire[31]) );
  XOR U386 ( .A(sreg[95]), .B(n348), .Z(n349) );
  XOR U387 ( .A(n355), .B(n356), .Z(n350) );
  XOR U388 ( .A(n357), .B(n348), .Z(n356) );
  XOR U389 ( .A(n358), .B(n359), .Z(n348) );
  NOR U390 ( .A(n360), .B(n361), .Z(n358) );
  AND U391 ( .A(b[0]), .B(a[31]), .Z(n357) );
  XOR U392 ( .A(n362), .B(n363), .Z(n355) );
  XOR U393 ( .A(n364), .B(n365), .Z(n363) );
  AND U394 ( .A(b[2]), .B(a[29]), .Z(n365) );
  AND U395 ( .A(a[28]), .B(b[3]), .Z(n364) );
  AND U396 ( .A(b[1]), .B(a[30]), .Z(n362) );
  XOR U397 ( .A(n361), .B(n360), .Z(swire[30]) );
  XOR U398 ( .A(sreg[94]), .B(n359), .Z(n360) );
  XOR U399 ( .A(n366), .B(n367), .Z(n361) );
  XOR U400 ( .A(n368), .B(n359), .Z(n367) );
  XOR U401 ( .A(n369), .B(n370), .Z(n359) );
  NOR U402 ( .A(n371), .B(n372), .Z(n369) );
  AND U403 ( .A(b[0]), .B(a[30]), .Z(n368) );
  XOR U404 ( .A(n373), .B(n374), .Z(n366) );
  XOR U405 ( .A(n375), .B(n376), .Z(n374) );
  AND U406 ( .A(b[2]), .B(a[28]), .Z(n376) );
  AND U407 ( .A(a[27]), .B(b[3]), .Z(n375) );
  AND U408 ( .A(b[1]), .B(a[29]), .Z(n373) );
  XOR U409 ( .A(n372), .B(n371), .Z(swire[29]) );
  XOR U410 ( .A(sreg[93]), .B(n370), .Z(n371) );
  XOR U411 ( .A(n377), .B(n378), .Z(n372) );
  XOR U412 ( .A(n379), .B(n370), .Z(n378) );
  XOR U413 ( .A(n380), .B(n381), .Z(n370) );
  NOR U414 ( .A(n382), .B(n383), .Z(n380) );
  AND U415 ( .A(b[0]), .B(a[29]), .Z(n379) );
  XOR U416 ( .A(n384), .B(n385), .Z(n377) );
  XOR U417 ( .A(n386), .B(n387), .Z(n385) );
  AND U418 ( .A(b[2]), .B(a[27]), .Z(n387) );
  AND U419 ( .A(a[26]), .B(b[3]), .Z(n386) );
  AND U420 ( .A(b[1]), .B(a[28]), .Z(n384) );
  XOR U421 ( .A(n383), .B(n382), .Z(swire[28]) );
  XOR U422 ( .A(sreg[92]), .B(n381), .Z(n382) );
  XOR U423 ( .A(n388), .B(n389), .Z(n383) );
  XOR U424 ( .A(n390), .B(n381), .Z(n389) );
  XOR U425 ( .A(n391), .B(n392), .Z(n381) );
  NOR U426 ( .A(n393), .B(n394), .Z(n391) );
  AND U427 ( .A(b[0]), .B(a[28]), .Z(n390) );
  XOR U428 ( .A(n395), .B(n396), .Z(n388) );
  XOR U429 ( .A(n397), .B(n398), .Z(n396) );
  AND U430 ( .A(b[2]), .B(a[26]), .Z(n398) );
  AND U431 ( .A(a[25]), .B(b[3]), .Z(n397) );
  AND U432 ( .A(b[1]), .B(a[27]), .Z(n395) );
  XOR U433 ( .A(n394), .B(n393), .Z(swire[27]) );
  XOR U434 ( .A(sreg[91]), .B(n392), .Z(n393) );
  XOR U435 ( .A(n399), .B(n400), .Z(n394) );
  XOR U436 ( .A(n401), .B(n392), .Z(n400) );
  XOR U437 ( .A(n402), .B(n403), .Z(n392) );
  NOR U438 ( .A(n404), .B(n405), .Z(n402) );
  AND U439 ( .A(b[0]), .B(a[27]), .Z(n401) );
  XOR U440 ( .A(n406), .B(n407), .Z(n399) );
  XOR U441 ( .A(n408), .B(n409), .Z(n407) );
  AND U442 ( .A(b[2]), .B(a[25]), .Z(n409) );
  AND U443 ( .A(a[24]), .B(b[3]), .Z(n408) );
  AND U444 ( .A(b[1]), .B(a[26]), .Z(n406) );
  XOR U445 ( .A(n405), .B(n404), .Z(swire[26]) );
  XOR U446 ( .A(sreg[90]), .B(n403), .Z(n404) );
  XOR U447 ( .A(n410), .B(n411), .Z(n405) );
  XOR U448 ( .A(n412), .B(n403), .Z(n411) );
  XOR U449 ( .A(n413), .B(n414), .Z(n403) );
  NOR U450 ( .A(n415), .B(n416), .Z(n413) );
  AND U451 ( .A(b[0]), .B(a[26]), .Z(n412) );
  XOR U452 ( .A(n417), .B(n418), .Z(n410) );
  XOR U453 ( .A(n419), .B(n420), .Z(n418) );
  AND U454 ( .A(b[2]), .B(a[24]), .Z(n420) );
  AND U455 ( .A(a[23]), .B(b[3]), .Z(n419) );
  AND U456 ( .A(b[1]), .B(a[25]), .Z(n417) );
  XOR U457 ( .A(n416), .B(n415), .Z(swire[25]) );
  XOR U458 ( .A(sreg[89]), .B(n414), .Z(n415) );
  XOR U459 ( .A(n421), .B(n422), .Z(n416) );
  XOR U460 ( .A(n423), .B(n414), .Z(n422) );
  XOR U461 ( .A(n424), .B(n425), .Z(n414) );
  NOR U462 ( .A(n426), .B(n427), .Z(n424) );
  AND U463 ( .A(b[0]), .B(a[25]), .Z(n423) );
  XOR U464 ( .A(n428), .B(n429), .Z(n421) );
  XOR U465 ( .A(n430), .B(n431), .Z(n429) );
  AND U466 ( .A(b[2]), .B(a[23]), .Z(n431) );
  AND U467 ( .A(a[22]), .B(b[3]), .Z(n430) );
  AND U468 ( .A(b[1]), .B(a[24]), .Z(n428) );
  XOR U469 ( .A(n427), .B(n426), .Z(swire[24]) );
  XOR U470 ( .A(sreg[88]), .B(n425), .Z(n426) );
  XOR U471 ( .A(n432), .B(n433), .Z(n427) );
  XOR U472 ( .A(n434), .B(n425), .Z(n433) );
  XOR U473 ( .A(n435), .B(n436), .Z(n425) );
  NOR U474 ( .A(n437), .B(n438), .Z(n435) );
  AND U475 ( .A(b[0]), .B(a[24]), .Z(n434) );
  XOR U476 ( .A(n439), .B(n440), .Z(n432) );
  XOR U477 ( .A(n441), .B(n442), .Z(n440) );
  AND U478 ( .A(b[2]), .B(a[22]), .Z(n442) );
  AND U479 ( .A(a[21]), .B(b[3]), .Z(n441) );
  AND U480 ( .A(b[1]), .B(a[23]), .Z(n439) );
  XOR U481 ( .A(n438), .B(n437), .Z(swire[23]) );
  XOR U482 ( .A(sreg[87]), .B(n436), .Z(n437) );
  XOR U483 ( .A(n443), .B(n444), .Z(n438) );
  XOR U484 ( .A(n445), .B(n436), .Z(n444) );
  XOR U485 ( .A(n446), .B(n447), .Z(n436) );
  NOR U486 ( .A(n448), .B(n449), .Z(n446) );
  AND U487 ( .A(b[0]), .B(a[23]), .Z(n445) );
  XOR U488 ( .A(n450), .B(n451), .Z(n443) );
  XOR U489 ( .A(n452), .B(n453), .Z(n451) );
  AND U490 ( .A(b[2]), .B(a[21]), .Z(n453) );
  AND U491 ( .A(a[20]), .B(b[3]), .Z(n452) );
  AND U492 ( .A(b[1]), .B(a[22]), .Z(n450) );
  XOR U493 ( .A(n449), .B(n448), .Z(swire[22]) );
  XOR U494 ( .A(sreg[86]), .B(n447), .Z(n448) );
  XOR U495 ( .A(n454), .B(n455), .Z(n449) );
  XOR U496 ( .A(n456), .B(n447), .Z(n455) );
  XOR U497 ( .A(n457), .B(n458), .Z(n447) );
  NOR U498 ( .A(n459), .B(n460), .Z(n457) );
  AND U499 ( .A(b[0]), .B(a[22]), .Z(n456) );
  XOR U500 ( .A(n461), .B(n462), .Z(n454) );
  XOR U501 ( .A(n463), .B(n464), .Z(n462) );
  AND U502 ( .A(b[2]), .B(a[20]), .Z(n464) );
  AND U503 ( .A(a[19]), .B(b[3]), .Z(n463) );
  AND U504 ( .A(b[1]), .B(a[21]), .Z(n461) );
  XOR U505 ( .A(n460), .B(n459), .Z(swire[21]) );
  XOR U506 ( .A(sreg[85]), .B(n458), .Z(n459) );
  XOR U507 ( .A(n465), .B(n466), .Z(n460) );
  XOR U508 ( .A(n467), .B(n458), .Z(n466) );
  XOR U509 ( .A(n468), .B(n469), .Z(n458) );
  NOR U510 ( .A(n470), .B(n471), .Z(n468) );
  AND U511 ( .A(b[0]), .B(a[21]), .Z(n467) );
  XOR U512 ( .A(n472), .B(n473), .Z(n465) );
  XOR U513 ( .A(n474), .B(n475), .Z(n473) );
  AND U514 ( .A(b[2]), .B(a[19]), .Z(n475) );
  AND U515 ( .A(a[18]), .B(b[3]), .Z(n474) );
  AND U516 ( .A(b[1]), .B(a[20]), .Z(n472) );
  XOR U517 ( .A(n471), .B(n470), .Z(swire[20]) );
  XOR U518 ( .A(sreg[84]), .B(n469), .Z(n470) );
  XOR U519 ( .A(n476), .B(n477), .Z(n471) );
  XOR U520 ( .A(n478), .B(n469), .Z(n477) );
  XOR U521 ( .A(n479), .B(n480), .Z(n469) );
  NOR U522 ( .A(n481), .B(n482), .Z(n479) );
  AND U523 ( .A(b[0]), .B(a[20]), .Z(n478) );
  XOR U524 ( .A(n483), .B(n484), .Z(n476) );
  XOR U525 ( .A(n485), .B(n486), .Z(n484) );
  AND U526 ( .A(b[2]), .B(a[18]), .Z(n486) );
  AND U527 ( .A(a[17]), .B(b[3]), .Z(n485) );
  AND U528 ( .A(b[1]), .B(a[19]), .Z(n483) );
  XOR U529 ( .A(n482), .B(n481), .Z(swire[19]) );
  XOR U530 ( .A(sreg[83]), .B(n480), .Z(n481) );
  XOR U531 ( .A(n487), .B(n488), .Z(n482) );
  XOR U532 ( .A(n489), .B(n480), .Z(n488) );
  XOR U533 ( .A(n490), .B(n491), .Z(n480) );
  NOR U534 ( .A(n492), .B(n493), .Z(n490) );
  AND U535 ( .A(b[0]), .B(a[19]), .Z(n489) );
  XOR U536 ( .A(n494), .B(n495), .Z(n487) );
  XOR U537 ( .A(n496), .B(n497), .Z(n495) );
  AND U538 ( .A(b[2]), .B(a[17]), .Z(n497) );
  AND U539 ( .A(a[16]), .B(b[3]), .Z(n496) );
  AND U540 ( .A(b[1]), .B(a[18]), .Z(n494) );
  XOR U541 ( .A(n493), .B(n492), .Z(swire[18]) );
  XOR U542 ( .A(sreg[82]), .B(n491), .Z(n492) );
  XOR U543 ( .A(n498), .B(n499), .Z(n493) );
  XOR U544 ( .A(n500), .B(n491), .Z(n499) );
  XOR U545 ( .A(n501), .B(n502), .Z(n491) );
  NOR U546 ( .A(n503), .B(n504), .Z(n501) );
  AND U547 ( .A(b[0]), .B(a[18]), .Z(n500) );
  XOR U548 ( .A(n505), .B(n506), .Z(n498) );
  XOR U549 ( .A(n507), .B(n508), .Z(n506) );
  AND U550 ( .A(b[2]), .B(a[16]), .Z(n508) );
  AND U551 ( .A(a[15]), .B(b[3]), .Z(n507) );
  AND U552 ( .A(b[1]), .B(a[17]), .Z(n505) );
  XOR U553 ( .A(n504), .B(n503), .Z(swire[17]) );
  XOR U554 ( .A(sreg[81]), .B(n502), .Z(n503) );
  XOR U555 ( .A(n509), .B(n510), .Z(n504) );
  XOR U556 ( .A(n511), .B(n502), .Z(n510) );
  XOR U557 ( .A(n512), .B(n513), .Z(n502) );
  NOR U558 ( .A(n514), .B(n515), .Z(n512) );
  AND U559 ( .A(b[0]), .B(a[17]), .Z(n511) );
  XOR U560 ( .A(n516), .B(n517), .Z(n509) );
  XOR U561 ( .A(n518), .B(n519), .Z(n517) );
  AND U562 ( .A(b[2]), .B(a[15]), .Z(n519) );
  AND U563 ( .A(a[14]), .B(b[3]), .Z(n518) );
  AND U564 ( .A(b[1]), .B(a[16]), .Z(n516) );
  XOR U565 ( .A(n515), .B(n514), .Z(swire[16]) );
  XOR U566 ( .A(sreg[80]), .B(n513), .Z(n514) );
  XOR U567 ( .A(n520), .B(n521), .Z(n515) );
  XOR U568 ( .A(n522), .B(n513), .Z(n521) );
  XOR U569 ( .A(n523), .B(n524), .Z(n513) );
  NOR U570 ( .A(n525), .B(n526), .Z(n523) );
  AND U571 ( .A(b[0]), .B(a[16]), .Z(n522) );
  XOR U572 ( .A(n527), .B(n528), .Z(n520) );
  XOR U573 ( .A(n529), .B(n530), .Z(n528) );
  AND U574 ( .A(b[2]), .B(a[14]), .Z(n530) );
  AND U575 ( .A(a[13]), .B(b[3]), .Z(n529) );
  AND U576 ( .A(b[1]), .B(a[15]), .Z(n527) );
  XOR U577 ( .A(n526), .B(n525), .Z(swire[15]) );
  XOR U578 ( .A(sreg[79]), .B(n524), .Z(n525) );
  XOR U579 ( .A(n531), .B(n532), .Z(n526) );
  XOR U580 ( .A(n533), .B(n524), .Z(n532) );
  XOR U581 ( .A(n534), .B(n535), .Z(n524) );
  NOR U582 ( .A(n536), .B(n537), .Z(n534) );
  AND U583 ( .A(b[0]), .B(a[15]), .Z(n533) );
  XOR U584 ( .A(n538), .B(n539), .Z(n531) );
  XOR U585 ( .A(n540), .B(n541), .Z(n539) );
  AND U586 ( .A(b[2]), .B(a[13]), .Z(n541) );
  AND U587 ( .A(a[12]), .B(b[3]), .Z(n540) );
  AND U588 ( .A(b[1]), .B(a[14]), .Z(n538) );
  XOR U589 ( .A(n537), .B(n536), .Z(swire[14]) );
  XOR U590 ( .A(sreg[78]), .B(n535), .Z(n536) );
  XOR U591 ( .A(n542), .B(n543), .Z(n537) );
  XOR U592 ( .A(n544), .B(n535), .Z(n543) );
  XOR U593 ( .A(n545), .B(n546), .Z(n535) );
  NOR U594 ( .A(n547), .B(n548), .Z(n545) );
  AND U595 ( .A(b[0]), .B(a[14]), .Z(n544) );
  XOR U596 ( .A(n549), .B(n550), .Z(n542) );
  XOR U597 ( .A(n551), .B(n552), .Z(n550) );
  AND U598 ( .A(b[2]), .B(a[12]), .Z(n552) );
  AND U599 ( .A(a[11]), .B(b[3]), .Z(n551) );
  AND U600 ( .A(b[1]), .B(a[13]), .Z(n549) );
  XOR U601 ( .A(n548), .B(n547), .Z(swire[13]) );
  XOR U602 ( .A(sreg[77]), .B(n546), .Z(n547) );
  XOR U603 ( .A(n553), .B(n554), .Z(n548) );
  XOR U604 ( .A(n555), .B(n546), .Z(n554) );
  XOR U605 ( .A(n556), .B(n557), .Z(n546) );
  NOR U606 ( .A(n558), .B(n559), .Z(n556) );
  AND U607 ( .A(b[0]), .B(a[13]), .Z(n555) );
  XOR U608 ( .A(n560), .B(n561), .Z(n553) );
  XOR U609 ( .A(n562), .B(n563), .Z(n561) );
  AND U610 ( .A(b[2]), .B(a[11]), .Z(n563) );
  AND U611 ( .A(a[10]), .B(b[3]), .Z(n562) );
  AND U612 ( .A(b[1]), .B(a[12]), .Z(n560) );
  XOR U613 ( .A(n559), .B(n558), .Z(swire[12]) );
  XOR U614 ( .A(sreg[76]), .B(n557), .Z(n558) );
  XOR U615 ( .A(n564), .B(n565), .Z(n559) );
  XOR U616 ( .A(n566), .B(n557), .Z(n565) );
  XOR U617 ( .A(n567), .B(n568), .Z(n557) );
  NOR U618 ( .A(n569), .B(n570), .Z(n567) );
  AND U619 ( .A(b[0]), .B(a[12]), .Z(n566) );
  XOR U620 ( .A(n571), .B(n572), .Z(n564) );
  XOR U621 ( .A(n573), .B(n574), .Z(n572) );
  AND U622 ( .A(b[2]), .B(a[10]), .Z(n574) );
  AND U623 ( .A(a[9]), .B(b[3]), .Z(n573) );
  AND U624 ( .A(b[1]), .B(a[11]), .Z(n571) );
  XOR U625 ( .A(n570), .B(n569), .Z(swire[11]) );
  XOR U626 ( .A(sreg[75]), .B(n568), .Z(n569) );
  XOR U627 ( .A(n575), .B(n576), .Z(n570) );
  XOR U628 ( .A(n577), .B(n568), .Z(n576) );
  XOR U629 ( .A(n578), .B(n579), .Z(n568) );
  NOR U630 ( .A(n580), .B(n581), .Z(n578) );
  AND U631 ( .A(b[0]), .B(a[11]), .Z(n577) );
  XOR U632 ( .A(n582), .B(n583), .Z(n575) );
  XOR U633 ( .A(n584), .B(n585), .Z(n583) );
  AND U634 ( .A(b[2]), .B(a[9]), .Z(n585) );
  AND U635 ( .A(a[8]), .B(b[3]), .Z(n584) );
  AND U636 ( .A(b[1]), .B(a[10]), .Z(n582) );
  XOR U637 ( .A(n581), .B(n580), .Z(swire[10]) );
  XOR U638 ( .A(sreg[74]), .B(n579), .Z(n580) );
  XOR U639 ( .A(n586), .B(n587), .Z(n581) );
  XOR U640 ( .A(n588), .B(n579), .Z(n587) );
  XOR U641 ( .A(n589), .B(n590), .Z(n579) );
  NOR U642 ( .A(n2), .B(n1), .Z(n589) );
  XOR U643 ( .A(sreg[73]), .B(n590), .Z(n1) );
  XOR U644 ( .A(n591), .B(n592), .Z(n2) );
  XOR U645 ( .A(n593), .B(n590), .Z(n592) );
  XOR U646 ( .A(n594), .B(n595), .Z(n590) );
  NOR U647 ( .A(n4), .B(n3), .Z(n594) );
  XOR U648 ( .A(n596), .B(n597), .Z(n3) );
  XOR U649 ( .A(n598), .B(n595), .Z(n597) );
  AND U650 ( .A(b[0]), .B(a[8]), .Z(n598) );
  XOR U651 ( .A(n599), .B(n600), .Z(n596) );
  XOR U652 ( .A(n601), .B(n602), .Z(n600) );
  AND U653 ( .A(a[5]), .B(b[3]), .Z(n602) );
  AND U654 ( .A(a[7]), .B(b[1]), .Z(n601) );
  AND U655 ( .A(b[2]), .B(a[6]), .Z(n599) );
  XOR U656 ( .A(sreg[72]), .B(n595), .Z(n4) );
  XOR U657 ( .A(n603), .B(n604), .Z(n595) );
  NOR U658 ( .A(n6), .B(n5), .Z(n603) );
  XOR U659 ( .A(n605), .B(n606), .Z(n5) );
  XOR U660 ( .A(n607), .B(n604), .Z(n606) );
  AND U661 ( .A(a[7]), .B(b[0]), .Z(n607) );
  XOR U662 ( .A(n608), .B(n609), .Z(n605) );
  XOR U663 ( .A(n610), .B(n611), .Z(n609) );
  AND U664 ( .A(a[5]), .B(b[2]), .Z(n611) );
  AND U665 ( .A(a[4]), .B(b[3]), .Z(n610) );
  AND U666 ( .A(b[1]), .B(a[6]), .Z(n608) );
  XOR U667 ( .A(sreg[71]), .B(n604), .Z(n6) );
  XOR U668 ( .A(n612), .B(n613), .Z(n604) );
  NOR U669 ( .A(n8), .B(n7), .Z(n612) );
  XOR U670 ( .A(n614), .B(n615), .Z(n7) );
  XOR U671 ( .A(n616), .B(n613), .Z(n615) );
  AND U672 ( .A(b[0]), .B(a[6]), .Z(n616) );
  XOR U673 ( .A(n617), .B(n618), .Z(n614) );
  XOR U674 ( .A(n619), .B(n620), .Z(n618) );
  AND U675 ( .A(a[3]), .B(b[3]), .Z(n620) );
  AND U676 ( .A(b[2]), .B(a[4]), .Z(n619) );
  AND U677 ( .A(a[5]), .B(b[1]), .Z(n617) );
  XOR U678 ( .A(sreg[70]), .B(n613), .Z(n8) );
  XOR U679 ( .A(n621), .B(n622), .Z(n613) );
  NOR U680 ( .A(n44), .B(n43), .Z(n621) );
  XOR U681 ( .A(n623), .B(n624), .Z(n43) );
  XOR U682 ( .A(n625), .B(n622), .Z(n624) );
  AND U683 ( .A(b[0]), .B(a[5]), .Z(n625) );
  XOR U684 ( .A(n626), .B(n627), .Z(n623) );
  XOR U685 ( .A(n628), .B(n629), .Z(n627) );
  AND U686 ( .A(a[2]), .B(b[3]), .Z(n629) );
  AND U687 ( .A(a[4]), .B(b[1]), .Z(n628) );
  AND U688 ( .A(b[2]), .B(a[3]), .Z(n626) );
  XOR U689 ( .A(sreg[69]), .B(n622), .Z(n44) );
  XOR U690 ( .A(n630), .B(n631), .Z(n622) );
  NOR U691 ( .A(n156), .B(n155), .Z(n630) );
  XOR U692 ( .A(n632), .B(n633), .Z(n155) );
  XOR U693 ( .A(n634), .B(n631), .Z(n633) );
  AND U694 ( .A(b[0]), .B(a[4]), .Z(n634) );
  XOR U695 ( .A(n635), .B(n636), .Z(n632) );
  XOR U696 ( .A(n637), .B(n638), .Z(n636) );
  AND U697 ( .A(b[2]), .B(a[2]), .Z(n638) );
  AND U698 ( .A(a[1]), .B(b[3]), .Z(n637) );
  AND U699 ( .A(a[3]), .B(b[1]), .Z(n635) );
  XOR U700 ( .A(sreg[68]), .B(n631), .Z(n156) );
  XOR U701 ( .A(n639), .B(n640), .Z(n631) );
  NOR U702 ( .A(n641), .B(n642), .Z(n639) );
  AND U703 ( .A(b[0]), .B(a[9]), .Z(n593) );
  XOR U704 ( .A(n643), .B(n644), .Z(n591) );
  XOR U705 ( .A(n645), .B(n646), .Z(n644) );
  AND U706 ( .A(a[6]), .B(b[3]), .Z(n646) );
  AND U707 ( .A(a[7]), .B(b[2]), .Z(n645) );
  AND U708 ( .A(b[1]), .B(a[8]), .Z(n643) );
  AND U709 ( .A(b[0]), .B(a[10]), .Z(n588) );
  XOR U710 ( .A(n647), .B(n648), .Z(n586) );
  XOR U711 ( .A(n649), .B(n650), .Z(n648) );
  AND U712 ( .A(b[2]), .B(a[8]), .Z(n650) );
  AND U713 ( .A(a[7]), .B(b[3]), .Z(n649) );
  AND U714 ( .A(b[1]), .B(a[9]), .Z(n647) );
  XOR U715 ( .A(n642), .B(n641), .Z(c[63]) );
  XOR U716 ( .A(sreg[67]), .B(n640), .Z(n641) );
  XOR U717 ( .A(n651), .B(n652), .Z(n642) );
  XOR U718 ( .A(n653), .B(n640), .Z(n652) );
  XOR U719 ( .A(n654), .B(n655), .Z(n640) );
  NOR U720 ( .A(n656), .B(n657), .Z(n654) );
  AND U721 ( .A(b[0]), .B(a[3]), .Z(n653) );
  XOR U722 ( .A(n658), .B(n659), .Z(n651) );
  XOR U723 ( .A(n660), .B(n661), .Z(n659) );
  AND U724 ( .A(b[2]), .B(a[1]), .Z(n661) );
  AND U725 ( .A(a[0]), .B(b[3]), .Z(n660) );
  AND U726 ( .A(a[2]), .B(b[1]), .Z(n658) );
  XOR U727 ( .A(n657), .B(n656), .Z(c[62]) );
  XOR U728 ( .A(sreg[66]), .B(n655), .Z(n656) );
  XOR U729 ( .A(n662), .B(n663), .Z(n657) );
  XOR U730 ( .A(n665), .B(n666), .Z(n655) );
  NAND U731 ( .A(n667), .B(n668), .Z(n666) );
  AND U732 ( .A(b[0]), .B(a[2]), .Z(n664) );
  XOR U733 ( .A(n669), .B(n670), .Z(n662) );
  AND U734 ( .A(a[1]), .B(b[1]), .Z(n670) );
  AND U735 ( .A(b[2]), .B(a[0]), .Z(n669) );
  XOR U736 ( .A(n667), .B(n668), .Z(c[61]) );
  XOR U737 ( .A(sreg[65]), .B(n665), .Z(n668) );
  XNOR U738 ( .A(n665), .B(n671), .Z(n667) );
  XOR U739 ( .A(n672), .B(n673), .Z(n671) );
  NAND U740 ( .A(b[0]), .B(a[1]), .Z(n673) );
  AND U741 ( .A(a[0]), .B(b[1]), .Z(n672) );
  ANDN U742 ( .B(sreg[64]), .A(n674), .Z(n665) );
  XNOR U743 ( .A(sreg[64]), .B(n674), .Z(c[60]) );
  NAND U744 ( .A(a[0]), .B(b[0]), .Z(n674) );
endmodule

