
module hamming_N160_CC2 ( clk, rst, x, y, o );
  input [79:0] x;
  input [79:0] y;
  output [7:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526;
  wire   [7:0] oglobal;

  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  NAND U83 ( .A(n191), .B(n190), .Z(n1) );
  NAND U84 ( .A(n188), .B(n189), .Z(n2) );
  AND U85 ( .A(n1), .B(n2), .Z(n386) );
  NAND U86 ( .A(n398), .B(n399), .Z(n3) );
  XOR U87 ( .A(n398), .B(n399), .Z(n4) );
  NANDN U88 ( .A(n397), .B(n4), .Z(n5) );
  NAND U89 ( .A(n3), .B(n5), .Z(n468) );
  XOR U90 ( .A(n259), .B(n257), .Z(n6) );
  NANDN U91 ( .A(n258), .B(n6), .Z(n7) );
  NAND U92 ( .A(n259), .B(n257), .Z(n8) );
  AND U93 ( .A(n7), .B(n8), .Z(n422) );
  NAND U94 ( .A(n201), .B(n202), .Z(n9) );
  XOR U95 ( .A(n201), .B(n202), .Z(n10) );
  NANDN U96 ( .A(n200), .B(n10), .Z(n11) );
  NAND U97 ( .A(n9), .B(n11), .Z(n427) );
  NAND U98 ( .A(n440), .B(n442), .Z(n12) );
  XOR U99 ( .A(n440), .B(n442), .Z(n13) );
  NAND U100 ( .A(n13), .B(n441), .Z(n14) );
  NAND U101 ( .A(n12), .B(n14), .Z(n497) );
  XOR U102 ( .A(n338), .B(n336), .Z(n15) );
  NANDN U103 ( .A(n337), .B(n15), .Z(n16) );
  NAND U104 ( .A(n338), .B(n336), .Z(n17) );
  AND U105 ( .A(n16), .B(n17), .Z(n373) );
  XOR U106 ( .A(n304), .B(n302), .Z(n18) );
  NANDN U107 ( .A(n303), .B(n18), .Z(n19) );
  NAND U108 ( .A(n304), .B(n302), .Z(n20) );
  AND U109 ( .A(n19), .B(n20), .Z(n365) );
  NAND U110 ( .A(n221), .B(n222), .Z(n21) );
  XOR U111 ( .A(n221), .B(n222), .Z(n22) );
  NANDN U112 ( .A(n220), .B(n22), .Z(n23) );
  NAND U113 ( .A(n21), .B(n23), .Z(n378) );
  NAND U114 ( .A(n341), .B(n342), .Z(n24) );
  XOR U115 ( .A(n341), .B(n342), .Z(n25) );
  NANDN U116 ( .A(n340), .B(n25), .Z(n26) );
  NAND U117 ( .A(n24), .B(n26), .Z(n358) );
  NAND U118 ( .A(n426), .B(n427), .Z(n27) );
  XOR U119 ( .A(n426), .B(n427), .Z(n28) );
  NANDN U120 ( .A(n425), .B(n28), .Z(n29) );
  NAND U121 ( .A(n27), .B(n29), .Z(n460) );
  XOR U122 ( .A(n354), .B(n355), .Z(n30) );
  NANDN U123 ( .A(n356), .B(n30), .Z(n31) );
  NAND U124 ( .A(n354), .B(n355), .Z(n32) );
  AND U125 ( .A(n31), .B(n32), .Z(n455) );
  NAND U126 ( .A(n464), .B(n465), .Z(n33) );
  XOR U127 ( .A(n464), .B(n465), .Z(n34) );
  NANDN U128 ( .A(n463), .B(n34), .Z(n35) );
  NAND U129 ( .A(n33), .B(n35), .Z(n492) );
  NAND U130 ( .A(n497), .B(n499), .Z(n36) );
  XOR U131 ( .A(n497), .B(n499), .Z(n37) );
  NAND U132 ( .A(n37), .B(n498), .Z(n38) );
  NAND U133 ( .A(n36), .B(n38), .Z(n509) );
  NAND U134 ( .A(n210), .B(n209), .Z(n39) );
  NAND U135 ( .A(n207), .B(n208), .Z(n40) );
  AND U136 ( .A(n39), .B(n40), .Z(n398) );
  NAND U137 ( .A(n392), .B(n393), .Z(n41) );
  XOR U138 ( .A(n392), .B(n393), .Z(n42) );
  NANDN U139 ( .A(n391), .B(n42), .Z(n43) );
  NAND U140 ( .A(n41), .B(n43), .Z(n470) );
  NAND U141 ( .A(n386), .B(n387), .Z(n44) );
  XOR U142 ( .A(n386), .B(n387), .Z(n45) );
  NANDN U143 ( .A(n385), .B(n45), .Z(n46) );
  NAND U144 ( .A(n44), .B(n46), .Z(n466) );
  XOR U145 ( .A(oglobal[1]), .B(n389), .Z(n47) );
  XNOR U146 ( .A(n390), .B(n47), .Z(n374) );
  NAND U147 ( .A(n421), .B(n423), .Z(n48) );
  XOR U148 ( .A(n421), .B(n423), .Z(n49) );
  NAND U149 ( .A(n49), .B(n422), .Z(n50) );
  NAND U150 ( .A(n48), .B(n50), .Z(n465) );
  NAND U151 ( .A(n403), .B(n404), .Z(n51) );
  XOR U152 ( .A(n403), .B(n404), .Z(n52) );
  NANDN U153 ( .A(n402), .B(n52), .Z(n53) );
  NAND U154 ( .A(n51), .B(n53), .Z(n451) );
  NAND U155 ( .A(n179), .B(n180), .Z(n54) );
  XOR U156 ( .A(n179), .B(n180), .Z(n55) );
  NANDN U157 ( .A(n178), .B(n55), .Z(n56) );
  NAND U158 ( .A(n54), .B(n56), .Z(n354) );
  XNOR U159 ( .A(n435), .B(n434), .Z(n348) );
  NAND U160 ( .A(n473), .B(n474), .Z(n57) );
  XOR U161 ( .A(n473), .B(n474), .Z(n58) );
  NANDN U162 ( .A(n472), .B(n58), .Z(n59) );
  NAND U163 ( .A(n57), .B(n59), .Z(n485) );
  NAND U164 ( .A(n501), .B(n503), .Z(n60) );
  XOR U165 ( .A(n501), .B(n503), .Z(n61) );
  NAND U166 ( .A(n61), .B(n502), .Z(n62) );
  NAND U167 ( .A(n60), .B(n62), .Z(n505) );
  NAND U168 ( .A(n509), .B(n510), .Z(n63) );
  XOR U169 ( .A(n509), .B(n510), .Z(n64) );
  NANDN U170 ( .A(n508), .B(n64), .Z(n65) );
  NAND U171 ( .A(n63), .B(n65), .Z(n515) );
  XOR U172 ( .A(n382), .B(n383), .Z(n66) );
  NANDN U173 ( .A(n384), .B(n66), .Z(n67) );
  NAND U174 ( .A(n382), .B(n383), .Z(n68) );
  AND U175 ( .A(n67), .B(n68), .Z(n467) );
  NAND U176 ( .A(n419), .B(n420), .Z(n69) );
  XOR U177 ( .A(n419), .B(n420), .Z(n70) );
  NANDN U178 ( .A(n418), .B(n70), .Z(n71) );
  NAND U179 ( .A(n69), .B(n71), .Z(n464) );
  XOR U180 ( .A(oglobal[1]), .B(n389), .Z(n72) );
  NANDN U181 ( .A(n390), .B(n72), .Z(n73) );
  NAND U182 ( .A(oglobal[1]), .B(n389), .Z(n74) );
  AND U183 ( .A(n73), .B(n74), .Z(n445) );
  NAND U184 ( .A(n468), .B(n470), .Z(n75) );
  XOR U185 ( .A(n468), .B(n470), .Z(n76) );
  NAND U186 ( .A(n76), .B(n469), .Z(n77) );
  NAND U187 ( .A(n75), .B(n77), .Z(n486) );
  NAND U188 ( .A(n263), .B(n264), .Z(n78) );
  XOR U189 ( .A(n263), .B(n264), .Z(n79) );
  NANDN U190 ( .A(n262), .B(n79), .Z(n80) );
  NAND U191 ( .A(n78), .B(n80), .Z(n433) );
  XOR U192 ( .A(n452), .B(n450), .Z(n81) );
  NANDN U193 ( .A(n451), .B(n81), .Z(n82) );
  NAND U194 ( .A(n452), .B(n450), .Z(n83) );
  AND U195 ( .A(n82), .B(n83), .Z(n498) );
  NAND U196 ( .A(n430), .B(n431), .Z(n84) );
  XOR U197 ( .A(n430), .B(n431), .Z(n85) );
  NANDN U198 ( .A(n429), .B(n85), .Z(n86) );
  NAND U199 ( .A(n84), .B(n86), .Z(n473) );
  XOR U200 ( .A(n175), .B(n177), .Z(n87) );
  XNOR U201 ( .A(n176), .B(n87), .Z(n345) );
  XNOR U202 ( .A(n457), .B(n456), .Z(n479) );
  NAND U203 ( .A(n506), .B(n507), .Z(n88) );
  XOR U204 ( .A(n506), .B(n507), .Z(n89) );
  NANDN U205 ( .A(n505), .B(n89), .Z(n90) );
  NAND U206 ( .A(n88), .B(n90), .Z(n513) );
  NAND U207 ( .A(n206), .B(n205), .Z(n91) );
  NAND U208 ( .A(n203), .B(n204), .Z(n92) );
  AND U209 ( .A(n91), .B(n92), .Z(n399) );
  NAND U210 ( .A(n395), .B(n396), .Z(n93) );
  XOR U211 ( .A(n395), .B(n396), .Z(n94) );
  NANDN U212 ( .A(n394), .B(n94), .Z(n95) );
  NAND U213 ( .A(n93), .B(n95), .Z(n469) );
  XNOR U214 ( .A(n313), .B(n312), .Z(n314) );
  XNOR U215 ( .A(n307), .B(n306), .Z(n308) );
  NAND U216 ( .A(n160), .B(n159), .Z(n96) );
  NAND U217 ( .A(n157), .B(n158), .Z(n97) );
  AND U218 ( .A(n96), .B(n97), .Z(n393) );
  NAND U219 ( .A(n249), .B(n250), .Z(n98) );
  XOR U220 ( .A(n249), .B(n250), .Z(n99) );
  NANDN U221 ( .A(n248), .B(n99), .Z(n100) );
  NAND U222 ( .A(n98), .B(n100), .Z(n421) );
  NAND U223 ( .A(n467), .B(n466), .Z(n101) );
  XOR U224 ( .A(n467), .B(n466), .Z(n102) );
  NANDN U225 ( .A(oglobal[2]), .B(n102), .Z(n103) );
  NAND U226 ( .A(n101), .B(n103), .Z(n488) );
  NAND U227 ( .A(n379), .B(n380), .Z(n104) );
  XOR U228 ( .A(n379), .B(n380), .Z(n105) );
  NAND U229 ( .A(n105), .B(n378), .Z(n106) );
  NAND U230 ( .A(n104), .B(n106), .Z(n441) );
  XOR U231 ( .A(n358), .B(n357), .Z(n107) );
  XNOR U232 ( .A(n360), .B(n107), .Z(n432) );
  NAND U233 ( .A(n461), .B(n462), .Z(n108) );
  XOR U234 ( .A(n461), .B(n462), .Z(n109) );
  NAND U235 ( .A(n109), .B(n460), .Z(n110) );
  NAND U236 ( .A(n108), .B(n110), .Z(n494) );
  XOR U237 ( .A(n177), .B(n175), .Z(n111) );
  NANDN U238 ( .A(n176), .B(n111), .Z(n112) );
  NAND U239 ( .A(n177), .B(n175), .Z(n113) );
  AND U240 ( .A(n112), .B(n113), .Z(n356) );
  XOR U241 ( .A(n343), .B(n344), .Z(n114) );
  NANDN U242 ( .A(n345), .B(n114), .Z(n115) );
  NAND U243 ( .A(n343), .B(n344), .Z(n116) );
  AND U244 ( .A(n115), .B(n116), .Z(n349) );
  NAND U245 ( .A(n483), .B(n485), .Z(n117) );
  XOR U246 ( .A(n483), .B(n485), .Z(n118) );
  NAND U247 ( .A(n118), .B(n484), .Z(n119) );
  NAND U248 ( .A(n117), .B(n119), .Z(n506) );
  NAND U249 ( .A(n520), .B(n521), .Z(n525) );
  XOR U250 ( .A(x[13]), .B(y[13]), .Z(n196) );
  XOR U251 ( .A(x[9]), .B(y[9]), .Z(n193) );
  XOR U252 ( .A(x[11]), .B(y[11]), .Z(n192) );
  XOR U253 ( .A(n193), .B(n192), .Z(n195) );
  XOR U254 ( .A(n196), .B(n195), .Z(n259) );
  XOR U255 ( .A(x[25]), .B(y[25]), .Z(n298) );
  XOR U256 ( .A(x[21]), .B(y[21]), .Z(n295) );
  XNOR U257 ( .A(x[23]), .B(y[23]), .Z(n296) );
  XNOR U258 ( .A(n295), .B(n296), .Z(n297) );
  XNOR U259 ( .A(n298), .B(n297), .Z(n258) );
  XOR U260 ( .A(x[19]), .B(y[19]), .Z(n292) );
  XOR U261 ( .A(x[15]), .B(y[15]), .Z(n289) );
  XNOR U262 ( .A(x[17]), .B(y[17]), .Z(n290) );
  XNOR U263 ( .A(n289), .B(n290), .Z(n291) );
  XOR U264 ( .A(n292), .B(n291), .Z(n257) );
  XOR U265 ( .A(n258), .B(n257), .Z(n120) );
  XOR U266 ( .A(n259), .B(n120), .Z(n177) );
  XOR U267 ( .A(x[7]), .B(y[7]), .Z(n184) );
  XOR U268 ( .A(x[5]), .B(y[5]), .Z(n182) );
  XNOR U269 ( .A(x[3]), .B(y[3]), .Z(n183) );
  XOR U270 ( .A(n182), .B(n183), .Z(n185) );
  XOR U271 ( .A(n184), .B(n185), .Z(n340) );
  XOR U272 ( .A(x[4]), .B(y[4]), .Z(n237) );
  XOR U273 ( .A(x[6]), .B(y[6]), .Z(n235) );
  XNOR U274 ( .A(x[8]), .B(y[8]), .Z(n236) );
  XOR U275 ( .A(n235), .B(n236), .Z(n238) );
  XNOR U276 ( .A(n237), .B(n238), .Z(n342) );
  XOR U277 ( .A(x[1]), .B(y[1]), .Z(n231) );
  XOR U278 ( .A(x[0]), .B(y[0]), .Z(n229) );
  XNOR U279 ( .A(x[2]), .B(y[2]), .Z(n230) );
  XOR U280 ( .A(n229), .B(n230), .Z(n232) );
  XNOR U281 ( .A(n231), .B(n232), .Z(n341) );
  XNOR U282 ( .A(n342), .B(n341), .Z(n121) );
  XOR U283 ( .A(n340), .B(n121), .Z(n176) );
  XOR U284 ( .A(x[64]), .B(y[64]), .Z(n147) );
  XOR U285 ( .A(x[66]), .B(y[66]), .Z(n144) );
  XNOR U286 ( .A(x[68]), .B(y[68]), .Z(n145) );
  XNOR U287 ( .A(n144), .B(n145), .Z(n146) );
  XOR U288 ( .A(n147), .B(n146), .Z(n338) );
  XOR U289 ( .A(x[58]), .B(y[58]), .Z(n164) );
  XOR U290 ( .A(x[60]), .B(y[60]), .Z(n161) );
  XNOR U291 ( .A(x[62]), .B(y[62]), .Z(n162) );
  XNOR U292 ( .A(n161), .B(n162), .Z(n163) );
  XNOR U293 ( .A(n164), .B(n163), .Z(n337) );
  XOR U294 ( .A(x[70]), .B(y[70]), .Z(n243) );
  XNOR U295 ( .A(x[72]), .B(y[72]), .Z(n241) );
  XNOR U296 ( .A(oglobal[0]), .B(n241), .Z(n242) );
  XOR U297 ( .A(n243), .B(n242), .Z(n336) );
  XOR U298 ( .A(n337), .B(n336), .Z(n122) );
  XOR U299 ( .A(n338), .B(n122), .Z(n175) );
  XOR U300 ( .A(x[22]), .B(y[22]), .Z(n170) );
  XOR U301 ( .A(x[24]), .B(y[24]), .Z(n167) );
  XNOR U302 ( .A(x[26]), .B(y[26]), .Z(n168) );
  XNOR U303 ( .A(n167), .B(n168), .Z(n169) );
  XNOR U304 ( .A(n170), .B(n169), .Z(n202) );
  XOR U305 ( .A(x[10]), .B(y[10]), .Z(n153) );
  XOR U306 ( .A(x[12]), .B(y[12]), .Z(n150) );
  XNOR U307 ( .A(x[14]), .B(y[14]), .Z(n151) );
  XNOR U308 ( .A(n150), .B(n151), .Z(n152) );
  XNOR U309 ( .A(n153), .B(n152), .Z(n201) );
  XOR U310 ( .A(x[16]), .B(y[16]), .Z(n141) );
  XOR U311 ( .A(x[18]), .B(y[18]), .Z(n138) );
  XNOR U312 ( .A(x[20]), .B(y[20]), .Z(n139) );
  XNOR U313 ( .A(n138), .B(n139), .Z(n140) );
  XOR U314 ( .A(n141), .B(n140), .Z(n200) );
  XOR U315 ( .A(n201), .B(n200), .Z(n123) );
  XNOR U316 ( .A(n202), .B(n123), .Z(n264) );
  XOR U317 ( .A(x[40]), .B(y[40]), .Z(n206) );
  XOR U318 ( .A(x[42]), .B(y[42]), .Z(n204) );
  XOR U319 ( .A(x[44]), .B(y[44]), .Z(n203) );
  XOR U320 ( .A(n204), .B(n203), .Z(n205) );
  XNOR U321 ( .A(n206), .B(n205), .Z(n253) );
  XOR U322 ( .A(x[28]), .B(y[28]), .Z(n160) );
  XOR U323 ( .A(x[30]), .B(y[30]), .Z(n158) );
  XOR U324 ( .A(x[32]), .B(y[32]), .Z(n157) );
  XOR U325 ( .A(n158), .B(n157), .Z(n159) );
  XNOR U326 ( .A(n160), .B(n159), .Z(n252) );
  XOR U327 ( .A(x[34]), .B(y[34]), .Z(n215) );
  XOR U328 ( .A(x[36]), .B(y[36]), .Z(n212) );
  XOR U329 ( .A(x[38]), .B(y[38]), .Z(n211) );
  XOR U330 ( .A(n212), .B(n211), .Z(n214) );
  XOR U331 ( .A(n215), .B(n214), .Z(n251) );
  XOR U332 ( .A(n252), .B(n251), .Z(n124) );
  XNOR U333 ( .A(n253), .B(n124), .Z(n263) );
  XOR U334 ( .A(x[52]), .B(y[52]), .Z(n210) );
  XOR U335 ( .A(x[54]), .B(y[54]), .Z(n208) );
  XOR U336 ( .A(x[56]), .B(y[56]), .Z(n207) );
  XOR U337 ( .A(n208), .B(n207), .Z(n209) );
  XNOR U338 ( .A(n210), .B(n209), .Z(n250) );
  XOR U339 ( .A(x[46]), .B(y[46]), .Z(n135) );
  XOR U340 ( .A(x[48]), .B(y[48]), .Z(n132) );
  XNOR U341 ( .A(x[50]), .B(y[50]), .Z(n133) );
  XNOR U342 ( .A(n132), .B(n133), .Z(n134) );
  XNOR U343 ( .A(n135), .B(n134), .Z(n249) );
  XOR U344 ( .A(x[74]), .B(y[74]), .Z(n191) );
  XOR U345 ( .A(x[76]), .B(y[76]), .Z(n189) );
  XOR U346 ( .A(x[78]), .B(y[78]), .Z(n188) );
  XOR U347 ( .A(n189), .B(n188), .Z(n190) );
  XOR U348 ( .A(n191), .B(n190), .Z(n248) );
  XOR U349 ( .A(n249), .B(n248), .Z(n125) );
  XOR U350 ( .A(n250), .B(n125), .Z(n262) );
  XOR U351 ( .A(n263), .B(n262), .Z(n126) );
  XOR U352 ( .A(n264), .B(n126), .Z(n343) );
  XOR U353 ( .A(x[63]), .B(y[63]), .Z(n315) );
  XOR U354 ( .A(x[61]), .B(y[61]), .Z(n312) );
  XNOR U355 ( .A(x[71]), .B(y[71]), .Z(n313) );
  XNOR U356 ( .A(n315), .B(n314), .Z(n304) );
  XOR U357 ( .A(x[55]), .B(y[55]), .Z(n332) );
  XOR U358 ( .A(x[75]), .B(y[75]), .Z(n330) );
  XNOR U359 ( .A(x[53]), .B(y[53]), .Z(n331) );
  XOR U360 ( .A(n330), .B(n331), .Z(n333) );
  XOR U361 ( .A(n332), .B(n333), .Z(n302) );
  XOR U362 ( .A(x[59]), .B(y[59]), .Z(n309) );
  XOR U363 ( .A(x[57]), .B(y[57]), .Z(n306) );
  XNOR U364 ( .A(x[73]), .B(y[73]), .Z(n307) );
  XOR U365 ( .A(n309), .B(n308), .Z(n303) );
  XOR U366 ( .A(n302), .B(n303), .Z(n127) );
  XNOR U367 ( .A(n304), .B(n127), .Z(n180) );
  XOR U368 ( .A(x[37]), .B(y[37]), .Z(n274) );
  XOR U369 ( .A(x[35]), .B(y[35]), .Z(n271) );
  XNOR U370 ( .A(x[33]), .B(y[33]), .Z(n272) );
  XNOR U371 ( .A(n271), .B(n272), .Z(n273) );
  XNOR U372 ( .A(n274), .B(n273), .Z(n225) );
  XOR U373 ( .A(x[31]), .B(y[31]), .Z(n286) );
  XOR U374 ( .A(x[27]), .B(y[27]), .Z(n283) );
  XNOR U375 ( .A(x[29]), .B(y[29]), .Z(n284) );
  XNOR U376 ( .A(n283), .B(n284), .Z(n285) );
  XNOR U377 ( .A(n286), .B(n285), .Z(n224) );
  XOR U378 ( .A(x[43]), .B(y[43]), .Z(n280) );
  XOR U379 ( .A(x[41]), .B(y[41]), .Z(n277) );
  XNOR U380 ( .A(x[39]), .B(y[39]), .Z(n278) );
  XNOR U381 ( .A(n277), .B(n278), .Z(n279) );
  XOR U382 ( .A(n280), .B(n279), .Z(n223) );
  XOR U383 ( .A(n224), .B(n223), .Z(n128) );
  XNOR U384 ( .A(n225), .B(n128), .Z(n179) );
  XOR U385 ( .A(x[47]), .B(y[47]), .Z(n268) );
  XOR U386 ( .A(x[79]), .B(y[79]), .Z(n265) );
  XNOR U387 ( .A(x[45]), .B(y[45]), .Z(n266) );
  XNOR U388 ( .A(n265), .B(n266), .Z(n267) );
  XNOR U389 ( .A(n268), .B(n267), .Z(n222) );
  XOR U390 ( .A(x[67]), .B(y[67]), .Z(n321) );
  XOR U391 ( .A(x[69]), .B(y[69]), .Z(n318) );
  XNOR U392 ( .A(x[65]), .B(y[65]), .Z(n319) );
  XNOR U393 ( .A(n318), .B(n319), .Z(n320) );
  XNOR U394 ( .A(n321), .B(n320), .Z(n221) );
  XOR U395 ( .A(x[51]), .B(y[51]), .Z(n327) );
  XOR U396 ( .A(x[77]), .B(y[77]), .Z(n324) );
  XNOR U397 ( .A(x[49]), .B(y[49]), .Z(n325) );
  XNOR U398 ( .A(n324), .B(n325), .Z(n326) );
  XOR U399 ( .A(n327), .B(n326), .Z(n220) );
  XOR U400 ( .A(n221), .B(n220), .Z(n129) );
  XOR U401 ( .A(n222), .B(n129), .Z(n178) );
  XOR U402 ( .A(n179), .B(n178), .Z(n130) );
  XOR U403 ( .A(n180), .B(n130), .Z(n344) );
  XOR U404 ( .A(n343), .B(n344), .Z(n131) );
  XNOR U405 ( .A(n345), .B(n131), .Z(o[0]) );
  NANDN U406 ( .A(n133), .B(n132), .Z(n137) );
  NAND U407 ( .A(n135), .B(n134), .Z(n136) );
  NAND U408 ( .A(n137), .B(n136), .Z(n418) );
  NANDN U409 ( .A(n139), .B(n138), .Z(n143) );
  NAND U410 ( .A(n141), .B(n140), .Z(n142) );
  AND U411 ( .A(n143), .B(n142), .Z(n396) );
  NANDN U412 ( .A(n145), .B(n144), .Z(n149) );
  NAND U413 ( .A(n147), .B(n146), .Z(n148) );
  AND U414 ( .A(n149), .B(n148), .Z(n395) );
  NANDN U415 ( .A(n151), .B(n150), .Z(n155) );
  NAND U416 ( .A(n153), .B(n152), .Z(n154) );
  NAND U417 ( .A(n155), .B(n154), .Z(n394) );
  XOR U418 ( .A(n395), .B(n394), .Z(n156) );
  XNOR U419 ( .A(n396), .B(n156), .Z(n420) );
  NANDN U420 ( .A(n162), .B(n161), .Z(n166) );
  NAND U421 ( .A(n164), .B(n163), .Z(n165) );
  AND U422 ( .A(n166), .B(n165), .Z(n392) );
  NANDN U423 ( .A(n168), .B(n167), .Z(n172) );
  NAND U424 ( .A(n170), .B(n169), .Z(n171) );
  NAND U425 ( .A(n172), .B(n171), .Z(n391) );
  XOR U426 ( .A(n392), .B(n391), .Z(n173) );
  XNOR U427 ( .A(n393), .B(n173), .Z(n419) );
  XNOR U428 ( .A(n420), .B(n419), .Z(n174) );
  XOR U429 ( .A(n418), .B(n174), .Z(n355) );
  XNOR U430 ( .A(n356), .B(n354), .Z(n181) );
  XOR U431 ( .A(n355), .B(n181), .Z(n350) );
  NANDN U432 ( .A(n183), .B(n182), .Z(n187) );
  NANDN U433 ( .A(n185), .B(n184), .Z(n186) );
  AND U434 ( .A(n187), .B(n186), .Z(n387) );
  IV U435 ( .A(n192), .Z(n194) );
  NANDN U436 ( .A(n194), .B(n193), .Z(n198) );
  NAND U437 ( .A(n196), .B(n195), .Z(n197) );
  NAND U438 ( .A(n198), .B(n197), .Z(n385) );
  XOR U439 ( .A(n386), .B(n385), .Z(n199) );
  XOR U440 ( .A(n387), .B(n199), .Z(n425) );
  IV U441 ( .A(n211), .Z(n213) );
  NANDN U442 ( .A(n213), .B(n212), .Z(n217) );
  NAND U443 ( .A(n215), .B(n214), .Z(n216) );
  NAND U444 ( .A(n217), .B(n216), .Z(n397) );
  XOR U445 ( .A(n398), .B(n397), .Z(n218) );
  XNOR U446 ( .A(n399), .B(n218), .Z(n426) );
  XNOR U447 ( .A(n427), .B(n426), .Z(n219) );
  XOR U448 ( .A(n425), .B(n219), .Z(n430) );
  NANDN U449 ( .A(n224), .B(n223), .Z(n228) );
  ANDN U450 ( .B(n224), .A(n223), .Z(n226) );
  OR U451 ( .A(n226), .B(n225), .Z(n227) );
  AND U452 ( .A(n228), .B(n227), .Z(n380) );
  NANDN U453 ( .A(n230), .B(n229), .Z(n234) );
  NANDN U454 ( .A(n232), .B(n231), .Z(n233) );
  NAND U455 ( .A(n234), .B(n233), .Z(n383) );
  NANDN U456 ( .A(n236), .B(n235), .Z(n240) );
  NANDN U457 ( .A(n238), .B(n237), .Z(n239) );
  AND U458 ( .A(n240), .B(n239), .Z(n384) );
  NANDN U459 ( .A(n241), .B(oglobal[0]), .Z(n245) );
  NAND U460 ( .A(n243), .B(n242), .Z(n244) );
  NAND U461 ( .A(n245), .B(n244), .Z(n382) );
  XOR U462 ( .A(n384), .B(n382), .Z(n246) );
  XOR U463 ( .A(n383), .B(n246), .Z(n379) );
  XNOR U464 ( .A(n380), .B(n379), .Z(n247) );
  XNOR U465 ( .A(n378), .B(n247), .Z(n431) );
  NANDN U466 ( .A(n252), .B(n251), .Z(n256) );
  ANDN U467 ( .B(n252), .A(n251), .Z(n254) );
  OR U468 ( .A(n254), .B(n253), .Z(n255) );
  AND U469 ( .A(n256), .B(n255), .Z(n423) );
  XNOR U470 ( .A(n423), .B(n422), .Z(n260) );
  XOR U471 ( .A(n421), .B(n260), .Z(n429) );
  XOR U472 ( .A(n431), .B(n429), .Z(n261) );
  XOR U473 ( .A(n430), .B(n261), .Z(n434) );
  NANDN U474 ( .A(n266), .B(n265), .Z(n270) );
  NAND U475 ( .A(n268), .B(n267), .Z(n269) );
  AND U476 ( .A(n270), .B(n269), .Z(n411) );
  NANDN U477 ( .A(n272), .B(n271), .Z(n276) );
  NAND U478 ( .A(n274), .B(n273), .Z(n275) );
  NAND U479 ( .A(n276), .B(n275), .Z(n412) );
  XNOR U480 ( .A(n411), .B(n412), .Z(n413) );
  NANDN U481 ( .A(n278), .B(n277), .Z(n282) );
  NAND U482 ( .A(n280), .B(n279), .Z(n281) );
  NAND U483 ( .A(n282), .B(n281), .Z(n414) );
  XOR U484 ( .A(n413), .B(n414), .Z(n366) );
  NANDN U485 ( .A(n284), .B(n283), .Z(n288) );
  NAND U486 ( .A(n286), .B(n285), .Z(n287) );
  NAND U487 ( .A(n288), .B(n287), .Z(n402) );
  NANDN U488 ( .A(n290), .B(n289), .Z(n294) );
  NAND U489 ( .A(n292), .B(n291), .Z(n293) );
  AND U490 ( .A(n294), .B(n293), .Z(n404) );
  NANDN U491 ( .A(n296), .B(n295), .Z(n300) );
  NAND U492 ( .A(n298), .B(n297), .Z(n299) );
  AND U493 ( .A(n300), .B(n299), .Z(n403) );
  XNOR U494 ( .A(n404), .B(n403), .Z(n301) );
  XOR U495 ( .A(n402), .B(n301), .Z(n368) );
  XNOR U496 ( .A(n368), .B(n365), .Z(n305) );
  XOR U497 ( .A(n366), .B(n305), .Z(n360) );
  NANDN U498 ( .A(n307), .B(n306), .Z(n311) );
  NAND U499 ( .A(n309), .B(n308), .Z(n310) );
  NAND U500 ( .A(n311), .B(n310), .Z(n389) );
  NANDN U501 ( .A(n313), .B(n312), .Z(n317) );
  NAND U502 ( .A(n315), .B(n314), .Z(n316) );
  AND U503 ( .A(n317), .B(n316), .Z(n390) );
  NANDN U504 ( .A(n319), .B(n318), .Z(n323) );
  NAND U505 ( .A(n321), .B(n320), .Z(n322) );
  AND U506 ( .A(n323), .B(n322), .Z(n405) );
  NANDN U507 ( .A(n325), .B(n324), .Z(n329) );
  NAND U508 ( .A(n327), .B(n326), .Z(n328) );
  NAND U509 ( .A(n329), .B(n328), .Z(n406) );
  XNOR U510 ( .A(n405), .B(n406), .Z(n407) );
  NANDN U511 ( .A(n331), .B(n330), .Z(n335) );
  NANDN U512 ( .A(n333), .B(n332), .Z(n334) );
  NAND U513 ( .A(n335), .B(n334), .Z(n408) );
  XOR U514 ( .A(n407), .B(n408), .Z(n372) );
  XOR U515 ( .A(n372), .B(n373), .Z(n339) );
  XNOR U516 ( .A(n374), .B(n339), .Z(n359) );
  IV U517 ( .A(n359), .Z(n357) );
  XOR U518 ( .A(n433), .B(n432), .Z(n435) );
  IV U519 ( .A(n348), .Z(n347) );
  XOR U520 ( .A(n347), .B(n349), .Z(n346) );
  XNOR U521 ( .A(n350), .B(n346), .Z(o[1]) );
  OR U522 ( .A(n349), .B(n347), .Z(n353) );
  ANDN U523 ( .B(n349), .A(n348), .Z(n351) );
  OR U524 ( .A(n351), .B(n350), .Z(n352) );
  AND U525 ( .A(n353), .B(n352), .Z(n477) );
  NANDN U526 ( .A(n357), .B(n358), .Z(n363) );
  NOR U527 ( .A(n359), .B(n358), .Z(n361) );
  NANDN U528 ( .A(n361), .B(n360), .Z(n362) );
  AND U529 ( .A(n363), .B(n362), .Z(n454) );
  XNOR U530 ( .A(n455), .B(n454), .Z(n456) );
  IV U531 ( .A(n366), .Z(n364) );
  NANDN U532 ( .A(n364), .B(n365), .Z(n370) );
  NOR U533 ( .A(n366), .B(n365), .Z(n367) );
  OR U534 ( .A(n368), .B(n367), .Z(n369) );
  AND U535 ( .A(n370), .B(n369), .Z(n440) );
  IV U536 ( .A(n372), .Z(n371) );
  OR U537 ( .A(n373), .B(n371), .Z(n377) );
  ANDN U538 ( .B(n373), .A(n372), .Z(n375) );
  NANDN U539 ( .A(n375), .B(n374), .Z(n376) );
  AND U540 ( .A(n377), .B(n376), .Z(n442) );
  XNOR U541 ( .A(n442), .B(n441), .Z(n381) );
  XOR U542 ( .A(n440), .B(n381), .Z(n457) );
  XOR U543 ( .A(n467), .B(n466), .Z(n388) );
  XNOR U544 ( .A(oglobal[2]), .B(n388), .Z(n446) );
  XNOR U545 ( .A(n469), .B(n468), .Z(n400) );
  XOR U546 ( .A(n470), .B(n400), .Z(n444) );
  XOR U547 ( .A(n445), .B(n444), .Z(n401) );
  XNOR U548 ( .A(n446), .B(n401), .Z(n462) );
  NANDN U549 ( .A(n406), .B(n405), .Z(n410) );
  NANDN U550 ( .A(n408), .B(n407), .Z(n409) );
  AND U551 ( .A(n410), .B(n409), .Z(n452) );
  NANDN U552 ( .A(n412), .B(n411), .Z(n416) );
  NANDN U553 ( .A(n414), .B(n413), .Z(n415) );
  AND U554 ( .A(n416), .B(n415), .Z(n450) );
  XNOR U555 ( .A(n452), .B(n450), .Z(n417) );
  XOR U556 ( .A(n451), .B(n417), .Z(n463) );
  XNOR U557 ( .A(n464), .B(n465), .Z(n424) );
  XOR U558 ( .A(n463), .B(n424), .Z(n461) );
  XNOR U559 ( .A(n461), .B(n460), .Z(n428) );
  XNOR U560 ( .A(n462), .B(n428), .Z(n474) );
  NANDN U561 ( .A(n433), .B(n432), .Z(n437) );
  NANDN U562 ( .A(n435), .B(n434), .Z(n436) );
  NAND U563 ( .A(n437), .B(n436), .Z(n472) );
  XOR U564 ( .A(n473), .B(n472), .Z(n438) );
  XOR U565 ( .A(n474), .B(n438), .Z(n476) );
  IV U566 ( .A(n476), .Z(n475) );
  XOR U567 ( .A(n479), .B(n475), .Z(n439) );
  XNOR U568 ( .A(n477), .B(n439), .Z(o[2]) );
  IV U569 ( .A(n444), .Z(n443) );
  OR U570 ( .A(n445), .B(n443), .Z(n449) );
  ANDN U571 ( .B(n445), .A(n444), .Z(n447) );
  OR U572 ( .A(n447), .B(n446), .Z(n448) );
  AND U573 ( .A(n449), .B(n448), .Z(n499) );
  XNOR U574 ( .A(n499), .B(n498), .Z(n453) );
  XOR U575 ( .A(n497), .B(n453), .Z(n503) );
  NANDN U576 ( .A(n455), .B(n454), .Z(n459) );
  NANDN U577 ( .A(n457), .B(n456), .Z(n458) );
  AND U578 ( .A(n459), .B(n458), .Z(n502) );
  XNOR U579 ( .A(n486), .B(oglobal[3]), .Z(n487) );
  XNOR U580 ( .A(n488), .B(n487), .Z(n491) );
  XNOR U581 ( .A(n492), .B(n491), .Z(n493) );
  XNOR U582 ( .A(n494), .B(n493), .Z(n501) );
  XNOR U583 ( .A(n502), .B(n501), .Z(n471) );
  XOR U584 ( .A(n503), .B(n471), .Z(n483) );
  OR U585 ( .A(n477), .B(n475), .Z(n481) );
  ANDN U586 ( .B(n477), .A(n476), .Z(n478) );
  OR U587 ( .A(n479), .B(n478), .Z(n480) );
  AND U588 ( .A(n481), .B(n480), .Z(n484) );
  XNOR U589 ( .A(n485), .B(n484), .Z(n482) );
  XOR U590 ( .A(n483), .B(n482), .Z(o[3]) );
  NANDN U591 ( .A(n486), .B(oglobal[3]), .Z(n490) );
  NANDN U592 ( .A(n488), .B(n487), .Z(n489) );
  NAND U593 ( .A(n490), .B(n489), .Z(n511) );
  XOR U594 ( .A(oglobal[4]), .B(n511), .Z(n508) );
  NANDN U595 ( .A(n492), .B(n491), .Z(n496) );
  NANDN U596 ( .A(n494), .B(n493), .Z(n495) );
  AND U597 ( .A(n496), .B(n495), .Z(n510) );
  XNOR U598 ( .A(n510), .B(n509), .Z(n500) );
  XOR U599 ( .A(n508), .B(n500), .Z(n507) );
  XNOR U600 ( .A(n507), .B(n505), .Z(n504) );
  XNOR U601 ( .A(n506), .B(n504), .Z(o[4]) );
  AND U602 ( .A(oglobal[4]), .B(n511), .Z(n518) );
  XOR U603 ( .A(n518), .B(oglobal[5]), .Z(n514) );
  XNOR U604 ( .A(n515), .B(n514), .Z(n512) );
  XNOR U605 ( .A(n513), .B(n512), .Z(o[5]) );
  NANDN U606 ( .A(n513), .B(n514), .Z(n517) );
  NANDN U607 ( .A(n514), .B(n513), .Z(n516) );
  ANDN U608 ( .B(n516), .A(n515), .Z(n521) );
  ANDN U609 ( .B(n517), .A(n521), .Z(n519) );
  AND U610 ( .A(n518), .B(oglobal[5]), .Z(n520) );
  ANDN U611 ( .B(n519), .A(n520), .Z(n523) );
  NANDN U612 ( .A(n523), .B(n525), .Z(n522) );
  XNOR U613 ( .A(oglobal[6]), .B(n522), .Z(o[6]) );
  NANDN U614 ( .A(n523), .B(oglobal[6]), .Z(n524) );
  AND U615 ( .A(n525), .B(n524), .Z(n526) );
  XNOR U616 ( .A(oglobal[7]), .B(n526), .Z(o[7]) );
endmodule

