
module MUX_N256_0 ( A, B, S, O );
  input [255:0] A;
  input [255:0] B;
  output [255:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[50]), .B(n109), .Z(O[50]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U166 ( .A(A[4]), .B(n111), .Z(O[4]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U169 ( .A(A[49]), .B(n113), .Z(O[49]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U172 ( .A(A[48]), .B(n115), .Z(O[48]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U175 ( .A(A[47]), .B(n117), .Z(O[47]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U178 ( .A(A[46]), .B(n119), .Z(O[46]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U181 ( .A(A[45]), .B(n121), .Z(O[45]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U184 ( .A(A[44]), .B(n123), .Z(O[44]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U187 ( .A(A[43]), .B(n125), .Z(O[43]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U190 ( .A(A[42]), .B(n127), .Z(O[42]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U193 ( .A(A[41]), .B(n129), .Z(O[41]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U196 ( .A(A[40]), .B(n131), .Z(O[40]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U199 ( .A(A[3]), .B(n133), .Z(O[3]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U202 ( .A(A[39]), .B(n135), .Z(O[39]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U205 ( .A(A[38]), .B(n137), .Z(O[38]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U208 ( .A(A[37]), .B(n139), .Z(O[37]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U211 ( .A(A[36]), .B(n141), .Z(O[36]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U214 ( .A(A[35]), .B(n143), .Z(O[35]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U217 ( .A(A[34]), .B(n145), .Z(O[34]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U220 ( .A(A[33]), .B(n147), .Z(O[33]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U223 ( .A(A[32]), .B(n149), .Z(O[32]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U226 ( .A(A[31]), .B(n151), .Z(O[31]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U229 ( .A(A[30]), .B(n153), .Z(O[30]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U232 ( .A(A[2]), .B(n155), .Z(O[2]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U235 ( .A(A[29]), .B(n157), .Z(O[29]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U238 ( .A(A[28]), .B(n159), .Z(O[28]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U241 ( .A(A[27]), .B(n161), .Z(O[27]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U244 ( .A(A[26]), .B(n163), .Z(O[26]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U247 ( .A(A[25]), .B(n165), .Z(O[25]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U250 ( .A(A[255]), .B(n167), .Z(O[255]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[255]), .B(A[255]), .Z(n168) );
  XOR U253 ( .A(A[254]), .B(n169), .Z(O[254]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[254]), .B(A[254]), .Z(n170) );
  XOR U256 ( .A(A[253]), .B(n171), .Z(O[253]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[253]), .B(A[253]), .Z(n172) );
  XOR U259 ( .A(A[252]), .B(n173), .Z(O[252]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[252]), .B(A[252]), .Z(n174) );
  XOR U262 ( .A(A[251]), .B(n175), .Z(O[251]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[251]), .B(A[251]), .Z(n176) );
  XOR U265 ( .A(A[250]), .B(n177), .Z(O[250]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[250]), .B(A[250]), .Z(n178) );
  XOR U268 ( .A(A[24]), .B(n179), .Z(O[24]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[24]), .B(A[24]), .Z(n180) );
  XOR U271 ( .A(A[249]), .B(n181), .Z(O[249]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[249]), .B(A[249]), .Z(n182) );
  XOR U274 ( .A(A[248]), .B(n183), .Z(O[248]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[248]), .B(A[248]), .Z(n184) );
  XOR U277 ( .A(A[247]), .B(n185), .Z(O[247]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[247]), .B(A[247]), .Z(n186) );
  XOR U280 ( .A(A[246]), .B(n187), .Z(O[246]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[246]), .B(A[246]), .Z(n188) );
  XOR U283 ( .A(A[245]), .B(n189), .Z(O[245]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[245]), .B(A[245]), .Z(n190) );
  XOR U286 ( .A(A[244]), .B(n191), .Z(O[244]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[244]), .B(A[244]), .Z(n192) );
  XOR U289 ( .A(A[243]), .B(n193), .Z(O[243]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[243]), .B(A[243]), .Z(n194) );
  XOR U292 ( .A(A[242]), .B(n195), .Z(O[242]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[242]), .B(A[242]), .Z(n196) );
  XOR U295 ( .A(A[241]), .B(n197), .Z(O[241]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[241]), .B(A[241]), .Z(n198) );
  XOR U298 ( .A(A[240]), .B(n199), .Z(O[240]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[240]), .B(A[240]), .Z(n200) );
  XOR U301 ( .A(A[23]), .B(n201), .Z(O[23]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[23]), .B(A[23]), .Z(n202) );
  XOR U304 ( .A(A[239]), .B(n203), .Z(O[239]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[239]), .B(A[239]), .Z(n204) );
  XOR U307 ( .A(A[238]), .B(n205), .Z(O[238]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[238]), .B(A[238]), .Z(n206) );
  XOR U310 ( .A(A[237]), .B(n207), .Z(O[237]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[237]), .B(A[237]), .Z(n208) );
  XOR U313 ( .A(A[236]), .B(n209), .Z(O[236]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[236]), .B(A[236]), .Z(n210) );
  XOR U316 ( .A(A[235]), .B(n211), .Z(O[235]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[235]), .B(A[235]), .Z(n212) );
  XOR U319 ( .A(A[234]), .B(n213), .Z(O[234]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[234]), .B(A[234]), .Z(n214) );
  XOR U322 ( .A(A[233]), .B(n215), .Z(O[233]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[233]), .B(A[233]), .Z(n216) );
  XOR U325 ( .A(A[232]), .B(n217), .Z(O[232]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[232]), .B(A[232]), .Z(n218) );
  XOR U328 ( .A(A[231]), .B(n219), .Z(O[231]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[231]), .B(A[231]), .Z(n220) );
  XOR U331 ( .A(A[230]), .B(n221), .Z(O[230]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[230]), .B(A[230]), .Z(n222) );
  XOR U334 ( .A(A[22]), .B(n223), .Z(O[22]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[22]), .B(A[22]), .Z(n224) );
  XOR U337 ( .A(A[229]), .B(n225), .Z(O[229]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n226) );
  XOR U340 ( .A(A[228]), .B(n227), .Z(O[228]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[228]), .B(A[228]), .Z(n228) );
  XOR U343 ( .A(A[227]), .B(n229), .Z(O[227]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[227]), .B(A[227]), .Z(n230) );
  XOR U346 ( .A(A[226]), .B(n231), .Z(O[226]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[226]), .B(A[226]), .Z(n232) );
  XOR U349 ( .A(A[225]), .B(n233), .Z(O[225]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[225]), .B(A[225]), .Z(n234) );
  XOR U352 ( .A(A[224]), .B(n235), .Z(O[224]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[224]), .B(A[224]), .Z(n236) );
  XOR U355 ( .A(A[223]), .B(n237), .Z(O[223]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[223]), .B(A[223]), .Z(n238) );
  XOR U358 ( .A(A[222]), .B(n239), .Z(O[222]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[222]), .B(A[222]), .Z(n240) );
  XOR U361 ( .A(A[221]), .B(n241), .Z(O[221]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[221]), .B(A[221]), .Z(n242) );
  XOR U364 ( .A(A[220]), .B(n243), .Z(O[220]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[220]), .B(A[220]), .Z(n244) );
  XOR U367 ( .A(A[21]), .B(n245), .Z(O[21]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[21]), .B(A[21]), .Z(n246) );
  XOR U370 ( .A(A[219]), .B(n247), .Z(O[219]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[219]), .B(A[219]), .Z(n248) );
  XOR U373 ( .A(A[218]), .B(n249), .Z(O[218]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[218]), .B(A[218]), .Z(n250) );
  XOR U376 ( .A(A[217]), .B(n251), .Z(O[217]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[217]), .B(A[217]), .Z(n252) );
  XOR U379 ( .A(A[216]), .B(n253), .Z(O[216]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[216]), .B(A[216]), .Z(n254) );
  XOR U382 ( .A(A[215]), .B(n255), .Z(O[215]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[215]), .B(A[215]), .Z(n256) );
  XOR U385 ( .A(A[214]), .B(n257), .Z(O[214]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[214]), .B(A[214]), .Z(n258) );
  XOR U388 ( .A(A[213]), .B(n259), .Z(O[213]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[213]), .B(A[213]), .Z(n260) );
  XOR U391 ( .A(A[212]), .B(n261), .Z(O[212]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[212]), .B(A[212]), .Z(n262) );
  XOR U394 ( .A(A[211]), .B(n263), .Z(O[211]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[211]), .B(A[211]), .Z(n264) );
  XOR U397 ( .A(A[210]), .B(n265), .Z(O[210]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[210]), .B(A[210]), .Z(n266) );
  XOR U400 ( .A(A[20]), .B(n267), .Z(O[20]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[20]), .B(A[20]), .Z(n268) );
  XOR U403 ( .A(A[209]), .B(n269), .Z(O[209]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[209]), .B(A[209]), .Z(n270) );
  XOR U406 ( .A(A[208]), .B(n271), .Z(O[208]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[208]), .B(A[208]), .Z(n272) );
  XOR U409 ( .A(A[207]), .B(n273), .Z(O[207]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[207]), .B(A[207]), .Z(n274) );
  XOR U412 ( .A(A[206]), .B(n275), .Z(O[206]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[206]), .B(A[206]), .Z(n276) );
  XOR U415 ( .A(A[205]), .B(n277), .Z(O[205]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[205]), .B(A[205]), .Z(n278) );
  XOR U418 ( .A(A[204]), .B(n279), .Z(O[204]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[204]), .B(A[204]), .Z(n280) );
  XOR U421 ( .A(A[203]), .B(n281), .Z(O[203]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[203]), .B(A[203]), .Z(n282) );
  XOR U424 ( .A(A[202]), .B(n283), .Z(O[202]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[202]), .B(A[202]), .Z(n284) );
  XOR U427 ( .A(A[201]), .B(n285), .Z(O[201]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[201]), .B(A[201]), .Z(n286) );
  XOR U430 ( .A(A[200]), .B(n287), .Z(O[200]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[200]), .B(A[200]), .Z(n288) );
  XOR U433 ( .A(A[1]), .B(n289), .Z(O[1]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[1]), .B(A[1]), .Z(n290) );
  XOR U436 ( .A(A[19]), .B(n291), .Z(O[19]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[19]), .B(A[19]), .Z(n292) );
  XOR U439 ( .A(A[199]), .B(n293), .Z(O[199]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[199]), .B(A[199]), .Z(n294) );
  XOR U442 ( .A(A[198]), .B(n295), .Z(O[198]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[198]), .B(A[198]), .Z(n296) );
  XOR U445 ( .A(A[197]), .B(n297), .Z(O[197]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[197]), .B(A[197]), .Z(n298) );
  XOR U448 ( .A(A[196]), .B(n299), .Z(O[196]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[196]), .B(A[196]), .Z(n300) );
  XOR U451 ( .A(A[195]), .B(n301), .Z(O[195]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[195]), .B(A[195]), .Z(n302) );
  XOR U454 ( .A(A[194]), .B(n303), .Z(O[194]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[194]), .B(A[194]), .Z(n304) );
  XOR U457 ( .A(A[193]), .B(n305), .Z(O[193]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[193]), .B(A[193]), .Z(n306) );
  XOR U460 ( .A(A[192]), .B(n307), .Z(O[192]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[192]), .B(A[192]), .Z(n308) );
  XOR U463 ( .A(A[191]), .B(n309), .Z(O[191]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[191]), .B(A[191]), .Z(n310) );
  XOR U466 ( .A(A[190]), .B(n311), .Z(O[190]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[190]), .B(A[190]), .Z(n312) );
  XOR U469 ( .A(A[18]), .B(n313), .Z(O[18]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[18]), .B(A[18]), .Z(n314) );
  XOR U472 ( .A(A[189]), .B(n315), .Z(O[189]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[189]), .B(A[189]), .Z(n316) );
  XOR U475 ( .A(A[188]), .B(n317), .Z(O[188]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[188]), .B(A[188]), .Z(n318) );
  XOR U478 ( .A(A[187]), .B(n319), .Z(O[187]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[187]), .B(A[187]), .Z(n320) );
  XOR U481 ( .A(A[186]), .B(n321), .Z(O[186]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[186]), .B(A[186]), .Z(n322) );
  XOR U484 ( .A(A[185]), .B(n323), .Z(O[185]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[185]), .B(A[185]), .Z(n324) );
  XOR U487 ( .A(A[184]), .B(n325), .Z(O[184]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[184]), .B(A[184]), .Z(n326) );
  XOR U490 ( .A(A[183]), .B(n327), .Z(O[183]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[183]), .B(A[183]), .Z(n328) );
  XOR U493 ( .A(A[182]), .B(n329), .Z(O[182]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[182]), .B(A[182]), .Z(n330) );
  XOR U496 ( .A(A[181]), .B(n331), .Z(O[181]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[181]), .B(A[181]), .Z(n332) );
  XOR U499 ( .A(A[180]), .B(n333), .Z(O[180]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[180]), .B(A[180]), .Z(n334) );
  XOR U502 ( .A(A[17]), .B(n335), .Z(O[17]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[17]), .B(A[17]), .Z(n336) );
  XOR U505 ( .A(A[179]), .B(n337), .Z(O[179]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[179]), .B(A[179]), .Z(n338) );
  XOR U508 ( .A(A[178]), .B(n339), .Z(O[178]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[178]), .B(A[178]), .Z(n340) );
  XOR U511 ( .A(A[177]), .B(n341), .Z(O[177]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[177]), .B(A[177]), .Z(n342) );
  XOR U514 ( .A(A[176]), .B(n343), .Z(O[176]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[176]), .B(A[176]), .Z(n344) );
  XOR U517 ( .A(A[175]), .B(n345), .Z(O[175]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[175]), .B(A[175]), .Z(n346) );
  XOR U520 ( .A(A[174]), .B(n347), .Z(O[174]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[174]), .B(A[174]), .Z(n348) );
  XOR U523 ( .A(A[173]), .B(n349), .Z(O[173]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[173]), .B(A[173]), .Z(n350) );
  XOR U526 ( .A(A[172]), .B(n351), .Z(O[172]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[172]), .B(A[172]), .Z(n352) );
  XOR U529 ( .A(A[171]), .B(n353), .Z(O[171]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[171]), .B(A[171]), .Z(n354) );
  XOR U532 ( .A(A[170]), .B(n355), .Z(O[170]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[170]), .B(A[170]), .Z(n356) );
  XOR U535 ( .A(A[16]), .B(n357), .Z(O[16]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[16]), .B(A[16]), .Z(n358) );
  XOR U538 ( .A(A[169]), .B(n359), .Z(O[169]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[169]), .B(A[169]), .Z(n360) );
  XOR U541 ( .A(A[168]), .B(n361), .Z(O[168]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[168]), .B(A[168]), .Z(n362) );
  XOR U544 ( .A(A[167]), .B(n363), .Z(O[167]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[167]), .B(A[167]), .Z(n364) );
  XOR U547 ( .A(A[166]), .B(n365), .Z(O[166]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[166]), .B(A[166]), .Z(n366) );
  XOR U550 ( .A(A[165]), .B(n367), .Z(O[165]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[165]), .B(A[165]), .Z(n368) );
  XOR U553 ( .A(A[164]), .B(n369), .Z(O[164]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[164]), .B(A[164]), .Z(n370) );
  XOR U556 ( .A(A[163]), .B(n371), .Z(O[163]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[163]), .B(A[163]), .Z(n372) );
  XOR U559 ( .A(A[162]), .B(n373), .Z(O[162]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[162]), .B(A[162]), .Z(n374) );
  XOR U562 ( .A(A[161]), .B(n375), .Z(O[161]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[161]), .B(A[161]), .Z(n376) );
  XOR U565 ( .A(A[160]), .B(n377), .Z(O[160]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[160]), .B(A[160]), .Z(n378) );
  XOR U568 ( .A(A[15]), .B(n379), .Z(O[15]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[15]), .B(A[15]), .Z(n380) );
  XOR U571 ( .A(A[159]), .B(n381), .Z(O[159]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[159]), .B(A[159]), .Z(n382) );
  XOR U574 ( .A(A[158]), .B(n383), .Z(O[158]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[158]), .B(A[158]), .Z(n384) );
  XOR U577 ( .A(A[157]), .B(n385), .Z(O[157]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[157]), .B(A[157]), .Z(n386) );
  XOR U580 ( .A(A[156]), .B(n387), .Z(O[156]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[156]), .B(A[156]), .Z(n388) );
  XOR U583 ( .A(A[155]), .B(n389), .Z(O[155]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[155]), .B(A[155]), .Z(n390) );
  XOR U586 ( .A(A[154]), .B(n391), .Z(O[154]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[154]), .B(A[154]), .Z(n392) );
  XOR U589 ( .A(A[153]), .B(n393), .Z(O[153]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[153]), .B(A[153]), .Z(n394) );
  XOR U592 ( .A(A[152]), .B(n395), .Z(O[152]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[152]), .B(A[152]), .Z(n396) );
  XOR U595 ( .A(A[151]), .B(n397), .Z(O[151]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[151]), .B(A[151]), .Z(n398) );
  XOR U598 ( .A(A[150]), .B(n399), .Z(O[150]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[150]), .B(A[150]), .Z(n400) );
  XOR U601 ( .A(A[14]), .B(n401), .Z(O[14]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[14]), .B(A[14]), .Z(n402) );
  XOR U604 ( .A(A[149]), .B(n403), .Z(O[149]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[149]), .B(A[149]), .Z(n404) );
  XOR U607 ( .A(A[148]), .B(n405), .Z(O[148]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[148]), .B(A[148]), .Z(n406) );
  XOR U610 ( .A(A[147]), .B(n407), .Z(O[147]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[147]), .B(A[147]), .Z(n408) );
  XOR U613 ( .A(A[146]), .B(n409), .Z(O[146]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[146]), .B(A[146]), .Z(n410) );
  XOR U616 ( .A(A[145]), .B(n411), .Z(O[145]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[145]), .B(A[145]), .Z(n412) );
  XOR U619 ( .A(A[144]), .B(n413), .Z(O[144]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[144]), .B(A[144]), .Z(n414) );
  XOR U622 ( .A(A[143]), .B(n415), .Z(O[143]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[143]), .B(A[143]), .Z(n416) );
  XOR U625 ( .A(A[142]), .B(n417), .Z(O[142]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[142]), .B(A[142]), .Z(n418) );
  XOR U628 ( .A(A[141]), .B(n419), .Z(O[141]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[141]), .B(A[141]), .Z(n420) );
  XOR U631 ( .A(A[140]), .B(n421), .Z(O[140]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[140]), .B(A[140]), .Z(n422) );
  XOR U634 ( .A(A[13]), .B(n423), .Z(O[13]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[13]), .B(A[13]), .Z(n424) );
  XOR U637 ( .A(A[139]), .B(n425), .Z(O[139]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[139]), .B(A[139]), .Z(n426) );
  XOR U640 ( .A(A[138]), .B(n427), .Z(O[138]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[138]), .B(A[138]), .Z(n428) );
  XOR U643 ( .A(A[137]), .B(n429), .Z(O[137]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[137]), .B(A[137]), .Z(n430) );
  XOR U646 ( .A(A[136]), .B(n431), .Z(O[136]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[136]), .B(A[136]), .Z(n432) );
  XOR U649 ( .A(A[135]), .B(n433), .Z(O[135]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[135]), .B(A[135]), .Z(n434) );
  XOR U652 ( .A(A[134]), .B(n435), .Z(O[134]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[134]), .B(A[134]), .Z(n436) );
  XOR U655 ( .A(A[133]), .B(n437), .Z(O[133]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[133]), .B(A[133]), .Z(n438) );
  XOR U658 ( .A(A[132]), .B(n439), .Z(O[132]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[132]), .B(A[132]), .Z(n440) );
  XOR U661 ( .A(A[131]), .B(n441), .Z(O[131]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[131]), .B(A[131]), .Z(n442) );
  XOR U664 ( .A(A[130]), .B(n443), .Z(O[130]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[130]), .B(A[130]), .Z(n444) );
  XOR U667 ( .A(A[12]), .B(n445), .Z(O[12]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[12]), .B(A[12]), .Z(n446) );
  XOR U670 ( .A(A[129]), .B(n447), .Z(O[129]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[129]), .B(A[129]), .Z(n448) );
  XOR U673 ( .A(A[128]), .B(n449), .Z(O[128]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[128]), .B(A[128]), .Z(n450) );
  XOR U676 ( .A(A[127]), .B(n451), .Z(O[127]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[127]), .B(A[127]), .Z(n452) );
  XOR U679 ( .A(A[126]), .B(n453), .Z(O[126]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[126]), .B(A[126]), .Z(n454) );
  XOR U682 ( .A(A[125]), .B(n455), .Z(O[125]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[125]), .B(A[125]), .Z(n456) );
  XOR U685 ( .A(A[124]), .B(n457), .Z(O[124]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[124]), .B(A[124]), .Z(n458) );
  XOR U688 ( .A(A[123]), .B(n459), .Z(O[123]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[123]), .B(A[123]), .Z(n460) );
  XOR U691 ( .A(A[122]), .B(n461), .Z(O[122]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[122]), .B(A[122]), .Z(n462) );
  XOR U694 ( .A(A[121]), .B(n463), .Z(O[121]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[121]), .B(A[121]), .Z(n464) );
  XOR U697 ( .A(A[120]), .B(n465), .Z(O[120]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[120]), .B(A[120]), .Z(n466) );
  XOR U700 ( .A(A[11]), .B(n467), .Z(O[11]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[11]), .B(A[11]), .Z(n468) );
  XOR U703 ( .A(A[119]), .B(n469), .Z(O[119]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[119]), .B(A[119]), .Z(n470) );
  XOR U706 ( .A(A[118]), .B(n471), .Z(O[118]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[118]), .B(A[118]), .Z(n472) );
  XOR U709 ( .A(A[117]), .B(n473), .Z(O[117]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[117]), .B(A[117]), .Z(n474) );
  XOR U712 ( .A(A[116]), .B(n475), .Z(O[116]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[116]), .B(A[116]), .Z(n476) );
  XOR U715 ( .A(A[115]), .B(n477), .Z(O[115]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[115]), .B(A[115]), .Z(n478) );
  XOR U718 ( .A(A[114]), .B(n479), .Z(O[114]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[114]), .B(A[114]), .Z(n480) );
  XOR U721 ( .A(A[113]), .B(n481), .Z(O[113]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[113]), .B(A[113]), .Z(n482) );
  XOR U724 ( .A(A[112]), .B(n483), .Z(O[112]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[112]), .B(A[112]), .Z(n484) );
  XOR U727 ( .A(A[111]), .B(n485), .Z(O[111]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[111]), .B(A[111]), .Z(n486) );
  XOR U730 ( .A(A[110]), .B(n487), .Z(O[110]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[110]), .B(A[110]), .Z(n488) );
  XOR U733 ( .A(A[10]), .B(n489), .Z(O[10]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[10]), .B(A[10]), .Z(n490) );
  XOR U736 ( .A(A[109]), .B(n491), .Z(O[109]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[109]), .B(A[109]), .Z(n492) );
  XOR U739 ( .A(A[108]), .B(n493), .Z(O[108]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[108]), .B(A[108]), .Z(n494) );
  XOR U742 ( .A(A[107]), .B(n495), .Z(O[107]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[107]), .B(A[107]), .Z(n496) );
  XOR U745 ( .A(A[106]), .B(n497), .Z(O[106]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[106]), .B(A[106]), .Z(n498) );
  XOR U748 ( .A(A[105]), .B(n499), .Z(O[105]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[105]), .B(A[105]), .Z(n500) );
  XOR U751 ( .A(A[104]), .B(n501), .Z(O[104]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[104]), .B(A[104]), .Z(n502) );
  XOR U754 ( .A(A[103]), .B(n503), .Z(O[103]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[103]), .B(A[103]), .Z(n504) );
  XOR U757 ( .A(A[102]), .B(n505), .Z(O[102]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[102]), .B(A[102]), .Z(n506) );
  XOR U760 ( .A(A[101]), .B(n507), .Z(O[101]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[101]), .B(A[101]), .Z(n508) );
  XOR U763 ( .A(A[100]), .B(n509), .Z(O[100]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[100]), .B(A[100]), .Z(n510) );
  XOR U766 ( .A(A[0]), .B(n511), .Z(O[0]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[0]), .B(A[0]), .Z(n512) );
endmodule


module MUX_N258_0 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_0 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_1033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_1034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  ANDN U1 ( .B(CI), .A(S), .Z(CO) );
  XOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_1035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_1289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N258 ( A, B, CI, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  input CI;
  output CO;

  wire   [257:1] C;

  FA_0 \FAINST[0].FA_  ( .A(1'b0), .B(B[0]), .CI(1'b0), .S(S[0]) );
  FA_1289 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(S[1]), .CO(C[2])
         );
  FA_1288 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_1287 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_1286 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_1285 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_1284 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_1283 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_1282 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_1281 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10]) );
  FA_1280 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_1279 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_1278 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_1277 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_1276 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_1275 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_1274 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_1273 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_1272 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_1271 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_1270 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_1269 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_1268 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_1267 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_1266 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_1265 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_1264 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_1263 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_1262 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_1261 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_1260 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_1259 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_1258 \FAINST[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_1257 \FAINST[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_1256 \FAINST[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_1255 \FAINST[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_1254 \FAINST[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_1253 \FAINST[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_1252 \FAINST[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_1251 \FAINST[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_1250 \FAINST[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_1249 \FAINST[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_1248 \FAINST[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_1247 \FAINST[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_1246 \FAINST[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_1245 \FAINST[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_1244 \FAINST[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_1243 \FAINST[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_1242 \FAINST[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_1241 \FAINST[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_1240 \FAINST[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_1239 \FAINST[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_1238 \FAINST[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_1237 \FAINST[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_1236 \FAINST[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_1235 \FAINST[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_1234 \FAINST[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_1233 \FAINST[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_1232 \FAINST[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_1231 \FAINST[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_1230 \FAINST[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_1229 \FAINST[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_1228 \FAINST[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_1227 \FAINST[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_1226 \FAINST[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_1225 \FAINST[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_1224 \FAINST[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_1223 \FAINST[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_1222 \FAINST[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_1221 \FAINST[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_1220 \FAINST[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_1219 \FAINST[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_1218 \FAINST[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_1217 \FAINST[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_1216 \FAINST[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_1215 \FAINST[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_1214 \FAINST[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_1213 \FAINST[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_1212 \FAINST[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_1211 \FAINST[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_1210 \FAINST[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_1209 \FAINST[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_1208 \FAINST[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_1207 \FAINST[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_1206 \FAINST[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_1205 \FAINST[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_1204 \FAINST[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_1203 \FAINST[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_1202 \FAINST[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_1201 \FAINST[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_1200 \FAINST[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_1199 \FAINST[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_1198 \FAINST[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_1197 \FAINST[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_1196 \FAINST[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_1195 \FAINST[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_1194 \FAINST[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_1193 \FAINST[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_1192 \FAINST[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_1191 \FAINST[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_1190 \FAINST[100].FA_  ( .A(A[100]), .B(B[100]), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_1189 \FAINST[101].FA_  ( .A(A[101]), .B(B[101]), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_1188 \FAINST[102].FA_  ( .A(A[102]), .B(B[102]), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_1187 \FAINST[103].FA_  ( .A(A[103]), .B(B[103]), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_1186 \FAINST[104].FA_  ( .A(A[104]), .B(B[104]), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_1185 \FAINST[105].FA_  ( .A(A[105]), .B(B[105]), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_1184 \FAINST[106].FA_  ( .A(A[106]), .B(B[106]), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_1183 \FAINST[107].FA_  ( .A(A[107]), .B(B[107]), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_1182 \FAINST[108].FA_  ( .A(A[108]), .B(B[108]), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_1181 \FAINST[109].FA_  ( .A(A[109]), .B(B[109]), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_1180 \FAINST[110].FA_  ( .A(A[110]), .B(B[110]), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_1179 \FAINST[111].FA_  ( .A(A[111]), .B(B[111]), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_1178 \FAINST[112].FA_  ( .A(A[112]), .B(B[112]), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_1177 \FAINST[113].FA_  ( .A(A[113]), .B(B[113]), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_1176 \FAINST[114].FA_  ( .A(A[114]), .B(B[114]), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_1175 \FAINST[115].FA_  ( .A(A[115]), .B(B[115]), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_1174 \FAINST[116].FA_  ( .A(A[116]), .B(B[116]), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_1173 \FAINST[117].FA_  ( .A(A[117]), .B(B[117]), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_1172 \FAINST[118].FA_  ( .A(A[118]), .B(B[118]), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_1171 \FAINST[119].FA_  ( .A(A[119]), .B(B[119]), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_1170 \FAINST[120].FA_  ( .A(A[120]), .B(B[120]), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_1169 \FAINST[121].FA_  ( .A(A[121]), .B(B[121]), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_1168 \FAINST[122].FA_  ( .A(A[122]), .B(B[122]), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_1167 \FAINST[123].FA_  ( .A(A[123]), .B(B[123]), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_1166 \FAINST[124].FA_  ( .A(A[124]), .B(B[124]), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_1165 \FAINST[125].FA_  ( .A(A[125]), .B(B[125]), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_1164 \FAINST[126].FA_  ( .A(A[126]), .B(B[126]), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_1163 \FAINST[127].FA_  ( .A(A[127]), .B(B[127]), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_1162 \FAINST[128].FA_  ( .A(A[128]), .B(B[128]), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_1161 \FAINST[129].FA_  ( .A(A[129]), .B(B[129]), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_1160 \FAINST[130].FA_  ( .A(A[130]), .B(B[130]), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_1159 \FAINST[131].FA_  ( .A(A[131]), .B(B[131]), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_1158 \FAINST[132].FA_  ( .A(A[132]), .B(B[132]), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_1157 \FAINST[133].FA_  ( .A(A[133]), .B(B[133]), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_1156 \FAINST[134].FA_  ( .A(A[134]), .B(B[134]), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_1155 \FAINST[135].FA_  ( .A(A[135]), .B(B[135]), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_1154 \FAINST[136].FA_  ( .A(A[136]), .B(B[136]), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_1153 \FAINST[137].FA_  ( .A(A[137]), .B(B[137]), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_1152 \FAINST[138].FA_  ( .A(A[138]), .B(B[138]), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_1151 \FAINST[139].FA_  ( .A(A[139]), .B(B[139]), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_1150 \FAINST[140].FA_  ( .A(A[140]), .B(B[140]), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_1149 \FAINST[141].FA_  ( .A(A[141]), .B(B[141]), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_1148 \FAINST[142].FA_  ( .A(A[142]), .B(B[142]), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_1147 \FAINST[143].FA_  ( .A(A[143]), .B(B[143]), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_1146 \FAINST[144].FA_  ( .A(A[144]), .B(B[144]), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_1145 \FAINST[145].FA_  ( .A(A[145]), .B(B[145]), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_1144 \FAINST[146].FA_  ( .A(A[146]), .B(B[146]), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_1143 \FAINST[147].FA_  ( .A(A[147]), .B(B[147]), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_1142 \FAINST[148].FA_  ( .A(A[148]), .B(B[148]), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_1141 \FAINST[149].FA_  ( .A(A[149]), .B(B[149]), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_1140 \FAINST[150].FA_  ( .A(A[150]), .B(B[150]), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_1139 \FAINST[151].FA_  ( .A(A[151]), .B(B[151]), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_1138 \FAINST[152].FA_  ( .A(A[152]), .B(B[152]), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_1137 \FAINST[153].FA_  ( .A(A[153]), .B(B[153]), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_1136 \FAINST[154].FA_  ( .A(A[154]), .B(B[154]), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_1135 \FAINST[155].FA_  ( .A(A[155]), .B(B[155]), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_1134 \FAINST[156].FA_  ( .A(A[156]), .B(B[156]), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_1133 \FAINST[157].FA_  ( .A(A[157]), .B(B[157]), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_1132 \FAINST[158].FA_  ( .A(A[158]), .B(B[158]), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_1131 \FAINST[159].FA_  ( .A(A[159]), .B(B[159]), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_1130 \FAINST[160].FA_  ( .A(A[160]), .B(B[160]), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_1129 \FAINST[161].FA_  ( .A(A[161]), .B(B[161]), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_1128 \FAINST[162].FA_  ( .A(A[162]), .B(B[162]), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_1127 \FAINST[163].FA_  ( .A(A[163]), .B(B[163]), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_1126 \FAINST[164].FA_  ( .A(A[164]), .B(B[164]), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_1125 \FAINST[165].FA_  ( .A(A[165]), .B(B[165]), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_1124 \FAINST[166].FA_  ( .A(A[166]), .B(B[166]), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_1123 \FAINST[167].FA_  ( .A(A[167]), .B(B[167]), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_1122 \FAINST[168].FA_  ( .A(A[168]), .B(B[168]), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_1121 \FAINST[169].FA_  ( .A(A[169]), .B(B[169]), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_1120 \FAINST[170].FA_  ( .A(A[170]), .B(B[170]), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_1119 \FAINST[171].FA_  ( .A(A[171]), .B(B[171]), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_1118 \FAINST[172].FA_  ( .A(A[172]), .B(B[172]), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_1117 \FAINST[173].FA_  ( .A(A[173]), .B(B[173]), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_1116 \FAINST[174].FA_  ( .A(A[174]), .B(B[174]), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_1115 \FAINST[175].FA_  ( .A(A[175]), .B(B[175]), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_1114 \FAINST[176].FA_  ( .A(A[176]), .B(B[176]), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_1113 \FAINST[177].FA_  ( .A(A[177]), .B(B[177]), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_1112 \FAINST[178].FA_  ( .A(A[178]), .B(B[178]), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_1111 \FAINST[179].FA_  ( .A(A[179]), .B(B[179]), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_1110 \FAINST[180].FA_  ( .A(A[180]), .B(B[180]), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_1109 \FAINST[181].FA_  ( .A(A[181]), .B(B[181]), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_1108 \FAINST[182].FA_  ( .A(A[182]), .B(B[182]), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_1107 \FAINST[183].FA_  ( .A(A[183]), .B(B[183]), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_1106 \FAINST[184].FA_  ( .A(A[184]), .B(B[184]), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_1105 \FAINST[185].FA_  ( .A(A[185]), .B(B[185]), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_1104 \FAINST[186].FA_  ( .A(A[186]), .B(B[186]), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_1103 \FAINST[187].FA_  ( .A(A[187]), .B(B[187]), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_1102 \FAINST[188].FA_  ( .A(A[188]), .B(B[188]), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_1101 \FAINST[189].FA_  ( .A(A[189]), .B(B[189]), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_1100 \FAINST[190].FA_  ( .A(A[190]), .B(B[190]), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_1099 \FAINST[191].FA_  ( .A(A[191]), .B(B[191]), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_1098 \FAINST[192].FA_  ( .A(A[192]), .B(B[192]), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_1097 \FAINST[193].FA_  ( .A(A[193]), .B(B[193]), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_1096 \FAINST[194].FA_  ( .A(A[194]), .B(B[194]), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_1095 \FAINST[195].FA_  ( .A(A[195]), .B(B[195]), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_1094 \FAINST[196].FA_  ( .A(A[196]), .B(B[196]), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_1093 \FAINST[197].FA_  ( .A(A[197]), .B(B[197]), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_1092 \FAINST[198].FA_  ( .A(A[198]), .B(B[198]), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_1091 \FAINST[199].FA_  ( .A(A[199]), .B(B[199]), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_1090 \FAINST[200].FA_  ( .A(A[200]), .B(B[200]), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_1089 \FAINST[201].FA_  ( .A(A[201]), .B(B[201]), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_1088 \FAINST[202].FA_  ( .A(A[202]), .B(B[202]), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_1087 \FAINST[203].FA_  ( .A(A[203]), .B(B[203]), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_1086 \FAINST[204].FA_  ( .A(A[204]), .B(B[204]), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_1085 \FAINST[205].FA_  ( .A(A[205]), .B(B[205]), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_1084 \FAINST[206].FA_  ( .A(A[206]), .B(B[206]), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_1083 \FAINST[207].FA_  ( .A(A[207]), .B(B[207]), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_1082 \FAINST[208].FA_  ( .A(A[208]), .B(B[208]), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_1081 \FAINST[209].FA_  ( .A(A[209]), .B(B[209]), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_1080 \FAINST[210].FA_  ( .A(A[210]), .B(B[210]), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_1079 \FAINST[211].FA_  ( .A(A[211]), .B(B[211]), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_1078 \FAINST[212].FA_  ( .A(A[212]), .B(B[212]), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_1077 \FAINST[213].FA_  ( .A(A[213]), .B(B[213]), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_1076 \FAINST[214].FA_  ( .A(A[214]), .B(B[214]), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_1075 \FAINST[215].FA_  ( .A(A[215]), .B(B[215]), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_1074 \FAINST[216].FA_  ( .A(A[216]), .B(B[216]), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_1073 \FAINST[217].FA_  ( .A(A[217]), .B(B[217]), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_1072 \FAINST[218].FA_  ( .A(A[218]), .B(B[218]), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_1071 \FAINST[219].FA_  ( .A(A[219]), .B(B[219]), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_1070 \FAINST[220].FA_  ( .A(A[220]), .B(B[220]), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_1069 \FAINST[221].FA_  ( .A(A[221]), .B(B[221]), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_1068 \FAINST[222].FA_  ( .A(A[222]), .B(B[222]), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_1067 \FAINST[223].FA_  ( .A(A[223]), .B(B[223]), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_1066 \FAINST[224].FA_  ( .A(A[224]), .B(B[224]), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_1065 \FAINST[225].FA_  ( .A(A[225]), .B(B[225]), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_1064 \FAINST[226].FA_  ( .A(A[226]), .B(B[226]), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_1063 \FAINST[227].FA_  ( .A(A[227]), .B(B[227]), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_1062 \FAINST[228].FA_  ( .A(A[228]), .B(B[228]), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_1061 \FAINST[229].FA_  ( .A(A[229]), .B(B[229]), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_1060 \FAINST[230].FA_  ( .A(A[230]), .B(B[230]), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_1059 \FAINST[231].FA_  ( .A(A[231]), .B(B[231]), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_1058 \FAINST[232].FA_  ( .A(A[232]), .B(B[232]), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_1057 \FAINST[233].FA_  ( .A(A[233]), .B(B[233]), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_1056 \FAINST[234].FA_  ( .A(A[234]), .B(B[234]), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_1055 \FAINST[235].FA_  ( .A(A[235]), .B(B[235]), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_1054 \FAINST[236].FA_  ( .A(A[236]), .B(B[236]), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_1053 \FAINST[237].FA_  ( .A(A[237]), .B(B[237]), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_1052 \FAINST[238].FA_  ( .A(A[238]), .B(B[238]), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_1051 \FAINST[239].FA_  ( .A(A[239]), .B(B[239]), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_1050 \FAINST[240].FA_  ( .A(A[240]), .B(B[240]), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_1049 \FAINST[241].FA_  ( .A(A[241]), .B(B[241]), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_1048 \FAINST[242].FA_  ( .A(A[242]), .B(B[242]), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_1047 \FAINST[243].FA_  ( .A(A[243]), .B(B[243]), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_1046 \FAINST[244].FA_  ( .A(A[244]), .B(B[244]), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_1045 \FAINST[245].FA_  ( .A(A[245]), .B(B[245]), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_1044 \FAINST[246].FA_  ( .A(A[246]), .B(B[246]), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_1043 \FAINST[247].FA_  ( .A(A[247]), .B(B[247]), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_1042 \FAINST[248].FA_  ( .A(A[248]), .B(B[248]), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_1041 \FAINST[249].FA_  ( .A(A[249]), .B(B[249]), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_1040 \FAINST[250].FA_  ( .A(A[250]), .B(B[250]), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_1039 \FAINST[251].FA_  ( .A(A[251]), .B(B[251]), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_1038 \FAINST[252].FA_  ( .A(A[252]), .B(B[252]), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_1037 \FAINST[253].FA_  ( .A(A[253]), .B(B[253]), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_1036 \FAINST[254].FA_  ( .A(A[254]), .B(B[254]), .CI(C[254]), .S(S[254]), 
        .CO(C[255]) );
  FA_1035 \FAINST[255].FA_  ( .A(A[255]), .B(B[255]), .CI(C[255]), .S(S[255]), 
        .CO(C[256]) );
  FA_1034 \FAINST[256].FA_  ( .A(A[256]), .B(1'b0), .CI(C[256]), .S(S[256]), 
        .CO(C[257]) );
  FA_1033 \FAINST[257].FA_  ( .A(A[257]), .B(1'b0), .CI(C[257]), .S(S[257]) );
endmodule


module FA_775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_1032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N258_0 ( A, B, O );
  input [257:0] A;
  input [257:0] B;
  output O;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258;
  wire   [257:1] C;

  FA_1032 \FAINST[0].FA_  ( .A(A[0]), .B(n258), .CI(1'b1), .CO(C[1]) );
  FA_1031 \FAINST[1].FA_  ( .A(A[1]), .B(n257), .CI(C[1]), .CO(C[2]) );
  FA_1030 \FAINST[2].FA_  ( .A(A[2]), .B(n256), .CI(C[2]), .CO(C[3]) );
  FA_1029 \FAINST[3].FA_  ( .A(A[3]), .B(n255), .CI(C[3]), .CO(C[4]) );
  FA_1028 \FAINST[4].FA_  ( .A(A[4]), .B(n254), .CI(C[4]), .CO(C[5]) );
  FA_1027 \FAINST[5].FA_  ( .A(A[5]), .B(n253), .CI(C[5]), .CO(C[6]) );
  FA_1026 \FAINST[6].FA_  ( .A(A[6]), .B(n252), .CI(C[6]), .CO(C[7]) );
  FA_1025 \FAINST[7].FA_  ( .A(A[7]), .B(n251), .CI(C[7]), .CO(C[8]) );
  FA_1024 \FAINST[8].FA_  ( .A(A[8]), .B(n250), .CI(C[8]), .CO(C[9]) );
  FA_1023 \FAINST[9].FA_  ( .A(A[9]), .B(n249), .CI(C[9]), .CO(C[10]) );
  FA_1022 \FAINST[10].FA_  ( .A(A[10]), .B(n248), .CI(C[10]), .CO(C[11]) );
  FA_1021 \FAINST[11].FA_  ( .A(A[11]), .B(n247), .CI(C[11]), .CO(C[12]) );
  FA_1020 \FAINST[12].FA_  ( .A(A[12]), .B(n246), .CI(C[12]), .CO(C[13]) );
  FA_1019 \FAINST[13].FA_  ( .A(A[13]), .B(n245), .CI(C[13]), .CO(C[14]) );
  FA_1018 \FAINST[14].FA_  ( .A(A[14]), .B(n244), .CI(C[14]), .CO(C[15]) );
  FA_1017 \FAINST[15].FA_  ( .A(A[15]), .B(n243), .CI(C[15]), .CO(C[16]) );
  FA_1016 \FAINST[16].FA_  ( .A(A[16]), .B(n242), .CI(C[16]), .CO(C[17]) );
  FA_1015 \FAINST[17].FA_  ( .A(A[17]), .B(n241), .CI(C[17]), .CO(C[18]) );
  FA_1014 \FAINST[18].FA_  ( .A(A[18]), .B(n240), .CI(C[18]), .CO(C[19]) );
  FA_1013 \FAINST[19].FA_  ( .A(A[19]), .B(n239), .CI(C[19]), .CO(C[20]) );
  FA_1012 \FAINST[20].FA_  ( .A(A[20]), .B(n238), .CI(C[20]), .CO(C[21]) );
  FA_1011 \FAINST[21].FA_  ( .A(A[21]), .B(n237), .CI(C[21]), .CO(C[22]) );
  FA_1010 \FAINST[22].FA_  ( .A(A[22]), .B(n236), .CI(C[22]), .CO(C[23]) );
  FA_1009 \FAINST[23].FA_  ( .A(A[23]), .B(n235), .CI(C[23]), .CO(C[24]) );
  FA_1008 \FAINST[24].FA_  ( .A(A[24]), .B(n234), .CI(C[24]), .CO(C[25]) );
  FA_1007 \FAINST[25].FA_  ( .A(A[25]), .B(n233), .CI(C[25]), .CO(C[26]) );
  FA_1006 \FAINST[26].FA_  ( .A(A[26]), .B(n232), .CI(C[26]), .CO(C[27]) );
  FA_1005 \FAINST[27].FA_  ( .A(A[27]), .B(n231), .CI(C[27]), .CO(C[28]) );
  FA_1004 \FAINST[28].FA_  ( .A(A[28]), .B(n230), .CI(C[28]), .CO(C[29]) );
  FA_1003 \FAINST[29].FA_  ( .A(A[29]), .B(n229), .CI(C[29]), .CO(C[30]) );
  FA_1002 \FAINST[30].FA_  ( .A(A[30]), .B(n228), .CI(C[30]), .CO(C[31]) );
  FA_1001 \FAINST[31].FA_  ( .A(A[31]), .B(n227), .CI(C[31]), .CO(C[32]) );
  FA_1000 \FAINST[32].FA_  ( .A(A[32]), .B(n226), .CI(C[32]), .CO(C[33]) );
  FA_999 \FAINST[33].FA_  ( .A(A[33]), .B(n225), .CI(C[33]), .CO(C[34]) );
  FA_998 \FAINST[34].FA_  ( .A(A[34]), .B(n224), .CI(C[34]), .CO(C[35]) );
  FA_997 \FAINST[35].FA_  ( .A(A[35]), .B(n223), .CI(C[35]), .CO(C[36]) );
  FA_996 \FAINST[36].FA_  ( .A(A[36]), .B(n222), .CI(C[36]), .CO(C[37]) );
  FA_995 \FAINST[37].FA_  ( .A(A[37]), .B(n221), .CI(C[37]), .CO(C[38]) );
  FA_994 \FAINST[38].FA_  ( .A(A[38]), .B(n220), .CI(C[38]), .CO(C[39]) );
  FA_993 \FAINST[39].FA_  ( .A(A[39]), .B(n219), .CI(C[39]), .CO(C[40]) );
  FA_992 \FAINST[40].FA_  ( .A(A[40]), .B(n218), .CI(C[40]), .CO(C[41]) );
  FA_991 \FAINST[41].FA_  ( .A(A[41]), .B(n217), .CI(C[41]), .CO(C[42]) );
  FA_990 \FAINST[42].FA_  ( .A(A[42]), .B(n216), .CI(C[42]), .CO(C[43]) );
  FA_989 \FAINST[43].FA_  ( .A(A[43]), .B(n215), .CI(C[43]), .CO(C[44]) );
  FA_988 \FAINST[44].FA_  ( .A(A[44]), .B(n214), .CI(C[44]), .CO(C[45]) );
  FA_987 \FAINST[45].FA_  ( .A(A[45]), .B(n213), .CI(C[45]), .CO(C[46]) );
  FA_986 \FAINST[46].FA_  ( .A(A[46]), .B(n212), .CI(C[46]), .CO(C[47]) );
  FA_985 \FAINST[47].FA_  ( .A(A[47]), .B(n211), .CI(C[47]), .CO(C[48]) );
  FA_984 \FAINST[48].FA_  ( .A(A[48]), .B(n210), .CI(C[48]), .CO(C[49]) );
  FA_983 \FAINST[49].FA_  ( .A(A[49]), .B(n209), .CI(C[49]), .CO(C[50]) );
  FA_982 \FAINST[50].FA_  ( .A(A[50]), .B(n208), .CI(C[50]), .CO(C[51]) );
  FA_981 \FAINST[51].FA_  ( .A(A[51]), .B(n207), .CI(C[51]), .CO(C[52]) );
  FA_980 \FAINST[52].FA_  ( .A(A[52]), .B(n206), .CI(C[52]), .CO(C[53]) );
  FA_979 \FAINST[53].FA_  ( .A(A[53]), .B(n205), .CI(C[53]), .CO(C[54]) );
  FA_978 \FAINST[54].FA_  ( .A(A[54]), .B(n204), .CI(C[54]), .CO(C[55]) );
  FA_977 \FAINST[55].FA_  ( .A(A[55]), .B(n203), .CI(C[55]), .CO(C[56]) );
  FA_976 \FAINST[56].FA_  ( .A(A[56]), .B(n202), .CI(C[56]), .CO(C[57]) );
  FA_975 \FAINST[57].FA_  ( .A(A[57]), .B(n201), .CI(C[57]), .CO(C[58]) );
  FA_974 \FAINST[58].FA_  ( .A(A[58]), .B(n200), .CI(C[58]), .CO(C[59]) );
  FA_973 \FAINST[59].FA_  ( .A(A[59]), .B(n199), .CI(C[59]), .CO(C[60]) );
  FA_972 \FAINST[60].FA_  ( .A(A[60]), .B(n198), .CI(C[60]), .CO(C[61]) );
  FA_971 \FAINST[61].FA_  ( .A(A[61]), .B(n197), .CI(C[61]), .CO(C[62]) );
  FA_970 \FAINST[62].FA_  ( .A(A[62]), .B(n196), .CI(C[62]), .CO(C[63]) );
  FA_969 \FAINST[63].FA_  ( .A(A[63]), .B(n195), .CI(C[63]), .CO(C[64]) );
  FA_968 \FAINST[64].FA_  ( .A(A[64]), .B(n194), .CI(C[64]), .CO(C[65]) );
  FA_967 \FAINST[65].FA_  ( .A(A[65]), .B(n193), .CI(C[65]), .CO(C[66]) );
  FA_966 \FAINST[66].FA_  ( .A(A[66]), .B(n192), .CI(C[66]), .CO(C[67]) );
  FA_965 \FAINST[67].FA_  ( .A(A[67]), .B(n191), .CI(C[67]), .CO(C[68]) );
  FA_964 \FAINST[68].FA_  ( .A(A[68]), .B(n190), .CI(C[68]), .CO(C[69]) );
  FA_963 \FAINST[69].FA_  ( .A(A[69]), .B(n189), .CI(C[69]), .CO(C[70]) );
  FA_962 \FAINST[70].FA_  ( .A(A[70]), .B(n188), .CI(C[70]), .CO(C[71]) );
  FA_961 \FAINST[71].FA_  ( .A(A[71]), .B(n187), .CI(C[71]), .CO(C[72]) );
  FA_960 \FAINST[72].FA_  ( .A(A[72]), .B(n186), .CI(C[72]), .CO(C[73]) );
  FA_959 \FAINST[73].FA_  ( .A(A[73]), .B(n185), .CI(C[73]), .CO(C[74]) );
  FA_958 \FAINST[74].FA_  ( .A(A[74]), .B(n184), .CI(C[74]), .CO(C[75]) );
  FA_957 \FAINST[75].FA_  ( .A(A[75]), .B(n183), .CI(C[75]), .CO(C[76]) );
  FA_956 \FAINST[76].FA_  ( .A(A[76]), .B(n182), .CI(C[76]), .CO(C[77]) );
  FA_955 \FAINST[77].FA_  ( .A(A[77]), .B(n181), .CI(C[77]), .CO(C[78]) );
  FA_954 \FAINST[78].FA_  ( .A(A[78]), .B(n180), .CI(C[78]), .CO(C[79]) );
  FA_953 \FAINST[79].FA_  ( .A(A[79]), .B(n179), .CI(C[79]), .CO(C[80]) );
  FA_952 \FAINST[80].FA_  ( .A(A[80]), .B(n178), .CI(C[80]), .CO(C[81]) );
  FA_951 \FAINST[81].FA_  ( .A(A[81]), .B(n177), .CI(C[81]), .CO(C[82]) );
  FA_950 \FAINST[82].FA_  ( .A(A[82]), .B(n176), .CI(C[82]), .CO(C[83]) );
  FA_949 \FAINST[83].FA_  ( .A(A[83]), .B(n175), .CI(C[83]), .CO(C[84]) );
  FA_948 \FAINST[84].FA_  ( .A(A[84]), .B(n174), .CI(C[84]), .CO(C[85]) );
  FA_947 \FAINST[85].FA_  ( .A(A[85]), .B(n173), .CI(C[85]), .CO(C[86]) );
  FA_946 \FAINST[86].FA_  ( .A(A[86]), .B(n172), .CI(C[86]), .CO(C[87]) );
  FA_945 \FAINST[87].FA_  ( .A(A[87]), .B(n171), .CI(C[87]), .CO(C[88]) );
  FA_944 \FAINST[88].FA_  ( .A(A[88]), .B(n170), .CI(C[88]), .CO(C[89]) );
  FA_943 \FAINST[89].FA_  ( .A(A[89]), .B(n169), .CI(C[89]), .CO(C[90]) );
  FA_942 \FAINST[90].FA_  ( .A(A[90]), .B(n168), .CI(C[90]), .CO(C[91]) );
  FA_941 \FAINST[91].FA_  ( .A(A[91]), .B(n167), .CI(C[91]), .CO(C[92]) );
  FA_940 \FAINST[92].FA_  ( .A(A[92]), .B(n166), .CI(C[92]), .CO(C[93]) );
  FA_939 \FAINST[93].FA_  ( .A(A[93]), .B(n165), .CI(C[93]), .CO(C[94]) );
  FA_938 \FAINST[94].FA_  ( .A(A[94]), .B(n164), .CI(C[94]), .CO(C[95]) );
  FA_937 \FAINST[95].FA_  ( .A(A[95]), .B(n163), .CI(C[95]), .CO(C[96]) );
  FA_936 \FAINST[96].FA_  ( .A(A[96]), .B(n162), .CI(C[96]), .CO(C[97]) );
  FA_935 \FAINST[97].FA_  ( .A(A[97]), .B(n161), .CI(C[97]), .CO(C[98]) );
  FA_934 \FAINST[98].FA_  ( .A(A[98]), .B(n160), .CI(C[98]), .CO(C[99]) );
  FA_933 \FAINST[99].FA_  ( .A(A[99]), .B(n159), .CI(C[99]), .CO(C[100]) );
  FA_932 \FAINST[100].FA_  ( .A(A[100]), .B(n158), .CI(C[100]), .CO(C[101]) );
  FA_931 \FAINST[101].FA_  ( .A(A[101]), .B(n157), .CI(C[101]), .CO(C[102]) );
  FA_930 \FAINST[102].FA_  ( .A(A[102]), .B(n156), .CI(C[102]), .CO(C[103]) );
  FA_929 \FAINST[103].FA_  ( .A(A[103]), .B(n155), .CI(C[103]), .CO(C[104]) );
  FA_928 \FAINST[104].FA_  ( .A(A[104]), .B(n154), .CI(C[104]), .CO(C[105]) );
  FA_927 \FAINST[105].FA_  ( .A(A[105]), .B(n153), .CI(C[105]), .CO(C[106]) );
  FA_926 \FAINST[106].FA_  ( .A(A[106]), .B(n152), .CI(C[106]), .CO(C[107]) );
  FA_925 \FAINST[107].FA_  ( .A(A[107]), .B(n151), .CI(C[107]), .CO(C[108]) );
  FA_924 \FAINST[108].FA_  ( .A(A[108]), .B(n150), .CI(C[108]), .CO(C[109]) );
  FA_923 \FAINST[109].FA_  ( .A(A[109]), .B(n149), .CI(C[109]), .CO(C[110]) );
  FA_922 \FAINST[110].FA_  ( .A(A[110]), .B(n148), .CI(C[110]), .CO(C[111]) );
  FA_921 \FAINST[111].FA_  ( .A(A[111]), .B(n147), .CI(C[111]), .CO(C[112]) );
  FA_920 \FAINST[112].FA_  ( .A(A[112]), .B(n146), .CI(C[112]), .CO(C[113]) );
  FA_919 \FAINST[113].FA_  ( .A(A[113]), .B(n145), .CI(C[113]), .CO(C[114]) );
  FA_918 \FAINST[114].FA_  ( .A(A[114]), .B(n144), .CI(C[114]), .CO(C[115]) );
  FA_917 \FAINST[115].FA_  ( .A(A[115]), .B(n143), .CI(C[115]), .CO(C[116]) );
  FA_916 \FAINST[116].FA_  ( .A(A[116]), .B(n142), .CI(C[116]), .CO(C[117]) );
  FA_915 \FAINST[117].FA_  ( .A(A[117]), .B(n141), .CI(C[117]), .CO(C[118]) );
  FA_914 \FAINST[118].FA_  ( .A(A[118]), .B(n140), .CI(C[118]), .CO(C[119]) );
  FA_913 \FAINST[119].FA_  ( .A(A[119]), .B(n139), .CI(C[119]), .CO(C[120]) );
  FA_912 \FAINST[120].FA_  ( .A(A[120]), .B(n138), .CI(C[120]), .CO(C[121]) );
  FA_911 \FAINST[121].FA_  ( .A(A[121]), .B(n137), .CI(C[121]), .CO(C[122]) );
  FA_910 \FAINST[122].FA_  ( .A(A[122]), .B(n136), .CI(C[122]), .CO(C[123]) );
  FA_909 \FAINST[123].FA_  ( .A(A[123]), .B(n135), .CI(C[123]), .CO(C[124]) );
  FA_908 \FAINST[124].FA_  ( .A(A[124]), .B(n134), .CI(C[124]), .CO(C[125]) );
  FA_907 \FAINST[125].FA_  ( .A(A[125]), .B(n133), .CI(C[125]), .CO(C[126]) );
  FA_906 \FAINST[126].FA_  ( .A(A[126]), .B(n132), .CI(C[126]), .CO(C[127]) );
  FA_905 \FAINST[127].FA_  ( .A(A[127]), .B(n131), .CI(C[127]), .CO(C[128]) );
  FA_904 \FAINST[128].FA_  ( .A(A[128]), .B(n130), .CI(C[128]), .CO(C[129]) );
  FA_903 \FAINST[129].FA_  ( .A(A[129]), .B(n129), .CI(C[129]), .CO(C[130]) );
  FA_902 \FAINST[130].FA_  ( .A(A[130]), .B(n128), .CI(C[130]), .CO(C[131]) );
  FA_901 \FAINST[131].FA_  ( .A(A[131]), .B(n127), .CI(C[131]), .CO(C[132]) );
  FA_900 \FAINST[132].FA_  ( .A(A[132]), .B(n126), .CI(C[132]), .CO(C[133]) );
  FA_899 \FAINST[133].FA_  ( .A(A[133]), .B(n125), .CI(C[133]), .CO(C[134]) );
  FA_898 \FAINST[134].FA_  ( .A(A[134]), .B(n124), .CI(C[134]), .CO(C[135]) );
  FA_897 \FAINST[135].FA_  ( .A(A[135]), .B(n123), .CI(C[135]), .CO(C[136]) );
  FA_896 \FAINST[136].FA_  ( .A(A[136]), .B(n122), .CI(C[136]), .CO(C[137]) );
  FA_895 \FAINST[137].FA_  ( .A(A[137]), .B(n121), .CI(C[137]), .CO(C[138]) );
  FA_894 \FAINST[138].FA_  ( .A(A[138]), .B(n120), .CI(C[138]), .CO(C[139]) );
  FA_893 \FAINST[139].FA_  ( .A(A[139]), .B(n119), .CI(C[139]), .CO(C[140]) );
  FA_892 \FAINST[140].FA_  ( .A(A[140]), .B(n118), .CI(C[140]), .CO(C[141]) );
  FA_891 \FAINST[141].FA_  ( .A(A[141]), .B(n117), .CI(C[141]), .CO(C[142]) );
  FA_890 \FAINST[142].FA_  ( .A(A[142]), .B(n116), .CI(C[142]), .CO(C[143]) );
  FA_889 \FAINST[143].FA_  ( .A(A[143]), .B(n115), .CI(C[143]), .CO(C[144]) );
  FA_888 \FAINST[144].FA_  ( .A(A[144]), .B(n114), .CI(C[144]), .CO(C[145]) );
  FA_887 \FAINST[145].FA_  ( .A(A[145]), .B(n113), .CI(C[145]), .CO(C[146]) );
  FA_886 \FAINST[146].FA_  ( .A(A[146]), .B(n112), .CI(C[146]), .CO(C[147]) );
  FA_885 \FAINST[147].FA_  ( .A(A[147]), .B(n111), .CI(C[147]), .CO(C[148]) );
  FA_884 \FAINST[148].FA_  ( .A(A[148]), .B(n110), .CI(C[148]), .CO(C[149]) );
  FA_883 \FAINST[149].FA_  ( .A(A[149]), .B(n109), .CI(C[149]), .CO(C[150]) );
  FA_882 \FAINST[150].FA_  ( .A(A[150]), .B(n108), .CI(C[150]), .CO(C[151]) );
  FA_881 \FAINST[151].FA_  ( .A(A[151]), .B(n107), .CI(C[151]), .CO(C[152]) );
  FA_880 \FAINST[152].FA_  ( .A(A[152]), .B(n106), .CI(C[152]), .CO(C[153]) );
  FA_879 \FAINST[153].FA_  ( .A(A[153]), .B(n105), .CI(C[153]), .CO(C[154]) );
  FA_878 \FAINST[154].FA_  ( .A(A[154]), .B(n104), .CI(C[154]), .CO(C[155]) );
  FA_877 \FAINST[155].FA_  ( .A(A[155]), .B(n103), .CI(C[155]), .CO(C[156]) );
  FA_876 \FAINST[156].FA_  ( .A(A[156]), .B(n102), .CI(C[156]), .CO(C[157]) );
  FA_875 \FAINST[157].FA_  ( .A(A[157]), .B(n101), .CI(C[157]), .CO(C[158]) );
  FA_874 \FAINST[158].FA_  ( .A(A[158]), .B(n100), .CI(C[158]), .CO(C[159]) );
  FA_873 \FAINST[159].FA_  ( .A(A[159]), .B(n99), .CI(C[159]), .CO(C[160]) );
  FA_872 \FAINST[160].FA_  ( .A(A[160]), .B(n98), .CI(C[160]), .CO(C[161]) );
  FA_871 \FAINST[161].FA_  ( .A(A[161]), .B(n97), .CI(C[161]), .CO(C[162]) );
  FA_870 \FAINST[162].FA_  ( .A(A[162]), .B(n96), .CI(C[162]), .CO(C[163]) );
  FA_869 \FAINST[163].FA_  ( .A(A[163]), .B(n95), .CI(C[163]), .CO(C[164]) );
  FA_868 \FAINST[164].FA_  ( .A(A[164]), .B(n94), .CI(C[164]), .CO(C[165]) );
  FA_867 \FAINST[165].FA_  ( .A(A[165]), .B(n93), .CI(C[165]), .CO(C[166]) );
  FA_866 \FAINST[166].FA_  ( .A(A[166]), .B(n92), .CI(C[166]), .CO(C[167]) );
  FA_865 \FAINST[167].FA_  ( .A(A[167]), .B(n91), .CI(C[167]), .CO(C[168]) );
  FA_864 \FAINST[168].FA_  ( .A(A[168]), .B(n90), .CI(C[168]), .CO(C[169]) );
  FA_863 \FAINST[169].FA_  ( .A(A[169]), .B(n89), .CI(C[169]), .CO(C[170]) );
  FA_862 \FAINST[170].FA_  ( .A(A[170]), .B(n88), .CI(C[170]), .CO(C[171]) );
  FA_861 \FAINST[171].FA_  ( .A(A[171]), .B(n87), .CI(C[171]), .CO(C[172]) );
  FA_860 \FAINST[172].FA_  ( .A(A[172]), .B(n86), .CI(C[172]), .CO(C[173]) );
  FA_859 \FAINST[173].FA_  ( .A(A[173]), .B(n85), .CI(C[173]), .CO(C[174]) );
  FA_858 \FAINST[174].FA_  ( .A(A[174]), .B(n84), .CI(C[174]), .CO(C[175]) );
  FA_857 \FAINST[175].FA_  ( .A(A[175]), .B(n83), .CI(C[175]), .CO(C[176]) );
  FA_856 \FAINST[176].FA_  ( .A(A[176]), .B(n82), .CI(C[176]), .CO(C[177]) );
  FA_855 \FAINST[177].FA_  ( .A(A[177]), .B(n81), .CI(C[177]), .CO(C[178]) );
  FA_854 \FAINST[178].FA_  ( .A(A[178]), .B(n80), .CI(C[178]), .CO(C[179]) );
  FA_853 \FAINST[179].FA_  ( .A(A[179]), .B(n79), .CI(C[179]), .CO(C[180]) );
  FA_852 \FAINST[180].FA_  ( .A(A[180]), .B(n78), .CI(C[180]), .CO(C[181]) );
  FA_851 \FAINST[181].FA_  ( .A(A[181]), .B(n77), .CI(C[181]), .CO(C[182]) );
  FA_850 \FAINST[182].FA_  ( .A(A[182]), .B(n76), .CI(C[182]), .CO(C[183]) );
  FA_849 \FAINST[183].FA_  ( .A(A[183]), .B(n75), .CI(C[183]), .CO(C[184]) );
  FA_848 \FAINST[184].FA_  ( .A(A[184]), .B(n74), .CI(C[184]), .CO(C[185]) );
  FA_847 \FAINST[185].FA_  ( .A(A[185]), .B(n73), .CI(C[185]), .CO(C[186]) );
  FA_846 \FAINST[186].FA_  ( .A(A[186]), .B(n72), .CI(C[186]), .CO(C[187]) );
  FA_845 \FAINST[187].FA_  ( .A(A[187]), .B(n71), .CI(C[187]), .CO(C[188]) );
  FA_844 \FAINST[188].FA_  ( .A(A[188]), .B(n70), .CI(C[188]), .CO(C[189]) );
  FA_843 \FAINST[189].FA_  ( .A(A[189]), .B(n69), .CI(C[189]), .CO(C[190]) );
  FA_842 \FAINST[190].FA_  ( .A(A[190]), .B(n68), .CI(C[190]), .CO(C[191]) );
  FA_841 \FAINST[191].FA_  ( .A(A[191]), .B(n67), .CI(C[191]), .CO(C[192]) );
  FA_840 \FAINST[192].FA_  ( .A(A[192]), .B(n66), .CI(C[192]), .CO(C[193]) );
  FA_839 \FAINST[193].FA_  ( .A(A[193]), .B(n65), .CI(C[193]), .CO(C[194]) );
  FA_838 \FAINST[194].FA_  ( .A(A[194]), .B(n64), .CI(C[194]), .CO(C[195]) );
  FA_837 \FAINST[195].FA_  ( .A(A[195]), .B(n63), .CI(C[195]), .CO(C[196]) );
  FA_836 \FAINST[196].FA_  ( .A(A[196]), .B(n62), .CI(C[196]), .CO(C[197]) );
  FA_835 \FAINST[197].FA_  ( .A(A[197]), .B(n61), .CI(C[197]), .CO(C[198]) );
  FA_834 \FAINST[198].FA_  ( .A(A[198]), .B(n60), .CI(C[198]), .CO(C[199]) );
  FA_833 \FAINST[199].FA_  ( .A(A[199]), .B(n59), .CI(C[199]), .CO(C[200]) );
  FA_832 \FAINST[200].FA_  ( .A(A[200]), .B(n58), .CI(C[200]), .CO(C[201]) );
  FA_831 \FAINST[201].FA_  ( .A(A[201]), .B(n57), .CI(C[201]), .CO(C[202]) );
  FA_830 \FAINST[202].FA_  ( .A(A[202]), .B(n56), .CI(C[202]), .CO(C[203]) );
  FA_829 \FAINST[203].FA_  ( .A(A[203]), .B(n55), .CI(C[203]), .CO(C[204]) );
  FA_828 \FAINST[204].FA_  ( .A(A[204]), .B(n54), .CI(C[204]), .CO(C[205]) );
  FA_827 \FAINST[205].FA_  ( .A(A[205]), .B(n53), .CI(C[205]), .CO(C[206]) );
  FA_826 \FAINST[206].FA_  ( .A(A[206]), .B(n52), .CI(C[206]), .CO(C[207]) );
  FA_825 \FAINST[207].FA_  ( .A(A[207]), .B(n51), .CI(C[207]), .CO(C[208]) );
  FA_824 \FAINST[208].FA_  ( .A(A[208]), .B(n50), .CI(C[208]), .CO(C[209]) );
  FA_823 \FAINST[209].FA_  ( .A(A[209]), .B(n49), .CI(C[209]), .CO(C[210]) );
  FA_822 \FAINST[210].FA_  ( .A(A[210]), .B(n48), .CI(C[210]), .CO(C[211]) );
  FA_821 \FAINST[211].FA_  ( .A(A[211]), .B(n47), .CI(C[211]), .CO(C[212]) );
  FA_820 \FAINST[212].FA_  ( .A(A[212]), .B(n46), .CI(C[212]), .CO(C[213]) );
  FA_819 \FAINST[213].FA_  ( .A(A[213]), .B(n45), .CI(C[213]), .CO(C[214]) );
  FA_818 \FAINST[214].FA_  ( .A(A[214]), .B(n44), .CI(C[214]), .CO(C[215]) );
  FA_817 \FAINST[215].FA_  ( .A(A[215]), .B(n43), .CI(C[215]), .CO(C[216]) );
  FA_816 \FAINST[216].FA_  ( .A(A[216]), .B(n42), .CI(C[216]), .CO(C[217]) );
  FA_815 \FAINST[217].FA_  ( .A(A[217]), .B(n41), .CI(C[217]), .CO(C[218]) );
  FA_814 \FAINST[218].FA_  ( .A(A[218]), .B(n40), .CI(C[218]), .CO(C[219]) );
  FA_813 \FAINST[219].FA_  ( .A(A[219]), .B(n39), .CI(C[219]), .CO(C[220]) );
  FA_812 \FAINST[220].FA_  ( .A(A[220]), .B(n38), .CI(C[220]), .CO(C[221]) );
  FA_811 \FAINST[221].FA_  ( .A(A[221]), .B(n37), .CI(C[221]), .CO(C[222]) );
  FA_810 \FAINST[222].FA_  ( .A(A[222]), .B(n36), .CI(C[222]), .CO(C[223]) );
  FA_809 \FAINST[223].FA_  ( .A(A[223]), .B(n35), .CI(C[223]), .CO(C[224]) );
  FA_808 \FAINST[224].FA_  ( .A(A[224]), .B(n34), .CI(C[224]), .CO(C[225]) );
  FA_807 \FAINST[225].FA_  ( .A(A[225]), .B(n33), .CI(C[225]), .CO(C[226]) );
  FA_806 \FAINST[226].FA_  ( .A(A[226]), .B(n32), .CI(C[226]), .CO(C[227]) );
  FA_805 \FAINST[227].FA_  ( .A(A[227]), .B(n31), .CI(C[227]), .CO(C[228]) );
  FA_804 \FAINST[228].FA_  ( .A(A[228]), .B(n30), .CI(C[228]), .CO(C[229]) );
  FA_803 \FAINST[229].FA_  ( .A(A[229]), .B(n29), .CI(C[229]), .CO(C[230]) );
  FA_802 \FAINST[230].FA_  ( .A(A[230]), .B(n28), .CI(C[230]), .CO(C[231]) );
  FA_801 \FAINST[231].FA_  ( .A(A[231]), .B(n27), .CI(C[231]), .CO(C[232]) );
  FA_800 \FAINST[232].FA_  ( .A(A[232]), .B(n26), .CI(C[232]), .CO(C[233]) );
  FA_799 \FAINST[233].FA_  ( .A(A[233]), .B(n25), .CI(C[233]), .CO(C[234]) );
  FA_798 \FAINST[234].FA_  ( .A(A[234]), .B(n24), .CI(C[234]), .CO(C[235]) );
  FA_797 \FAINST[235].FA_  ( .A(A[235]), .B(n23), .CI(C[235]), .CO(C[236]) );
  FA_796 \FAINST[236].FA_  ( .A(A[236]), .B(n22), .CI(C[236]), .CO(C[237]) );
  FA_795 \FAINST[237].FA_  ( .A(A[237]), .B(n21), .CI(C[237]), .CO(C[238]) );
  FA_794 \FAINST[238].FA_  ( .A(A[238]), .B(n20), .CI(C[238]), .CO(C[239]) );
  FA_793 \FAINST[239].FA_  ( .A(A[239]), .B(n19), .CI(C[239]), .CO(C[240]) );
  FA_792 \FAINST[240].FA_  ( .A(A[240]), .B(n18), .CI(C[240]), .CO(C[241]) );
  FA_791 \FAINST[241].FA_  ( .A(A[241]), .B(n17), .CI(C[241]), .CO(C[242]) );
  FA_790 \FAINST[242].FA_  ( .A(A[242]), .B(n16), .CI(C[242]), .CO(C[243]) );
  FA_789 \FAINST[243].FA_  ( .A(A[243]), .B(n15), .CI(C[243]), .CO(C[244]) );
  FA_788 \FAINST[244].FA_  ( .A(A[244]), .B(n14), .CI(C[244]), .CO(C[245]) );
  FA_787 \FAINST[245].FA_  ( .A(A[245]), .B(n13), .CI(C[245]), .CO(C[246]) );
  FA_786 \FAINST[246].FA_  ( .A(A[246]), .B(n12), .CI(C[246]), .CO(C[247]) );
  FA_785 \FAINST[247].FA_  ( .A(A[247]), .B(n11), .CI(C[247]), .CO(C[248]) );
  FA_784 \FAINST[248].FA_  ( .A(A[248]), .B(n10), .CI(C[248]), .CO(C[249]) );
  FA_783 \FAINST[249].FA_  ( .A(A[249]), .B(n9), .CI(C[249]), .CO(C[250]) );
  FA_782 \FAINST[250].FA_  ( .A(A[250]), .B(n8), .CI(C[250]), .CO(C[251]) );
  FA_781 \FAINST[251].FA_  ( .A(A[251]), .B(n7), .CI(C[251]), .CO(C[252]) );
  FA_780 \FAINST[252].FA_  ( .A(A[252]), .B(n6), .CI(C[252]), .CO(C[253]) );
  FA_779 \FAINST[253].FA_  ( .A(A[253]), .B(n5), .CI(C[253]), .CO(C[254]) );
  FA_778 \FAINST[254].FA_  ( .A(A[254]), .B(n4), .CI(C[254]), .CO(C[255]) );
  FA_777 \FAINST[255].FA_  ( .A(A[255]), .B(n3), .CI(C[255]), .CO(C[256]) );
  FA_776 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .CO(C[257]) );
  FA_775 \FAINST[257].FA_  ( .A(A[257]), .B(1'b1), .CI(C[257]), .CO(O) );
  IV U2 ( .A(B[159]), .Z(n99) );
  IV U3 ( .A(B[160]), .Z(n98) );
  IV U4 ( .A(B[161]), .Z(n97) );
  IV U5 ( .A(B[162]), .Z(n96) );
  IV U6 ( .A(B[163]), .Z(n95) );
  IV U7 ( .A(B[164]), .Z(n94) );
  IV U8 ( .A(B[165]), .Z(n93) );
  IV U9 ( .A(B[166]), .Z(n92) );
  IV U10 ( .A(B[167]), .Z(n91) );
  IV U11 ( .A(B[168]), .Z(n90) );
  IV U12 ( .A(B[249]), .Z(n9) );
  IV U13 ( .A(B[169]), .Z(n89) );
  IV U14 ( .A(B[170]), .Z(n88) );
  IV U15 ( .A(B[171]), .Z(n87) );
  IV U16 ( .A(B[172]), .Z(n86) );
  IV U17 ( .A(B[173]), .Z(n85) );
  IV U18 ( .A(B[174]), .Z(n84) );
  IV U19 ( .A(B[175]), .Z(n83) );
  IV U20 ( .A(B[176]), .Z(n82) );
  IV U21 ( .A(B[177]), .Z(n81) );
  IV U22 ( .A(B[178]), .Z(n80) );
  IV U23 ( .A(B[250]), .Z(n8) );
  IV U24 ( .A(B[179]), .Z(n79) );
  IV U25 ( .A(B[180]), .Z(n78) );
  IV U26 ( .A(B[181]), .Z(n77) );
  IV U27 ( .A(B[182]), .Z(n76) );
  IV U28 ( .A(B[183]), .Z(n75) );
  IV U29 ( .A(B[184]), .Z(n74) );
  IV U30 ( .A(B[185]), .Z(n73) );
  IV U31 ( .A(B[186]), .Z(n72) );
  IV U32 ( .A(B[187]), .Z(n71) );
  IV U33 ( .A(B[188]), .Z(n70) );
  IV U34 ( .A(B[251]), .Z(n7) );
  IV U35 ( .A(B[189]), .Z(n69) );
  IV U36 ( .A(B[190]), .Z(n68) );
  IV U37 ( .A(B[191]), .Z(n67) );
  IV U38 ( .A(B[192]), .Z(n66) );
  IV U39 ( .A(B[193]), .Z(n65) );
  IV U40 ( .A(B[194]), .Z(n64) );
  IV U41 ( .A(B[195]), .Z(n63) );
  IV U42 ( .A(B[196]), .Z(n62) );
  IV U43 ( .A(B[197]), .Z(n61) );
  IV U44 ( .A(B[198]), .Z(n60) );
  IV U45 ( .A(B[252]), .Z(n6) );
  IV U46 ( .A(B[199]), .Z(n59) );
  IV U47 ( .A(B[200]), .Z(n58) );
  IV U48 ( .A(B[201]), .Z(n57) );
  IV U49 ( .A(B[202]), .Z(n56) );
  IV U50 ( .A(B[203]), .Z(n55) );
  IV U51 ( .A(B[204]), .Z(n54) );
  IV U52 ( .A(B[205]), .Z(n53) );
  IV U53 ( .A(B[206]), .Z(n52) );
  IV U54 ( .A(B[207]), .Z(n51) );
  IV U55 ( .A(B[208]), .Z(n50) );
  IV U56 ( .A(B[253]), .Z(n5) );
  IV U57 ( .A(B[209]), .Z(n49) );
  IV U58 ( .A(B[210]), .Z(n48) );
  IV U59 ( .A(B[211]), .Z(n47) );
  IV U60 ( .A(B[212]), .Z(n46) );
  IV U61 ( .A(B[213]), .Z(n45) );
  IV U62 ( .A(B[214]), .Z(n44) );
  IV U63 ( .A(B[215]), .Z(n43) );
  IV U64 ( .A(B[216]), .Z(n42) );
  IV U65 ( .A(B[217]), .Z(n41) );
  IV U66 ( .A(B[218]), .Z(n40) );
  IV U67 ( .A(B[254]), .Z(n4) );
  IV U68 ( .A(B[219]), .Z(n39) );
  IV U69 ( .A(B[220]), .Z(n38) );
  IV U70 ( .A(B[221]), .Z(n37) );
  IV U71 ( .A(B[222]), .Z(n36) );
  IV U72 ( .A(B[223]), .Z(n35) );
  IV U73 ( .A(B[224]), .Z(n34) );
  IV U74 ( .A(B[225]), .Z(n33) );
  IV U75 ( .A(B[226]), .Z(n32) );
  IV U76 ( .A(B[227]), .Z(n31) );
  IV U77 ( .A(B[228]), .Z(n30) );
  IV U78 ( .A(B[255]), .Z(n3) );
  IV U79 ( .A(B[229]), .Z(n29) );
  IV U80 ( .A(B[230]), .Z(n28) );
  IV U81 ( .A(B[231]), .Z(n27) );
  IV U82 ( .A(B[232]), .Z(n26) );
  IV U83 ( .A(B[0]), .Z(n258) );
  IV U84 ( .A(B[1]), .Z(n257) );
  IV U85 ( .A(B[2]), .Z(n256) );
  IV U86 ( .A(B[3]), .Z(n255) );
  IV U87 ( .A(B[4]), .Z(n254) );
  IV U88 ( .A(B[5]), .Z(n253) );
  IV U89 ( .A(B[6]), .Z(n252) );
  IV U90 ( .A(B[7]), .Z(n251) );
  IV U91 ( .A(B[8]), .Z(n250) );
  IV U92 ( .A(B[233]), .Z(n25) );
  IV U93 ( .A(B[9]), .Z(n249) );
  IV U94 ( .A(B[10]), .Z(n248) );
  IV U95 ( .A(B[11]), .Z(n247) );
  IV U96 ( .A(B[12]), .Z(n246) );
  IV U97 ( .A(B[13]), .Z(n245) );
  IV U98 ( .A(B[14]), .Z(n244) );
  IV U99 ( .A(B[15]), .Z(n243) );
  IV U100 ( .A(B[16]), .Z(n242) );
  IV U101 ( .A(B[17]), .Z(n241) );
  IV U102 ( .A(B[18]), .Z(n240) );
  IV U103 ( .A(B[234]), .Z(n24) );
  IV U104 ( .A(B[19]), .Z(n239) );
  IV U105 ( .A(B[20]), .Z(n238) );
  IV U106 ( .A(B[21]), .Z(n237) );
  IV U107 ( .A(B[22]), .Z(n236) );
  IV U108 ( .A(B[23]), .Z(n235) );
  IV U109 ( .A(B[24]), .Z(n234) );
  IV U110 ( .A(B[25]), .Z(n233) );
  IV U111 ( .A(B[26]), .Z(n232) );
  IV U112 ( .A(B[27]), .Z(n231) );
  IV U113 ( .A(B[28]), .Z(n230) );
  IV U114 ( .A(B[235]), .Z(n23) );
  IV U115 ( .A(B[29]), .Z(n229) );
  IV U116 ( .A(B[30]), .Z(n228) );
  IV U117 ( .A(B[31]), .Z(n227) );
  IV U118 ( .A(B[32]), .Z(n226) );
  IV U119 ( .A(B[33]), .Z(n225) );
  IV U120 ( .A(B[34]), .Z(n224) );
  IV U121 ( .A(B[35]), .Z(n223) );
  IV U122 ( .A(B[36]), .Z(n222) );
  IV U123 ( .A(B[37]), .Z(n221) );
  IV U124 ( .A(B[38]), .Z(n220) );
  IV U125 ( .A(B[236]), .Z(n22) );
  IV U126 ( .A(B[39]), .Z(n219) );
  IV U127 ( .A(B[40]), .Z(n218) );
  IV U128 ( .A(B[41]), .Z(n217) );
  IV U129 ( .A(B[42]), .Z(n216) );
  IV U130 ( .A(B[43]), .Z(n215) );
  IV U131 ( .A(B[44]), .Z(n214) );
  IV U132 ( .A(B[45]), .Z(n213) );
  IV U133 ( .A(B[46]), .Z(n212) );
  IV U134 ( .A(B[47]), .Z(n211) );
  IV U135 ( .A(B[48]), .Z(n210) );
  IV U136 ( .A(B[237]), .Z(n21) );
  IV U137 ( .A(B[49]), .Z(n209) );
  IV U138 ( .A(B[50]), .Z(n208) );
  IV U139 ( .A(B[51]), .Z(n207) );
  IV U140 ( .A(B[52]), .Z(n206) );
  IV U141 ( .A(B[53]), .Z(n205) );
  IV U142 ( .A(B[54]), .Z(n204) );
  IV U143 ( .A(B[55]), .Z(n203) );
  IV U144 ( .A(B[56]), .Z(n202) );
  IV U145 ( .A(B[57]), .Z(n201) );
  IV U146 ( .A(B[58]), .Z(n200) );
  IV U147 ( .A(B[238]), .Z(n20) );
  IV U148 ( .A(B[59]), .Z(n199) );
  IV U149 ( .A(B[60]), .Z(n198) );
  IV U150 ( .A(B[61]), .Z(n197) );
  IV U151 ( .A(B[62]), .Z(n196) );
  IV U152 ( .A(B[63]), .Z(n195) );
  IV U153 ( .A(B[64]), .Z(n194) );
  IV U154 ( .A(B[65]), .Z(n193) );
  IV U155 ( .A(B[66]), .Z(n192) );
  IV U156 ( .A(B[67]), .Z(n191) );
  IV U157 ( .A(B[68]), .Z(n190) );
  IV U158 ( .A(B[239]), .Z(n19) );
  IV U159 ( .A(B[69]), .Z(n189) );
  IV U160 ( .A(B[70]), .Z(n188) );
  IV U161 ( .A(B[71]), .Z(n187) );
  IV U162 ( .A(B[72]), .Z(n186) );
  IV U163 ( .A(B[73]), .Z(n185) );
  IV U164 ( .A(B[74]), .Z(n184) );
  IV U165 ( .A(B[75]), .Z(n183) );
  IV U166 ( .A(B[76]), .Z(n182) );
  IV U167 ( .A(B[77]), .Z(n181) );
  IV U168 ( .A(B[78]), .Z(n180) );
  IV U169 ( .A(B[240]), .Z(n18) );
  IV U170 ( .A(B[79]), .Z(n179) );
  IV U171 ( .A(B[80]), .Z(n178) );
  IV U172 ( .A(B[81]), .Z(n177) );
  IV U173 ( .A(B[82]), .Z(n176) );
  IV U174 ( .A(B[83]), .Z(n175) );
  IV U175 ( .A(B[84]), .Z(n174) );
  IV U176 ( .A(B[85]), .Z(n173) );
  IV U177 ( .A(B[86]), .Z(n172) );
  IV U178 ( .A(B[87]), .Z(n171) );
  IV U179 ( .A(B[88]), .Z(n170) );
  IV U180 ( .A(B[241]), .Z(n17) );
  IV U181 ( .A(B[89]), .Z(n169) );
  IV U182 ( .A(B[90]), .Z(n168) );
  IV U183 ( .A(B[91]), .Z(n167) );
  IV U184 ( .A(B[92]), .Z(n166) );
  IV U185 ( .A(B[93]), .Z(n165) );
  IV U186 ( .A(B[94]), .Z(n164) );
  IV U187 ( .A(B[95]), .Z(n163) );
  IV U188 ( .A(B[96]), .Z(n162) );
  IV U189 ( .A(B[97]), .Z(n161) );
  IV U190 ( .A(B[98]), .Z(n160) );
  IV U191 ( .A(B[242]), .Z(n16) );
  IV U192 ( .A(B[99]), .Z(n159) );
  IV U193 ( .A(B[100]), .Z(n158) );
  IV U194 ( .A(B[101]), .Z(n157) );
  IV U195 ( .A(B[102]), .Z(n156) );
  IV U196 ( .A(B[103]), .Z(n155) );
  IV U197 ( .A(B[104]), .Z(n154) );
  IV U198 ( .A(B[105]), .Z(n153) );
  IV U199 ( .A(B[106]), .Z(n152) );
  IV U200 ( .A(B[107]), .Z(n151) );
  IV U201 ( .A(B[108]), .Z(n150) );
  IV U202 ( .A(B[243]), .Z(n15) );
  IV U203 ( .A(B[109]), .Z(n149) );
  IV U204 ( .A(B[110]), .Z(n148) );
  IV U205 ( .A(B[111]), .Z(n147) );
  IV U206 ( .A(B[112]), .Z(n146) );
  IV U207 ( .A(B[113]), .Z(n145) );
  IV U208 ( .A(B[114]), .Z(n144) );
  IV U209 ( .A(B[115]), .Z(n143) );
  IV U210 ( .A(B[116]), .Z(n142) );
  IV U211 ( .A(B[117]), .Z(n141) );
  IV U212 ( .A(B[118]), .Z(n140) );
  IV U213 ( .A(B[244]), .Z(n14) );
  IV U214 ( .A(B[119]), .Z(n139) );
  IV U215 ( .A(B[120]), .Z(n138) );
  IV U216 ( .A(B[121]), .Z(n137) );
  IV U217 ( .A(B[122]), .Z(n136) );
  IV U218 ( .A(B[123]), .Z(n135) );
  IV U219 ( .A(B[124]), .Z(n134) );
  IV U220 ( .A(B[125]), .Z(n133) );
  IV U221 ( .A(B[126]), .Z(n132) );
  IV U222 ( .A(B[127]), .Z(n131) );
  IV U223 ( .A(B[128]), .Z(n130) );
  IV U224 ( .A(B[245]), .Z(n13) );
  IV U225 ( .A(B[129]), .Z(n129) );
  IV U226 ( .A(B[130]), .Z(n128) );
  IV U227 ( .A(B[131]), .Z(n127) );
  IV U228 ( .A(B[132]), .Z(n126) );
  IV U229 ( .A(B[133]), .Z(n125) );
  IV U230 ( .A(B[134]), .Z(n124) );
  IV U231 ( .A(B[135]), .Z(n123) );
  IV U232 ( .A(B[136]), .Z(n122) );
  IV U233 ( .A(B[137]), .Z(n121) );
  IV U234 ( .A(B[138]), .Z(n120) );
  IV U235 ( .A(B[246]), .Z(n12) );
  IV U236 ( .A(B[139]), .Z(n119) );
  IV U237 ( .A(B[140]), .Z(n118) );
  IV U238 ( .A(B[141]), .Z(n117) );
  IV U239 ( .A(B[142]), .Z(n116) );
  IV U240 ( .A(B[143]), .Z(n115) );
  IV U241 ( .A(B[144]), .Z(n114) );
  IV U242 ( .A(B[145]), .Z(n113) );
  IV U243 ( .A(B[146]), .Z(n112) );
  IV U244 ( .A(B[147]), .Z(n111) );
  IV U245 ( .A(B[148]), .Z(n110) );
  IV U246 ( .A(B[247]), .Z(n11) );
  IV U247 ( .A(B[149]), .Z(n109) );
  IV U248 ( .A(B[150]), .Z(n108) );
  IV U249 ( .A(B[151]), .Z(n107) );
  IV U250 ( .A(B[152]), .Z(n106) );
  IV U251 ( .A(B[153]), .Z(n105) );
  IV U252 ( .A(B[154]), .Z(n104) );
  IV U253 ( .A(B[155]), .Z(n103) );
  IV U254 ( .A(B[156]), .Z(n102) );
  IV U255 ( .A(B[157]), .Z(n101) );
  IV U256 ( .A(B[158]), .Z(n100) );
  IV U257 ( .A(B[248]), .Z(n10) );
endmodule


module FA_517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  NANDN U1 ( .A(CI), .B(S), .Z(CO) );
  XNOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N258_0 ( A, B, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258;
  wire   [257:1] C;

  FA_774 \FAINST[0].FA_  ( .A(A[0]), .B(n258), .CI(1'b1), .S(S[0]), .CO(C[1])
         );
  FA_773 \FAINST[1].FA_  ( .A(A[1]), .B(n257), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_772 \FAINST[2].FA_  ( .A(A[2]), .B(n256), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_771 \FAINST[3].FA_  ( .A(A[3]), .B(n255), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_770 \FAINST[4].FA_  ( .A(A[4]), .B(n254), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_769 \FAINST[5].FA_  ( .A(A[5]), .B(n253), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_768 \FAINST[6].FA_  ( .A(A[6]), .B(n252), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_767 \FAINST[7].FA_  ( .A(A[7]), .B(n251), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_766 \FAINST[8].FA_  ( .A(A[8]), .B(n250), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_765 \FAINST[9].FA_  ( .A(A[9]), .B(n249), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_764 \FAINST[10].FA_  ( .A(A[10]), .B(n248), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_763 \FAINST[11].FA_  ( .A(A[11]), .B(n247), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_762 \FAINST[12].FA_  ( .A(A[12]), .B(n246), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_761 \FAINST[13].FA_  ( .A(A[13]), .B(n245), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_760 \FAINST[14].FA_  ( .A(A[14]), .B(n244), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_759 \FAINST[15].FA_  ( .A(A[15]), .B(n243), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_758 \FAINST[16].FA_  ( .A(A[16]), .B(n242), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_757 \FAINST[17].FA_  ( .A(A[17]), .B(n241), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_756 \FAINST[18].FA_  ( .A(A[18]), .B(n240), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_755 \FAINST[19].FA_  ( .A(A[19]), .B(n239), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_754 \FAINST[20].FA_  ( .A(A[20]), .B(n238), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_753 \FAINST[21].FA_  ( .A(A[21]), .B(n237), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_752 \FAINST[22].FA_  ( .A(A[22]), .B(n236), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_751 \FAINST[23].FA_  ( .A(A[23]), .B(n235), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_750 \FAINST[24].FA_  ( .A(A[24]), .B(n234), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_749 \FAINST[25].FA_  ( .A(A[25]), .B(n233), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_748 \FAINST[26].FA_  ( .A(A[26]), .B(n232), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_747 \FAINST[27].FA_  ( .A(A[27]), .B(n231), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_746 \FAINST[28].FA_  ( .A(A[28]), .B(n230), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_745 \FAINST[29].FA_  ( .A(A[29]), .B(n229), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_744 \FAINST[30].FA_  ( .A(A[30]), .B(n228), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_743 \FAINST[31].FA_  ( .A(A[31]), .B(n227), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_742 \FAINST[32].FA_  ( .A(A[32]), .B(n226), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_741 \FAINST[33].FA_  ( .A(A[33]), .B(n225), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_740 \FAINST[34].FA_  ( .A(A[34]), .B(n224), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_739 \FAINST[35].FA_  ( .A(A[35]), .B(n223), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_738 \FAINST[36].FA_  ( .A(A[36]), .B(n222), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_737 \FAINST[37].FA_  ( .A(A[37]), .B(n221), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_736 \FAINST[38].FA_  ( .A(A[38]), .B(n220), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_735 \FAINST[39].FA_  ( .A(A[39]), .B(n219), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_734 \FAINST[40].FA_  ( .A(A[40]), .B(n218), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_733 \FAINST[41].FA_  ( .A(A[41]), .B(n217), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_732 \FAINST[42].FA_  ( .A(A[42]), .B(n216), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_731 \FAINST[43].FA_  ( .A(A[43]), .B(n215), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_730 \FAINST[44].FA_  ( .A(A[44]), .B(n214), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_729 \FAINST[45].FA_  ( .A(A[45]), .B(n213), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_728 \FAINST[46].FA_  ( .A(A[46]), .B(n212), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_727 \FAINST[47].FA_  ( .A(A[47]), .B(n211), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_726 \FAINST[48].FA_  ( .A(A[48]), .B(n210), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_725 \FAINST[49].FA_  ( .A(A[49]), .B(n209), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_724 \FAINST[50].FA_  ( .A(A[50]), .B(n208), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_723 \FAINST[51].FA_  ( .A(A[51]), .B(n207), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_722 \FAINST[52].FA_  ( .A(A[52]), .B(n206), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_721 \FAINST[53].FA_  ( .A(A[53]), .B(n205), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_720 \FAINST[54].FA_  ( .A(A[54]), .B(n204), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_719 \FAINST[55].FA_  ( .A(A[55]), .B(n203), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_718 \FAINST[56].FA_  ( .A(A[56]), .B(n202), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_717 \FAINST[57].FA_  ( .A(A[57]), .B(n201), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_716 \FAINST[58].FA_  ( .A(A[58]), .B(n200), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_715 \FAINST[59].FA_  ( .A(A[59]), .B(n199), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_714 \FAINST[60].FA_  ( .A(A[60]), .B(n198), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_713 \FAINST[61].FA_  ( .A(A[61]), .B(n197), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_712 \FAINST[62].FA_  ( .A(A[62]), .B(n196), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_711 \FAINST[63].FA_  ( .A(A[63]), .B(n195), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_710 \FAINST[64].FA_  ( .A(A[64]), .B(n194), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_709 \FAINST[65].FA_  ( .A(A[65]), .B(n193), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_708 \FAINST[66].FA_  ( .A(A[66]), .B(n192), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_707 \FAINST[67].FA_  ( .A(A[67]), .B(n191), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_706 \FAINST[68].FA_  ( .A(A[68]), .B(n190), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_705 \FAINST[69].FA_  ( .A(A[69]), .B(n189), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_704 \FAINST[70].FA_  ( .A(A[70]), .B(n188), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_703 \FAINST[71].FA_  ( .A(A[71]), .B(n187), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_702 \FAINST[72].FA_  ( .A(A[72]), .B(n186), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_701 \FAINST[73].FA_  ( .A(A[73]), .B(n185), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_700 \FAINST[74].FA_  ( .A(A[74]), .B(n184), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_699 \FAINST[75].FA_  ( .A(A[75]), .B(n183), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_698 \FAINST[76].FA_  ( .A(A[76]), .B(n182), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_697 \FAINST[77].FA_  ( .A(A[77]), .B(n181), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_696 \FAINST[78].FA_  ( .A(A[78]), .B(n180), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_695 \FAINST[79].FA_  ( .A(A[79]), .B(n179), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_694 \FAINST[80].FA_  ( .A(A[80]), .B(n178), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_693 \FAINST[81].FA_  ( .A(A[81]), .B(n177), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_692 \FAINST[82].FA_  ( .A(A[82]), .B(n176), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_691 \FAINST[83].FA_  ( .A(A[83]), .B(n175), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_690 \FAINST[84].FA_  ( .A(A[84]), .B(n174), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_689 \FAINST[85].FA_  ( .A(A[85]), .B(n173), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_688 \FAINST[86].FA_  ( .A(A[86]), .B(n172), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_687 \FAINST[87].FA_  ( .A(A[87]), .B(n171), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_686 \FAINST[88].FA_  ( .A(A[88]), .B(n170), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_685 \FAINST[89].FA_  ( .A(A[89]), .B(n169), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_684 \FAINST[90].FA_  ( .A(A[90]), .B(n168), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_683 \FAINST[91].FA_  ( .A(A[91]), .B(n167), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_682 \FAINST[92].FA_  ( .A(A[92]), .B(n166), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_681 \FAINST[93].FA_  ( .A(A[93]), .B(n165), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_680 \FAINST[94].FA_  ( .A(A[94]), .B(n164), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_679 \FAINST[95].FA_  ( .A(A[95]), .B(n163), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_678 \FAINST[96].FA_  ( .A(A[96]), .B(n162), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_677 \FAINST[97].FA_  ( .A(A[97]), .B(n161), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_676 \FAINST[98].FA_  ( .A(A[98]), .B(n160), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_675 \FAINST[99].FA_  ( .A(A[99]), .B(n159), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_674 \FAINST[100].FA_  ( .A(A[100]), .B(n158), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_673 \FAINST[101].FA_  ( .A(A[101]), .B(n157), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_672 \FAINST[102].FA_  ( .A(A[102]), .B(n156), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_671 \FAINST[103].FA_  ( .A(A[103]), .B(n155), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_670 \FAINST[104].FA_  ( .A(A[104]), .B(n154), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_669 \FAINST[105].FA_  ( .A(A[105]), .B(n153), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_668 \FAINST[106].FA_  ( .A(A[106]), .B(n152), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_667 \FAINST[107].FA_  ( .A(A[107]), .B(n151), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_666 \FAINST[108].FA_  ( .A(A[108]), .B(n150), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_665 \FAINST[109].FA_  ( .A(A[109]), .B(n149), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_664 \FAINST[110].FA_  ( .A(A[110]), .B(n148), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_663 \FAINST[111].FA_  ( .A(A[111]), .B(n147), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_662 \FAINST[112].FA_  ( .A(A[112]), .B(n146), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_661 \FAINST[113].FA_  ( .A(A[113]), .B(n145), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_660 \FAINST[114].FA_  ( .A(A[114]), .B(n144), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_659 \FAINST[115].FA_  ( .A(A[115]), .B(n143), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_658 \FAINST[116].FA_  ( .A(A[116]), .B(n142), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_657 \FAINST[117].FA_  ( .A(A[117]), .B(n141), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_656 \FAINST[118].FA_  ( .A(A[118]), .B(n140), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_655 \FAINST[119].FA_  ( .A(A[119]), .B(n139), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_654 \FAINST[120].FA_  ( .A(A[120]), .B(n138), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_653 \FAINST[121].FA_  ( .A(A[121]), .B(n137), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_652 \FAINST[122].FA_  ( .A(A[122]), .B(n136), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_651 \FAINST[123].FA_  ( .A(A[123]), .B(n135), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_650 \FAINST[124].FA_  ( .A(A[124]), .B(n134), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_649 \FAINST[125].FA_  ( .A(A[125]), .B(n133), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_648 \FAINST[126].FA_  ( .A(A[126]), .B(n132), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_647 \FAINST[127].FA_  ( .A(A[127]), .B(n131), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_646 \FAINST[128].FA_  ( .A(A[128]), .B(n130), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_645 \FAINST[129].FA_  ( .A(A[129]), .B(n129), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_644 \FAINST[130].FA_  ( .A(A[130]), .B(n128), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_643 \FAINST[131].FA_  ( .A(A[131]), .B(n127), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_642 \FAINST[132].FA_  ( .A(A[132]), .B(n126), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_641 \FAINST[133].FA_  ( .A(A[133]), .B(n125), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_640 \FAINST[134].FA_  ( .A(A[134]), .B(n124), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_639 \FAINST[135].FA_  ( .A(A[135]), .B(n123), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_638 \FAINST[136].FA_  ( .A(A[136]), .B(n122), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_637 \FAINST[137].FA_  ( .A(A[137]), .B(n121), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_636 \FAINST[138].FA_  ( .A(A[138]), .B(n120), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_635 \FAINST[139].FA_  ( .A(A[139]), .B(n119), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_634 \FAINST[140].FA_  ( .A(A[140]), .B(n118), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_633 \FAINST[141].FA_  ( .A(A[141]), .B(n117), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_632 \FAINST[142].FA_  ( .A(A[142]), .B(n116), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_631 \FAINST[143].FA_  ( .A(A[143]), .B(n115), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_630 \FAINST[144].FA_  ( .A(A[144]), .B(n114), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_629 \FAINST[145].FA_  ( .A(A[145]), .B(n113), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_628 \FAINST[146].FA_  ( .A(A[146]), .B(n112), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_627 \FAINST[147].FA_  ( .A(A[147]), .B(n111), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_626 \FAINST[148].FA_  ( .A(A[148]), .B(n110), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_625 \FAINST[149].FA_  ( .A(A[149]), .B(n109), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_624 \FAINST[150].FA_  ( .A(A[150]), .B(n108), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_623 \FAINST[151].FA_  ( .A(A[151]), .B(n107), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_622 \FAINST[152].FA_  ( .A(A[152]), .B(n106), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_621 \FAINST[153].FA_  ( .A(A[153]), .B(n105), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_620 \FAINST[154].FA_  ( .A(A[154]), .B(n104), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_619 \FAINST[155].FA_  ( .A(A[155]), .B(n103), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_618 \FAINST[156].FA_  ( .A(A[156]), .B(n102), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_617 \FAINST[157].FA_  ( .A(A[157]), .B(n101), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_616 \FAINST[158].FA_  ( .A(A[158]), .B(n100), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_615 \FAINST[159].FA_  ( .A(A[159]), .B(n99), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_614 \FAINST[160].FA_  ( .A(A[160]), .B(n98), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_613 \FAINST[161].FA_  ( .A(A[161]), .B(n97), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_612 \FAINST[162].FA_  ( .A(A[162]), .B(n96), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_611 \FAINST[163].FA_  ( .A(A[163]), .B(n95), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_610 \FAINST[164].FA_  ( .A(A[164]), .B(n94), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_609 \FAINST[165].FA_  ( .A(A[165]), .B(n93), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_608 \FAINST[166].FA_  ( .A(A[166]), .B(n92), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_607 \FAINST[167].FA_  ( .A(A[167]), .B(n91), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_606 \FAINST[168].FA_  ( .A(A[168]), .B(n90), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_605 \FAINST[169].FA_  ( .A(A[169]), .B(n89), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_604 \FAINST[170].FA_  ( .A(A[170]), .B(n88), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_603 \FAINST[171].FA_  ( .A(A[171]), .B(n87), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_602 \FAINST[172].FA_  ( .A(A[172]), .B(n86), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_601 \FAINST[173].FA_  ( .A(A[173]), .B(n85), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_600 \FAINST[174].FA_  ( .A(A[174]), .B(n84), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_599 \FAINST[175].FA_  ( .A(A[175]), .B(n83), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_598 \FAINST[176].FA_  ( .A(A[176]), .B(n82), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_597 \FAINST[177].FA_  ( .A(A[177]), .B(n81), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_596 \FAINST[178].FA_  ( .A(A[178]), .B(n80), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_595 \FAINST[179].FA_  ( .A(A[179]), .B(n79), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_594 \FAINST[180].FA_  ( .A(A[180]), .B(n78), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_593 \FAINST[181].FA_  ( .A(A[181]), .B(n77), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_592 \FAINST[182].FA_  ( .A(A[182]), .B(n76), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_591 \FAINST[183].FA_  ( .A(A[183]), .B(n75), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_590 \FAINST[184].FA_  ( .A(A[184]), .B(n74), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_589 \FAINST[185].FA_  ( .A(A[185]), .B(n73), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_588 \FAINST[186].FA_  ( .A(A[186]), .B(n72), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_587 \FAINST[187].FA_  ( .A(A[187]), .B(n71), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_586 \FAINST[188].FA_  ( .A(A[188]), .B(n70), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_585 \FAINST[189].FA_  ( .A(A[189]), .B(n69), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_584 \FAINST[190].FA_  ( .A(A[190]), .B(n68), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_583 \FAINST[191].FA_  ( .A(A[191]), .B(n67), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_582 \FAINST[192].FA_  ( .A(A[192]), .B(n66), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_581 \FAINST[193].FA_  ( .A(A[193]), .B(n65), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_580 \FAINST[194].FA_  ( .A(A[194]), .B(n64), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_579 \FAINST[195].FA_  ( .A(A[195]), .B(n63), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_578 \FAINST[196].FA_  ( .A(A[196]), .B(n62), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_577 \FAINST[197].FA_  ( .A(A[197]), .B(n61), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_576 \FAINST[198].FA_  ( .A(A[198]), .B(n60), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_575 \FAINST[199].FA_  ( .A(A[199]), .B(n59), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_574 \FAINST[200].FA_  ( .A(A[200]), .B(n58), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_573 \FAINST[201].FA_  ( .A(A[201]), .B(n57), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_572 \FAINST[202].FA_  ( .A(A[202]), .B(n56), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_571 \FAINST[203].FA_  ( .A(A[203]), .B(n55), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_570 \FAINST[204].FA_  ( .A(A[204]), .B(n54), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_569 \FAINST[205].FA_  ( .A(A[205]), .B(n53), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_568 \FAINST[206].FA_  ( .A(A[206]), .B(n52), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_567 \FAINST[207].FA_  ( .A(A[207]), .B(n51), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_566 \FAINST[208].FA_  ( .A(A[208]), .B(n50), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_565 \FAINST[209].FA_  ( .A(A[209]), .B(n49), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_564 \FAINST[210].FA_  ( .A(A[210]), .B(n48), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_563 \FAINST[211].FA_  ( .A(A[211]), .B(n47), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_562 \FAINST[212].FA_  ( .A(A[212]), .B(n46), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_561 \FAINST[213].FA_  ( .A(A[213]), .B(n45), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_560 \FAINST[214].FA_  ( .A(A[214]), .B(n44), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_559 \FAINST[215].FA_  ( .A(A[215]), .B(n43), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_558 \FAINST[216].FA_  ( .A(A[216]), .B(n42), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_557 \FAINST[217].FA_  ( .A(A[217]), .B(n41), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_556 \FAINST[218].FA_  ( .A(A[218]), .B(n40), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_555 \FAINST[219].FA_  ( .A(A[219]), .B(n39), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_554 \FAINST[220].FA_  ( .A(A[220]), .B(n38), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_553 \FAINST[221].FA_  ( .A(A[221]), .B(n37), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_552 \FAINST[222].FA_  ( .A(A[222]), .B(n36), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_551 \FAINST[223].FA_  ( .A(A[223]), .B(n35), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_550 \FAINST[224].FA_  ( .A(A[224]), .B(n34), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_549 \FAINST[225].FA_  ( .A(A[225]), .B(n33), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_548 \FAINST[226].FA_  ( .A(A[226]), .B(n32), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_547 \FAINST[227].FA_  ( .A(A[227]), .B(n31), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_546 \FAINST[228].FA_  ( .A(A[228]), .B(n30), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_545 \FAINST[229].FA_  ( .A(A[229]), .B(n29), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_544 \FAINST[230].FA_  ( .A(A[230]), .B(n28), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_543 \FAINST[231].FA_  ( .A(A[231]), .B(n27), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_542 \FAINST[232].FA_  ( .A(A[232]), .B(n26), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_541 \FAINST[233].FA_  ( .A(A[233]), .B(n25), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_540 \FAINST[234].FA_  ( .A(A[234]), .B(n24), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_539 \FAINST[235].FA_  ( .A(A[235]), .B(n23), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_538 \FAINST[236].FA_  ( .A(A[236]), .B(n22), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_537 \FAINST[237].FA_  ( .A(A[237]), .B(n21), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_536 \FAINST[238].FA_  ( .A(A[238]), .B(n20), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_535 \FAINST[239].FA_  ( .A(A[239]), .B(n19), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_534 \FAINST[240].FA_  ( .A(A[240]), .B(n18), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_533 \FAINST[241].FA_  ( .A(A[241]), .B(n17), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_532 \FAINST[242].FA_  ( .A(A[242]), .B(n16), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_531 \FAINST[243].FA_  ( .A(A[243]), .B(n15), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_530 \FAINST[244].FA_  ( .A(A[244]), .B(n14), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_529 \FAINST[245].FA_  ( .A(A[245]), .B(n13), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_528 \FAINST[246].FA_  ( .A(A[246]), .B(n12), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_527 \FAINST[247].FA_  ( .A(A[247]), .B(n11), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_526 \FAINST[248].FA_  ( .A(A[248]), .B(n10), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_525 \FAINST[249].FA_  ( .A(A[249]), .B(n9), .CI(C[249]), .S(S[249]), .CO(
        C[250]) );
  FA_524 \FAINST[250].FA_  ( .A(A[250]), .B(n8), .CI(C[250]), .S(S[250]), .CO(
        C[251]) );
  FA_523 \FAINST[251].FA_  ( .A(A[251]), .B(n7), .CI(C[251]), .S(S[251]), .CO(
        C[252]) );
  FA_522 \FAINST[252].FA_  ( .A(A[252]), .B(n6), .CI(C[252]), .S(S[252]), .CO(
        C[253]) );
  FA_521 \FAINST[253].FA_  ( .A(A[253]), .B(n5), .CI(C[253]), .S(S[253]), .CO(
        C[254]) );
  FA_520 \FAINST[254].FA_  ( .A(A[254]), .B(n4), .CI(C[254]), .S(S[254]), .CO(
        C[255]) );
  FA_519 \FAINST[255].FA_  ( .A(A[255]), .B(n3), .CI(C[255]), .S(S[255]), .CO(
        C[256]) );
  FA_518 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .S(S[256]), 
        .CO(C[257]) );
  FA_517 \FAINST[257].FA_  ( .A(A[257]), .B(1'b1), .CI(C[257]), .S(S[257]) );
  IV U2 ( .A(B[159]), .Z(n99) );
  IV U3 ( .A(B[160]), .Z(n98) );
  IV U4 ( .A(B[161]), .Z(n97) );
  IV U5 ( .A(B[162]), .Z(n96) );
  IV U6 ( .A(B[163]), .Z(n95) );
  IV U7 ( .A(B[164]), .Z(n94) );
  IV U8 ( .A(B[165]), .Z(n93) );
  IV U9 ( .A(B[166]), .Z(n92) );
  IV U10 ( .A(B[167]), .Z(n91) );
  IV U11 ( .A(B[168]), .Z(n90) );
  IV U12 ( .A(B[249]), .Z(n9) );
  IV U13 ( .A(B[169]), .Z(n89) );
  IV U14 ( .A(B[170]), .Z(n88) );
  IV U15 ( .A(B[171]), .Z(n87) );
  IV U16 ( .A(B[172]), .Z(n86) );
  IV U17 ( .A(B[173]), .Z(n85) );
  IV U18 ( .A(B[174]), .Z(n84) );
  IV U19 ( .A(B[175]), .Z(n83) );
  IV U20 ( .A(B[176]), .Z(n82) );
  IV U21 ( .A(B[177]), .Z(n81) );
  IV U22 ( .A(B[178]), .Z(n80) );
  IV U23 ( .A(B[250]), .Z(n8) );
  IV U24 ( .A(B[179]), .Z(n79) );
  IV U25 ( .A(B[180]), .Z(n78) );
  IV U26 ( .A(B[181]), .Z(n77) );
  IV U27 ( .A(B[182]), .Z(n76) );
  IV U28 ( .A(B[183]), .Z(n75) );
  IV U29 ( .A(B[184]), .Z(n74) );
  IV U30 ( .A(B[185]), .Z(n73) );
  IV U31 ( .A(B[186]), .Z(n72) );
  IV U32 ( .A(B[187]), .Z(n71) );
  IV U33 ( .A(B[188]), .Z(n70) );
  IV U34 ( .A(B[251]), .Z(n7) );
  IV U35 ( .A(B[189]), .Z(n69) );
  IV U36 ( .A(B[190]), .Z(n68) );
  IV U37 ( .A(B[191]), .Z(n67) );
  IV U38 ( .A(B[192]), .Z(n66) );
  IV U39 ( .A(B[193]), .Z(n65) );
  IV U40 ( .A(B[194]), .Z(n64) );
  IV U41 ( .A(B[195]), .Z(n63) );
  IV U42 ( .A(B[196]), .Z(n62) );
  IV U43 ( .A(B[197]), .Z(n61) );
  IV U44 ( .A(B[198]), .Z(n60) );
  IV U45 ( .A(B[252]), .Z(n6) );
  IV U46 ( .A(B[199]), .Z(n59) );
  IV U47 ( .A(B[200]), .Z(n58) );
  IV U48 ( .A(B[201]), .Z(n57) );
  IV U49 ( .A(B[202]), .Z(n56) );
  IV U50 ( .A(B[203]), .Z(n55) );
  IV U51 ( .A(B[204]), .Z(n54) );
  IV U52 ( .A(B[205]), .Z(n53) );
  IV U53 ( .A(B[206]), .Z(n52) );
  IV U54 ( .A(B[207]), .Z(n51) );
  IV U55 ( .A(B[208]), .Z(n50) );
  IV U56 ( .A(B[253]), .Z(n5) );
  IV U57 ( .A(B[209]), .Z(n49) );
  IV U58 ( .A(B[210]), .Z(n48) );
  IV U59 ( .A(B[211]), .Z(n47) );
  IV U60 ( .A(B[212]), .Z(n46) );
  IV U61 ( .A(B[213]), .Z(n45) );
  IV U62 ( .A(B[214]), .Z(n44) );
  IV U63 ( .A(B[215]), .Z(n43) );
  IV U64 ( .A(B[216]), .Z(n42) );
  IV U65 ( .A(B[217]), .Z(n41) );
  IV U66 ( .A(B[218]), .Z(n40) );
  IV U67 ( .A(B[254]), .Z(n4) );
  IV U68 ( .A(B[219]), .Z(n39) );
  IV U69 ( .A(B[220]), .Z(n38) );
  IV U70 ( .A(B[221]), .Z(n37) );
  IV U71 ( .A(B[222]), .Z(n36) );
  IV U72 ( .A(B[223]), .Z(n35) );
  IV U73 ( .A(B[224]), .Z(n34) );
  IV U74 ( .A(B[225]), .Z(n33) );
  IV U75 ( .A(B[226]), .Z(n32) );
  IV U76 ( .A(B[227]), .Z(n31) );
  IV U77 ( .A(B[228]), .Z(n30) );
  IV U78 ( .A(B[255]), .Z(n3) );
  IV U79 ( .A(B[229]), .Z(n29) );
  IV U80 ( .A(B[230]), .Z(n28) );
  IV U81 ( .A(B[231]), .Z(n27) );
  IV U82 ( .A(B[232]), .Z(n26) );
  IV U83 ( .A(B[0]), .Z(n258) );
  IV U84 ( .A(B[1]), .Z(n257) );
  IV U85 ( .A(B[2]), .Z(n256) );
  IV U86 ( .A(B[3]), .Z(n255) );
  IV U87 ( .A(B[4]), .Z(n254) );
  IV U88 ( .A(B[5]), .Z(n253) );
  IV U89 ( .A(B[6]), .Z(n252) );
  IV U90 ( .A(B[7]), .Z(n251) );
  IV U91 ( .A(B[8]), .Z(n250) );
  IV U92 ( .A(B[233]), .Z(n25) );
  IV U93 ( .A(B[9]), .Z(n249) );
  IV U94 ( .A(B[10]), .Z(n248) );
  IV U95 ( .A(B[11]), .Z(n247) );
  IV U96 ( .A(B[12]), .Z(n246) );
  IV U97 ( .A(B[13]), .Z(n245) );
  IV U98 ( .A(B[14]), .Z(n244) );
  IV U99 ( .A(B[15]), .Z(n243) );
  IV U100 ( .A(B[16]), .Z(n242) );
  IV U101 ( .A(B[17]), .Z(n241) );
  IV U102 ( .A(B[18]), .Z(n240) );
  IV U103 ( .A(B[234]), .Z(n24) );
  IV U104 ( .A(B[19]), .Z(n239) );
  IV U105 ( .A(B[20]), .Z(n238) );
  IV U106 ( .A(B[21]), .Z(n237) );
  IV U107 ( .A(B[22]), .Z(n236) );
  IV U108 ( .A(B[23]), .Z(n235) );
  IV U109 ( .A(B[24]), .Z(n234) );
  IV U110 ( .A(B[25]), .Z(n233) );
  IV U111 ( .A(B[26]), .Z(n232) );
  IV U112 ( .A(B[27]), .Z(n231) );
  IV U113 ( .A(B[28]), .Z(n230) );
  IV U114 ( .A(B[235]), .Z(n23) );
  IV U115 ( .A(B[29]), .Z(n229) );
  IV U116 ( .A(B[30]), .Z(n228) );
  IV U117 ( .A(B[31]), .Z(n227) );
  IV U118 ( .A(B[32]), .Z(n226) );
  IV U119 ( .A(B[33]), .Z(n225) );
  IV U120 ( .A(B[34]), .Z(n224) );
  IV U121 ( .A(B[35]), .Z(n223) );
  IV U122 ( .A(B[36]), .Z(n222) );
  IV U123 ( .A(B[37]), .Z(n221) );
  IV U124 ( .A(B[38]), .Z(n220) );
  IV U125 ( .A(B[236]), .Z(n22) );
  IV U126 ( .A(B[39]), .Z(n219) );
  IV U127 ( .A(B[40]), .Z(n218) );
  IV U128 ( .A(B[41]), .Z(n217) );
  IV U129 ( .A(B[42]), .Z(n216) );
  IV U130 ( .A(B[43]), .Z(n215) );
  IV U131 ( .A(B[44]), .Z(n214) );
  IV U132 ( .A(B[45]), .Z(n213) );
  IV U133 ( .A(B[46]), .Z(n212) );
  IV U134 ( .A(B[47]), .Z(n211) );
  IV U135 ( .A(B[48]), .Z(n210) );
  IV U136 ( .A(B[237]), .Z(n21) );
  IV U137 ( .A(B[49]), .Z(n209) );
  IV U138 ( .A(B[50]), .Z(n208) );
  IV U139 ( .A(B[51]), .Z(n207) );
  IV U140 ( .A(B[52]), .Z(n206) );
  IV U141 ( .A(B[53]), .Z(n205) );
  IV U142 ( .A(B[54]), .Z(n204) );
  IV U143 ( .A(B[55]), .Z(n203) );
  IV U144 ( .A(B[56]), .Z(n202) );
  IV U145 ( .A(B[57]), .Z(n201) );
  IV U146 ( .A(B[58]), .Z(n200) );
  IV U147 ( .A(B[238]), .Z(n20) );
  IV U148 ( .A(B[59]), .Z(n199) );
  IV U149 ( .A(B[60]), .Z(n198) );
  IV U150 ( .A(B[61]), .Z(n197) );
  IV U151 ( .A(B[62]), .Z(n196) );
  IV U152 ( .A(B[63]), .Z(n195) );
  IV U153 ( .A(B[64]), .Z(n194) );
  IV U154 ( .A(B[65]), .Z(n193) );
  IV U155 ( .A(B[66]), .Z(n192) );
  IV U156 ( .A(B[67]), .Z(n191) );
  IV U157 ( .A(B[68]), .Z(n190) );
  IV U158 ( .A(B[239]), .Z(n19) );
  IV U159 ( .A(B[69]), .Z(n189) );
  IV U160 ( .A(B[70]), .Z(n188) );
  IV U161 ( .A(B[71]), .Z(n187) );
  IV U162 ( .A(B[72]), .Z(n186) );
  IV U163 ( .A(B[73]), .Z(n185) );
  IV U164 ( .A(B[74]), .Z(n184) );
  IV U165 ( .A(B[75]), .Z(n183) );
  IV U166 ( .A(B[76]), .Z(n182) );
  IV U167 ( .A(B[77]), .Z(n181) );
  IV U168 ( .A(B[78]), .Z(n180) );
  IV U169 ( .A(B[240]), .Z(n18) );
  IV U170 ( .A(B[79]), .Z(n179) );
  IV U171 ( .A(B[80]), .Z(n178) );
  IV U172 ( .A(B[81]), .Z(n177) );
  IV U173 ( .A(B[82]), .Z(n176) );
  IV U174 ( .A(B[83]), .Z(n175) );
  IV U175 ( .A(B[84]), .Z(n174) );
  IV U176 ( .A(B[85]), .Z(n173) );
  IV U177 ( .A(B[86]), .Z(n172) );
  IV U178 ( .A(B[87]), .Z(n171) );
  IV U179 ( .A(B[88]), .Z(n170) );
  IV U180 ( .A(B[241]), .Z(n17) );
  IV U181 ( .A(B[89]), .Z(n169) );
  IV U182 ( .A(B[90]), .Z(n168) );
  IV U183 ( .A(B[91]), .Z(n167) );
  IV U184 ( .A(B[92]), .Z(n166) );
  IV U185 ( .A(B[93]), .Z(n165) );
  IV U186 ( .A(B[94]), .Z(n164) );
  IV U187 ( .A(B[95]), .Z(n163) );
  IV U188 ( .A(B[96]), .Z(n162) );
  IV U189 ( .A(B[97]), .Z(n161) );
  IV U190 ( .A(B[98]), .Z(n160) );
  IV U191 ( .A(B[242]), .Z(n16) );
  IV U192 ( .A(B[99]), .Z(n159) );
  IV U193 ( .A(B[100]), .Z(n158) );
  IV U194 ( .A(B[101]), .Z(n157) );
  IV U195 ( .A(B[102]), .Z(n156) );
  IV U196 ( .A(B[103]), .Z(n155) );
  IV U197 ( .A(B[104]), .Z(n154) );
  IV U198 ( .A(B[105]), .Z(n153) );
  IV U199 ( .A(B[106]), .Z(n152) );
  IV U200 ( .A(B[107]), .Z(n151) );
  IV U201 ( .A(B[108]), .Z(n150) );
  IV U202 ( .A(B[243]), .Z(n15) );
  IV U203 ( .A(B[109]), .Z(n149) );
  IV U204 ( .A(B[110]), .Z(n148) );
  IV U205 ( .A(B[111]), .Z(n147) );
  IV U206 ( .A(B[112]), .Z(n146) );
  IV U207 ( .A(B[113]), .Z(n145) );
  IV U208 ( .A(B[114]), .Z(n144) );
  IV U209 ( .A(B[115]), .Z(n143) );
  IV U210 ( .A(B[116]), .Z(n142) );
  IV U211 ( .A(B[117]), .Z(n141) );
  IV U212 ( .A(B[118]), .Z(n140) );
  IV U213 ( .A(B[244]), .Z(n14) );
  IV U214 ( .A(B[119]), .Z(n139) );
  IV U215 ( .A(B[120]), .Z(n138) );
  IV U216 ( .A(B[121]), .Z(n137) );
  IV U217 ( .A(B[122]), .Z(n136) );
  IV U218 ( .A(B[123]), .Z(n135) );
  IV U219 ( .A(B[124]), .Z(n134) );
  IV U220 ( .A(B[125]), .Z(n133) );
  IV U221 ( .A(B[126]), .Z(n132) );
  IV U222 ( .A(B[127]), .Z(n131) );
  IV U223 ( .A(B[128]), .Z(n130) );
  IV U224 ( .A(B[245]), .Z(n13) );
  IV U225 ( .A(B[129]), .Z(n129) );
  IV U226 ( .A(B[130]), .Z(n128) );
  IV U227 ( .A(B[131]), .Z(n127) );
  IV U228 ( .A(B[132]), .Z(n126) );
  IV U229 ( .A(B[133]), .Z(n125) );
  IV U230 ( .A(B[134]), .Z(n124) );
  IV U231 ( .A(B[135]), .Z(n123) );
  IV U232 ( .A(B[136]), .Z(n122) );
  IV U233 ( .A(B[137]), .Z(n121) );
  IV U234 ( .A(B[138]), .Z(n120) );
  IV U235 ( .A(B[246]), .Z(n12) );
  IV U236 ( .A(B[139]), .Z(n119) );
  IV U237 ( .A(B[140]), .Z(n118) );
  IV U238 ( .A(B[141]), .Z(n117) );
  IV U239 ( .A(B[142]), .Z(n116) );
  IV U240 ( .A(B[143]), .Z(n115) );
  IV U241 ( .A(B[144]), .Z(n114) );
  IV U242 ( .A(B[145]), .Z(n113) );
  IV U243 ( .A(B[146]), .Z(n112) );
  IV U244 ( .A(B[147]), .Z(n111) );
  IV U245 ( .A(B[148]), .Z(n110) );
  IV U246 ( .A(B[247]), .Z(n11) );
  IV U247 ( .A(B[149]), .Z(n109) );
  IV U248 ( .A(B[150]), .Z(n108) );
  IV U249 ( .A(B[151]), .Z(n107) );
  IV U250 ( .A(B[152]), .Z(n106) );
  IV U251 ( .A(B[153]), .Z(n105) );
  IV U252 ( .A(B[154]), .Z(n104) );
  IV U253 ( .A(B[155]), .Z(n103) );
  IV U254 ( .A(B[156]), .Z(n102) );
  IV U255 ( .A(B[157]), .Z(n101) );
  IV U256 ( .A(B[158]), .Z(n100) );
  IV U257 ( .A(B[248]), .Z(n10) );
endmodule


module MUX_N258_1 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N258_2 ( A, B, S, O );
  input [257:0] A;
  input [257:0] B;
  output [257:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U56 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U57 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U58 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U59 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U60 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U61 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U62 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U63 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U64 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U65 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U66 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U67 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U68 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U69 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U70 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U71 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U72 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U73 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U74 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U75 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U76 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U77 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U78 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U79 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U80 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U81 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U82 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U83 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U84 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U85 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U86 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U87 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U88 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U89 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U90 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U91 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U92 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U93 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U94 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U95 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U96 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U97 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U98 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U99 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U100 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U101 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U102 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U103 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U104 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U105 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U106 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U107 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U108 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U109 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U110 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U111 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U112 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U113 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U114 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U115 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U116 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U117 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U118 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U119 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U120 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U121 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U122 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U123 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U124 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U125 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U126 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U127 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U128 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U129 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U130 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U131 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U132 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U133 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U134 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U135 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U136 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U137 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U138 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U139 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U140 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U141 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U142 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U143 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U144 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U145 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U146 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U147 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U148 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U149 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U150 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U151 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U152 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U153 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U154 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U155 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U156 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U157 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U158 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U159 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U160 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U161 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U162 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U163 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U164 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U165 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U166 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U167 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U168 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U169 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U170 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U171 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U172 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U173 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U174 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U175 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U176 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U177 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U178 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U179 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U180 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U181 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U182 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U183 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U184 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U185 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U186 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U187 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U188 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U189 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U190 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U191 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U192 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U193 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U194 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U195 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U196 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U197 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U198 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U199 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U200 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U201 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U202 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U203 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U204 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U205 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U206 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U207 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U208 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U209 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U210 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U211 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U212 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U213 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U214 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U215 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U216 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U217 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U218 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U219 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U220 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U221 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U222 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U223 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U224 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U225 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U226 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U227 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U228 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U229 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U230 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U231 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U232 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U233 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U234 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U235 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U236 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U237 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U238 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U239 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U240 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U241 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U242 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U243 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U244 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U245 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U246 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U247 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U248 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U249 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U250 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U251 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U252 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U253 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U254 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U255 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U256 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N258_1 ( A, B, O );
  input [257:0] A;
  input [257:0] B;
  output O;
  wire   n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517;
  wire   [257:1] C;

  FA_516 \FAINST[0].FA_  ( .A(A[0]), .B(n260), .CI(1'b1), .CO(C[1]) );
  FA_515 \FAINST[1].FA_  ( .A(A[1]), .B(n261), .CI(C[1]), .CO(C[2]) );
  FA_514 \FAINST[2].FA_  ( .A(A[2]), .B(n262), .CI(C[2]), .CO(C[3]) );
  FA_513 \FAINST[3].FA_  ( .A(A[3]), .B(n263), .CI(C[3]), .CO(C[4]) );
  FA_512 \FAINST[4].FA_  ( .A(A[4]), .B(n264), .CI(C[4]), .CO(C[5]) );
  FA_511 \FAINST[5].FA_  ( .A(A[5]), .B(n265), .CI(C[5]), .CO(C[6]) );
  FA_510 \FAINST[6].FA_  ( .A(A[6]), .B(n266), .CI(C[6]), .CO(C[7]) );
  FA_509 \FAINST[7].FA_  ( .A(A[7]), .B(n267), .CI(C[7]), .CO(C[8]) );
  FA_508 \FAINST[8].FA_  ( .A(A[8]), .B(n268), .CI(C[8]), .CO(C[9]) );
  FA_507 \FAINST[9].FA_  ( .A(A[9]), .B(n269), .CI(C[9]), .CO(C[10]) );
  FA_506 \FAINST[10].FA_  ( .A(A[10]), .B(n270), .CI(C[10]), .CO(C[11]) );
  FA_505 \FAINST[11].FA_  ( .A(A[11]), .B(n271), .CI(C[11]), .CO(C[12]) );
  FA_504 \FAINST[12].FA_  ( .A(A[12]), .B(n272), .CI(C[12]), .CO(C[13]) );
  FA_503 \FAINST[13].FA_  ( .A(A[13]), .B(n273), .CI(C[13]), .CO(C[14]) );
  FA_502 \FAINST[14].FA_  ( .A(A[14]), .B(n274), .CI(C[14]), .CO(C[15]) );
  FA_501 \FAINST[15].FA_  ( .A(A[15]), .B(n275), .CI(C[15]), .CO(C[16]) );
  FA_500 \FAINST[16].FA_  ( .A(A[16]), .B(n276), .CI(C[16]), .CO(C[17]) );
  FA_499 \FAINST[17].FA_  ( .A(A[17]), .B(n277), .CI(C[17]), .CO(C[18]) );
  FA_498 \FAINST[18].FA_  ( .A(A[18]), .B(n278), .CI(C[18]), .CO(C[19]) );
  FA_497 \FAINST[19].FA_  ( .A(A[19]), .B(n279), .CI(C[19]), .CO(C[20]) );
  FA_496 \FAINST[20].FA_  ( .A(A[20]), .B(n280), .CI(C[20]), .CO(C[21]) );
  FA_495 \FAINST[21].FA_  ( .A(A[21]), .B(n281), .CI(C[21]), .CO(C[22]) );
  FA_494 \FAINST[22].FA_  ( .A(A[22]), .B(n282), .CI(C[22]), .CO(C[23]) );
  FA_493 \FAINST[23].FA_  ( .A(A[23]), .B(n283), .CI(C[23]), .CO(C[24]) );
  FA_492 \FAINST[24].FA_  ( .A(A[24]), .B(n284), .CI(C[24]), .CO(C[25]) );
  FA_491 \FAINST[25].FA_  ( .A(A[25]), .B(n285), .CI(C[25]), .CO(C[26]) );
  FA_490 \FAINST[26].FA_  ( .A(A[26]), .B(n286), .CI(C[26]), .CO(C[27]) );
  FA_489 \FAINST[27].FA_  ( .A(A[27]), .B(n287), .CI(C[27]), .CO(C[28]) );
  FA_488 \FAINST[28].FA_  ( .A(A[28]), .B(n288), .CI(C[28]), .CO(C[29]) );
  FA_487 \FAINST[29].FA_  ( .A(A[29]), .B(n289), .CI(C[29]), .CO(C[30]) );
  FA_486 \FAINST[30].FA_  ( .A(A[30]), .B(n290), .CI(C[30]), .CO(C[31]) );
  FA_485 \FAINST[31].FA_  ( .A(A[31]), .B(n291), .CI(C[31]), .CO(C[32]) );
  FA_484 \FAINST[32].FA_  ( .A(A[32]), .B(n292), .CI(C[32]), .CO(C[33]) );
  FA_483 \FAINST[33].FA_  ( .A(A[33]), .B(n293), .CI(C[33]), .CO(C[34]) );
  FA_482 \FAINST[34].FA_  ( .A(A[34]), .B(n294), .CI(C[34]), .CO(C[35]) );
  FA_481 \FAINST[35].FA_  ( .A(A[35]), .B(n295), .CI(C[35]), .CO(C[36]) );
  FA_480 \FAINST[36].FA_  ( .A(A[36]), .B(n296), .CI(C[36]), .CO(C[37]) );
  FA_479 \FAINST[37].FA_  ( .A(A[37]), .B(n297), .CI(C[37]), .CO(C[38]) );
  FA_478 \FAINST[38].FA_  ( .A(A[38]), .B(n298), .CI(C[38]), .CO(C[39]) );
  FA_477 \FAINST[39].FA_  ( .A(A[39]), .B(n299), .CI(C[39]), .CO(C[40]) );
  FA_476 \FAINST[40].FA_  ( .A(A[40]), .B(n300), .CI(C[40]), .CO(C[41]) );
  FA_475 \FAINST[41].FA_  ( .A(A[41]), .B(n301), .CI(C[41]), .CO(C[42]) );
  FA_474 \FAINST[42].FA_  ( .A(A[42]), .B(n302), .CI(C[42]), .CO(C[43]) );
  FA_473 \FAINST[43].FA_  ( .A(A[43]), .B(n303), .CI(C[43]), .CO(C[44]) );
  FA_472 \FAINST[44].FA_  ( .A(A[44]), .B(n304), .CI(C[44]), .CO(C[45]) );
  FA_471 \FAINST[45].FA_  ( .A(A[45]), .B(n305), .CI(C[45]), .CO(C[46]) );
  FA_470 \FAINST[46].FA_  ( .A(A[46]), .B(n306), .CI(C[46]), .CO(C[47]) );
  FA_469 \FAINST[47].FA_  ( .A(A[47]), .B(n307), .CI(C[47]), .CO(C[48]) );
  FA_468 \FAINST[48].FA_  ( .A(A[48]), .B(n308), .CI(C[48]), .CO(C[49]) );
  FA_467 \FAINST[49].FA_  ( .A(A[49]), .B(n309), .CI(C[49]), .CO(C[50]) );
  FA_466 \FAINST[50].FA_  ( .A(A[50]), .B(n310), .CI(C[50]), .CO(C[51]) );
  FA_465 \FAINST[51].FA_  ( .A(A[51]), .B(n311), .CI(C[51]), .CO(C[52]) );
  FA_464 \FAINST[52].FA_  ( .A(A[52]), .B(n312), .CI(C[52]), .CO(C[53]) );
  FA_463 \FAINST[53].FA_  ( .A(A[53]), .B(n313), .CI(C[53]), .CO(C[54]) );
  FA_462 \FAINST[54].FA_  ( .A(A[54]), .B(n314), .CI(C[54]), .CO(C[55]) );
  FA_461 \FAINST[55].FA_  ( .A(A[55]), .B(n315), .CI(C[55]), .CO(C[56]) );
  FA_460 \FAINST[56].FA_  ( .A(A[56]), .B(n316), .CI(C[56]), .CO(C[57]) );
  FA_459 \FAINST[57].FA_  ( .A(A[57]), .B(n317), .CI(C[57]), .CO(C[58]) );
  FA_458 \FAINST[58].FA_  ( .A(A[58]), .B(n318), .CI(C[58]), .CO(C[59]) );
  FA_457 \FAINST[59].FA_  ( .A(A[59]), .B(n319), .CI(C[59]), .CO(C[60]) );
  FA_456 \FAINST[60].FA_  ( .A(A[60]), .B(n320), .CI(C[60]), .CO(C[61]) );
  FA_455 \FAINST[61].FA_  ( .A(A[61]), .B(n321), .CI(C[61]), .CO(C[62]) );
  FA_454 \FAINST[62].FA_  ( .A(A[62]), .B(n322), .CI(C[62]), .CO(C[63]) );
  FA_453 \FAINST[63].FA_  ( .A(A[63]), .B(n323), .CI(C[63]), .CO(C[64]) );
  FA_452 \FAINST[64].FA_  ( .A(A[64]), .B(n324), .CI(C[64]), .CO(C[65]) );
  FA_451 \FAINST[65].FA_  ( .A(A[65]), .B(n325), .CI(C[65]), .CO(C[66]) );
  FA_450 \FAINST[66].FA_  ( .A(A[66]), .B(n326), .CI(C[66]), .CO(C[67]) );
  FA_449 \FAINST[67].FA_  ( .A(A[67]), .B(n327), .CI(C[67]), .CO(C[68]) );
  FA_448 \FAINST[68].FA_  ( .A(A[68]), .B(n328), .CI(C[68]), .CO(C[69]) );
  FA_447 \FAINST[69].FA_  ( .A(A[69]), .B(n329), .CI(C[69]), .CO(C[70]) );
  FA_446 \FAINST[70].FA_  ( .A(A[70]), .B(n330), .CI(C[70]), .CO(C[71]) );
  FA_445 \FAINST[71].FA_  ( .A(A[71]), .B(n331), .CI(C[71]), .CO(C[72]) );
  FA_444 \FAINST[72].FA_  ( .A(A[72]), .B(n332), .CI(C[72]), .CO(C[73]) );
  FA_443 \FAINST[73].FA_  ( .A(A[73]), .B(n333), .CI(C[73]), .CO(C[74]) );
  FA_442 \FAINST[74].FA_  ( .A(A[74]), .B(n334), .CI(C[74]), .CO(C[75]) );
  FA_441 \FAINST[75].FA_  ( .A(A[75]), .B(n335), .CI(C[75]), .CO(C[76]) );
  FA_440 \FAINST[76].FA_  ( .A(A[76]), .B(n336), .CI(C[76]), .CO(C[77]) );
  FA_439 \FAINST[77].FA_  ( .A(A[77]), .B(n337), .CI(C[77]), .CO(C[78]) );
  FA_438 \FAINST[78].FA_  ( .A(A[78]), .B(n338), .CI(C[78]), .CO(C[79]) );
  FA_437 \FAINST[79].FA_  ( .A(A[79]), .B(n339), .CI(C[79]), .CO(C[80]) );
  FA_436 \FAINST[80].FA_  ( .A(A[80]), .B(n340), .CI(C[80]), .CO(C[81]) );
  FA_435 \FAINST[81].FA_  ( .A(A[81]), .B(n341), .CI(C[81]), .CO(C[82]) );
  FA_434 \FAINST[82].FA_  ( .A(A[82]), .B(n342), .CI(C[82]), .CO(C[83]) );
  FA_433 \FAINST[83].FA_  ( .A(A[83]), .B(n343), .CI(C[83]), .CO(C[84]) );
  FA_432 \FAINST[84].FA_  ( .A(A[84]), .B(n344), .CI(C[84]), .CO(C[85]) );
  FA_431 \FAINST[85].FA_  ( .A(A[85]), .B(n345), .CI(C[85]), .CO(C[86]) );
  FA_430 \FAINST[86].FA_  ( .A(A[86]), .B(n346), .CI(C[86]), .CO(C[87]) );
  FA_429 \FAINST[87].FA_  ( .A(A[87]), .B(n347), .CI(C[87]), .CO(C[88]) );
  FA_428 \FAINST[88].FA_  ( .A(A[88]), .B(n348), .CI(C[88]), .CO(C[89]) );
  FA_427 \FAINST[89].FA_  ( .A(A[89]), .B(n349), .CI(C[89]), .CO(C[90]) );
  FA_426 \FAINST[90].FA_  ( .A(A[90]), .B(n350), .CI(C[90]), .CO(C[91]) );
  FA_425 \FAINST[91].FA_  ( .A(A[91]), .B(n351), .CI(C[91]), .CO(C[92]) );
  FA_424 \FAINST[92].FA_  ( .A(A[92]), .B(n352), .CI(C[92]), .CO(C[93]) );
  FA_423 \FAINST[93].FA_  ( .A(A[93]), .B(n353), .CI(C[93]), .CO(C[94]) );
  FA_422 \FAINST[94].FA_  ( .A(A[94]), .B(n354), .CI(C[94]), .CO(C[95]) );
  FA_421 \FAINST[95].FA_  ( .A(A[95]), .B(n355), .CI(C[95]), .CO(C[96]) );
  FA_420 \FAINST[96].FA_  ( .A(A[96]), .B(n356), .CI(C[96]), .CO(C[97]) );
  FA_419 \FAINST[97].FA_  ( .A(A[97]), .B(n357), .CI(C[97]), .CO(C[98]) );
  FA_418 \FAINST[98].FA_  ( .A(A[98]), .B(n358), .CI(C[98]), .CO(C[99]) );
  FA_417 \FAINST[99].FA_  ( .A(A[99]), .B(n359), .CI(C[99]), .CO(C[100]) );
  FA_416 \FAINST[100].FA_  ( .A(A[100]), .B(n360), .CI(C[100]), .CO(C[101]) );
  FA_415 \FAINST[101].FA_  ( .A(A[101]), .B(n361), .CI(C[101]), .CO(C[102]) );
  FA_414 \FAINST[102].FA_  ( .A(A[102]), .B(n362), .CI(C[102]), .CO(C[103]) );
  FA_413 \FAINST[103].FA_  ( .A(A[103]), .B(n363), .CI(C[103]), .CO(C[104]) );
  FA_412 \FAINST[104].FA_  ( .A(A[104]), .B(n364), .CI(C[104]), .CO(C[105]) );
  FA_411 \FAINST[105].FA_  ( .A(A[105]), .B(n365), .CI(C[105]), .CO(C[106]) );
  FA_410 \FAINST[106].FA_  ( .A(A[106]), .B(n366), .CI(C[106]), .CO(C[107]) );
  FA_409 \FAINST[107].FA_  ( .A(A[107]), .B(n367), .CI(C[107]), .CO(C[108]) );
  FA_408 \FAINST[108].FA_  ( .A(A[108]), .B(n368), .CI(C[108]), .CO(C[109]) );
  FA_407 \FAINST[109].FA_  ( .A(A[109]), .B(n369), .CI(C[109]), .CO(C[110]) );
  FA_406 \FAINST[110].FA_  ( .A(A[110]), .B(n370), .CI(C[110]), .CO(C[111]) );
  FA_405 \FAINST[111].FA_  ( .A(A[111]), .B(n371), .CI(C[111]), .CO(C[112]) );
  FA_404 \FAINST[112].FA_  ( .A(A[112]), .B(n372), .CI(C[112]), .CO(C[113]) );
  FA_403 \FAINST[113].FA_  ( .A(A[113]), .B(n373), .CI(C[113]), .CO(C[114]) );
  FA_402 \FAINST[114].FA_  ( .A(A[114]), .B(n374), .CI(C[114]), .CO(C[115]) );
  FA_401 \FAINST[115].FA_  ( .A(A[115]), .B(n375), .CI(C[115]), .CO(C[116]) );
  FA_400 \FAINST[116].FA_  ( .A(A[116]), .B(n376), .CI(C[116]), .CO(C[117]) );
  FA_399 \FAINST[117].FA_  ( .A(A[117]), .B(n377), .CI(C[117]), .CO(C[118]) );
  FA_398 \FAINST[118].FA_  ( .A(A[118]), .B(n378), .CI(C[118]), .CO(C[119]) );
  FA_397 \FAINST[119].FA_  ( .A(A[119]), .B(n379), .CI(C[119]), .CO(C[120]) );
  FA_396 \FAINST[120].FA_  ( .A(A[120]), .B(n380), .CI(C[120]), .CO(C[121]) );
  FA_395 \FAINST[121].FA_  ( .A(A[121]), .B(n381), .CI(C[121]), .CO(C[122]) );
  FA_394 \FAINST[122].FA_  ( .A(A[122]), .B(n382), .CI(C[122]), .CO(C[123]) );
  FA_393 \FAINST[123].FA_  ( .A(A[123]), .B(n383), .CI(C[123]), .CO(C[124]) );
  FA_392 \FAINST[124].FA_  ( .A(A[124]), .B(n384), .CI(C[124]), .CO(C[125]) );
  FA_391 \FAINST[125].FA_  ( .A(A[125]), .B(n385), .CI(C[125]), .CO(C[126]) );
  FA_390 \FAINST[126].FA_  ( .A(A[126]), .B(n386), .CI(C[126]), .CO(C[127]) );
  FA_389 \FAINST[127].FA_  ( .A(A[127]), .B(n387), .CI(C[127]), .CO(C[128]) );
  FA_388 \FAINST[128].FA_  ( .A(A[128]), .B(n388), .CI(C[128]), .CO(C[129]) );
  FA_387 \FAINST[129].FA_  ( .A(A[129]), .B(n389), .CI(C[129]), .CO(C[130]) );
  FA_386 \FAINST[130].FA_  ( .A(A[130]), .B(n390), .CI(C[130]), .CO(C[131]) );
  FA_385 \FAINST[131].FA_  ( .A(A[131]), .B(n391), .CI(C[131]), .CO(C[132]) );
  FA_384 \FAINST[132].FA_  ( .A(A[132]), .B(n392), .CI(C[132]), .CO(C[133]) );
  FA_383 \FAINST[133].FA_  ( .A(A[133]), .B(n393), .CI(C[133]), .CO(C[134]) );
  FA_382 \FAINST[134].FA_  ( .A(A[134]), .B(n394), .CI(C[134]), .CO(C[135]) );
  FA_381 \FAINST[135].FA_  ( .A(A[135]), .B(n395), .CI(C[135]), .CO(C[136]) );
  FA_380 \FAINST[136].FA_  ( .A(A[136]), .B(n396), .CI(C[136]), .CO(C[137]) );
  FA_379 \FAINST[137].FA_  ( .A(A[137]), .B(n397), .CI(C[137]), .CO(C[138]) );
  FA_378 \FAINST[138].FA_  ( .A(A[138]), .B(n398), .CI(C[138]), .CO(C[139]) );
  FA_377 \FAINST[139].FA_  ( .A(A[139]), .B(n399), .CI(C[139]), .CO(C[140]) );
  FA_376 \FAINST[140].FA_  ( .A(A[140]), .B(n400), .CI(C[140]), .CO(C[141]) );
  FA_375 \FAINST[141].FA_  ( .A(A[141]), .B(n401), .CI(C[141]), .CO(C[142]) );
  FA_374 \FAINST[142].FA_  ( .A(A[142]), .B(n402), .CI(C[142]), .CO(C[143]) );
  FA_373 \FAINST[143].FA_  ( .A(A[143]), .B(n403), .CI(C[143]), .CO(C[144]) );
  FA_372 \FAINST[144].FA_  ( .A(A[144]), .B(n404), .CI(C[144]), .CO(C[145]) );
  FA_371 \FAINST[145].FA_  ( .A(A[145]), .B(n405), .CI(C[145]), .CO(C[146]) );
  FA_370 \FAINST[146].FA_  ( .A(A[146]), .B(n406), .CI(C[146]), .CO(C[147]) );
  FA_369 \FAINST[147].FA_  ( .A(A[147]), .B(n407), .CI(C[147]), .CO(C[148]) );
  FA_368 \FAINST[148].FA_  ( .A(A[148]), .B(n408), .CI(C[148]), .CO(C[149]) );
  FA_367 \FAINST[149].FA_  ( .A(A[149]), .B(n409), .CI(C[149]), .CO(C[150]) );
  FA_366 \FAINST[150].FA_  ( .A(A[150]), .B(n410), .CI(C[150]), .CO(C[151]) );
  FA_365 \FAINST[151].FA_  ( .A(A[151]), .B(n411), .CI(C[151]), .CO(C[152]) );
  FA_364 \FAINST[152].FA_  ( .A(A[152]), .B(n412), .CI(C[152]), .CO(C[153]) );
  FA_363 \FAINST[153].FA_  ( .A(A[153]), .B(n413), .CI(C[153]), .CO(C[154]) );
  FA_362 \FAINST[154].FA_  ( .A(A[154]), .B(n414), .CI(C[154]), .CO(C[155]) );
  FA_361 \FAINST[155].FA_  ( .A(A[155]), .B(n415), .CI(C[155]), .CO(C[156]) );
  FA_360 \FAINST[156].FA_  ( .A(A[156]), .B(n416), .CI(C[156]), .CO(C[157]) );
  FA_359 \FAINST[157].FA_  ( .A(A[157]), .B(n417), .CI(C[157]), .CO(C[158]) );
  FA_358 \FAINST[158].FA_  ( .A(A[158]), .B(n418), .CI(C[158]), .CO(C[159]) );
  FA_357 \FAINST[159].FA_  ( .A(A[159]), .B(n419), .CI(C[159]), .CO(C[160]) );
  FA_356 \FAINST[160].FA_  ( .A(A[160]), .B(n420), .CI(C[160]), .CO(C[161]) );
  FA_355 \FAINST[161].FA_  ( .A(A[161]), .B(n421), .CI(C[161]), .CO(C[162]) );
  FA_354 \FAINST[162].FA_  ( .A(A[162]), .B(n422), .CI(C[162]), .CO(C[163]) );
  FA_353 \FAINST[163].FA_  ( .A(A[163]), .B(n423), .CI(C[163]), .CO(C[164]) );
  FA_352 \FAINST[164].FA_  ( .A(A[164]), .B(n424), .CI(C[164]), .CO(C[165]) );
  FA_351 \FAINST[165].FA_  ( .A(A[165]), .B(n425), .CI(C[165]), .CO(C[166]) );
  FA_350 \FAINST[166].FA_  ( .A(A[166]), .B(n426), .CI(C[166]), .CO(C[167]) );
  FA_349 \FAINST[167].FA_  ( .A(A[167]), .B(n427), .CI(C[167]), .CO(C[168]) );
  FA_348 \FAINST[168].FA_  ( .A(A[168]), .B(n428), .CI(C[168]), .CO(C[169]) );
  FA_347 \FAINST[169].FA_  ( .A(A[169]), .B(n429), .CI(C[169]), .CO(C[170]) );
  FA_346 \FAINST[170].FA_  ( .A(A[170]), .B(n430), .CI(C[170]), .CO(C[171]) );
  FA_345 \FAINST[171].FA_  ( .A(A[171]), .B(n431), .CI(C[171]), .CO(C[172]) );
  FA_344 \FAINST[172].FA_  ( .A(A[172]), .B(n432), .CI(C[172]), .CO(C[173]) );
  FA_343 \FAINST[173].FA_  ( .A(A[173]), .B(n433), .CI(C[173]), .CO(C[174]) );
  FA_342 \FAINST[174].FA_  ( .A(A[174]), .B(n434), .CI(C[174]), .CO(C[175]) );
  FA_341 \FAINST[175].FA_  ( .A(A[175]), .B(n435), .CI(C[175]), .CO(C[176]) );
  FA_340 \FAINST[176].FA_  ( .A(A[176]), .B(n436), .CI(C[176]), .CO(C[177]) );
  FA_339 \FAINST[177].FA_  ( .A(A[177]), .B(n437), .CI(C[177]), .CO(C[178]) );
  FA_338 \FAINST[178].FA_  ( .A(A[178]), .B(n438), .CI(C[178]), .CO(C[179]) );
  FA_337 \FAINST[179].FA_  ( .A(A[179]), .B(n439), .CI(C[179]), .CO(C[180]) );
  FA_336 \FAINST[180].FA_  ( .A(A[180]), .B(n440), .CI(C[180]), .CO(C[181]) );
  FA_335 \FAINST[181].FA_  ( .A(A[181]), .B(n441), .CI(C[181]), .CO(C[182]) );
  FA_334 \FAINST[182].FA_  ( .A(A[182]), .B(n442), .CI(C[182]), .CO(C[183]) );
  FA_333 \FAINST[183].FA_  ( .A(A[183]), .B(n443), .CI(C[183]), .CO(C[184]) );
  FA_332 \FAINST[184].FA_  ( .A(A[184]), .B(n444), .CI(C[184]), .CO(C[185]) );
  FA_331 \FAINST[185].FA_  ( .A(A[185]), .B(n445), .CI(C[185]), .CO(C[186]) );
  FA_330 \FAINST[186].FA_  ( .A(A[186]), .B(n446), .CI(C[186]), .CO(C[187]) );
  FA_329 \FAINST[187].FA_  ( .A(A[187]), .B(n447), .CI(C[187]), .CO(C[188]) );
  FA_328 \FAINST[188].FA_  ( .A(A[188]), .B(n448), .CI(C[188]), .CO(C[189]) );
  FA_327 \FAINST[189].FA_  ( .A(A[189]), .B(n449), .CI(C[189]), .CO(C[190]) );
  FA_326 \FAINST[190].FA_  ( .A(A[190]), .B(n450), .CI(C[190]), .CO(C[191]) );
  FA_325 \FAINST[191].FA_  ( .A(A[191]), .B(n451), .CI(C[191]), .CO(C[192]) );
  FA_324 \FAINST[192].FA_  ( .A(A[192]), .B(n452), .CI(C[192]), .CO(C[193]) );
  FA_323 \FAINST[193].FA_  ( .A(A[193]), .B(n453), .CI(C[193]), .CO(C[194]) );
  FA_322 \FAINST[194].FA_  ( .A(A[194]), .B(n454), .CI(C[194]), .CO(C[195]) );
  FA_321 \FAINST[195].FA_  ( .A(A[195]), .B(n455), .CI(C[195]), .CO(C[196]) );
  FA_320 \FAINST[196].FA_  ( .A(A[196]), .B(n456), .CI(C[196]), .CO(C[197]) );
  FA_319 \FAINST[197].FA_  ( .A(A[197]), .B(n457), .CI(C[197]), .CO(C[198]) );
  FA_318 \FAINST[198].FA_  ( .A(A[198]), .B(n458), .CI(C[198]), .CO(C[199]) );
  FA_317 \FAINST[199].FA_  ( .A(A[199]), .B(n459), .CI(C[199]), .CO(C[200]) );
  FA_316 \FAINST[200].FA_  ( .A(A[200]), .B(n460), .CI(C[200]), .CO(C[201]) );
  FA_315 \FAINST[201].FA_  ( .A(A[201]), .B(n461), .CI(C[201]), .CO(C[202]) );
  FA_314 \FAINST[202].FA_  ( .A(A[202]), .B(n462), .CI(C[202]), .CO(C[203]) );
  FA_313 \FAINST[203].FA_  ( .A(A[203]), .B(n463), .CI(C[203]), .CO(C[204]) );
  FA_312 \FAINST[204].FA_  ( .A(A[204]), .B(n464), .CI(C[204]), .CO(C[205]) );
  FA_311 \FAINST[205].FA_  ( .A(A[205]), .B(n465), .CI(C[205]), .CO(C[206]) );
  FA_310 \FAINST[206].FA_  ( .A(A[206]), .B(n466), .CI(C[206]), .CO(C[207]) );
  FA_309 \FAINST[207].FA_  ( .A(A[207]), .B(n467), .CI(C[207]), .CO(C[208]) );
  FA_308 \FAINST[208].FA_  ( .A(A[208]), .B(n468), .CI(C[208]), .CO(C[209]) );
  FA_307 \FAINST[209].FA_  ( .A(A[209]), .B(n469), .CI(C[209]), .CO(C[210]) );
  FA_306 \FAINST[210].FA_  ( .A(A[210]), .B(n470), .CI(C[210]), .CO(C[211]) );
  FA_305 \FAINST[211].FA_  ( .A(A[211]), .B(n471), .CI(C[211]), .CO(C[212]) );
  FA_304 \FAINST[212].FA_  ( .A(A[212]), .B(n472), .CI(C[212]), .CO(C[213]) );
  FA_303 \FAINST[213].FA_  ( .A(A[213]), .B(n473), .CI(C[213]), .CO(C[214]) );
  FA_302 \FAINST[214].FA_  ( .A(A[214]), .B(n474), .CI(C[214]), .CO(C[215]) );
  FA_301 \FAINST[215].FA_  ( .A(A[215]), .B(n475), .CI(C[215]), .CO(C[216]) );
  FA_300 \FAINST[216].FA_  ( .A(A[216]), .B(n476), .CI(C[216]), .CO(C[217]) );
  FA_299 \FAINST[217].FA_  ( .A(A[217]), .B(n477), .CI(C[217]), .CO(C[218]) );
  FA_298 \FAINST[218].FA_  ( .A(A[218]), .B(n478), .CI(C[218]), .CO(C[219]) );
  FA_297 \FAINST[219].FA_  ( .A(A[219]), .B(n479), .CI(C[219]), .CO(C[220]) );
  FA_296 \FAINST[220].FA_  ( .A(A[220]), .B(n480), .CI(C[220]), .CO(C[221]) );
  FA_295 \FAINST[221].FA_  ( .A(A[221]), .B(n481), .CI(C[221]), .CO(C[222]) );
  FA_294 \FAINST[222].FA_  ( .A(A[222]), .B(n482), .CI(C[222]), .CO(C[223]) );
  FA_293 \FAINST[223].FA_  ( .A(A[223]), .B(n483), .CI(C[223]), .CO(C[224]) );
  FA_292 \FAINST[224].FA_  ( .A(A[224]), .B(n484), .CI(C[224]), .CO(C[225]) );
  FA_291 \FAINST[225].FA_  ( .A(A[225]), .B(n485), .CI(C[225]), .CO(C[226]) );
  FA_290 \FAINST[226].FA_  ( .A(A[226]), .B(n486), .CI(C[226]), .CO(C[227]) );
  FA_289 \FAINST[227].FA_  ( .A(A[227]), .B(n487), .CI(C[227]), .CO(C[228]) );
  FA_288 \FAINST[228].FA_  ( .A(A[228]), .B(n488), .CI(C[228]), .CO(C[229]) );
  FA_287 \FAINST[229].FA_  ( .A(A[229]), .B(n489), .CI(C[229]), .CO(C[230]) );
  FA_286 \FAINST[230].FA_  ( .A(A[230]), .B(n490), .CI(C[230]), .CO(C[231]) );
  FA_285 \FAINST[231].FA_  ( .A(A[231]), .B(n491), .CI(C[231]), .CO(C[232]) );
  FA_284 \FAINST[232].FA_  ( .A(A[232]), .B(n492), .CI(C[232]), .CO(C[233]) );
  FA_283 \FAINST[233].FA_  ( .A(A[233]), .B(n493), .CI(C[233]), .CO(C[234]) );
  FA_282 \FAINST[234].FA_  ( .A(A[234]), .B(n494), .CI(C[234]), .CO(C[235]) );
  FA_281 \FAINST[235].FA_  ( .A(A[235]), .B(n495), .CI(C[235]), .CO(C[236]) );
  FA_280 \FAINST[236].FA_  ( .A(A[236]), .B(n496), .CI(C[236]), .CO(C[237]) );
  FA_279 \FAINST[237].FA_  ( .A(A[237]), .B(n497), .CI(C[237]), .CO(C[238]) );
  FA_278 \FAINST[238].FA_  ( .A(A[238]), .B(n498), .CI(C[238]), .CO(C[239]) );
  FA_277 \FAINST[239].FA_  ( .A(A[239]), .B(n499), .CI(C[239]), .CO(C[240]) );
  FA_276 \FAINST[240].FA_  ( .A(A[240]), .B(n500), .CI(C[240]), .CO(C[241]) );
  FA_275 \FAINST[241].FA_  ( .A(A[241]), .B(n501), .CI(C[241]), .CO(C[242]) );
  FA_274 \FAINST[242].FA_  ( .A(A[242]), .B(n502), .CI(C[242]), .CO(C[243]) );
  FA_273 \FAINST[243].FA_  ( .A(A[243]), .B(n503), .CI(C[243]), .CO(C[244]) );
  FA_272 \FAINST[244].FA_  ( .A(A[244]), .B(n504), .CI(C[244]), .CO(C[245]) );
  FA_271 \FAINST[245].FA_  ( .A(A[245]), .B(n505), .CI(C[245]), .CO(C[246]) );
  FA_270 \FAINST[246].FA_  ( .A(A[246]), .B(n506), .CI(C[246]), .CO(C[247]) );
  FA_269 \FAINST[247].FA_  ( .A(A[247]), .B(n507), .CI(C[247]), .CO(C[248]) );
  FA_268 \FAINST[248].FA_  ( .A(A[248]), .B(n508), .CI(C[248]), .CO(C[249]) );
  FA_267 \FAINST[249].FA_  ( .A(A[249]), .B(n509), .CI(C[249]), .CO(C[250]) );
  FA_266 \FAINST[250].FA_  ( .A(A[250]), .B(n510), .CI(C[250]), .CO(C[251]) );
  FA_265 \FAINST[251].FA_  ( .A(A[251]), .B(n511), .CI(C[251]), .CO(C[252]) );
  FA_264 \FAINST[252].FA_  ( .A(A[252]), .B(n512), .CI(C[252]), .CO(C[253]) );
  FA_263 \FAINST[253].FA_  ( .A(A[253]), .B(n513), .CI(C[253]), .CO(C[254]) );
  FA_262 \FAINST[254].FA_  ( .A(A[254]), .B(n514), .CI(C[254]), .CO(C[255]) );
  FA_261 \FAINST[255].FA_  ( .A(A[255]), .B(n515), .CI(C[255]), .CO(C[256]) );
  FA_260 \FAINST[256].FA_  ( .A(1'b0), .B(n516), .CI(C[256]), .CO(C[257]) );
  FA_259 \FAINST[257].FA_  ( .A(1'b0), .B(n517), .CI(C[257]), .CO(O) );
  IV U2 ( .A(B[159]), .Z(n419) );
  IV U3 ( .A(B[160]), .Z(n420) );
  IV U4 ( .A(B[161]), .Z(n421) );
  IV U5 ( .A(B[162]), .Z(n422) );
  IV U6 ( .A(B[163]), .Z(n423) );
  IV U7 ( .A(B[164]), .Z(n424) );
  IV U8 ( .A(B[165]), .Z(n425) );
  IV U9 ( .A(B[166]), .Z(n426) );
  IV U10 ( .A(B[167]), .Z(n427) );
  IV U11 ( .A(B[168]), .Z(n428) );
  IV U12 ( .A(B[249]), .Z(n509) );
  IV U13 ( .A(B[169]), .Z(n429) );
  IV U14 ( .A(B[170]), .Z(n430) );
  IV U15 ( .A(B[171]), .Z(n431) );
  IV U16 ( .A(B[172]), .Z(n432) );
  IV U17 ( .A(B[173]), .Z(n433) );
  IV U18 ( .A(B[174]), .Z(n434) );
  IV U19 ( .A(B[175]), .Z(n435) );
  IV U20 ( .A(B[176]), .Z(n436) );
  IV U21 ( .A(B[177]), .Z(n437) );
  IV U22 ( .A(B[178]), .Z(n438) );
  IV U23 ( .A(B[250]), .Z(n510) );
  IV U24 ( .A(B[179]), .Z(n439) );
  IV U25 ( .A(B[180]), .Z(n440) );
  IV U26 ( .A(B[181]), .Z(n441) );
  IV U27 ( .A(B[182]), .Z(n442) );
  IV U28 ( .A(B[183]), .Z(n443) );
  IV U29 ( .A(B[184]), .Z(n444) );
  IV U30 ( .A(B[185]), .Z(n445) );
  IV U31 ( .A(B[186]), .Z(n446) );
  IV U32 ( .A(B[187]), .Z(n447) );
  IV U33 ( .A(B[188]), .Z(n448) );
  IV U34 ( .A(B[251]), .Z(n511) );
  IV U35 ( .A(B[189]), .Z(n449) );
  IV U36 ( .A(B[190]), .Z(n450) );
  IV U37 ( .A(B[191]), .Z(n451) );
  IV U38 ( .A(B[192]), .Z(n452) );
  IV U39 ( .A(B[193]), .Z(n453) );
  IV U40 ( .A(B[194]), .Z(n454) );
  IV U41 ( .A(B[195]), .Z(n455) );
  IV U42 ( .A(B[196]), .Z(n456) );
  IV U43 ( .A(B[197]), .Z(n457) );
  IV U44 ( .A(B[198]), .Z(n458) );
  IV U45 ( .A(B[252]), .Z(n512) );
  IV U46 ( .A(B[199]), .Z(n459) );
  IV U47 ( .A(B[200]), .Z(n460) );
  IV U48 ( .A(B[201]), .Z(n461) );
  IV U49 ( .A(B[202]), .Z(n462) );
  IV U50 ( .A(B[203]), .Z(n463) );
  IV U51 ( .A(B[204]), .Z(n464) );
  IV U52 ( .A(B[205]), .Z(n465) );
  IV U53 ( .A(B[206]), .Z(n466) );
  IV U54 ( .A(B[207]), .Z(n467) );
  IV U55 ( .A(B[208]), .Z(n468) );
  IV U56 ( .A(B[253]), .Z(n513) );
  IV U57 ( .A(B[209]), .Z(n469) );
  IV U58 ( .A(B[210]), .Z(n470) );
  IV U59 ( .A(B[211]), .Z(n471) );
  IV U60 ( .A(B[212]), .Z(n472) );
  IV U61 ( .A(B[213]), .Z(n473) );
  IV U62 ( .A(B[214]), .Z(n474) );
  IV U63 ( .A(B[215]), .Z(n475) );
  IV U64 ( .A(B[216]), .Z(n476) );
  IV U65 ( .A(B[217]), .Z(n477) );
  IV U66 ( .A(B[218]), .Z(n478) );
  IV U67 ( .A(B[254]), .Z(n514) );
  IV U68 ( .A(B[219]), .Z(n479) );
  IV U69 ( .A(B[220]), .Z(n480) );
  IV U70 ( .A(B[221]), .Z(n481) );
  IV U71 ( .A(B[222]), .Z(n482) );
  IV U72 ( .A(B[223]), .Z(n483) );
  IV U73 ( .A(B[224]), .Z(n484) );
  IV U74 ( .A(B[225]), .Z(n485) );
  IV U75 ( .A(B[226]), .Z(n486) );
  IV U76 ( .A(B[227]), .Z(n487) );
  IV U77 ( .A(B[228]), .Z(n488) );
  IV U78 ( .A(B[255]), .Z(n515) );
  IV U79 ( .A(B[229]), .Z(n489) );
  IV U80 ( .A(B[230]), .Z(n490) );
  IV U81 ( .A(B[231]), .Z(n491) );
  IV U82 ( .A(B[232]), .Z(n492) );
  IV U83 ( .A(B[0]), .Z(n260) );
  IV U84 ( .A(B[1]), .Z(n261) );
  IV U85 ( .A(B[2]), .Z(n262) );
  IV U86 ( .A(B[3]), .Z(n263) );
  IV U87 ( .A(B[4]), .Z(n264) );
  IV U88 ( .A(B[5]), .Z(n265) );
  IV U89 ( .A(B[6]), .Z(n266) );
  IV U90 ( .A(B[7]), .Z(n267) );
  IV U91 ( .A(B[8]), .Z(n268) );
  IV U92 ( .A(B[233]), .Z(n493) );
  IV U93 ( .A(B[9]), .Z(n269) );
  IV U94 ( .A(B[10]), .Z(n270) );
  IV U95 ( .A(B[11]), .Z(n271) );
  IV U96 ( .A(B[12]), .Z(n272) );
  IV U97 ( .A(B[13]), .Z(n273) );
  IV U98 ( .A(B[14]), .Z(n274) );
  IV U99 ( .A(B[15]), .Z(n275) );
  IV U100 ( .A(B[16]), .Z(n276) );
  IV U101 ( .A(B[17]), .Z(n277) );
  IV U102 ( .A(B[18]), .Z(n278) );
  IV U103 ( .A(B[234]), .Z(n494) );
  IV U104 ( .A(B[19]), .Z(n279) );
  IV U105 ( .A(B[20]), .Z(n280) );
  IV U106 ( .A(B[21]), .Z(n281) );
  IV U107 ( .A(B[22]), .Z(n282) );
  IV U108 ( .A(B[23]), .Z(n283) );
  IV U109 ( .A(B[24]), .Z(n284) );
  IV U110 ( .A(B[25]), .Z(n285) );
  IV U111 ( .A(B[26]), .Z(n286) );
  IV U112 ( .A(B[27]), .Z(n287) );
  IV U113 ( .A(B[28]), .Z(n288) );
  IV U114 ( .A(B[235]), .Z(n495) );
  IV U115 ( .A(B[29]), .Z(n289) );
  IV U116 ( .A(B[30]), .Z(n290) );
  IV U117 ( .A(B[31]), .Z(n291) );
  IV U118 ( .A(B[32]), .Z(n292) );
  IV U119 ( .A(B[33]), .Z(n293) );
  IV U120 ( .A(B[34]), .Z(n294) );
  IV U121 ( .A(B[35]), .Z(n295) );
  IV U122 ( .A(B[36]), .Z(n296) );
  IV U123 ( .A(B[37]), .Z(n297) );
  IV U124 ( .A(B[38]), .Z(n298) );
  IV U125 ( .A(B[236]), .Z(n496) );
  IV U126 ( .A(B[39]), .Z(n299) );
  IV U127 ( .A(B[40]), .Z(n300) );
  IV U128 ( .A(B[41]), .Z(n301) );
  IV U129 ( .A(B[42]), .Z(n302) );
  IV U130 ( .A(B[43]), .Z(n303) );
  IV U131 ( .A(B[44]), .Z(n304) );
  IV U132 ( .A(B[45]), .Z(n305) );
  IV U133 ( .A(B[46]), .Z(n306) );
  IV U134 ( .A(B[47]), .Z(n307) );
  IV U135 ( .A(B[48]), .Z(n308) );
  IV U136 ( .A(B[237]), .Z(n497) );
  IV U137 ( .A(B[49]), .Z(n309) );
  IV U138 ( .A(B[50]), .Z(n310) );
  IV U139 ( .A(B[51]), .Z(n311) );
  IV U140 ( .A(B[52]), .Z(n312) );
  IV U141 ( .A(B[53]), .Z(n313) );
  IV U142 ( .A(B[54]), .Z(n314) );
  IV U143 ( .A(B[55]), .Z(n315) );
  IV U144 ( .A(B[56]), .Z(n316) );
  IV U145 ( .A(B[57]), .Z(n317) );
  IV U146 ( .A(B[58]), .Z(n318) );
  IV U147 ( .A(B[238]), .Z(n498) );
  IV U148 ( .A(B[256]), .Z(n516) );
  IV U149 ( .A(B[59]), .Z(n319) );
  IV U150 ( .A(B[60]), .Z(n320) );
  IV U151 ( .A(B[61]), .Z(n321) );
  IV U152 ( .A(B[62]), .Z(n322) );
  IV U153 ( .A(B[63]), .Z(n323) );
  IV U154 ( .A(B[64]), .Z(n324) );
  IV U155 ( .A(B[65]), .Z(n325) );
  IV U156 ( .A(B[66]), .Z(n326) );
  IV U157 ( .A(B[67]), .Z(n327) );
  IV U158 ( .A(B[68]), .Z(n328) );
  IV U159 ( .A(B[239]), .Z(n499) );
  IV U160 ( .A(B[69]), .Z(n329) );
  IV U161 ( .A(B[70]), .Z(n330) );
  IV U162 ( .A(B[71]), .Z(n331) );
  IV U163 ( .A(B[72]), .Z(n332) );
  IV U164 ( .A(B[73]), .Z(n333) );
  IV U165 ( .A(B[74]), .Z(n334) );
  IV U166 ( .A(B[75]), .Z(n335) );
  IV U167 ( .A(B[76]), .Z(n336) );
  IV U168 ( .A(B[77]), .Z(n337) );
  IV U169 ( .A(B[78]), .Z(n338) );
  IV U170 ( .A(B[240]), .Z(n500) );
  IV U171 ( .A(B[79]), .Z(n339) );
  IV U172 ( .A(B[80]), .Z(n340) );
  IV U173 ( .A(B[81]), .Z(n341) );
  IV U174 ( .A(B[82]), .Z(n342) );
  IV U175 ( .A(B[83]), .Z(n343) );
  IV U176 ( .A(B[84]), .Z(n344) );
  IV U177 ( .A(B[85]), .Z(n345) );
  IV U178 ( .A(B[86]), .Z(n346) );
  IV U179 ( .A(B[87]), .Z(n347) );
  IV U180 ( .A(B[88]), .Z(n348) );
  IV U181 ( .A(B[241]), .Z(n501) );
  IV U182 ( .A(B[89]), .Z(n349) );
  IV U183 ( .A(B[90]), .Z(n350) );
  IV U184 ( .A(B[91]), .Z(n351) );
  IV U185 ( .A(B[92]), .Z(n352) );
  IV U186 ( .A(B[93]), .Z(n353) );
  IV U187 ( .A(B[94]), .Z(n354) );
  IV U188 ( .A(B[95]), .Z(n355) );
  IV U189 ( .A(B[96]), .Z(n356) );
  IV U190 ( .A(B[97]), .Z(n357) );
  IV U191 ( .A(B[98]), .Z(n358) );
  IV U192 ( .A(B[242]), .Z(n502) );
  IV U193 ( .A(B[99]), .Z(n359) );
  IV U194 ( .A(B[100]), .Z(n360) );
  IV U195 ( .A(B[101]), .Z(n361) );
  IV U196 ( .A(B[102]), .Z(n362) );
  IV U197 ( .A(B[103]), .Z(n363) );
  IV U198 ( .A(B[104]), .Z(n364) );
  IV U199 ( .A(B[105]), .Z(n365) );
  IV U200 ( .A(B[106]), .Z(n366) );
  IV U201 ( .A(B[107]), .Z(n367) );
  IV U202 ( .A(B[108]), .Z(n368) );
  IV U203 ( .A(B[243]), .Z(n503) );
  IV U204 ( .A(B[109]), .Z(n369) );
  IV U205 ( .A(B[110]), .Z(n370) );
  IV U206 ( .A(B[111]), .Z(n371) );
  IV U207 ( .A(B[112]), .Z(n372) );
  IV U208 ( .A(B[113]), .Z(n373) );
  IV U209 ( .A(B[114]), .Z(n374) );
  IV U210 ( .A(B[115]), .Z(n375) );
  IV U211 ( .A(B[116]), .Z(n376) );
  IV U212 ( .A(B[117]), .Z(n377) );
  IV U213 ( .A(B[118]), .Z(n378) );
  IV U214 ( .A(B[244]), .Z(n504) );
  IV U215 ( .A(B[119]), .Z(n379) );
  IV U216 ( .A(B[120]), .Z(n380) );
  IV U217 ( .A(B[121]), .Z(n381) );
  IV U218 ( .A(B[122]), .Z(n382) );
  IV U219 ( .A(B[123]), .Z(n383) );
  IV U220 ( .A(B[124]), .Z(n384) );
  IV U221 ( .A(B[125]), .Z(n385) );
  IV U222 ( .A(B[126]), .Z(n386) );
  IV U223 ( .A(B[127]), .Z(n387) );
  IV U224 ( .A(B[128]), .Z(n388) );
  IV U225 ( .A(B[245]), .Z(n505) );
  IV U226 ( .A(B[129]), .Z(n389) );
  IV U227 ( .A(B[130]), .Z(n390) );
  IV U228 ( .A(B[131]), .Z(n391) );
  IV U229 ( .A(B[132]), .Z(n392) );
  IV U230 ( .A(B[133]), .Z(n393) );
  IV U231 ( .A(B[134]), .Z(n394) );
  IV U232 ( .A(B[135]), .Z(n395) );
  IV U233 ( .A(B[136]), .Z(n396) );
  IV U234 ( .A(B[137]), .Z(n397) );
  IV U235 ( .A(B[138]), .Z(n398) );
  IV U236 ( .A(B[246]), .Z(n506) );
  IV U237 ( .A(B[139]), .Z(n399) );
  IV U238 ( .A(B[140]), .Z(n400) );
  IV U239 ( .A(B[141]), .Z(n401) );
  IV U240 ( .A(B[142]), .Z(n402) );
  IV U241 ( .A(B[143]), .Z(n403) );
  IV U242 ( .A(B[144]), .Z(n404) );
  IV U243 ( .A(B[145]), .Z(n405) );
  IV U244 ( .A(B[146]), .Z(n406) );
  IV U245 ( .A(B[147]), .Z(n407) );
  IV U246 ( .A(B[148]), .Z(n408) );
  IV U247 ( .A(B[247]), .Z(n507) );
  IV U248 ( .A(B[149]), .Z(n409) );
  IV U249 ( .A(B[150]), .Z(n410) );
  IV U250 ( .A(B[151]), .Z(n411) );
  IV U251 ( .A(B[152]), .Z(n412) );
  IV U252 ( .A(B[153]), .Z(n413) );
  IV U253 ( .A(B[154]), .Z(n414) );
  IV U254 ( .A(B[155]), .Z(n415) );
  IV U255 ( .A(B[156]), .Z(n416) );
  IV U256 ( .A(B[157]), .Z(n417) );
  IV U257 ( .A(B[158]), .Z(n418) );
  IV U258 ( .A(B[248]), .Z(n508) );
  IV U259 ( .A(B[257]), .Z(n517) );
endmodule


module FA_2 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_3 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_4 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_5 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_12 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_13 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_14 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_15 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_16 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_17 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_18 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_19 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_20 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_21 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_22 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_23 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_24 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_25 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_26 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_27 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_28 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_29 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_30 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_31 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_32 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_33 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_34 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_35 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_36 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_37 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_38 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_39 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_40 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_41 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_42 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_43 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_44 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_45 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_46 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_47 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_48 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_49 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_50 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_51 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_52 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_53 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_54 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_55 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_56 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_57 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_58 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_59 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_60 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_61 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_62 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_63 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_64 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_65 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_66 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_67 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_68 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_69 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_70 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_71 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_72 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_73 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_74 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_75 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_76 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_77 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_78 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_79 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_80 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_81 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_82 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_83 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_84 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_85 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_86 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_87 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_88 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_89 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_90 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_91 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_92 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_93 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_94 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_95 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_96 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_97 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_98 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_99 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N258_1 ( A, B, S, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] S;
  output CO;
  wire   n2, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512;
  wire   [257:1] C;

  FA_258 \FAINST[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(S[0]), .CO(C[1]) );
  FA_257 \FAINST[1].FA_  ( .A(A[1]), .B(n258), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_256 \FAINST[2].FA_  ( .A(A[2]), .B(n259), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_255 \FAINST[3].FA_  ( .A(A[3]), .B(n260), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_254 \FAINST[4].FA_  ( .A(A[4]), .B(n261), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_253 \FAINST[5].FA_  ( .A(A[5]), .B(n262), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_252 \FAINST[6].FA_  ( .A(A[6]), .B(n263), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_251 \FAINST[7].FA_  ( .A(A[7]), .B(n264), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_250 \FAINST[8].FA_  ( .A(A[8]), .B(n265), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_249 \FAINST[9].FA_  ( .A(A[9]), .B(n266), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_248 \FAINST[10].FA_  ( .A(A[10]), .B(n267), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_247 \FAINST[11].FA_  ( .A(A[11]), .B(n268), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_246 \FAINST[12].FA_  ( .A(A[12]), .B(n269), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_245 \FAINST[13].FA_  ( .A(A[13]), .B(n270), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_244 \FAINST[14].FA_  ( .A(A[14]), .B(n271), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_243 \FAINST[15].FA_  ( .A(A[15]), .B(n272), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_242 \FAINST[16].FA_  ( .A(A[16]), .B(n273), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_241 \FAINST[17].FA_  ( .A(A[17]), .B(n274), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_240 \FAINST[18].FA_  ( .A(A[18]), .B(n275), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_239 \FAINST[19].FA_  ( .A(A[19]), .B(n276), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_238 \FAINST[20].FA_  ( .A(A[20]), .B(n277), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_237 \FAINST[21].FA_  ( .A(A[21]), .B(n278), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_236 \FAINST[22].FA_  ( .A(A[22]), .B(n279), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_235 \FAINST[23].FA_  ( .A(A[23]), .B(n280), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_234 \FAINST[24].FA_  ( .A(A[24]), .B(n281), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_233 \FAINST[25].FA_  ( .A(A[25]), .B(n282), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_232 \FAINST[26].FA_  ( .A(A[26]), .B(n283), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_231 \FAINST[27].FA_  ( .A(A[27]), .B(n284), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_230 \FAINST[28].FA_  ( .A(A[28]), .B(n285), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_229 \FAINST[29].FA_  ( .A(A[29]), .B(n286), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_228 \FAINST[30].FA_  ( .A(A[30]), .B(n287), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_227 \FAINST[31].FA_  ( .A(A[31]), .B(n288), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_226 \FAINST[32].FA_  ( .A(A[32]), .B(n289), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_225 \FAINST[33].FA_  ( .A(A[33]), .B(n290), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_224 \FAINST[34].FA_  ( .A(A[34]), .B(n291), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_223 \FAINST[35].FA_  ( .A(A[35]), .B(n292), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_222 \FAINST[36].FA_  ( .A(A[36]), .B(n293), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_221 \FAINST[37].FA_  ( .A(A[37]), .B(n294), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_220 \FAINST[38].FA_  ( .A(A[38]), .B(n295), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_219 \FAINST[39].FA_  ( .A(A[39]), .B(n296), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_218 \FAINST[40].FA_  ( .A(A[40]), .B(n297), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_217 \FAINST[41].FA_  ( .A(A[41]), .B(n298), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_216 \FAINST[42].FA_  ( .A(A[42]), .B(n299), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_215 \FAINST[43].FA_  ( .A(A[43]), .B(n300), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_214 \FAINST[44].FA_  ( .A(A[44]), .B(n301), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_213 \FAINST[45].FA_  ( .A(A[45]), .B(n302), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_212 \FAINST[46].FA_  ( .A(A[46]), .B(n303), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_211 \FAINST[47].FA_  ( .A(A[47]), .B(n304), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_210 \FAINST[48].FA_  ( .A(A[48]), .B(n305), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_209 \FAINST[49].FA_  ( .A(A[49]), .B(n306), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_208 \FAINST[50].FA_  ( .A(A[50]), .B(n307), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_207 \FAINST[51].FA_  ( .A(A[51]), .B(n308), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_206 \FAINST[52].FA_  ( .A(A[52]), .B(n309), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_205 \FAINST[53].FA_  ( .A(A[53]), .B(n310), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_204 \FAINST[54].FA_  ( .A(A[54]), .B(n311), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_203 \FAINST[55].FA_  ( .A(A[55]), .B(n312), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_202 \FAINST[56].FA_  ( .A(A[56]), .B(n313), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_201 \FAINST[57].FA_  ( .A(A[57]), .B(n314), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_200 \FAINST[58].FA_  ( .A(A[58]), .B(n315), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_199 \FAINST[59].FA_  ( .A(A[59]), .B(n316), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_198 \FAINST[60].FA_  ( .A(A[60]), .B(n317), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_197 \FAINST[61].FA_  ( .A(A[61]), .B(n318), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_196 \FAINST[62].FA_  ( .A(A[62]), .B(n319), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_195 \FAINST[63].FA_  ( .A(A[63]), .B(n320), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_194 \FAINST[64].FA_  ( .A(A[64]), .B(n321), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_193 \FAINST[65].FA_  ( .A(A[65]), .B(n322), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_192 \FAINST[66].FA_  ( .A(A[66]), .B(n323), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_191 \FAINST[67].FA_  ( .A(A[67]), .B(n324), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_190 \FAINST[68].FA_  ( .A(A[68]), .B(n325), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_189 \FAINST[69].FA_  ( .A(A[69]), .B(n326), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_188 \FAINST[70].FA_  ( .A(A[70]), .B(n327), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_187 \FAINST[71].FA_  ( .A(A[71]), .B(n328), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_186 \FAINST[72].FA_  ( .A(A[72]), .B(n329), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_185 \FAINST[73].FA_  ( .A(A[73]), .B(n330), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_184 \FAINST[74].FA_  ( .A(A[74]), .B(n331), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_183 \FAINST[75].FA_  ( .A(A[75]), .B(n332), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_182 \FAINST[76].FA_  ( .A(A[76]), .B(n333), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_181 \FAINST[77].FA_  ( .A(A[77]), .B(n334), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_180 \FAINST[78].FA_  ( .A(A[78]), .B(n335), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_179 \FAINST[79].FA_  ( .A(A[79]), .B(n336), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_178 \FAINST[80].FA_  ( .A(A[80]), .B(n337), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_177 \FAINST[81].FA_  ( .A(A[81]), .B(n338), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_176 \FAINST[82].FA_  ( .A(A[82]), .B(n339), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_175 \FAINST[83].FA_  ( .A(A[83]), .B(n340), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_174 \FAINST[84].FA_  ( .A(A[84]), .B(n341), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_173 \FAINST[85].FA_  ( .A(A[85]), .B(n342), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_172 \FAINST[86].FA_  ( .A(A[86]), .B(n343), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_171 \FAINST[87].FA_  ( .A(A[87]), .B(n344), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_170 \FAINST[88].FA_  ( .A(A[88]), .B(n345), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_169 \FAINST[89].FA_  ( .A(A[89]), .B(n346), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_168 \FAINST[90].FA_  ( .A(A[90]), .B(n347), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_167 \FAINST[91].FA_  ( .A(A[91]), .B(n348), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_166 \FAINST[92].FA_  ( .A(A[92]), .B(n349), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_165 \FAINST[93].FA_  ( .A(A[93]), .B(n350), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_164 \FAINST[94].FA_  ( .A(A[94]), .B(n351), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_163 \FAINST[95].FA_  ( .A(A[95]), .B(n352), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_162 \FAINST[96].FA_  ( .A(A[96]), .B(n353), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_161 \FAINST[97].FA_  ( .A(A[97]), .B(n354), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_160 \FAINST[98].FA_  ( .A(A[98]), .B(n355), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_159 \FAINST[99].FA_  ( .A(A[99]), .B(n356), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_158 \FAINST[100].FA_  ( .A(A[100]), .B(n357), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_157 \FAINST[101].FA_  ( .A(A[101]), .B(n358), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_156 \FAINST[102].FA_  ( .A(A[102]), .B(n359), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_155 \FAINST[103].FA_  ( .A(A[103]), .B(n360), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_154 \FAINST[104].FA_  ( .A(A[104]), .B(n361), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_153 \FAINST[105].FA_  ( .A(A[105]), .B(n362), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_152 \FAINST[106].FA_  ( .A(A[106]), .B(n363), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_151 \FAINST[107].FA_  ( .A(A[107]), .B(n364), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_150 \FAINST[108].FA_  ( .A(A[108]), .B(n365), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_149 \FAINST[109].FA_  ( .A(A[109]), .B(n366), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_148 \FAINST[110].FA_  ( .A(A[110]), .B(n367), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_147 \FAINST[111].FA_  ( .A(A[111]), .B(n368), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_146 \FAINST[112].FA_  ( .A(A[112]), .B(n369), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_145 \FAINST[113].FA_  ( .A(A[113]), .B(n370), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_144 \FAINST[114].FA_  ( .A(A[114]), .B(n371), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_143 \FAINST[115].FA_  ( .A(A[115]), .B(n372), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_142 \FAINST[116].FA_  ( .A(A[116]), .B(n373), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_141 \FAINST[117].FA_  ( .A(A[117]), .B(n374), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_140 \FAINST[118].FA_  ( .A(A[118]), .B(n375), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_139 \FAINST[119].FA_  ( .A(A[119]), .B(n376), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_138 \FAINST[120].FA_  ( .A(A[120]), .B(n377), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_137 \FAINST[121].FA_  ( .A(A[121]), .B(n378), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_136 \FAINST[122].FA_  ( .A(A[122]), .B(n379), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_135 \FAINST[123].FA_  ( .A(A[123]), .B(n380), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_134 \FAINST[124].FA_  ( .A(A[124]), .B(n381), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_133 \FAINST[125].FA_  ( .A(A[125]), .B(n382), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_132 \FAINST[126].FA_  ( .A(A[126]), .B(n383), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_131 \FAINST[127].FA_  ( .A(A[127]), .B(n384), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_130 \FAINST[128].FA_  ( .A(A[128]), .B(n385), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_129 \FAINST[129].FA_  ( .A(A[129]), .B(n386), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_128 \FAINST[130].FA_  ( .A(A[130]), .B(n387), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_127 \FAINST[131].FA_  ( .A(A[131]), .B(n388), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_126 \FAINST[132].FA_  ( .A(A[132]), .B(n389), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_125 \FAINST[133].FA_  ( .A(A[133]), .B(n390), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_124 \FAINST[134].FA_  ( .A(A[134]), .B(n391), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_123 \FAINST[135].FA_  ( .A(A[135]), .B(n392), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_122 \FAINST[136].FA_  ( .A(A[136]), .B(n393), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_121 \FAINST[137].FA_  ( .A(A[137]), .B(n394), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_120 \FAINST[138].FA_  ( .A(A[138]), .B(n395), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_119 \FAINST[139].FA_  ( .A(A[139]), .B(n396), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_118 \FAINST[140].FA_  ( .A(A[140]), .B(n397), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_117 \FAINST[141].FA_  ( .A(A[141]), .B(n398), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_116 \FAINST[142].FA_  ( .A(A[142]), .B(n399), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_115 \FAINST[143].FA_  ( .A(A[143]), .B(n400), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_114 \FAINST[144].FA_  ( .A(A[144]), .B(n401), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_113 \FAINST[145].FA_  ( .A(A[145]), .B(n402), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_112 \FAINST[146].FA_  ( .A(A[146]), .B(n403), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_111 \FAINST[147].FA_  ( .A(A[147]), .B(n404), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_110 \FAINST[148].FA_  ( .A(A[148]), .B(n405), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_109 \FAINST[149].FA_  ( .A(A[149]), .B(n406), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_108 \FAINST[150].FA_  ( .A(A[150]), .B(n407), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_107 \FAINST[151].FA_  ( .A(A[151]), .B(n408), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_106 \FAINST[152].FA_  ( .A(A[152]), .B(n409), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_105 \FAINST[153].FA_  ( .A(A[153]), .B(n410), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_104 \FAINST[154].FA_  ( .A(A[154]), .B(n411), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_103 \FAINST[155].FA_  ( .A(A[155]), .B(n412), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_102 \FAINST[156].FA_  ( .A(A[156]), .B(n413), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_101 \FAINST[157].FA_  ( .A(A[157]), .B(n414), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_100 \FAINST[158].FA_  ( .A(A[158]), .B(n415), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_99 \FAINST[159].FA_  ( .A(A[159]), .B(n416), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_98 \FAINST[160].FA_  ( .A(A[160]), .B(n417), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_97 \FAINST[161].FA_  ( .A(A[161]), .B(n418), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_96 \FAINST[162].FA_  ( .A(A[162]), .B(n419), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_95 \FAINST[163].FA_  ( .A(A[163]), .B(n420), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_94 \FAINST[164].FA_  ( .A(A[164]), .B(n421), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_93 \FAINST[165].FA_  ( .A(A[165]), .B(n422), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_92 \FAINST[166].FA_  ( .A(A[166]), .B(n423), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_91 \FAINST[167].FA_  ( .A(A[167]), .B(n424), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_90 \FAINST[168].FA_  ( .A(A[168]), .B(n425), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_89 \FAINST[169].FA_  ( .A(A[169]), .B(n426), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_88 \FAINST[170].FA_  ( .A(A[170]), .B(n427), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_87 \FAINST[171].FA_  ( .A(A[171]), .B(n428), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_86 \FAINST[172].FA_  ( .A(A[172]), .B(n429), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_85 \FAINST[173].FA_  ( .A(A[173]), .B(n430), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_84 \FAINST[174].FA_  ( .A(A[174]), .B(n431), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_83 \FAINST[175].FA_  ( .A(A[175]), .B(n432), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_82 \FAINST[176].FA_  ( .A(A[176]), .B(n433), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_81 \FAINST[177].FA_  ( .A(A[177]), .B(n434), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_80 \FAINST[178].FA_  ( .A(A[178]), .B(n435), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_79 \FAINST[179].FA_  ( .A(A[179]), .B(n436), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_78 \FAINST[180].FA_  ( .A(A[180]), .B(n437), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_77 \FAINST[181].FA_  ( .A(A[181]), .B(n438), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_76 \FAINST[182].FA_  ( .A(A[182]), .B(n439), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_75 \FAINST[183].FA_  ( .A(A[183]), .B(n440), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_74 \FAINST[184].FA_  ( .A(A[184]), .B(n441), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_73 \FAINST[185].FA_  ( .A(A[185]), .B(n442), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_72 \FAINST[186].FA_  ( .A(A[186]), .B(n443), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_71 \FAINST[187].FA_  ( .A(A[187]), .B(n444), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_70 \FAINST[188].FA_  ( .A(A[188]), .B(n445), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_69 \FAINST[189].FA_  ( .A(A[189]), .B(n446), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_68 \FAINST[190].FA_  ( .A(A[190]), .B(n447), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_67 \FAINST[191].FA_  ( .A(A[191]), .B(n448), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_66 \FAINST[192].FA_  ( .A(A[192]), .B(n449), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_65 \FAINST[193].FA_  ( .A(A[193]), .B(n450), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_64 \FAINST[194].FA_  ( .A(A[194]), .B(n451), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_63 \FAINST[195].FA_  ( .A(A[195]), .B(n452), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_62 \FAINST[196].FA_  ( .A(A[196]), .B(n453), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_61 \FAINST[197].FA_  ( .A(A[197]), .B(n454), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_60 \FAINST[198].FA_  ( .A(A[198]), .B(n455), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_59 \FAINST[199].FA_  ( .A(A[199]), .B(n456), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_58 \FAINST[200].FA_  ( .A(A[200]), .B(n457), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_57 \FAINST[201].FA_  ( .A(A[201]), .B(n458), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_56 \FAINST[202].FA_  ( .A(A[202]), .B(n459), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_55 \FAINST[203].FA_  ( .A(A[203]), .B(n460), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_54 \FAINST[204].FA_  ( .A(A[204]), .B(n461), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_53 \FAINST[205].FA_  ( .A(A[205]), .B(n462), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_52 \FAINST[206].FA_  ( .A(A[206]), .B(n463), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_51 \FAINST[207].FA_  ( .A(A[207]), .B(n464), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_50 \FAINST[208].FA_  ( .A(A[208]), .B(n465), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_49 \FAINST[209].FA_  ( .A(A[209]), .B(n466), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_48 \FAINST[210].FA_  ( .A(A[210]), .B(n467), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_47 \FAINST[211].FA_  ( .A(A[211]), .B(n468), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_46 \FAINST[212].FA_  ( .A(A[212]), .B(n469), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_45 \FAINST[213].FA_  ( .A(A[213]), .B(n470), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_44 \FAINST[214].FA_  ( .A(A[214]), .B(n471), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_43 \FAINST[215].FA_  ( .A(A[215]), .B(n472), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_42 \FAINST[216].FA_  ( .A(A[216]), .B(n473), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_41 \FAINST[217].FA_  ( .A(A[217]), .B(n474), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_40 \FAINST[218].FA_  ( .A(A[218]), .B(n475), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_39 \FAINST[219].FA_  ( .A(A[219]), .B(n476), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_38 \FAINST[220].FA_  ( .A(A[220]), .B(n477), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_37 \FAINST[221].FA_  ( .A(A[221]), .B(n478), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_36 \FAINST[222].FA_  ( .A(A[222]), .B(n479), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_35 \FAINST[223].FA_  ( .A(A[223]), .B(n480), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_34 \FAINST[224].FA_  ( .A(A[224]), .B(n481), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_33 \FAINST[225].FA_  ( .A(A[225]), .B(n482), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_32 \FAINST[226].FA_  ( .A(A[226]), .B(n483), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_31 \FAINST[227].FA_  ( .A(A[227]), .B(n484), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_30 \FAINST[228].FA_  ( .A(A[228]), .B(n485), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_29 \FAINST[229].FA_  ( .A(A[229]), .B(n486), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_28 \FAINST[230].FA_  ( .A(A[230]), .B(n487), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_27 \FAINST[231].FA_  ( .A(A[231]), .B(n488), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_26 \FAINST[232].FA_  ( .A(A[232]), .B(n489), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_25 \FAINST[233].FA_  ( .A(A[233]), .B(n490), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_24 \FAINST[234].FA_  ( .A(A[234]), .B(n491), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_23 \FAINST[235].FA_  ( .A(A[235]), .B(n492), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_22 \FAINST[236].FA_  ( .A(A[236]), .B(n493), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_21 \FAINST[237].FA_  ( .A(A[237]), .B(n494), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_20 \FAINST[238].FA_  ( .A(A[238]), .B(n495), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_19 \FAINST[239].FA_  ( .A(A[239]), .B(n496), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_18 \FAINST[240].FA_  ( .A(A[240]), .B(n497), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_17 \FAINST[241].FA_  ( .A(A[241]), .B(n498), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_16 \FAINST[242].FA_  ( .A(A[242]), .B(n499), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_15 \FAINST[243].FA_  ( .A(A[243]), .B(n500), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_14 \FAINST[244].FA_  ( .A(A[244]), .B(n501), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_13 \FAINST[245].FA_  ( .A(A[245]), .B(n502), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_12 \FAINST[246].FA_  ( .A(A[246]), .B(n503), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_11 \FAINST[247].FA_  ( .A(A[247]), .B(n504), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_10 \FAINST[248].FA_  ( .A(A[248]), .B(n505), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_9 \FAINST[249].FA_  ( .A(A[249]), .B(n506), .CI(C[249]), .S(S[249]), .CO(
        C[250]) );
  FA_8 \FAINST[250].FA_  ( .A(A[250]), .B(n507), .CI(C[250]), .S(S[250]), .CO(
        C[251]) );
  FA_7 \FAINST[251].FA_  ( .A(A[251]), .B(n508), .CI(C[251]), .S(S[251]), .CO(
        C[252]) );
  FA_6 \FAINST[252].FA_  ( .A(A[252]), .B(n509), .CI(C[252]), .S(S[252]), .CO(
        C[253]) );
  FA_5 \FAINST[253].FA_  ( .A(A[253]), .B(n510), .CI(C[253]), .S(S[253]), .CO(
        C[254]) );
  FA_4 \FAINST[254].FA_  ( .A(A[254]), .B(n511), .CI(C[254]), .S(S[254]), .CO(
        C[255]) );
  FA_3 \FAINST[255].FA_  ( .A(A[255]), .B(n512), .CI(C[255]), .S(S[255]), .CO(
        C[256]) );
  FA_2 \FAINST[256].FA_  ( .A(A[256]), .B(1'b1), .CI(C[256]), .S(S[256]) );
  IV U2 ( .A(B[159]), .Z(n416) );
  IV U3 ( .A(B[160]), .Z(n417) );
  IV U4 ( .A(B[161]), .Z(n418) );
  IV U5 ( .A(B[162]), .Z(n419) );
  IV U6 ( .A(B[163]), .Z(n420) );
  IV U7 ( .A(B[164]), .Z(n421) );
  IV U8 ( .A(B[165]), .Z(n422) );
  IV U9 ( .A(B[166]), .Z(n423) );
  IV U10 ( .A(B[167]), .Z(n424) );
  IV U11 ( .A(B[168]), .Z(n425) );
  IV U12 ( .A(B[249]), .Z(n506) );
  IV U13 ( .A(B[169]), .Z(n426) );
  IV U14 ( .A(B[170]), .Z(n427) );
  IV U15 ( .A(B[171]), .Z(n428) );
  IV U16 ( .A(B[172]), .Z(n429) );
  IV U17 ( .A(B[173]), .Z(n430) );
  IV U18 ( .A(B[174]), .Z(n431) );
  IV U19 ( .A(B[175]), .Z(n432) );
  IV U20 ( .A(B[176]), .Z(n433) );
  IV U21 ( .A(B[177]), .Z(n434) );
  IV U22 ( .A(B[178]), .Z(n435) );
  IV U23 ( .A(B[250]), .Z(n507) );
  IV U24 ( .A(B[179]), .Z(n436) );
  IV U25 ( .A(B[180]), .Z(n437) );
  IV U26 ( .A(B[181]), .Z(n438) );
  IV U27 ( .A(B[182]), .Z(n439) );
  IV U28 ( .A(B[183]), .Z(n440) );
  IV U29 ( .A(B[184]), .Z(n441) );
  IV U30 ( .A(B[185]), .Z(n442) );
  IV U31 ( .A(B[186]), .Z(n443) );
  IV U32 ( .A(B[187]), .Z(n444) );
  IV U33 ( .A(B[188]), .Z(n445) );
  IV U34 ( .A(B[251]), .Z(n508) );
  IV U35 ( .A(B[189]), .Z(n446) );
  IV U36 ( .A(B[190]), .Z(n447) );
  IV U37 ( .A(B[191]), .Z(n448) );
  IV U38 ( .A(B[192]), .Z(n449) );
  IV U39 ( .A(B[193]), .Z(n450) );
  IV U40 ( .A(B[194]), .Z(n451) );
  IV U41 ( .A(B[195]), .Z(n452) );
  IV U42 ( .A(B[196]), .Z(n453) );
  IV U43 ( .A(B[197]), .Z(n454) );
  IV U44 ( .A(B[198]), .Z(n455) );
  IV U45 ( .A(B[252]), .Z(n509) );
  IV U46 ( .A(B[199]), .Z(n456) );
  IV U47 ( .A(B[200]), .Z(n457) );
  IV U48 ( .A(B[201]), .Z(n458) );
  IV U49 ( .A(B[202]), .Z(n459) );
  IV U50 ( .A(B[203]), .Z(n460) );
  IV U51 ( .A(B[204]), .Z(n461) );
  IV U52 ( .A(B[205]), .Z(n462) );
  IV U53 ( .A(B[206]), .Z(n463) );
  IV U54 ( .A(B[207]), .Z(n464) );
  IV U55 ( .A(B[208]), .Z(n465) );
  IV U56 ( .A(B[253]), .Z(n510) );
  IV U57 ( .A(B[209]), .Z(n466) );
  IV U58 ( .A(B[210]), .Z(n467) );
  IV U59 ( .A(B[211]), .Z(n468) );
  IV U60 ( .A(B[212]), .Z(n469) );
  IV U61 ( .A(B[213]), .Z(n470) );
  IV U62 ( .A(B[214]), .Z(n471) );
  IV U63 ( .A(B[215]), .Z(n472) );
  IV U64 ( .A(B[216]), .Z(n473) );
  IV U65 ( .A(B[217]), .Z(n474) );
  IV U66 ( .A(B[218]), .Z(n475) );
  IV U67 ( .A(B[254]), .Z(n511) );
  IV U68 ( .A(B[219]), .Z(n476) );
  IV U69 ( .A(B[220]), .Z(n477) );
  IV U70 ( .A(B[221]), .Z(n478) );
  IV U71 ( .A(B[222]), .Z(n479) );
  IV U72 ( .A(B[223]), .Z(n480) );
  IV U73 ( .A(B[224]), .Z(n481) );
  IV U74 ( .A(B[225]), .Z(n482) );
  IV U75 ( .A(B[226]), .Z(n483) );
  IV U76 ( .A(B[227]), .Z(n484) );
  IV U77 ( .A(B[228]), .Z(n485) );
  IV U78 ( .A(B[255]), .Z(n512) );
  IV U79 ( .A(B[229]), .Z(n486) );
  IV U80 ( .A(B[230]), .Z(n487) );
  IV U81 ( .A(B[231]), .Z(n488) );
  IV U82 ( .A(B[232]), .Z(n489) );
  IV U83 ( .A(B[0]), .Z(n2) );
  IV U84 ( .A(B[1]), .Z(n258) );
  IV U85 ( .A(B[2]), .Z(n259) );
  IV U86 ( .A(B[3]), .Z(n260) );
  IV U87 ( .A(B[4]), .Z(n261) );
  IV U88 ( .A(B[5]), .Z(n262) );
  IV U89 ( .A(B[6]), .Z(n263) );
  IV U90 ( .A(B[7]), .Z(n264) );
  IV U91 ( .A(B[8]), .Z(n265) );
  IV U92 ( .A(B[233]), .Z(n490) );
  IV U93 ( .A(B[9]), .Z(n266) );
  IV U94 ( .A(B[10]), .Z(n267) );
  IV U95 ( .A(B[11]), .Z(n268) );
  IV U96 ( .A(B[12]), .Z(n269) );
  IV U97 ( .A(B[13]), .Z(n270) );
  IV U98 ( .A(B[14]), .Z(n271) );
  IV U99 ( .A(B[15]), .Z(n272) );
  IV U100 ( .A(B[16]), .Z(n273) );
  IV U101 ( .A(B[17]), .Z(n274) );
  IV U102 ( .A(B[18]), .Z(n275) );
  IV U103 ( .A(B[234]), .Z(n491) );
  IV U104 ( .A(B[19]), .Z(n276) );
  IV U105 ( .A(B[20]), .Z(n277) );
  IV U106 ( .A(B[21]), .Z(n278) );
  IV U107 ( .A(B[22]), .Z(n279) );
  IV U108 ( .A(B[23]), .Z(n280) );
  IV U109 ( .A(B[24]), .Z(n281) );
  IV U110 ( .A(B[25]), .Z(n282) );
  IV U111 ( .A(B[26]), .Z(n283) );
  IV U112 ( .A(B[27]), .Z(n284) );
  IV U113 ( .A(B[28]), .Z(n285) );
  IV U114 ( .A(B[235]), .Z(n492) );
  IV U115 ( .A(B[29]), .Z(n286) );
  IV U116 ( .A(B[30]), .Z(n287) );
  IV U117 ( .A(B[31]), .Z(n288) );
  IV U118 ( .A(B[32]), .Z(n289) );
  IV U119 ( .A(B[33]), .Z(n290) );
  IV U120 ( .A(B[34]), .Z(n291) );
  IV U121 ( .A(B[35]), .Z(n292) );
  IV U122 ( .A(B[36]), .Z(n293) );
  IV U123 ( .A(B[37]), .Z(n294) );
  IV U124 ( .A(B[38]), .Z(n295) );
  IV U125 ( .A(B[236]), .Z(n493) );
  IV U126 ( .A(B[39]), .Z(n296) );
  IV U127 ( .A(B[40]), .Z(n297) );
  IV U128 ( .A(B[41]), .Z(n298) );
  IV U129 ( .A(B[42]), .Z(n299) );
  IV U130 ( .A(B[43]), .Z(n300) );
  IV U131 ( .A(B[44]), .Z(n301) );
  IV U132 ( .A(B[45]), .Z(n302) );
  IV U133 ( .A(B[46]), .Z(n303) );
  IV U134 ( .A(B[47]), .Z(n304) );
  IV U135 ( .A(B[48]), .Z(n305) );
  IV U136 ( .A(B[237]), .Z(n494) );
  IV U137 ( .A(B[49]), .Z(n306) );
  IV U138 ( .A(B[50]), .Z(n307) );
  IV U139 ( .A(B[51]), .Z(n308) );
  IV U140 ( .A(B[52]), .Z(n309) );
  IV U141 ( .A(B[53]), .Z(n310) );
  IV U142 ( .A(B[54]), .Z(n311) );
  IV U143 ( .A(B[55]), .Z(n312) );
  IV U144 ( .A(B[56]), .Z(n313) );
  IV U145 ( .A(B[57]), .Z(n314) );
  IV U146 ( .A(B[58]), .Z(n315) );
  IV U147 ( .A(B[238]), .Z(n495) );
  IV U148 ( .A(B[59]), .Z(n316) );
  IV U149 ( .A(B[60]), .Z(n317) );
  IV U150 ( .A(B[61]), .Z(n318) );
  IV U151 ( .A(B[62]), .Z(n319) );
  IV U152 ( .A(B[63]), .Z(n320) );
  IV U153 ( .A(B[64]), .Z(n321) );
  IV U154 ( .A(B[65]), .Z(n322) );
  IV U155 ( .A(B[66]), .Z(n323) );
  IV U156 ( .A(B[67]), .Z(n324) );
  IV U157 ( .A(B[68]), .Z(n325) );
  IV U158 ( .A(B[239]), .Z(n496) );
  IV U159 ( .A(B[69]), .Z(n326) );
  IV U160 ( .A(B[70]), .Z(n327) );
  IV U161 ( .A(B[71]), .Z(n328) );
  IV U162 ( .A(B[72]), .Z(n329) );
  IV U163 ( .A(B[73]), .Z(n330) );
  IV U164 ( .A(B[74]), .Z(n331) );
  IV U165 ( .A(B[75]), .Z(n332) );
  IV U166 ( .A(B[76]), .Z(n333) );
  IV U167 ( .A(B[77]), .Z(n334) );
  IV U168 ( .A(B[78]), .Z(n335) );
  IV U169 ( .A(B[240]), .Z(n497) );
  IV U170 ( .A(B[79]), .Z(n336) );
  IV U171 ( .A(B[80]), .Z(n337) );
  IV U172 ( .A(B[81]), .Z(n338) );
  IV U173 ( .A(B[82]), .Z(n339) );
  IV U174 ( .A(B[83]), .Z(n340) );
  IV U175 ( .A(B[84]), .Z(n341) );
  IV U176 ( .A(B[85]), .Z(n342) );
  IV U177 ( .A(B[86]), .Z(n343) );
  IV U178 ( .A(B[87]), .Z(n344) );
  IV U179 ( .A(B[88]), .Z(n345) );
  IV U180 ( .A(B[241]), .Z(n498) );
  IV U181 ( .A(B[89]), .Z(n346) );
  IV U182 ( .A(B[90]), .Z(n347) );
  IV U183 ( .A(B[91]), .Z(n348) );
  IV U184 ( .A(B[92]), .Z(n349) );
  IV U185 ( .A(B[93]), .Z(n350) );
  IV U186 ( .A(B[94]), .Z(n351) );
  IV U187 ( .A(B[95]), .Z(n352) );
  IV U188 ( .A(B[96]), .Z(n353) );
  IV U189 ( .A(B[97]), .Z(n354) );
  IV U190 ( .A(B[98]), .Z(n355) );
  IV U191 ( .A(B[242]), .Z(n499) );
  IV U192 ( .A(B[99]), .Z(n356) );
  IV U193 ( .A(B[100]), .Z(n357) );
  IV U194 ( .A(B[101]), .Z(n358) );
  IV U195 ( .A(B[102]), .Z(n359) );
  IV U196 ( .A(B[103]), .Z(n360) );
  IV U197 ( .A(B[104]), .Z(n361) );
  IV U198 ( .A(B[105]), .Z(n362) );
  IV U199 ( .A(B[106]), .Z(n363) );
  IV U200 ( .A(B[107]), .Z(n364) );
  IV U201 ( .A(B[108]), .Z(n365) );
  IV U202 ( .A(B[243]), .Z(n500) );
  IV U203 ( .A(B[109]), .Z(n366) );
  IV U204 ( .A(B[110]), .Z(n367) );
  IV U205 ( .A(B[111]), .Z(n368) );
  IV U206 ( .A(B[112]), .Z(n369) );
  IV U207 ( .A(B[113]), .Z(n370) );
  IV U208 ( .A(B[114]), .Z(n371) );
  IV U209 ( .A(B[115]), .Z(n372) );
  IV U210 ( .A(B[116]), .Z(n373) );
  IV U211 ( .A(B[117]), .Z(n374) );
  IV U212 ( .A(B[118]), .Z(n375) );
  IV U213 ( .A(B[244]), .Z(n501) );
  IV U214 ( .A(B[119]), .Z(n376) );
  IV U215 ( .A(B[120]), .Z(n377) );
  IV U216 ( .A(B[121]), .Z(n378) );
  IV U217 ( .A(B[122]), .Z(n379) );
  IV U218 ( .A(B[123]), .Z(n380) );
  IV U219 ( .A(B[124]), .Z(n381) );
  IV U220 ( .A(B[125]), .Z(n382) );
  IV U221 ( .A(B[126]), .Z(n383) );
  IV U222 ( .A(B[127]), .Z(n384) );
  IV U223 ( .A(B[128]), .Z(n385) );
  IV U224 ( .A(B[245]), .Z(n502) );
  IV U225 ( .A(B[129]), .Z(n386) );
  IV U226 ( .A(B[130]), .Z(n387) );
  IV U227 ( .A(B[131]), .Z(n388) );
  IV U228 ( .A(B[132]), .Z(n389) );
  IV U229 ( .A(B[133]), .Z(n390) );
  IV U230 ( .A(B[134]), .Z(n391) );
  IV U231 ( .A(B[135]), .Z(n392) );
  IV U232 ( .A(B[136]), .Z(n393) );
  IV U233 ( .A(B[137]), .Z(n394) );
  IV U234 ( .A(B[138]), .Z(n395) );
  IV U235 ( .A(B[246]), .Z(n503) );
  IV U236 ( .A(B[139]), .Z(n396) );
  IV U237 ( .A(B[140]), .Z(n397) );
  IV U238 ( .A(B[141]), .Z(n398) );
  IV U239 ( .A(B[142]), .Z(n399) );
  IV U240 ( .A(B[143]), .Z(n400) );
  IV U241 ( .A(B[144]), .Z(n401) );
  IV U242 ( .A(B[145]), .Z(n402) );
  IV U243 ( .A(B[146]), .Z(n403) );
  IV U244 ( .A(B[147]), .Z(n404) );
  IV U245 ( .A(B[148]), .Z(n405) );
  IV U246 ( .A(B[247]), .Z(n504) );
  IV U247 ( .A(B[149]), .Z(n406) );
  IV U248 ( .A(B[150]), .Z(n407) );
  IV U249 ( .A(B[151]), .Z(n408) );
  IV U250 ( .A(B[152]), .Z(n409) );
  IV U251 ( .A(B[153]), .Z(n410) );
  IV U252 ( .A(B[154]), .Z(n411) );
  IV U253 ( .A(B[155]), .Z(n412) );
  IV U254 ( .A(B[156]), .Z(n413) );
  IV U255 ( .A(B[157]), .Z(n414) );
  IV U256 ( .A(B[158]), .Z(n415) );
  IV U257 ( .A(B[248]), .Z(n505) );
endmodule


module modmult_step_N256 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   c1, c2, n1;
  wire   [257:0] w1;
  wire   [257:0] w2;
  wire   [257:0] w3;
  wire   [257:0] z2;
  wire   [257:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  MUX_N258_0 MUX_1 ( .A({1'b0, 1'b0, y}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(xregN_1), .O({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, w1[255:0]}) );
  MUX_N258_2 MUX_2 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(c1), .O({SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        w2[255:0]}) );
  MUX_N258_1 MUX_3 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .S(n1), .O({SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        w3[255:0]}) );
  ADD_N258 ADD_1 ( .A({zin[256:0], 1'b0}), .B({1'b0, 1'b0, w1[255:0]}), .CI(
        1'b0), .S(z2) );
  COMP_N258_0 COMP_1 ( .A(z2), .B({1'b0, 1'b0, n}), .O(c1) );
  SUB_N258_0 SUB_1 ( .A(z2), .B({1'b0, 1'b0, w2[255:0]}), .S(z3) );
  COMP_N258_1 COMP_2 ( .A({1'b0, 1'b0, n}), .B(z3), .O(c2) );
  SUB_N258_1 SUB_2 ( .A({1'b0, z3[256:0]}), .B({1'b0, 1'b0, w3[255:0]}), .S({
        SYNOPSYS_UNCONNECTED__6, zout[256:0]}) );
  IV U2 ( .A(c2), .Z(n1) );
endmodule


module modmult_N256_CC256 ( clk, rst, start, x, y, n, o );
  input [255:0] x;
  input [255:0] y;
  input [255:0] n;
  output [255:0] o;
  input clk, rst, start;
  wire   \zout[0][256] , \zin[0][256] , \zin[0][255] , \zin[0][254] ,
         \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] ,
         \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] ,
         \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] ,
         \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] ,
         \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] ,
         \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] ,
         \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] ,
         \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] ,
         \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] ,
         \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] ,
         \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] ,
         \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] ,
         \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] ,
         \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] ,
         \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] ,
         \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] ,
         \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] ,
         \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] ,
         \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] ,
         \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] ,
         \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] ,
         \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] ,
         \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] ,
         \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] ,
         \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] ,
         \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] ,
         \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] ,
         \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] ,
         \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] ,
         \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] ,
         \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] ,
         \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] ,
         \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] ,
         \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] ,
         \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] ,
         \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] ,
         \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] ,
         \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] ,
         \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] ,
         \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] ,
         \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] ,
         \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] ,
         \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] ,
         \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] ,
         \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] ,
         \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] ,
         \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] ,
         \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] ,
         \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] ,
         \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] ,
         \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] ,
         \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] ,
         \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] ,
         \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] ,
         \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] ,
         \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] ,
         \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] ,
         \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] ,
         \zin[0][2] , \zin[0][1] , \zin[0][0] ;
  wire   [255:0] xin;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N256 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[255]), .y(y), .n(n), .zin({1'b0, \zin[0][256] , \zin[0][255] , \zin[0][254] , 
        \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] , 
        \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] , 
        \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] , 
        \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] , 
        \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] , 
        \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] , 
        \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] , 
        \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] , 
        \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] , 
        \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] , 
        \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] , 
        \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] , 
        \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] , 
        \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] , 
        \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] , 
        \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] , 
        \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] , 
        \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] , 
        \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] , 
        \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] , 
        \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] , 
        \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] , 
        \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] , 
        \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] , 
        \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] , 
        \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] , 
        \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] , 
        \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] , 
        \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] , 
        \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] , 
        \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] , 
        \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] , 
        \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] , 
        \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] , 
        \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] , 
        \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] , 
        \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] , 
        \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] , 
        \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] , \zin[0][97] , 
        \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] , \zin[0][92] , 
        \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] , \zin[0][87] , 
        \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] , \zin[0][82] , 
        \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] , \zin[0][77] , 
        \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] , \zin[0][72] , 
        \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] , \zin[0][67] , 
        \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] , \zin[0][62] , 
        \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] , \zin[0][57] , 
        \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] , \zin[0][52] , 
        \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] , \zin[0][47] , 
        \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] , \zin[0][42] , 
        \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] , \zin[0][37] , 
        \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] , \zin[0][32] , 
        \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] , \zin[0][27] , 
        \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] , \zin[0][22] , 
        \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] , \zin[0][17] , 
        \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] , \zin[0][12] , 
        \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] , \zin[0][7] , 
        \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] , \zin[0][2] , 
        \zin[0][1] , \zin[0][0] }), .zout({SYNOPSYS_UNCONNECTED__0, 
        \zout[0][256] , o}) );
  DFF \xreg_reg[0]  ( .D(1'b0), .CLK(clk), .RST(start), .I(x[0]), .Q(xin[0])
         );
  DFF \xreg_reg[1]  ( .D(xin[0]), .CLK(clk), .RST(start), .I(x[1]), .Q(xin[1])
         );
  DFF \xreg_reg[2]  ( .D(xin[1]), .CLK(clk), .RST(start), .I(x[2]), .Q(xin[2])
         );
  DFF \xreg_reg[3]  ( .D(xin[2]), .CLK(clk), .RST(start), .I(x[3]), .Q(xin[3])
         );
  DFF \xreg_reg[4]  ( .D(xin[3]), .CLK(clk), .RST(start), .I(x[4]), .Q(xin[4])
         );
  DFF \xreg_reg[5]  ( .D(xin[4]), .CLK(clk), .RST(start), .I(x[5]), .Q(xin[5])
         );
  DFF \xreg_reg[6]  ( .D(xin[5]), .CLK(clk), .RST(start), .I(x[6]), .Q(xin[6])
         );
  DFF \xreg_reg[7]  ( .D(xin[6]), .CLK(clk), .RST(start), .I(x[7]), .Q(xin[7])
         );
  DFF \xreg_reg[8]  ( .D(xin[7]), .CLK(clk), .RST(start), .I(x[8]), .Q(xin[8])
         );
  DFF \xreg_reg[9]  ( .D(xin[8]), .CLK(clk), .RST(start), .I(x[9]), .Q(xin[9])
         );
  DFF \xreg_reg[10]  ( .D(xin[9]), .CLK(clk), .RST(start), .I(x[10]), .Q(
        xin[10]) );
  DFF \xreg_reg[11]  ( .D(xin[10]), .CLK(clk), .RST(start), .I(x[11]), .Q(
        xin[11]) );
  DFF \xreg_reg[12]  ( .D(xin[11]), .CLK(clk), .RST(start), .I(x[12]), .Q(
        xin[12]) );
  DFF \xreg_reg[13]  ( .D(xin[12]), .CLK(clk), .RST(start), .I(x[13]), .Q(
        xin[13]) );
  DFF \xreg_reg[14]  ( .D(xin[13]), .CLK(clk), .RST(start), .I(x[14]), .Q(
        xin[14]) );
  DFF \xreg_reg[15]  ( .D(xin[14]), .CLK(clk), .RST(start), .I(x[15]), .Q(
        xin[15]) );
  DFF \xreg_reg[16]  ( .D(xin[15]), .CLK(clk), .RST(start), .I(x[16]), .Q(
        xin[16]) );
  DFF \xreg_reg[17]  ( .D(xin[16]), .CLK(clk), .RST(start), .I(x[17]), .Q(
        xin[17]) );
  DFF \xreg_reg[18]  ( .D(xin[17]), .CLK(clk), .RST(start), .I(x[18]), .Q(
        xin[18]) );
  DFF \xreg_reg[19]  ( .D(xin[18]), .CLK(clk), .RST(start), .I(x[19]), .Q(
        xin[19]) );
  DFF \xreg_reg[20]  ( .D(xin[19]), .CLK(clk), .RST(start), .I(x[20]), .Q(
        xin[20]) );
  DFF \xreg_reg[21]  ( .D(xin[20]), .CLK(clk), .RST(start), .I(x[21]), .Q(
        xin[21]) );
  DFF \xreg_reg[22]  ( .D(xin[21]), .CLK(clk), .RST(start), .I(x[22]), .Q(
        xin[22]) );
  DFF \xreg_reg[23]  ( .D(xin[22]), .CLK(clk), .RST(start), .I(x[23]), .Q(
        xin[23]) );
  DFF \xreg_reg[24]  ( .D(xin[23]), .CLK(clk), .RST(start), .I(x[24]), .Q(
        xin[24]) );
  DFF \xreg_reg[25]  ( .D(xin[24]), .CLK(clk), .RST(start), .I(x[25]), .Q(
        xin[25]) );
  DFF \xreg_reg[26]  ( .D(xin[25]), .CLK(clk), .RST(start), .I(x[26]), .Q(
        xin[26]) );
  DFF \xreg_reg[27]  ( .D(xin[26]), .CLK(clk), .RST(start), .I(x[27]), .Q(
        xin[27]) );
  DFF \xreg_reg[28]  ( .D(xin[27]), .CLK(clk), .RST(start), .I(x[28]), .Q(
        xin[28]) );
  DFF \xreg_reg[29]  ( .D(xin[28]), .CLK(clk), .RST(start), .I(x[29]), .Q(
        xin[29]) );
  DFF \xreg_reg[30]  ( .D(xin[29]), .CLK(clk), .RST(start), .I(x[30]), .Q(
        xin[30]) );
  DFF \xreg_reg[31]  ( .D(xin[30]), .CLK(clk), .RST(start), .I(x[31]), .Q(
        xin[31]) );
  DFF \xreg_reg[32]  ( .D(xin[31]), .CLK(clk), .RST(start), .I(x[32]), .Q(
        xin[32]) );
  DFF \xreg_reg[33]  ( .D(xin[32]), .CLK(clk), .RST(start), .I(x[33]), .Q(
        xin[33]) );
  DFF \xreg_reg[34]  ( .D(xin[33]), .CLK(clk), .RST(start), .I(x[34]), .Q(
        xin[34]) );
  DFF \xreg_reg[35]  ( .D(xin[34]), .CLK(clk), .RST(start), .I(x[35]), .Q(
        xin[35]) );
  DFF \xreg_reg[36]  ( .D(xin[35]), .CLK(clk), .RST(start), .I(x[36]), .Q(
        xin[36]) );
  DFF \xreg_reg[37]  ( .D(xin[36]), .CLK(clk), .RST(start), .I(x[37]), .Q(
        xin[37]) );
  DFF \xreg_reg[38]  ( .D(xin[37]), .CLK(clk), .RST(start), .I(x[38]), .Q(
        xin[38]) );
  DFF \xreg_reg[39]  ( .D(xin[38]), .CLK(clk), .RST(start), .I(x[39]), .Q(
        xin[39]) );
  DFF \xreg_reg[40]  ( .D(xin[39]), .CLK(clk), .RST(start), .I(x[40]), .Q(
        xin[40]) );
  DFF \xreg_reg[41]  ( .D(xin[40]), .CLK(clk), .RST(start), .I(x[41]), .Q(
        xin[41]) );
  DFF \xreg_reg[42]  ( .D(xin[41]), .CLK(clk), .RST(start), .I(x[42]), .Q(
        xin[42]) );
  DFF \xreg_reg[43]  ( .D(xin[42]), .CLK(clk), .RST(start), .I(x[43]), .Q(
        xin[43]) );
  DFF \xreg_reg[44]  ( .D(xin[43]), .CLK(clk), .RST(start), .I(x[44]), .Q(
        xin[44]) );
  DFF \xreg_reg[45]  ( .D(xin[44]), .CLK(clk), .RST(start), .I(x[45]), .Q(
        xin[45]) );
  DFF \xreg_reg[46]  ( .D(xin[45]), .CLK(clk), .RST(start), .I(x[46]), .Q(
        xin[46]) );
  DFF \xreg_reg[47]  ( .D(xin[46]), .CLK(clk), .RST(start), .I(x[47]), .Q(
        xin[47]) );
  DFF \xreg_reg[48]  ( .D(xin[47]), .CLK(clk), .RST(start), .I(x[48]), .Q(
        xin[48]) );
  DFF \xreg_reg[49]  ( .D(xin[48]), .CLK(clk), .RST(start), .I(x[49]), .Q(
        xin[49]) );
  DFF \xreg_reg[50]  ( .D(xin[49]), .CLK(clk), .RST(start), .I(x[50]), .Q(
        xin[50]) );
  DFF \xreg_reg[51]  ( .D(xin[50]), .CLK(clk), .RST(start), .I(x[51]), .Q(
        xin[51]) );
  DFF \xreg_reg[52]  ( .D(xin[51]), .CLK(clk), .RST(start), .I(x[52]), .Q(
        xin[52]) );
  DFF \xreg_reg[53]  ( .D(xin[52]), .CLK(clk), .RST(start), .I(x[53]), .Q(
        xin[53]) );
  DFF \xreg_reg[54]  ( .D(xin[53]), .CLK(clk), .RST(start), .I(x[54]), .Q(
        xin[54]) );
  DFF \xreg_reg[55]  ( .D(xin[54]), .CLK(clk), .RST(start), .I(x[55]), .Q(
        xin[55]) );
  DFF \xreg_reg[56]  ( .D(xin[55]), .CLK(clk), .RST(start), .I(x[56]), .Q(
        xin[56]) );
  DFF \xreg_reg[57]  ( .D(xin[56]), .CLK(clk), .RST(start), .I(x[57]), .Q(
        xin[57]) );
  DFF \xreg_reg[58]  ( .D(xin[57]), .CLK(clk), .RST(start), .I(x[58]), .Q(
        xin[58]) );
  DFF \xreg_reg[59]  ( .D(xin[58]), .CLK(clk), .RST(start), .I(x[59]), .Q(
        xin[59]) );
  DFF \xreg_reg[60]  ( .D(xin[59]), .CLK(clk), .RST(start), .I(x[60]), .Q(
        xin[60]) );
  DFF \xreg_reg[61]  ( .D(xin[60]), .CLK(clk), .RST(start), .I(x[61]), .Q(
        xin[61]) );
  DFF \xreg_reg[62]  ( .D(xin[61]), .CLK(clk), .RST(start), .I(x[62]), .Q(
        xin[62]) );
  DFF \xreg_reg[63]  ( .D(xin[62]), .CLK(clk), .RST(start), .I(x[63]), .Q(
        xin[63]) );
  DFF \xreg_reg[64]  ( .D(xin[63]), .CLK(clk), .RST(start), .I(x[64]), .Q(
        xin[64]) );
  DFF \xreg_reg[65]  ( .D(xin[64]), .CLK(clk), .RST(start), .I(x[65]), .Q(
        xin[65]) );
  DFF \xreg_reg[66]  ( .D(xin[65]), .CLK(clk), .RST(start), .I(x[66]), .Q(
        xin[66]) );
  DFF \xreg_reg[67]  ( .D(xin[66]), .CLK(clk), .RST(start), .I(x[67]), .Q(
        xin[67]) );
  DFF \xreg_reg[68]  ( .D(xin[67]), .CLK(clk), .RST(start), .I(x[68]), .Q(
        xin[68]) );
  DFF \xreg_reg[69]  ( .D(xin[68]), .CLK(clk), .RST(start), .I(x[69]), .Q(
        xin[69]) );
  DFF \xreg_reg[70]  ( .D(xin[69]), .CLK(clk), .RST(start), .I(x[70]), .Q(
        xin[70]) );
  DFF \xreg_reg[71]  ( .D(xin[70]), .CLK(clk), .RST(start), .I(x[71]), .Q(
        xin[71]) );
  DFF \xreg_reg[72]  ( .D(xin[71]), .CLK(clk), .RST(start), .I(x[72]), .Q(
        xin[72]) );
  DFF \xreg_reg[73]  ( .D(xin[72]), .CLK(clk), .RST(start), .I(x[73]), .Q(
        xin[73]) );
  DFF \xreg_reg[74]  ( .D(xin[73]), .CLK(clk), .RST(start), .I(x[74]), .Q(
        xin[74]) );
  DFF \xreg_reg[75]  ( .D(xin[74]), .CLK(clk), .RST(start), .I(x[75]), .Q(
        xin[75]) );
  DFF \xreg_reg[76]  ( .D(xin[75]), .CLK(clk), .RST(start), .I(x[76]), .Q(
        xin[76]) );
  DFF \xreg_reg[77]  ( .D(xin[76]), .CLK(clk), .RST(start), .I(x[77]), .Q(
        xin[77]) );
  DFF \xreg_reg[78]  ( .D(xin[77]), .CLK(clk), .RST(start), .I(x[78]), .Q(
        xin[78]) );
  DFF \xreg_reg[79]  ( .D(xin[78]), .CLK(clk), .RST(start), .I(x[79]), .Q(
        xin[79]) );
  DFF \xreg_reg[80]  ( .D(xin[79]), .CLK(clk), .RST(start), .I(x[80]), .Q(
        xin[80]) );
  DFF \xreg_reg[81]  ( .D(xin[80]), .CLK(clk), .RST(start), .I(x[81]), .Q(
        xin[81]) );
  DFF \xreg_reg[82]  ( .D(xin[81]), .CLK(clk), .RST(start), .I(x[82]), .Q(
        xin[82]) );
  DFF \xreg_reg[83]  ( .D(xin[82]), .CLK(clk), .RST(start), .I(x[83]), .Q(
        xin[83]) );
  DFF \xreg_reg[84]  ( .D(xin[83]), .CLK(clk), .RST(start), .I(x[84]), .Q(
        xin[84]) );
  DFF \xreg_reg[85]  ( .D(xin[84]), .CLK(clk), .RST(start), .I(x[85]), .Q(
        xin[85]) );
  DFF \xreg_reg[86]  ( .D(xin[85]), .CLK(clk), .RST(start), .I(x[86]), .Q(
        xin[86]) );
  DFF \xreg_reg[87]  ( .D(xin[86]), .CLK(clk), .RST(start), .I(x[87]), .Q(
        xin[87]) );
  DFF \xreg_reg[88]  ( .D(xin[87]), .CLK(clk), .RST(start), .I(x[88]), .Q(
        xin[88]) );
  DFF \xreg_reg[89]  ( .D(xin[88]), .CLK(clk), .RST(start), .I(x[89]), .Q(
        xin[89]) );
  DFF \xreg_reg[90]  ( .D(xin[89]), .CLK(clk), .RST(start), .I(x[90]), .Q(
        xin[90]) );
  DFF \xreg_reg[91]  ( .D(xin[90]), .CLK(clk), .RST(start), .I(x[91]), .Q(
        xin[91]) );
  DFF \xreg_reg[92]  ( .D(xin[91]), .CLK(clk), .RST(start), .I(x[92]), .Q(
        xin[92]) );
  DFF \xreg_reg[93]  ( .D(xin[92]), .CLK(clk), .RST(start), .I(x[93]), .Q(
        xin[93]) );
  DFF \xreg_reg[94]  ( .D(xin[93]), .CLK(clk), .RST(start), .I(x[94]), .Q(
        xin[94]) );
  DFF \xreg_reg[95]  ( .D(xin[94]), .CLK(clk), .RST(start), .I(x[95]), .Q(
        xin[95]) );
  DFF \xreg_reg[96]  ( .D(xin[95]), .CLK(clk), .RST(start), .I(x[96]), .Q(
        xin[96]) );
  DFF \xreg_reg[97]  ( .D(xin[96]), .CLK(clk), .RST(start), .I(x[97]), .Q(
        xin[97]) );
  DFF \xreg_reg[98]  ( .D(xin[97]), .CLK(clk), .RST(start), .I(x[98]), .Q(
        xin[98]) );
  DFF \xreg_reg[99]  ( .D(xin[98]), .CLK(clk), .RST(start), .I(x[99]), .Q(
        xin[99]) );
  DFF \xreg_reg[100]  ( .D(xin[99]), .CLK(clk), .RST(start), .I(x[100]), .Q(
        xin[100]) );
  DFF \xreg_reg[101]  ( .D(xin[100]), .CLK(clk), .RST(start), .I(x[101]), .Q(
        xin[101]) );
  DFF \xreg_reg[102]  ( .D(xin[101]), .CLK(clk), .RST(start), .I(x[102]), .Q(
        xin[102]) );
  DFF \xreg_reg[103]  ( .D(xin[102]), .CLK(clk), .RST(start), .I(x[103]), .Q(
        xin[103]) );
  DFF \xreg_reg[104]  ( .D(xin[103]), .CLK(clk), .RST(start), .I(x[104]), .Q(
        xin[104]) );
  DFF \xreg_reg[105]  ( .D(xin[104]), .CLK(clk), .RST(start), .I(x[105]), .Q(
        xin[105]) );
  DFF \xreg_reg[106]  ( .D(xin[105]), .CLK(clk), .RST(start), .I(x[106]), .Q(
        xin[106]) );
  DFF \xreg_reg[107]  ( .D(xin[106]), .CLK(clk), .RST(start), .I(x[107]), .Q(
        xin[107]) );
  DFF \xreg_reg[108]  ( .D(xin[107]), .CLK(clk), .RST(start), .I(x[108]), .Q(
        xin[108]) );
  DFF \xreg_reg[109]  ( .D(xin[108]), .CLK(clk), .RST(start), .I(x[109]), .Q(
        xin[109]) );
  DFF \xreg_reg[110]  ( .D(xin[109]), .CLK(clk), .RST(start), .I(x[110]), .Q(
        xin[110]) );
  DFF \xreg_reg[111]  ( .D(xin[110]), .CLK(clk), .RST(start), .I(x[111]), .Q(
        xin[111]) );
  DFF \xreg_reg[112]  ( .D(xin[111]), .CLK(clk), .RST(start), .I(x[112]), .Q(
        xin[112]) );
  DFF \xreg_reg[113]  ( .D(xin[112]), .CLK(clk), .RST(start), .I(x[113]), .Q(
        xin[113]) );
  DFF \xreg_reg[114]  ( .D(xin[113]), .CLK(clk), .RST(start), .I(x[114]), .Q(
        xin[114]) );
  DFF \xreg_reg[115]  ( .D(xin[114]), .CLK(clk), .RST(start), .I(x[115]), .Q(
        xin[115]) );
  DFF \xreg_reg[116]  ( .D(xin[115]), .CLK(clk), .RST(start), .I(x[116]), .Q(
        xin[116]) );
  DFF \xreg_reg[117]  ( .D(xin[116]), .CLK(clk), .RST(start), .I(x[117]), .Q(
        xin[117]) );
  DFF \xreg_reg[118]  ( .D(xin[117]), .CLK(clk), .RST(start), .I(x[118]), .Q(
        xin[118]) );
  DFF \xreg_reg[119]  ( .D(xin[118]), .CLK(clk), .RST(start), .I(x[119]), .Q(
        xin[119]) );
  DFF \xreg_reg[120]  ( .D(xin[119]), .CLK(clk), .RST(start), .I(x[120]), .Q(
        xin[120]) );
  DFF \xreg_reg[121]  ( .D(xin[120]), .CLK(clk), .RST(start), .I(x[121]), .Q(
        xin[121]) );
  DFF \xreg_reg[122]  ( .D(xin[121]), .CLK(clk), .RST(start), .I(x[122]), .Q(
        xin[122]) );
  DFF \xreg_reg[123]  ( .D(xin[122]), .CLK(clk), .RST(start), .I(x[123]), .Q(
        xin[123]) );
  DFF \xreg_reg[124]  ( .D(xin[123]), .CLK(clk), .RST(start), .I(x[124]), .Q(
        xin[124]) );
  DFF \xreg_reg[125]  ( .D(xin[124]), .CLK(clk), .RST(start), .I(x[125]), .Q(
        xin[125]) );
  DFF \xreg_reg[126]  ( .D(xin[125]), .CLK(clk), .RST(start), .I(x[126]), .Q(
        xin[126]) );
  DFF \xreg_reg[127]  ( .D(xin[126]), .CLK(clk), .RST(start), .I(x[127]), .Q(
        xin[127]) );
  DFF \xreg_reg[128]  ( .D(xin[127]), .CLK(clk), .RST(start), .I(x[128]), .Q(
        xin[128]) );
  DFF \xreg_reg[129]  ( .D(xin[128]), .CLK(clk), .RST(start), .I(x[129]), .Q(
        xin[129]) );
  DFF \xreg_reg[130]  ( .D(xin[129]), .CLK(clk), .RST(start), .I(x[130]), .Q(
        xin[130]) );
  DFF \xreg_reg[131]  ( .D(xin[130]), .CLK(clk), .RST(start), .I(x[131]), .Q(
        xin[131]) );
  DFF \xreg_reg[132]  ( .D(xin[131]), .CLK(clk), .RST(start), .I(x[132]), .Q(
        xin[132]) );
  DFF \xreg_reg[133]  ( .D(xin[132]), .CLK(clk), .RST(start), .I(x[133]), .Q(
        xin[133]) );
  DFF \xreg_reg[134]  ( .D(xin[133]), .CLK(clk), .RST(start), .I(x[134]), .Q(
        xin[134]) );
  DFF \xreg_reg[135]  ( .D(xin[134]), .CLK(clk), .RST(start), .I(x[135]), .Q(
        xin[135]) );
  DFF \xreg_reg[136]  ( .D(xin[135]), .CLK(clk), .RST(start), .I(x[136]), .Q(
        xin[136]) );
  DFF \xreg_reg[137]  ( .D(xin[136]), .CLK(clk), .RST(start), .I(x[137]), .Q(
        xin[137]) );
  DFF \xreg_reg[138]  ( .D(xin[137]), .CLK(clk), .RST(start), .I(x[138]), .Q(
        xin[138]) );
  DFF \xreg_reg[139]  ( .D(xin[138]), .CLK(clk), .RST(start), .I(x[139]), .Q(
        xin[139]) );
  DFF \xreg_reg[140]  ( .D(xin[139]), .CLK(clk), .RST(start), .I(x[140]), .Q(
        xin[140]) );
  DFF \xreg_reg[141]  ( .D(xin[140]), .CLK(clk), .RST(start), .I(x[141]), .Q(
        xin[141]) );
  DFF \xreg_reg[142]  ( .D(xin[141]), .CLK(clk), .RST(start), .I(x[142]), .Q(
        xin[142]) );
  DFF \xreg_reg[143]  ( .D(xin[142]), .CLK(clk), .RST(start), .I(x[143]), .Q(
        xin[143]) );
  DFF \xreg_reg[144]  ( .D(xin[143]), .CLK(clk), .RST(start), .I(x[144]), .Q(
        xin[144]) );
  DFF \xreg_reg[145]  ( .D(xin[144]), .CLK(clk), .RST(start), .I(x[145]), .Q(
        xin[145]) );
  DFF \xreg_reg[146]  ( .D(xin[145]), .CLK(clk), .RST(start), .I(x[146]), .Q(
        xin[146]) );
  DFF \xreg_reg[147]  ( .D(xin[146]), .CLK(clk), .RST(start), .I(x[147]), .Q(
        xin[147]) );
  DFF \xreg_reg[148]  ( .D(xin[147]), .CLK(clk), .RST(start), .I(x[148]), .Q(
        xin[148]) );
  DFF \xreg_reg[149]  ( .D(xin[148]), .CLK(clk), .RST(start), .I(x[149]), .Q(
        xin[149]) );
  DFF \xreg_reg[150]  ( .D(xin[149]), .CLK(clk), .RST(start), .I(x[150]), .Q(
        xin[150]) );
  DFF \xreg_reg[151]  ( .D(xin[150]), .CLK(clk), .RST(start), .I(x[151]), .Q(
        xin[151]) );
  DFF \xreg_reg[152]  ( .D(xin[151]), .CLK(clk), .RST(start), .I(x[152]), .Q(
        xin[152]) );
  DFF \xreg_reg[153]  ( .D(xin[152]), .CLK(clk), .RST(start), .I(x[153]), .Q(
        xin[153]) );
  DFF \xreg_reg[154]  ( .D(xin[153]), .CLK(clk), .RST(start), .I(x[154]), .Q(
        xin[154]) );
  DFF \xreg_reg[155]  ( .D(xin[154]), .CLK(clk), .RST(start), .I(x[155]), .Q(
        xin[155]) );
  DFF \xreg_reg[156]  ( .D(xin[155]), .CLK(clk), .RST(start), .I(x[156]), .Q(
        xin[156]) );
  DFF \xreg_reg[157]  ( .D(xin[156]), .CLK(clk), .RST(start), .I(x[157]), .Q(
        xin[157]) );
  DFF \xreg_reg[158]  ( .D(xin[157]), .CLK(clk), .RST(start), .I(x[158]), .Q(
        xin[158]) );
  DFF \xreg_reg[159]  ( .D(xin[158]), .CLK(clk), .RST(start), .I(x[159]), .Q(
        xin[159]) );
  DFF \xreg_reg[160]  ( .D(xin[159]), .CLK(clk), .RST(start), .I(x[160]), .Q(
        xin[160]) );
  DFF \xreg_reg[161]  ( .D(xin[160]), .CLK(clk), .RST(start), .I(x[161]), .Q(
        xin[161]) );
  DFF \xreg_reg[162]  ( .D(xin[161]), .CLK(clk), .RST(start), .I(x[162]), .Q(
        xin[162]) );
  DFF \xreg_reg[163]  ( .D(xin[162]), .CLK(clk), .RST(start), .I(x[163]), .Q(
        xin[163]) );
  DFF \xreg_reg[164]  ( .D(xin[163]), .CLK(clk), .RST(start), .I(x[164]), .Q(
        xin[164]) );
  DFF \xreg_reg[165]  ( .D(xin[164]), .CLK(clk), .RST(start), .I(x[165]), .Q(
        xin[165]) );
  DFF \xreg_reg[166]  ( .D(xin[165]), .CLK(clk), .RST(start), .I(x[166]), .Q(
        xin[166]) );
  DFF \xreg_reg[167]  ( .D(xin[166]), .CLK(clk), .RST(start), .I(x[167]), .Q(
        xin[167]) );
  DFF \xreg_reg[168]  ( .D(xin[167]), .CLK(clk), .RST(start), .I(x[168]), .Q(
        xin[168]) );
  DFF \xreg_reg[169]  ( .D(xin[168]), .CLK(clk), .RST(start), .I(x[169]), .Q(
        xin[169]) );
  DFF \xreg_reg[170]  ( .D(xin[169]), .CLK(clk), .RST(start), .I(x[170]), .Q(
        xin[170]) );
  DFF \xreg_reg[171]  ( .D(xin[170]), .CLK(clk), .RST(start), .I(x[171]), .Q(
        xin[171]) );
  DFF \xreg_reg[172]  ( .D(xin[171]), .CLK(clk), .RST(start), .I(x[172]), .Q(
        xin[172]) );
  DFF \xreg_reg[173]  ( .D(xin[172]), .CLK(clk), .RST(start), .I(x[173]), .Q(
        xin[173]) );
  DFF \xreg_reg[174]  ( .D(xin[173]), .CLK(clk), .RST(start), .I(x[174]), .Q(
        xin[174]) );
  DFF \xreg_reg[175]  ( .D(xin[174]), .CLK(clk), .RST(start), .I(x[175]), .Q(
        xin[175]) );
  DFF \xreg_reg[176]  ( .D(xin[175]), .CLK(clk), .RST(start), .I(x[176]), .Q(
        xin[176]) );
  DFF \xreg_reg[177]  ( .D(xin[176]), .CLK(clk), .RST(start), .I(x[177]), .Q(
        xin[177]) );
  DFF \xreg_reg[178]  ( .D(xin[177]), .CLK(clk), .RST(start), .I(x[178]), .Q(
        xin[178]) );
  DFF \xreg_reg[179]  ( .D(xin[178]), .CLK(clk), .RST(start), .I(x[179]), .Q(
        xin[179]) );
  DFF \xreg_reg[180]  ( .D(xin[179]), .CLK(clk), .RST(start), .I(x[180]), .Q(
        xin[180]) );
  DFF \xreg_reg[181]  ( .D(xin[180]), .CLK(clk), .RST(start), .I(x[181]), .Q(
        xin[181]) );
  DFF \xreg_reg[182]  ( .D(xin[181]), .CLK(clk), .RST(start), .I(x[182]), .Q(
        xin[182]) );
  DFF \xreg_reg[183]  ( .D(xin[182]), .CLK(clk), .RST(start), .I(x[183]), .Q(
        xin[183]) );
  DFF \xreg_reg[184]  ( .D(xin[183]), .CLK(clk), .RST(start), .I(x[184]), .Q(
        xin[184]) );
  DFF \xreg_reg[185]  ( .D(xin[184]), .CLK(clk), .RST(start), .I(x[185]), .Q(
        xin[185]) );
  DFF \xreg_reg[186]  ( .D(xin[185]), .CLK(clk), .RST(start), .I(x[186]), .Q(
        xin[186]) );
  DFF \xreg_reg[187]  ( .D(xin[186]), .CLK(clk), .RST(start), .I(x[187]), .Q(
        xin[187]) );
  DFF \xreg_reg[188]  ( .D(xin[187]), .CLK(clk), .RST(start), .I(x[188]), .Q(
        xin[188]) );
  DFF \xreg_reg[189]  ( .D(xin[188]), .CLK(clk), .RST(start), .I(x[189]), .Q(
        xin[189]) );
  DFF \xreg_reg[190]  ( .D(xin[189]), .CLK(clk), .RST(start), .I(x[190]), .Q(
        xin[190]) );
  DFF \xreg_reg[191]  ( .D(xin[190]), .CLK(clk), .RST(start), .I(x[191]), .Q(
        xin[191]) );
  DFF \xreg_reg[192]  ( .D(xin[191]), .CLK(clk), .RST(start), .I(x[192]), .Q(
        xin[192]) );
  DFF \xreg_reg[193]  ( .D(xin[192]), .CLK(clk), .RST(start), .I(x[193]), .Q(
        xin[193]) );
  DFF \xreg_reg[194]  ( .D(xin[193]), .CLK(clk), .RST(start), .I(x[194]), .Q(
        xin[194]) );
  DFF \xreg_reg[195]  ( .D(xin[194]), .CLK(clk), .RST(start), .I(x[195]), .Q(
        xin[195]) );
  DFF \xreg_reg[196]  ( .D(xin[195]), .CLK(clk), .RST(start), .I(x[196]), .Q(
        xin[196]) );
  DFF \xreg_reg[197]  ( .D(xin[196]), .CLK(clk), .RST(start), .I(x[197]), .Q(
        xin[197]) );
  DFF \xreg_reg[198]  ( .D(xin[197]), .CLK(clk), .RST(start), .I(x[198]), .Q(
        xin[198]) );
  DFF \xreg_reg[199]  ( .D(xin[198]), .CLK(clk), .RST(start), .I(x[199]), .Q(
        xin[199]) );
  DFF \xreg_reg[200]  ( .D(xin[199]), .CLK(clk), .RST(start), .I(x[200]), .Q(
        xin[200]) );
  DFF \xreg_reg[201]  ( .D(xin[200]), .CLK(clk), .RST(start), .I(x[201]), .Q(
        xin[201]) );
  DFF \xreg_reg[202]  ( .D(xin[201]), .CLK(clk), .RST(start), .I(x[202]), .Q(
        xin[202]) );
  DFF \xreg_reg[203]  ( .D(xin[202]), .CLK(clk), .RST(start), .I(x[203]), .Q(
        xin[203]) );
  DFF \xreg_reg[204]  ( .D(xin[203]), .CLK(clk), .RST(start), .I(x[204]), .Q(
        xin[204]) );
  DFF \xreg_reg[205]  ( .D(xin[204]), .CLK(clk), .RST(start), .I(x[205]), .Q(
        xin[205]) );
  DFF \xreg_reg[206]  ( .D(xin[205]), .CLK(clk), .RST(start), .I(x[206]), .Q(
        xin[206]) );
  DFF \xreg_reg[207]  ( .D(xin[206]), .CLK(clk), .RST(start), .I(x[207]), .Q(
        xin[207]) );
  DFF \xreg_reg[208]  ( .D(xin[207]), .CLK(clk), .RST(start), .I(x[208]), .Q(
        xin[208]) );
  DFF \xreg_reg[209]  ( .D(xin[208]), .CLK(clk), .RST(start), .I(x[209]), .Q(
        xin[209]) );
  DFF \xreg_reg[210]  ( .D(xin[209]), .CLK(clk), .RST(start), .I(x[210]), .Q(
        xin[210]) );
  DFF \xreg_reg[211]  ( .D(xin[210]), .CLK(clk), .RST(start), .I(x[211]), .Q(
        xin[211]) );
  DFF \xreg_reg[212]  ( .D(xin[211]), .CLK(clk), .RST(start), .I(x[212]), .Q(
        xin[212]) );
  DFF \xreg_reg[213]  ( .D(xin[212]), .CLK(clk), .RST(start), .I(x[213]), .Q(
        xin[213]) );
  DFF \xreg_reg[214]  ( .D(xin[213]), .CLK(clk), .RST(start), .I(x[214]), .Q(
        xin[214]) );
  DFF \xreg_reg[215]  ( .D(xin[214]), .CLK(clk), .RST(start), .I(x[215]), .Q(
        xin[215]) );
  DFF \xreg_reg[216]  ( .D(xin[215]), .CLK(clk), .RST(start), .I(x[216]), .Q(
        xin[216]) );
  DFF \xreg_reg[217]  ( .D(xin[216]), .CLK(clk), .RST(start), .I(x[217]), .Q(
        xin[217]) );
  DFF \xreg_reg[218]  ( .D(xin[217]), .CLK(clk), .RST(start), .I(x[218]), .Q(
        xin[218]) );
  DFF \xreg_reg[219]  ( .D(xin[218]), .CLK(clk), .RST(start), .I(x[219]), .Q(
        xin[219]) );
  DFF \xreg_reg[220]  ( .D(xin[219]), .CLK(clk), .RST(start), .I(x[220]), .Q(
        xin[220]) );
  DFF \xreg_reg[221]  ( .D(xin[220]), .CLK(clk), .RST(start), .I(x[221]), .Q(
        xin[221]) );
  DFF \xreg_reg[222]  ( .D(xin[221]), .CLK(clk), .RST(start), .I(x[222]), .Q(
        xin[222]) );
  DFF \xreg_reg[223]  ( .D(xin[222]), .CLK(clk), .RST(start), .I(x[223]), .Q(
        xin[223]) );
  DFF \xreg_reg[224]  ( .D(xin[223]), .CLK(clk), .RST(start), .I(x[224]), .Q(
        xin[224]) );
  DFF \xreg_reg[225]  ( .D(xin[224]), .CLK(clk), .RST(start), .I(x[225]), .Q(
        xin[225]) );
  DFF \xreg_reg[226]  ( .D(xin[225]), .CLK(clk), .RST(start), .I(x[226]), .Q(
        xin[226]) );
  DFF \xreg_reg[227]  ( .D(xin[226]), .CLK(clk), .RST(start), .I(x[227]), .Q(
        xin[227]) );
  DFF \xreg_reg[228]  ( .D(xin[227]), .CLK(clk), .RST(start), .I(x[228]), .Q(
        xin[228]) );
  DFF \xreg_reg[229]  ( .D(xin[228]), .CLK(clk), .RST(start), .I(x[229]), .Q(
        xin[229]) );
  DFF \xreg_reg[230]  ( .D(xin[229]), .CLK(clk), .RST(start), .I(x[230]), .Q(
        xin[230]) );
  DFF \xreg_reg[231]  ( .D(xin[230]), .CLK(clk), .RST(start), .I(x[231]), .Q(
        xin[231]) );
  DFF \xreg_reg[232]  ( .D(xin[231]), .CLK(clk), .RST(start), .I(x[232]), .Q(
        xin[232]) );
  DFF \xreg_reg[233]  ( .D(xin[232]), .CLK(clk), .RST(start), .I(x[233]), .Q(
        xin[233]) );
  DFF \xreg_reg[234]  ( .D(xin[233]), .CLK(clk), .RST(start), .I(x[234]), .Q(
        xin[234]) );
  DFF \xreg_reg[235]  ( .D(xin[234]), .CLK(clk), .RST(start), .I(x[235]), .Q(
        xin[235]) );
  DFF \xreg_reg[236]  ( .D(xin[235]), .CLK(clk), .RST(start), .I(x[236]), .Q(
        xin[236]) );
  DFF \xreg_reg[237]  ( .D(xin[236]), .CLK(clk), .RST(start), .I(x[237]), .Q(
        xin[237]) );
  DFF \xreg_reg[238]  ( .D(xin[237]), .CLK(clk), .RST(start), .I(x[238]), .Q(
        xin[238]) );
  DFF \xreg_reg[239]  ( .D(xin[238]), .CLK(clk), .RST(start), .I(x[239]), .Q(
        xin[239]) );
  DFF \xreg_reg[240]  ( .D(xin[239]), .CLK(clk), .RST(start), .I(x[240]), .Q(
        xin[240]) );
  DFF \xreg_reg[241]  ( .D(xin[240]), .CLK(clk), .RST(start), .I(x[241]), .Q(
        xin[241]) );
  DFF \xreg_reg[242]  ( .D(xin[241]), .CLK(clk), .RST(start), .I(x[242]), .Q(
        xin[242]) );
  DFF \xreg_reg[243]  ( .D(xin[242]), .CLK(clk), .RST(start), .I(x[243]), .Q(
        xin[243]) );
  DFF \xreg_reg[244]  ( .D(xin[243]), .CLK(clk), .RST(start), .I(x[244]), .Q(
        xin[244]) );
  DFF \xreg_reg[245]  ( .D(xin[244]), .CLK(clk), .RST(start), .I(x[245]), .Q(
        xin[245]) );
  DFF \xreg_reg[246]  ( .D(xin[245]), .CLK(clk), .RST(start), .I(x[246]), .Q(
        xin[246]) );
  DFF \xreg_reg[247]  ( .D(xin[246]), .CLK(clk), .RST(start), .I(x[247]), .Q(
        xin[247]) );
  DFF \xreg_reg[248]  ( .D(xin[247]), .CLK(clk), .RST(start), .I(x[248]), .Q(
        xin[248]) );
  DFF \xreg_reg[249]  ( .D(xin[248]), .CLK(clk), .RST(start), .I(x[249]), .Q(
        xin[249]) );
  DFF \xreg_reg[250]  ( .D(xin[249]), .CLK(clk), .RST(start), .I(x[250]), .Q(
        xin[250]) );
  DFF \xreg_reg[251]  ( .D(xin[250]), .CLK(clk), .RST(start), .I(x[251]), .Q(
        xin[251]) );
  DFF \xreg_reg[252]  ( .D(xin[251]), .CLK(clk), .RST(start), .I(x[252]), .Q(
        xin[252]) );
  DFF \xreg_reg[253]  ( .D(xin[252]), .CLK(clk), .RST(start), .I(x[253]), .Q(
        xin[253]) );
  DFF \xreg_reg[254]  ( .D(xin[253]), .CLK(clk), .RST(start), .I(x[254]), .Q(
        xin[254]) );
  DFF \xreg_reg[255]  ( .D(xin[254]), .CLK(clk), .RST(start), .I(x[255]), .Q(
        xin[255]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][0] ) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1] ) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][2] ) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][3] ) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][4] ) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][5] ) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][6] ) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][7] ) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][8] ) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][9] ) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][10] ) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][11] ) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][12] ) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][13] ) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][14] ) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][15] ) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][16] ) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][17] ) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][18] ) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][19] ) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][20] ) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][21] ) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][22] ) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][23] ) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][24] ) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][25] ) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][26] ) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][27] ) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][28] ) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][29] ) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][30] ) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][31] ) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][32] ) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][33] ) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][34] ) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][35] ) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][36] ) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][37] ) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][38] ) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][39] ) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][40] ) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][41] ) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][42] ) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][43] ) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][44] ) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][45] ) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][46] ) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][47] ) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][48] ) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][49] ) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][50] ) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][51] ) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][52] ) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][53] ) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][54] ) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][55] ) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][56] ) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][57] ) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][58] ) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][59] ) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][60] ) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][61] ) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][62] ) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][63] ) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][64] ) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][65] ) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][66] ) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][67] ) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][68] ) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][69] ) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][70] ) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][71] ) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][72] ) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][73] ) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][74] ) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][75] ) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][76] ) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][77] ) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][78] ) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][79] ) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][80] ) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][81] ) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][82] ) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][83] ) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][84] ) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][85] ) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][86] ) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][87] ) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][88] ) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][89] ) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][90] ) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][91] ) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][92] ) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][93] ) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][94] ) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][95] ) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][96] ) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][97] ) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][98] ) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][99] ) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][100] ) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][101] ) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][102] ) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][103] ) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][104] ) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][105] ) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][106] ) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][107] ) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][108] ) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][109] ) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][110] ) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][111] ) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][112] ) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][113] ) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][114] ) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][115] ) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][116] ) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][117] ) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][118] ) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][119] ) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][120] ) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][121] ) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][122] ) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][123] ) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][124] ) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][125] ) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][126] ) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][127] ) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][128] ) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][129] ) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][130] ) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][131] ) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][132] ) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][133] ) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][134] ) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][135] ) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][136] ) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][137] ) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][138] ) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][139] ) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][140] ) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][141] ) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][142] ) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][143] ) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][144] ) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][145] ) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][146] ) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][147] ) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][148] ) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][149] ) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][150] ) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][151] ) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][152] ) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][153] ) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][154] ) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][155] ) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][156] ) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][157] ) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][158] ) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][159] ) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][160] ) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][161] ) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][162] ) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][163] ) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][164] ) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][165] ) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][166] ) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][167] ) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][168] ) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][169] ) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][170] ) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][171] ) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][172] ) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][173] ) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][174] ) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][175] ) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][176] ) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][177] ) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][178] ) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][179] ) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][180] ) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][181] ) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][182] ) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][183] ) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][184] ) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][185] ) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][186] ) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][187] ) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][188] ) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][189] ) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][190] ) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][191] ) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][192] ) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][193] ) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][194] ) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][195] ) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][196] ) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][197] ) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][198] ) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][199] ) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][200] ) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][201] ) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][202] ) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][203] ) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][204] ) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][205] ) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][206] ) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][207] ) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][208] ) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][209] ) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][210] ) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][211] ) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][212] ) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][213] ) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][214] ) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][215] ) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][216] ) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][217] ) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][218] ) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][219] ) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][220] ) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][221] ) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][222] ) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][223] ) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][224] ) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][225] ) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][226] ) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][227] ) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][228] ) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][229] ) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][230] ) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][231] ) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][232] ) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][233] ) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][234] ) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][235] ) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][236] ) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][237] ) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][238] ) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][239] ) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][240] ) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][241] ) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][242] ) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][243] ) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][244] ) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][245] ) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][246] ) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][247] ) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][248] ) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][249] ) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][250] ) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][251] ) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][252] ) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][253] ) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][254] ) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][255] ) );
  DFF \zreg_reg[256]  ( .D(\zout[0][256] ), .CLK(clk), .RST(start), .I(1'b0), 
        .Q(\zin[0][256] ) );
endmodule


module MUX_N256_1 ( A, B, S, O );
  input [255:0] A;
  input [255:0] B;
  output [255:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[50]), .B(n109), .Z(O[50]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U166 ( .A(A[4]), .B(n111), .Z(O[4]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U169 ( .A(A[49]), .B(n113), .Z(O[49]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U172 ( .A(A[48]), .B(n115), .Z(O[48]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U175 ( .A(A[47]), .B(n117), .Z(O[47]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U178 ( .A(A[46]), .B(n119), .Z(O[46]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U181 ( .A(A[45]), .B(n121), .Z(O[45]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U184 ( .A(A[44]), .B(n123), .Z(O[44]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U187 ( .A(A[43]), .B(n125), .Z(O[43]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U190 ( .A(A[42]), .B(n127), .Z(O[42]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U193 ( .A(A[41]), .B(n129), .Z(O[41]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U196 ( .A(A[40]), .B(n131), .Z(O[40]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U199 ( .A(A[3]), .B(n133), .Z(O[3]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U202 ( .A(A[39]), .B(n135), .Z(O[39]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U205 ( .A(A[38]), .B(n137), .Z(O[38]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U208 ( .A(A[37]), .B(n139), .Z(O[37]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U211 ( .A(A[36]), .B(n141), .Z(O[36]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U214 ( .A(A[35]), .B(n143), .Z(O[35]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U217 ( .A(A[34]), .B(n145), .Z(O[34]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U220 ( .A(A[33]), .B(n147), .Z(O[33]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U223 ( .A(A[32]), .B(n149), .Z(O[32]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U226 ( .A(A[31]), .B(n151), .Z(O[31]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U229 ( .A(A[30]), .B(n153), .Z(O[30]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U232 ( .A(A[2]), .B(n155), .Z(O[2]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U235 ( .A(A[29]), .B(n157), .Z(O[29]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U238 ( .A(A[28]), .B(n159), .Z(O[28]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U241 ( .A(A[27]), .B(n161), .Z(O[27]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U244 ( .A(A[26]), .B(n163), .Z(O[26]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U247 ( .A(A[25]), .B(n165), .Z(O[25]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U250 ( .A(A[255]), .B(n167), .Z(O[255]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[255]), .B(A[255]), .Z(n168) );
  XOR U253 ( .A(A[254]), .B(n169), .Z(O[254]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[254]), .B(A[254]), .Z(n170) );
  XOR U256 ( .A(A[253]), .B(n171), .Z(O[253]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[253]), .B(A[253]), .Z(n172) );
  XOR U259 ( .A(A[252]), .B(n173), .Z(O[252]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[252]), .B(A[252]), .Z(n174) );
  XOR U262 ( .A(A[251]), .B(n175), .Z(O[251]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[251]), .B(A[251]), .Z(n176) );
  XOR U265 ( .A(A[250]), .B(n177), .Z(O[250]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[250]), .B(A[250]), .Z(n178) );
  XOR U268 ( .A(A[24]), .B(n179), .Z(O[24]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[24]), .B(A[24]), .Z(n180) );
  XOR U271 ( .A(A[249]), .B(n181), .Z(O[249]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[249]), .B(A[249]), .Z(n182) );
  XOR U274 ( .A(A[248]), .B(n183), .Z(O[248]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[248]), .B(A[248]), .Z(n184) );
  XOR U277 ( .A(A[247]), .B(n185), .Z(O[247]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[247]), .B(A[247]), .Z(n186) );
  XOR U280 ( .A(A[246]), .B(n187), .Z(O[246]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[246]), .B(A[246]), .Z(n188) );
  XOR U283 ( .A(A[245]), .B(n189), .Z(O[245]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[245]), .B(A[245]), .Z(n190) );
  XOR U286 ( .A(A[244]), .B(n191), .Z(O[244]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[244]), .B(A[244]), .Z(n192) );
  XOR U289 ( .A(A[243]), .B(n193), .Z(O[243]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[243]), .B(A[243]), .Z(n194) );
  XOR U292 ( .A(A[242]), .B(n195), .Z(O[242]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[242]), .B(A[242]), .Z(n196) );
  XOR U295 ( .A(A[241]), .B(n197), .Z(O[241]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[241]), .B(A[241]), .Z(n198) );
  XOR U298 ( .A(A[240]), .B(n199), .Z(O[240]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[240]), .B(A[240]), .Z(n200) );
  XOR U301 ( .A(A[23]), .B(n201), .Z(O[23]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[23]), .B(A[23]), .Z(n202) );
  XOR U304 ( .A(A[239]), .B(n203), .Z(O[239]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[239]), .B(A[239]), .Z(n204) );
  XOR U307 ( .A(A[238]), .B(n205), .Z(O[238]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[238]), .B(A[238]), .Z(n206) );
  XOR U310 ( .A(A[237]), .B(n207), .Z(O[237]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[237]), .B(A[237]), .Z(n208) );
  XOR U313 ( .A(A[236]), .B(n209), .Z(O[236]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[236]), .B(A[236]), .Z(n210) );
  XOR U316 ( .A(A[235]), .B(n211), .Z(O[235]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[235]), .B(A[235]), .Z(n212) );
  XOR U319 ( .A(A[234]), .B(n213), .Z(O[234]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[234]), .B(A[234]), .Z(n214) );
  XOR U322 ( .A(A[233]), .B(n215), .Z(O[233]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[233]), .B(A[233]), .Z(n216) );
  XOR U325 ( .A(A[232]), .B(n217), .Z(O[232]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[232]), .B(A[232]), .Z(n218) );
  XOR U328 ( .A(A[231]), .B(n219), .Z(O[231]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[231]), .B(A[231]), .Z(n220) );
  XOR U331 ( .A(A[230]), .B(n221), .Z(O[230]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[230]), .B(A[230]), .Z(n222) );
  XOR U334 ( .A(A[22]), .B(n223), .Z(O[22]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[22]), .B(A[22]), .Z(n224) );
  XOR U337 ( .A(A[229]), .B(n225), .Z(O[229]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n226) );
  XOR U340 ( .A(A[228]), .B(n227), .Z(O[228]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[228]), .B(A[228]), .Z(n228) );
  XOR U343 ( .A(A[227]), .B(n229), .Z(O[227]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[227]), .B(A[227]), .Z(n230) );
  XOR U346 ( .A(A[226]), .B(n231), .Z(O[226]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[226]), .B(A[226]), .Z(n232) );
  XOR U349 ( .A(A[225]), .B(n233), .Z(O[225]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[225]), .B(A[225]), .Z(n234) );
  XOR U352 ( .A(A[224]), .B(n235), .Z(O[224]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[224]), .B(A[224]), .Z(n236) );
  XOR U355 ( .A(A[223]), .B(n237), .Z(O[223]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[223]), .B(A[223]), .Z(n238) );
  XOR U358 ( .A(A[222]), .B(n239), .Z(O[222]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[222]), .B(A[222]), .Z(n240) );
  XOR U361 ( .A(A[221]), .B(n241), .Z(O[221]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[221]), .B(A[221]), .Z(n242) );
  XOR U364 ( .A(A[220]), .B(n243), .Z(O[220]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[220]), .B(A[220]), .Z(n244) );
  XOR U367 ( .A(A[21]), .B(n245), .Z(O[21]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[21]), .B(A[21]), .Z(n246) );
  XOR U370 ( .A(A[219]), .B(n247), .Z(O[219]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[219]), .B(A[219]), .Z(n248) );
  XOR U373 ( .A(A[218]), .B(n249), .Z(O[218]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[218]), .B(A[218]), .Z(n250) );
  XOR U376 ( .A(A[217]), .B(n251), .Z(O[217]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[217]), .B(A[217]), .Z(n252) );
  XOR U379 ( .A(A[216]), .B(n253), .Z(O[216]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[216]), .B(A[216]), .Z(n254) );
  XOR U382 ( .A(A[215]), .B(n255), .Z(O[215]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[215]), .B(A[215]), .Z(n256) );
  XOR U385 ( .A(A[214]), .B(n257), .Z(O[214]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[214]), .B(A[214]), .Z(n258) );
  XOR U388 ( .A(A[213]), .B(n259), .Z(O[213]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[213]), .B(A[213]), .Z(n260) );
  XOR U391 ( .A(A[212]), .B(n261), .Z(O[212]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[212]), .B(A[212]), .Z(n262) );
  XOR U394 ( .A(A[211]), .B(n263), .Z(O[211]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[211]), .B(A[211]), .Z(n264) );
  XOR U397 ( .A(A[210]), .B(n265), .Z(O[210]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[210]), .B(A[210]), .Z(n266) );
  XOR U400 ( .A(A[20]), .B(n267), .Z(O[20]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[20]), .B(A[20]), .Z(n268) );
  XOR U403 ( .A(A[209]), .B(n269), .Z(O[209]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[209]), .B(A[209]), .Z(n270) );
  XOR U406 ( .A(A[208]), .B(n271), .Z(O[208]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[208]), .B(A[208]), .Z(n272) );
  XOR U409 ( .A(A[207]), .B(n273), .Z(O[207]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[207]), .B(A[207]), .Z(n274) );
  XOR U412 ( .A(A[206]), .B(n275), .Z(O[206]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[206]), .B(A[206]), .Z(n276) );
  XOR U415 ( .A(A[205]), .B(n277), .Z(O[205]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[205]), .B(A[205]), .Z(n278) );
  XOR U418 ( .A(A[204]), .B(n279), .Z(O[204]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[204]), .B(A[204]), .Z(n280) );
  XOR U421 ( .A(A[203]), .B(n281), .Z(O[203]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[203]), .B(A[203]), .Z(n282) );
  XOR U424 ( .A(A[202]), .B(n283), .Z(O[202]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[202]), .B(A[202]), .Z(n284) );
  XOR U427 ( .A(A[201]), .B(n285), .Z(O[201]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[201]), .B(A[201]), .Z(n286) );
  XOR U430 ( .A(A[200]), .B(n287), .Z(O[200]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[200]), .B(A[200]), .Z(n288) );
  XOR U433 ( .A(A[1]), .B(n289), .Z(O[1]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[1]), .B(A[1]), .Z(n290) );
  XOR U436 ( .A(A[19]), .B(n291), .Z(O[19]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[19]), .B(A[19]), .Z(n292) );
  XOR U439 ( .A(A[199]), .B(n293), .Z(O[199]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[199]), .B(A[199]), .Z(n294) );
  XOR U442 ( .A(A[198]), .B(n295), .Z(O[198]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[198]), .B(A[198]), .Z(n296) );
  XOR U445 ( .A(A[197]), .B(n297), .Z(O[197]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[197]), .B(A[197]), .Z(n298) );
  XOR U448 ( .A(A[196]), .B(n299), .Z(O[196]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[196]), .B(A[196]), .Z(n300) );
  XOR U451 ( .A(A[195]), .B(n301), .Z(O[195]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[195]), .B(A[195]), .Z(n302) );
  XOR U454 ( .A(A[194]), .B(n303), .Z(O[194]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[194]), .B(A[194]), .Z(n304) );
  XOR U457 ( .A(A[193]), .B(n305), .Z(O[193]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[193]), .B(A[193]), .Z(n306) );
  XOR U460 ( .A(A[192]), .B(n307), .Z(O[192]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[192]), .B(A[192]), .Z(n308) );
  XOR U463 ( .A(A[191]), .B(n309), .Z(O[191]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[191]), .B(A[191]), .Z(n310) );
  XOR U466 ( .A(A[190]), .B(n311), .Z(O[190]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[190]), .B(A[190]), .Z(n312) );
  XOR U469 ( .A(A[18]), .B(n313), .Z(O[18]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[18]), .B(A[18]), .Z(n314) );
  XOR U472 ( .A(A[189]), .B(n315), .Z(O[189]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[189]), .B(A[189]), .Z(n316) );
  XOR U475 ( .A(A[188]), .B(n317), .Z(O[188]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[188]), .B(A[188]), .Z(n318) );
  XOR U478 ( .A(A[187]), .B(n319), .Z(O[187]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[187]), .B(A[187]), .Z(n320) );
  XOR U481 ( .A(A[186]), .B(n321), .Z(O[186]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[186]), .B(A[186]), .Z(n322) );
  XOR U484 ( .A(A[185]), .B(n323), .Z(O[185]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[185]), .B(A[185]), .Z(n324) );
  XOR U487 ( .A(A[184]), .B(n325), .Z(O[184]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[184]), .B(A[184]), .Z(n326) );
  XOR U490 ( .A(A[183]), .B(n327), .Z(O[183]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[183]), .B(A[183]), .Z(n328) );
  XOR U493 ( .A(A[182]), .B(n329), .Z(O[182]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[182]), .B(A[182]), .Z(n330) );
  XOR U496 ( .A(A[181]), .B(n331), .Z(O[181]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[181]), .B(A[181]), .Z(n332) );
  XOR U499 ( .A(A[180]), .B(n333), .Z(O[180]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[180]), .B(A[180]), .Z(n334) );
  XOR U502 ( .A(A[17]), .B(n335), .Z(O[17]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[17]), .B(A[17]), .Z(n336) );
  XOR U505 ( .A(A[179]), .B(n337), .Z(O[179]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[179]), .B(A[179]), .Z(n338) );
  XOR U508 ( .A(A[178]), .B(n339), .Z(O[178]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[178]), .B(A[178]), .Z(n340) );
  XOR U511 ( .A(A[177]), .B(n341), .Z(O[177]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[177]), .B(A[177]), .Z(n342) );
  XOR U514 ( .A(A[176]), .B(n343), .Z(O[176]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[176]), .B(A[176]), .Z(n344) );
  XOR U517 ( .A(A[175]), .B(n345), .Z(O[175]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[175]), .B(A[175]), .Z(n346) );
  XOR U520 ( .A(A[174]), .B(n347), .Z(O[174]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[174]), .B(A[174]), .Z(n348) );
  XOR U523 ( .A(A[173]), .B(n349), .Z(O[173]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[173]), .B(A[173]), .Z(n350) );
  XOR U526 ( .A(A[172]), .B(n351), .Z(O[172]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[172]), .B(A[172]), .Z(n352) );
  XOR U529 ( .A(A[171]), .B(n353), .Z(O[171]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[171]), .B(A[171]), .Z(n354) );
  XOR U532 ( .A(A[170]), .B(n355), .Z(O[170]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[170]), .B(A[170]), .Z(n356) );
  XOR U535 ( .A(A[16]), .B(n357), .Z(O[16]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[16]), .B(A[16]), .Z(n358) );
  XOR U538 ( .A(A[169]), .B(n359), .Z(O[169]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[169]), .B(A[169]), .Z(n360) );
  XOR U541 ( .A(A[168]), .B(n361), .Z(O[168]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[168]), .B(A[168]), .Z(n362) );
  XOR U544 ( .A(A[167]), .B(n363), .Z(O[167]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[167]), .B(A[167]), .Z(n364) );
  XOR U547 ( .A(A[166]), .B(n365), .Z(O[166]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[166]), .B(A[166]), .Z(n366) );
  XOR U550 ( .A(A[165]), .B(n367), .Z(O[165]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[165]), .B(A[165]), .Z(n368) );
  XOR U553 ( .A(A[164]), .B(n369), .Z(O[164]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[164]), .B(A[164]), .Z(n370) );
  XOR U556 ( .A(A[163]), .B(n371), .Z(O[163]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[163]), .B(A[163]), .Z(n372) );
  XOR U559 ( .A(A[162]), .B(n373), .Z(O[162]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[162]), .B(A[162]), .Z(n374) );
  XOR U562 ( .A(A[161]), .B(n375), .Z(O[161]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[161]), .B(A[161]), .Z(n376) );
  XOR U565 ( .A(A[160]), .B(n377), .Z(O[160]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[160]), .B(A[160]), .Z(n378) );
  XOR U568 ( .A(A[15]), .B(n379), .Z(O[15]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[15]), .B(A[15]), .Z(n380) );
  XOR U571 ( .A(A[159]), .B(n381), .Z(O[159]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[159]), .B(A[159]), .Z(n382) );
  XOR U574 ( .A(A[158]), .B(n383), .Z(O[158]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[158]), .B(A[158]), .Z(n384) );
  XOR U577 ( .A(A[157]), .B(n385), .Z(O[157]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[157]), .B(A[157]), .Z(n386) );
  XOR U580 ( .A(A[156]), .B(n387), .Z(O[156]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[156]), .B(A[156]), .Z(n388) );
  XOR U583 ( .A(A[155]), .B(n389), .Z(O[155]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[155]), .B(A[155]), .Z(n390) );
  XOR U586 ( .A(A[154]), .B(n391), .Z(O[154]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[154]), .B(A[154]), .Z(n392) );
  XOR U589 ( .A(A[153]), .B(n393), .Z(O[153]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[153]), .B(A[153]), .Z(n394) );
  XOR U592 ( .A(A[152]), .B(n395), .Z(O[152]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[152]), .B(A[152]), .Z(n396) );
  XOR U595 ( .A(A[151]), .B(n397), .Z(O[151]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[151]), .B(A[151]), .Z(n398) );
  XOR U598 ( .A(A[150]), .B(n399), .Z(O[150]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[150]), .B(A[150]), .Z(n400) );
  XOR U601 ( .A(A[14]), .B(n401), .Z(O[14]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[14]), .B(A[14]), .Z(n402) );
  XOR U604 ( .A(A[149]), .B(n403), .Z(O[149]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[149]), .B(A[149]), .Z(n404) );
  XOR U607 ( .A(A[148]), .B(n405), .Z(O[148]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[148]), .B(A[148]), .Z(n406) );
  XOR U610 ( .A(A[147]), .B(n407), .Z(O[147]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[147]), .B(A[147]), .Z(n408) );
  XOR U613 ( .A(A[146]), .B(n409), .Z(O[146]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[146]), .B(A[146]), .Z(n410) );
  XOR U616 ( .A(A[145]), .B(n411), .Z(O[145]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[145]), .B(A[145]), .Z(n412) );
  XOR U619 ( .A(A[144]), .B(n413), .Z(O[144]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[144]), .B(A[144]), .Z(n414) );
  XOR U622 ( .A(A[143]), .B(n415), .Z(O[143]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[143]), .B(A[143]), .Z(n416) );
  XOR U625 ( .A(A[142]), .B(n417), .Z(O[142]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[142]), .B(A[142]), .Z(n418) );
  XOR U628 ( .A(A[141]), .B(n419), .Z(O[141]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[141]), .B(A[141]), .Z(n420) );
  XOR U631 ( .A(A[140]), .B(n421), .Z(O[140]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[140]), .B(A[140]), .Z(n422) );
  XOR U634 ( .A(A[13]), .B(n423), .Z(O[13]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[13]), .B(A[13]), .Z(n424) );
  XOR U637 ( .A(A[139]), .B(n425), .Z(O[139]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[139]), .B(A[139]), .Z(n426) );
  XOR U640 ( .A(A[138]), .B(n427), .Z(O[138]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[138]), .B(A[138]), .Z(n428) );
  XOR U643 ( .A(A[137]), .B(n429), .Z(O[137]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[137]), .B(A[137]), .Z(n430) );
  XOR U646 ( .A(A[136]), .B(n431), .Z(O[136]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[136]), .B(A[136]), .Z(n432) );
  XOR U649 ( .A(A[135]), .B(n433), .Z(O[135]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[135]), .B(A[135]), .Z(n434) );
  XOR U652 ( .A(A[134]), .B(n435), .Z(O[134]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[134]), .B(A[134]), .Z(n436) );
  XOR U655 ( .A(A[133]), .B(n437), .Z(O[133]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[133]), .B(A[133]), .Z(n438) );
  XOR U658 ( .A(A[132]), .B(n439), .Z(O[132]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[132]), .B(A[132]), .Z(n440) );
  XOR U661 ( .A(A[131]), .B(n441), .Z(O[131]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[131]), .B(A[131]), .Z(n442) );
  XOR U664 ( .A(A[130]), .B(n443), .Z(O[130]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[130]), .B(A[130]), .Z(n444) );
  XOR U667 ( .A(A[12]), .B(n445), .Z(O[12]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[12]), .B(A[12]), .Z(n446) );
  XOR U670 ( .A(A[129]), .B(n447), .Z(O[129]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[129]), .B(A[129]), .Z(n448) );
  XOR U673 ( .A(A[128]), .B(n449), .Z(O[128]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[128]), .B(A[128]), .Z(n450) );
  XOR U676 ( .A(A[127]), .B(n451), .Z(O[127]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[127]), .B(A[127]), .Z(n452) );
  XOR U679 ( .A(A[126]), .B(n453), .Z(O[126]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[126]), .B(A[126]), .Z(n454) );
  XOR U682 ( .A(A[125]), .B(n455), .Z(O[125]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[125]), .B(A[125]), .Z(n456) );
  XOR U685 ( .A(A[124]), .B(n457), .Z(O[124]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[124]), .B(A[124]), .Z(n458) );
  XOR U688 ( .A(A[123]), .B(n459), .Z(O[123]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[123]), .B(A[123]), .Z(n460) );
  XOR U691 ( .A(A[122]), .B(n461), .Z(O[122]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[122]), .B(A[122]), .Z(n462) );
  XOR U694 ( .A(A[121]), .B(n463), .Z(O[121]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[121]), .B(A[121]), .Z(n464) );
  XOR U697 ( .A(A[120]), .B(n465), .Z(O[120]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[120]), .B(A[120]), .Z(n466) );
  XOR U700 ( .A(A[11]), .B(n467), .Z(O[11]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[11]), .B(A[11]), .Z(n468) );
  XOR U703 ( .A(A[119]), .B(n469), .Z(O[119]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[119]), .B(A[119]), .Z(n470) );
  XOR U706 ( .A(A[118]), .B(n471), .Z(O[118]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[118]), .B(A[118]), .Z(n472) );
  XOR U709 ( .A(A[117]), .B(n473), .Z(O[117]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[117]), .B(A[117]), .Z(n474) );
  XOR U712 ( .A(A[116]), .B(n475), .Z(O[116]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[116]), .B(A[116]), .Z(n476) );
  XOR U715 ( .A(A[115]), .B(n477), .Z(O[115]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[115]), .B(A[115]), .Z(n478) );
  XOR U718 ( .A(A[114]), .B(n479), .Z(O[114]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[114]), .B(A[114]), .Z(n480) );
  XOR U721 ( .A(A[113]), .B(n481), .Z(O[113]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[113]), .B(A[113]), .Z(n482) );
  XOR U724 ( .A(A[112]), .B(n483), .Z(O[112]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[112]), .B(A[112]), .Z(n484) );
  XOR U727 ( .A(A[111]), .B(n485), .Z(O[111]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[111]), .B(A[111]), .Z(n486) );
  XOR U730 ( .A(A[110]), .B(n487), .Z(O[110]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[110]), .B(A[110]), .Z(n488) );
  XOR U733 ( .A(A[10]), .B(n489), .Z(O[10]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[10]), .B(A[10]), .Z(n490) );
  XOR U736 ( .A(A[109]), .B(n491), .Z(O[109]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[109]), .B(A[109]), .Z(n492) );
  XOR U739 ( .A(A[108]), .B(n493), .Z(O[108]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[108]), .B(A[108]), .Z(n494) );
  XOR U742 ( .A(A[107]), .B(n495), .Z(O[107]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[107]), .B(A[107]), .Z(n496) );
  XOR U745 ( .A(A[106]), .B(n497), .Z(O[106]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[106]), .B(A[106]), .Z(n498) );
  XOR U748 ( .A(A[105]), .B(n499), .Z(O[105]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[105]), .B(A[105]), .Z(n500) );
  XOR U751 ( .A(A[104]), .B(n501), .Z(O[104]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[104]), .B(A[104]), .Z(n502) );
  XOR U754 ( .A(A[103]), .B(n503), .Z(O[103]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[103]), .B(A[103]), .Z(n504) );
  XOR U757 ( .A(A[102]), .B(n505), .Z(O[102]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[102]), .B(A[102]), .Z(n506) );
  XOR U760 ( .A(A[101]), .B(n507), .Z(O[101]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[101]), .B(A[101]), .Z(n508) );
  XOR U763 ( .A(A[100]), .B(n509), .Z(O[100]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[100]), .B(A[100]), .Z(n510) );
  XOR U766 ( .A(A[0]), .B(n511), .Z(O[0]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[0]), .B(A[0]), .Z(n512) );
endmodule


module MUX_N256_2 ( A, B, S, O );
  input [255:0] A;
  input [255:0] B;
  output [255:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510;

  XOR U1 ( .A(B[8]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(B[8]), .Z(n2) );
  XOR U4 ( .A(B[98]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(B[98]), .Z(n4) );
  XOR U7 ( .A(B[97]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(B[97]), .Z(n6) );
  XOR U10 ( .A(B[96]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(B[96]), .Z(n8) );
  XOR U13 ( .A(B[95]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(B[95]), .Z(n10) );
  XOR U16 ( .A(B[94]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(B[94]), .Z(n12) );
  XOR U19 ( .A(B[93]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(B[93]), .Z(n14) );
  XOR U22 ( .A(B[92]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(B[92]), .Z(n16) );
  XOR U25 ( .A(B[91]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(B[91]), .Z(n18) );
  XOR U28 ( .A(B[90]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(B[90]), .Z(n20) );
  XOR U31 ( .A(B[89]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(B[89]), .Z(n22) );
  XOR U34 ( .A(B[7]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(B[7]), .Z(n24) );
  XOR U37 ( .A(B[88]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(B[88]), .Z(n26) );
  XOR U40 ( .A(B[87]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(B[87]), .Z(n28) );
  XOR U43 ( .A(B[86]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(B[86]), .Z(n30) );
  XOR U46 ( .A(B[85]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(B[85]), .Z(n32) );
  XOR U49 ( .A(B[84]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(B[84]), .Z(n34) );
  XOR U52 ( .A(B[83]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(B[83]), .Z(n36) );
  XOR U55 ( .A(B[82]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(B[82]), .Z(n38) );
  XOR U58 ( .A(B[81]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(B[81]), .Z(n40) );
  XOR U61 ( .A(B[80]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(B[80]), .Z(n42) );
  XOR U64 ( .A(B[79]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(B[79]), .Z(n44) );
  XOR U67 ( .A(B[6]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(B[6]), .Z(n46) );
  XOR U70 ( .A(B[78]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(B[78]), .Z(n48) );
  XOR U73 ( .A(B[77]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(B[77]), .Z(n50) );
  XOR U76 ( .A(B[76]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(B[76]), .Z(n52) );
  XOR U79 ( .A(B[75]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(B[75]), .Z(n54) );
  XOR U82 ( .A(B[74]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(B[74]), .Z(n56) );
  XOR U85 ( .A(B[73]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(B[73]), .Z(n58) );
  XOR U88 ( .A(B[72]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(B[72]), .Z(n60) );
  XOR U91 ( .A(B[71]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(B[71]), .Z(n62) );
  XOR U94 ( .A(B[70]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(B[70]), .Z(n64) );
  XOR U97 ( .A(B[69]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(B[69]), .Z(n66) );
  XOR U100 ( .A(B[5]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(B[5]), .Z(n68) );
  XOR U103 ( .A(B[68]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(B[68]), .Z(n70) );
  XOR U106 ( .A(B[67]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(B[67]), .Z(n72) );
  XOR U109 ( .A(B[66]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(B[66]), .Z(n74) );
  XOR U112 ( .A(B[65]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(B[65]), .Z(n76) );
  XOR U115 ( .A(B[64]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(B[64]), .Z(n78) );
  XOR U118 ( .A(B[63]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(B[63]), .Z(n80) );
  XOR U121 ( .A(B[62]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(B[62]), .Z(n82) );
  XOR U124 ( .A(B[61]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(B[61]), .Z(n84) );
  XOR U127 ( .A(B[60]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(B[60]), .Z(n86) );
  XOR U130 ( .A(B[59]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(B[59]), .Z(n88) );
  XOR U133 ( .A(B[4]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(B[4]), .Z(n90) );
  XOR U136 ( .A(B[58]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(B[58]), .Z(n92) );
  XOR U139 ( .A(B[57]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(B[57]), .Z(n94) );
  XOR U142 ( .A(B[56]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(B[56]), .Z(n96) );
  XOR U145 ( .A(B[55]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(B[55]), .Z(n98) );
  XOR U148 ( .A(B[54]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(B[54]), .Z(n100) );
  XOR U151 ( .A(B[53]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(B[53]), .Z(n102) );
  XOR U154 ( .A(B[52]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(B[52]), .Z(n104) );
  XOR U157 ( .A(B[51]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(B[51]), .Z(n106) );
  XOR U160 ( .A(B[50]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(B[50]), .Z(n108) );
  XOR U163 ( .A(B[49]), .B(n109), .Z(O[50]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[50]), .B(B[49]), .Z(n110) );
  XOR U166 ( .A(B[3]), .B(n111), .Z(O[4]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[4]), .B(B[3]), .Z(n112) );
  XOR U169 ( .A(B[48]), .B(n113), .Z(O[49]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[49]), .B(B[48]), .Z(n114) );
  XOR U172 ( .A(B[47]), .B(n115), .Z(O[48]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[48]), .B(B[47]), .Z(n116) );
  XOR U175 ( .A(B[46]), .B(n117), .Z(O[47]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[47]), .B(B[46]), .Z(n118) );
  XOR U178 ( .A(B[45]), .B(n119), .Z(O[46]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[46]), .B(B[45]), .Z(n120) );
  XOR U181 ( .A(B[44]), .B(n121), .Z(O[45]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[45]), .B(B[44]), .Z(n122) );
  XOR U184 ( .A(B[43]), .B(n123), .Z(O[44]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[44]), .B(B[43]), .Z(n124) );
  XOR U187 ( .A(B[42]), .B(n125), .Z(O[43]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[43]), .B(B[42]), .Z(n126) );
  XOR U190 ( .A(B[41]), .B(n127), .Z(O[42]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[42]), .B(B[41]), .Z(n128) );
  XOR U193 ( .A(B[40]), .B(n129), .Z(O[41]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[41]), .B(B[40]), .Z(n130) );
  XOR U196 ( .A(B[39]), .B(n131), .Z(O[40]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[40]), .B(B[39]), .Z(n132) );
  XOR U199 ( .A(B[2]), .B(n133), .Z(O[3]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[3]), .B(B[2]), .Z(n134) );
  XOR U202 ( .A(B[38]), .B(n135), .Z(O[39]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[39]), .B(B[38]), .Z(n136) );
  XOR U205 ( .A(B[37]), .B(n137), .Z(O[38]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[38]), .B(B[37]), .Z(n138) );
  XOR U208 ( .A(B[36]), .B(n139), .Z(O[37]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[37]), .B(B[36]), .Z(n140) );
  XOR U211 ( .A(B[35]), .B(n141), .Z(O[36]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[36]), .B(B[35]), .Z(n142) );
  XOR U214 ( .A(B[34]), .B(n143), .Z(O[35]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[35]), .B(B[34]), .Z(n144) );
  XOR U217 ( .A(B[33]), .B(n145), .Z(O[34]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[34]), .B(B[33]), .Z(n146) );
  XOR U220 ( .A(B[32]), .B(n147), .Z(O[33]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[33]), .B(B[32]), .Z(n148) );
  XOR U223 ( .A(B[31]), .B(n149), .Z(O[32]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[32]), .B(B[31]), .Z(n150) );
  XOR U226 ( .A(B[30]), .B(n151), .Z(O[31]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[31]), .B(B[30]), .Z(n152) );
  XOR U229 ( .A(B[29]), .B(n153), .Z(O[30]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[30]), .B(B[29]), .Z(n154) );
  XOR U232 ( .A(B[1]), .B(n155), .Z(O[2]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[2]), .B(B[1]), .Z(n156) );
  XOR U235 ( .A(B[28]), .B(n157), .Z(O[29]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[29]), .B(B[28]), .Z(n158) );
  XOR U238 ( .A(B[27]), .B(n159), .Z(O[28]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[28]), .B(B[27]), .Z(n160) );
  XOR U241 ( .A(B[26]), .B(n161), .Z(O[27]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[27]), .B(B[26]), .Z(n162) );
  XOR U244 ( .A(B[25]), .B(n163), .Z(O[26]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[26]), .B(B[25]), .Z(n164) );
  XOR U247 ( .A(B[24]), .B(n165), .Z(O[25]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[25]), .B(B[24]), .Z(n166) );
  XOR U250 ( .A(B[254]), .B(n167), .Z(O[255]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[255]), .B(B[254]), .Z(n168) );
  XOR U253 ( .A(B[253]), .B(n169), .Z(O[254]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[254]), .B(B[253]), .Z(n170) );
  XOR U256 ( .A(B[252]), .B(n171), .Z(O[253]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[253]), .B(B[252]), .Z(n172) );
  XOR U259 ( .A(B[251]), .B(n173), .Z(O[252]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[252]), .B(B[251]), .Z(n174) );
  XOR U262 ( .A(B[250]), .B(n175), .Z(O[251]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[251]), .B(B[250]), .Z(n176) );
  XOR U265 ( .A(B[249]), .B(n177), .Z(O[250]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[250]), .B(B[249]), .Z(n178) );
  XOR U268 ( .A(B[23]), .B(n179), .Z(O[24]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[24]), .B(B[23]), .Z(n180) );
  XOR U271 ( .A(B[248]), .B(n181), .Z(O[249]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[249]), .B(B[248]), .Z(n182) );
  XOR U274 ( .A(B[247]), .B(n183), .Z(O[248]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[248]), .B(B[247]), .Z(n184) );
  XOR U277 ( .A(B[246]), .B(n185), .Z(O[247]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[247]), .B(B[246]), .Z(n186) );
  XOR U280 ( .A(B[245]), .B(n187), .Z(O[246]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[246]), .B(B[245]), .Z(n188) );
  XOR U283 ( .A(B[244]), .B(n189), .Z(O[245]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[245]), .B(B[244]), .Z(n190) );
  XOR U286 ( .A(B[243]), .B(n191), .Z(O[244]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[244]), .B(B[243]), .Z(n192) );
  XOR U289 ( .A(B[242]), .B(n193), .Z(O[243]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[243]), .B(B[242]), .Z(n194) );
  XOR U292 ( .A(B[241]), .B(n195), .Z(O[242]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[242]), .B(B[241]), .Z(n196) );
  XOR U295 ( .A(B[240]), .B(n197), .Z(O[241]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[241]), .B(B[240]), .Z(n198) );
  XOR U298 ( .A(B[239]), .B(n199), .Z(O[240]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[240]), .B(B[239]), .Z(n200) );
  XOR U301 ( .A(B[22]), .B(n201), .Z(O[23]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[23]), .B(B[22]), .Z(n202) );
  XOR U304 ( .A(B[238]), .B(n203), .Z(O[239]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[239]), .B(B[238]), .Z(n204) );
  XOR U307 ( .A(B[237]), .B(n205), .Z(O[238]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[238]), .B(B[237]), .Z(n206) );
  XOR U310 ( .A(B[236]), .B(n207), .Z(O[237]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[237]), .B(B[236]), .Z(n208) );
  XOR U313 ( .A(B[235]), .B(n209), .Z(O[236]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[236]), .B(B[235]), .Z(n210) );
  XOR U316 ( .A(B[234]), .B(n211), .Z(O[235]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[235]), .B(B[234]), .Z(n212) );
  XOR U319 ( .A(B[233]), .B(n213), .Z(O[234]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[234]), .B(B[233]), .Z(n214) );
  XOR U322 ( .A(B[232]), .B(n215), .Z(O[233]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[233]), .B(B[232]), .Z(n216) );
  XOR U325 ( .A(B[231]), .B(n217), .Z(O[232]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[232]), .B(B[231]), .Z(n218) );
  XOR U328 ( .A(B[230]), .B(n219), .Z(O[231]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[231]), .B(B[230]), .Z(n220) );
  XOR U331 ( .A(B[229]), .B(n221), .Z(O[230]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[230]), .B(B[229]), .Z(n222) );
  XOR U334 ( .A(B[21]), .B(n223), .Z(O[22]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[22]), .B(B[21]), .Z(n224) );
  XOR U337 ( .A(B[228]), .B(n225), .Z(O[229]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[229]), .B(B[228]), .Z(n226) );
  XOR U340 ( .A(B[227]), .B(n227), .Z(O[228]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[228]), .B(B[227]), .Z(n228) );
  XOR U343 ( .A(B[226]), .B(n229), .Z(O[227]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[227]), .B(B[226]), .Z(n230) );
  XOR U346 ( .A(B[225]), .B(n231), .Z(O[226]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[226]), .B(B[225]), .Z(n232) );
  XOR U349 ( .A(B[224]), .B(n233), .Z(O[225]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[225]), .B(B[224]), .Z(n234) );
  XOR U352 ( .A(B[223]), .B(n235), .Z(O[224]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[224]), .B(B[223]), .Z(n236) );
  XOR U355 ( .A(B[222]), .B(n237), .Z(O[223]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[223]), .B(B[222]), .Z(n238) );
  XOR U358 ( .A(B[221]), .B(n239), .Z(O[222]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[222]), .B(B[221]), .Z(n240) );
  XOR U361 ( .A(B[220]), .B(n241), .Z(O[221]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[221]), .B(B[220]), .Z(n242) );
  XOR U364 ( .A(B[219]), .B(n243), .Z(O[220]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[220]), .B(B[219]), .Z(n244) );
  XOR U367 ( .A(B[20]), .B(n245), .Z(O[21]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[21]), .B(B[20]), .Z(n246) );
  XOR U370 ( .A(B[218]), .B(n247), .Z(O[219]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[219]), .B(B[218]), .Z(n248) );
  XOR U373 ( .A(B[217]), .B(n249), .Z(O[218]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[218]), .B(B[217]), .Z(n250) );
  XOR U376 ( .A(B[216]), .B(n251), .Z(O[217]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[217]), .B(B[216]), .Z(n252) );
  XOR U379 ( .A(B[215]), .B(n253), .Z(O[216]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[216]), .B(B[215]), .Z(n254) );
  XOR U382 ( .A(B[214]), .B(n255), .Z(O[215]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[215]), .B(B[214]), .Z(n256) );
  XOR U385 ( .A(B[213]), .B(n257), .Z(O[214]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[214]), .B(B[213]), .Z(n258) );
  XOR U388 ( .A(B[212]), .B(n259), .Z(O[213]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[213]), .B(B[212]), .Z(n260) );
  XOR U391 ( .A(B[211]), .B(n261), .Z(O[212]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[212]), .B(B[211]), .Z(n262) );
  XOR U394 ( .A(B[210]), .B(n263), .Z(O[211]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[211]), .B(B[210]), .Z(n264) );
  XOR U397 ( .A(B[209]), .B(n265), .Z(O[210]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[210]), .B(B[209]), .Z(n266) );
  XOR U400 ( .A(B[19]), .B(n267), .Z(O[20]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[20]), .B(B[19]), .Z(n268) );
  XOR U403 ( .A(B[208]), .B(n269), .Z(O[209]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[209]), .B(B[208]), .Z(n270) );
  XOR U406 ( .A(B[207]), .B(n271), .Z(O[208]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[208]), .B(B[207]), .Z(n272) );
  XOR U409 ( .A(B[206]), .B(n273), .Z(O[207]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[207]), .B(B[206]), .Z(n274) );
  XOR U412 ( .A(B[205]), .B(n275), .Z(O[206]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[206]), .B(B[205]), .Z(n276) );
  XOR U415 ( .A(B[204]), .B(n277), .Z(O[205]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[205]), .B(B[204]), .Z(n278) );
  XOR U418 ( .A(B[203]), .B(n279), .Z(O[204]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[204]), .B(B[203]), .Z(n280) );
  XOR U421 ( .A(B[202]), .B(n281), .Z(O[203]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[203]), .B(B[202]), .Z(n282) );
  XOR U424 ( .A(B[201]), .B(n283), .Z(O[202]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[202]), .B(B[201]), .Z(n284) );
  XOR U427 ( .A(B[200]), .B(n285), .Z(O[201]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[201]), .B(B[200]), .Z(n286) );
  XOR U430 ( .A(B[199]), .B(n287), .Z(O[200]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[200]), .B(B[199]), .Z(n288) );
  XOR U433 ( .A(B[0]), .B(n289), .Z(O[1]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[1]), .B(B[0]), .Z(n290) );
  XOR U436 ( .A(B[18]), .B(n291), .Z(O[19]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[19]), .B(B[18]), .Z(n292) );
  XOR U439 ( .A(B[198]), .B(n293), .Z(O[199]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[199]), .B(B[198]), .Z(n294) );
  XOR U442 ( .A(B[197]), .B(n295), .Z(O[198]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[198]), .B(B[197]), .Z(n296) );
  XOR U445 ( .A(B[196]), .B(n297), .Z(O[197]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[197]), .B(B[196]), .Z(n298) );
  XOR U448 ( .A(B[195]), .B(n299), .Z(O[196]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[196]), .B(B[195]), .Z(n300) );
  XOR U451 ( .A(B[194]), .B(n301), .Z(O[195]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[195]), .B(B[194]), .Z(n302) );
  XOR U454 ( .A(B[193]), .B(n303), .Z(O[194]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[194]), .B(B[193]), .Z(n304) );
  XOR U457 ( .A(B[192]), .B(n305), .Z(O[193]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[193]), .B(B[192]), .Z(n306) );
  XOR U460 ( .A(B[191]), .B(n307), .Z(O[192]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[192]), .B(B[191]), .Z(n308) );
  XOR U463 ( .A(B[190]), .B(n309), .Z(O[191]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[191]), .B(B[190]), .Z(n310) );
  XOR U466 ( .A(B[189]), .B(n311), .Z(O[190]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[190]), .B(B[189]), .Z(n312) );
  XOR U469 ( .A(B[17]), .B(n313), .Z(O[18]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[18]), .B(B[17]), .Z(n314) );
  XOR U472 ( .A(B[188]), .B(n315), .Z(O[189]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[189]), .B(B[188]), .Z(n316) );
  XOR U475 ( .A(B[187]), .B(n317), .Z(O[188]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[188]), .B(B[187]), .Z(n318) );
  XOR U478 ( .A(B[186]), .B(n319), .Z(O[187]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[187]), .B(B[186]), .Z(n320) );
  XOR U481 ( .A(B[185]), .B(n321), .Z(O[186]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[186]), .B(B[185]), .Z(n322) );
  XOR U484 ( .A(B[184]), .B(n323), .Z(O[185]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[185]), .B(B[184]), .Z(n324) );
  XOR U487 ( .A(B[183]), .B(n325), .Z(O[184]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[184]), .B(B[183]), .Z(n326) );
  XOR U490 ( .A(B[182]), .B(n327), .Z(O[183]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[183]), .B(B[182]), .Z(n328) );
  XOR U493 ( .A(B[181]), .B(n329), .Z(O[182]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[182]), .B(B[181]), .Z(n330) );
  XOR U496 ( .A(B[180]), .B(n331), .Z(O[181]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[181]), .B(B[180]), .Z(n332) );
  XOR U499 ( .A(B[179]), .B(n333), .Z(O[180]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[180]), .B(B[179]), .Z(n334) );
  XOR U502 ( .A(B[16]), .B(n335), .Z(O[17]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[17]), .B(B[16]), .Z(n336) );
  XOR U505 ( .A(B[178]), .B(n337), .Z(O[179]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[179]), .B(B[178]), .Z(n338) );
  XOR U508 ( .A(B[177]), .B(n339), .Z(O[178]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[178]), .B(B[177]), .Z(n340) );
  XOR U511 ( .A(B[176]), .B(n341), .Z(O[177]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[177]), .B(B[176]), .Z(n342) );
  XOR U514 ( .A(B[175]), .B(n343), .Z(O[176]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[176]), .B(B[175]), .Z(n344) );
  XOR U517 ( .A(B[174]), .B(n345), .Z(O[175]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[175]), .B(B[174]), .Z(n346) );
  XOR U520 ( .A(B[173]), .B(n347), .Z(O[174]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[174]), .B(B[173]), .Z(n348) );
  XOR U523 ( .A(B[172]), .B(n349), .Z(O[173]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[173]), .B(B[172]), .Z(n350) );
  XOR U526 ( .A(B[171]), .B(n351), .Z(O[172]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[172]), .B(B[171]), .Z(n352) );
  XOR U529 ( .A(B[170]), .B(n353), .Z(O[171]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[171]), .B(B[170]), .Z(n354) );
  XOR U532 ( .A(B[169]), .B(n355), .Z(O[170]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[170]), .B(B[169]), .Z(n356) );
  XOR U535 ( .A(B[15]), .B(n357), .Z(O[16]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[16]), .B(B[15]), .Z(n358) );
  XOR U538 ( .A(B[168]), .B(n359), .Z(O[169]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[169]), .B(B[168]), .Z(n360) );
  XOR U541 ( .A(B[167]), .B(n361), .Z(O[168]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[168]), .B(B[167]), .Z(n362) );
  XOR U544 ( .A(B[166]), .B(n363), .Z(O[167]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[167]), .B(B[166]), .Z(n364) );
  XOR U547 ( .A(B[165]), .B(n365), .Z(O[166]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[166]), .B(B[165]), .Z(n366) );
  XOR U550 ( .A(B[164]), .B(n367), .Z(O[165]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[165]), .B(B[164]), .Z(n368) );
  XOR U553 ( .A(B[163]), .B(n369), .Z(O[164]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[164]), .B(B[163]), .Z(n370) );
  XOR U556 ( .A(B[162]), .B(n371), .Z(O[163]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[163]), .B(B[162]), .Z(n372) );
  XOR U559 ( .A(B[161]), .B(n373), .Z(O[162]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[162]), .B(B[161]), .Z(n374) );
  XOR U562 ( .A(B[160]), .B(n375), .Z(O[161]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[161]), .B(B[160]), .Z(n376) );
  XOR U565 ( .A(B[159]), .B(n377), .Z(O[160]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[160]), .B(B[159]), .Z(n378) );
  XOR U568 ( .A(B[14]), .B(n379), .Z(O[15]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[15]), .B(B[14]), .Z(n380) );
  XOR U571 ( .A(B[158]), .B(n381), .Z(O[159]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[159]), .B(B[158]), .Z(n382) );
  XOR U574 ( .A(B[157]), .B(n383), .Z(O[158]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[158]), .B(B[157]), .Z(n384) );
  XOR U577 ( .A(B[156]), .B(n385), .Z(O[157]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[157]), .B(B[156]), .Z(n386) );
  XOR U580 ( .A(B[155]), .B(n387), .Z(O[156]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[156]), .B(B[155]), .Z(n388) );
  XOR U583 ( .A(B[154]), .B(n389), .Z(O[155]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[155]), .B(B[154]), .Z(n390) );
  XOR U586 ( .A(B[153]), .B(n391), .Z(O[154]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[154]), .B(B[153]), .Z(n392) );
  XOR U589 ( .A(B[152]), .B(n393), .Z(O[153]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[153]), .B(B[152]), .Z(n394) );
  XOR U592 ( .A(B[151]), .B(n395), .Z(O[152]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[152]), .B(B[151]), .Z(n396) );
  XOR U595 ( .A(B[150]), .B(n397), .Z(O[151]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[151]), .B(B[150]), .Z(n398) );
  XOR U598 ( .A(B[149]), .B(n399), .Z(O[150]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[150]), .B(B[149]), .Z(n400) );
  XOR U601 ( .A(B[13]), .B(n401), .Z(O[14]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[14]), .B(B[13]), .Z(n402) );
  XOR U604 ( .A(B[148]), .B(n403), .Z(O[149]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[149]), .B(B[148]), .Z(n404) );
  XOR U607 ( .A(B[147]), .B(n405), .Z(O[148]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[148]), .B(B[147]), .Z(n406) );
  XOR U610 ( .A(B[146]), .B(n407), .Z(O[147]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[147]), .B(B[146]), .Z(n408) );
  XOR U613 ( .A(B[145]), .B(n409), .Z(O[146]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[146]), .B(B[145]), .Z(n410) );
  XOR U616 ( .A(B[144]), .B(n411), .Z(O[145]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[145]), .B(B[144]), .Z(n412) );
  XOR U619 ( .A(B[143]), .B(n413), .Z(O[144]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[144]), .B(B[143]), .Z(n414) );
  XOR U622 ( .A(B[142]), .B(n415), .Z(O[143]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[143]), .B(B[142]), .Z(n416) );
  XOR U625 ( .A(B[141]), .B(n417), .Z(O[142]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[142]), .B(B[141]), .Z(n418) );
  XOR U628 ( .A(B[140]), .B(n419), .Z(O[141]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[141]), .B(B[140]), .Z(n420) );
  XOR U631 ( .A(B[139]), .B(n421), .Z(O[140]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[140]), .B(B[139]), .Z(n422) );
  XOR U634 ( .A(B[12]), .B(n423), .Z(O[13]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[13]), .B(B[12]), .Z(n424) );
  XOR U637 ( .A(B[138]), .B(n425), .Z(O[139]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[139]), .B(B[138]), .Z(n426) );
  XOR U640 ( .A(B[137]), .B(n427), .Z(O[138]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[138]), .B(B[137]), .Z(n428) );
  XOR U643 ( .A(B[136]), .B(n429), .Z(O[137]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[137]), .B(B[136]), .Z(n430) );
  XOR U646 ( .A(B[135]), .B(n431), .Z(O[136]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[136]), .B(B[135]), .Z(n432) );
  XOR U649 ( .A(B[134]), .B(n433), .Z(O[135]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[135]), .B(B[134]), .Z(n434) );
  XOR U652 ( .A(B[133]), .B(n435), .Z(O[134]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[134]), .B(B[133]), .Z(n436) );
  XOR U655 ( .A(B[132]), .B(n437), .Z(O[133]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[133]), .B(B[132]), .Z(n438) );
  XOR U658 ( .A(B[131]), .B(n439), .Z(O[132]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[132]), .B(B[131]), .Z(n440) );
  XOR U661 ( .A(B[130]), .B(n441), .Z(O[131]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[131]), .B(B[130]), .Z(n442) );
  XOR U664 ( .A(B[129]), .B(n443), .Z(O[130]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[130]), .B(B[129]), .Z(n444) );
  XOR U667 ( .A(B[11]), .B(n445), .Z(O[12]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[12]), .B(B[11]), .Z(n446) );
  XOR U670 ( .A(B[128]), .B(n447), .Z(O[129]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[129]), .B(B[128]), .Z(n448) );
  XOR U673 ( .A(B[127]), .B(n449), .Z(O[128]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[128]), .B(B[127]), .Z(n450) );
  XOR U676 ( .A(B[126]), .B(n451), .Z(O[127]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[127]), .B(B[126]), .Z(n452) );
  XOR U679 ( .A(B[125]), .B(n453), .Z(O[126]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[126]), .B(B[125]), .Z(n454) );
  XOR U682 ( .A(B[124]), .B(n455), .Z(O[125]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[125]), .B(B[124]), .Z(n456) );
  XOR U685 ( .A(B[123]), .B(n457), .Z(O[124]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[124]), .B(B[123]), .Z(n458) );
  XOR U688 ( .A(B[122]), .B(n459), .Z(O[123]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[123]), .B(B[122]), .Z(n460) );
  XOR U691 ( .A(B[121]), .B(n461), .Z(O[122]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[122]), .B(B[121]), .Z(n462) );
  XOR U694 ( .A(B[120]), .B(n463), .Z(O[121]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[121]), .B(B[120]), .Z(n464) );
  XOR U697 ( .A(B[119]), .B(n465), .Z(O[120]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[120]), .B(B[119]), .Z(n466) );
  XOR U700 ( .A(B[10]), .B(n467), .Z(O[11]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[11]), .B(B[10]), .Z(n468) );
  XOR U703 ( .A(B[118]), .B(n469), .Z(O[119]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[119]), .B(B[118]), .Z(n470) );
  XOR U706 ( .A(B[117]), .B(n471), .Z(O[118]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[118]), .B(B[117]), .Z(n472) );
  XOR U709 ( .A(B[116]), .B(n473), .Z(O[117]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[117]), .B(B[116]), .Z(n474) );
  XOR U712 ( .A(B[115]), .B(n475), .Z(O[116]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[116]), .B(B[115]), .Z(n476) );
  XOR U715 ( .A(B[114]), .B(n477), .Z(O[115]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[115]), .B(B[114]), .Z(n478) );
  XOR U718 ( .A(B[113]), .B(n479), .Z(O[114]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[114]), .B(B[113]), .Z(n480) );
  XOR U721 ( .A(B[112]), .B(n481), .Z(O[113]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[113]), .B(B[112]), .Z(n482) );
  XOR U724 ( .A(B[111]), .B(n483), .Z(O[112]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[112]), .B(B[111]), .Z(n484) );
  XOR U727 ( .A(B[110]), .B(n485), .Z(O[111]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[111]), .B(B[110]), .Z(n486) );
  XOR U730 ( .A(B[109]), .B(n487), .Z(O[110]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[110]), .B(B[109]), .Z(n488) );
  XOR U733 ( .A(B[9]), .B(n489), .Z(O[10]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[9]), .B(B[10]), .Z(n490) );
  XOR U736 ( .A(B[108]), .B(n491), .Z(O[109]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[109]), .B(B[108]), .Z(n492) );
  XOR U739 ( .A(B[107]), .B(n493), .Z(O[108]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[108]), .B(B[107]), .Z(n494) );
  XOR U742 ( .A(B[106]), .B(n495), .Z(O[107]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[107]), .B(B[106]), .Z(n496) );
  XOR U745 ( .A(B[105]), .B(n497), .Z(O[106]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[106]), .B(B[105]), .Z(n498) );
  XOR U748 ( .A(B[104]), .B(n499), .Z(O[105]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[105]), .B(B[104]), .Z(n500) );
  XOR U751 ( .A(B[103]), .B(n501), .Z(O[104]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[104]), .B(B[103]), .Z(n502) );
  XOR U754 ( .A(B[102]), .B(n503), .Z(O[103]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[103]), .B(B[102]), .Z(n504) );
  XOR U757 ( .A(B[101]), .B(n505), .Z(O[102]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[102]), .B(B[101]), .Z(n506) );
  XOR U760 ( .A(B[100]), .B(n507), .Z(O[101]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[101]), .B(B[100]), .Z(n508) );
  XOR U763 ( .A(B[99]), .B(n509), .Z(O[100]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[99]), .B(B[100]), .Z(n510) );
  AND U766 ( .A(B[0]), .B(S), .Z(O[0]) );
endmodule


module modexp_2N_NN_N256_CC131072 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   _0_net_, first_one, mul_pow, n6, n8, n265, n266, n267, n268;
  wire   [255:0] start_in;
  wire   [255:0] ein;
  wire   [255:0] creg_next;
  wire   [255:0] o;
  wire   [255:0] ereg_next;
  wire   [255:0] y;

  MUX_N256_0 MUX_4 ( .A(o), .B(c), .S(_0_net_), .O(creg_next) );
  MUX_N256_2 MUX_6 ( .A({ein[254:0], 1'b0}), .B(ein), .S(mul_pow), .O(
        ereg_next) );
  MUX_N256_1 MUX_9 ( .A(m), .B(c), .S(mul_pow), .O(y) );
  modmult_N256_CC256 modmult_1 ( .clk(clk), .rst(1'b0), .start(start_in[0]), 
        .x(c), .y(y), .n(n), .o(o) );
  DFF \start_reg_reg[0]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[255]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e[0]), .Q(
        ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e[1]), .Q(
        ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e[2]), .Q(
        ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e[3]), .Q(
        ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e[4]), .Q(
        ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e[5]), .Q(
        ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e[6]), .Q(
        ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e[7]), .Q(
        ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e[8]), .Q(
        ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e[9]), .Q(
        ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(e[10]), .Q(
        ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(e[11]), .Q(
        ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(e[12]), .Q(
        ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(e[13]), .Q(
        ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(e[14]), .Q(
        ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(e[15]), .Q(
        ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(e[16]), .Q(
        ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(e[17]), .Q(
        ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(e[18]), .Q(
        ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(e[19]), .Q(
        ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(e[20]), .Q(
        ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(e[21]), .Q(
        ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(e[22]), .Q(
        ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(e[23]), .Q(
        ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(e[24]), .Q(
        ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(e[25]), .Q(
        ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(e[26]), .Q(
        ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(e[27]), .Q(
        ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(e[28]), .Q(
        ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(e[29]), .Q(
        ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(e[30]), .Q(
        ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(e[31]), .Q(
        ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(e[32]), .Q(
        ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(e[33]), .Q(
        ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(e[34]), .Q(
        ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(e[35]), .Q(
        ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(e[36]), .Q(
        ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(e[37]), .Q(
        ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(e[38]), .Q(
        ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(e[39]), .Q(
        ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(e[40]), .Q(
        ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(e[41]), .Q(
        ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(e[42]), .Q(
        ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(e[43]), .Q(
        ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(e[44]), .Q(
        ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(e[45]), .Q(
        ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(e[46]), .Q(
        ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(e[47]), .Q(
        ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(e[48]), .Q(
        ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(e[49]), .Q(
        ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(e[50]), .Q(
        ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(e[51]), .Q(
        ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(e[52]), .Q(
        ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(e[53]), .Q(
        ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(e[54]), .Q(
        ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(e[55]), .Q(
        ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(e[56]), .Q(
        ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(e[57]), .Q(
        ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(e[58]), .Q(
        ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(e[59]), .Q(
        ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(e[60]), .Q(
        ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(e[61]), .Q(
        ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(e[62]), .Q(
        ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(e[63]), .Q(
        ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(e[64]), .Q(
        ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(e[65]), .Q(
        ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(e[66]), .Q(
        ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(e[67]), .Q(
        ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(e[68]), .Q(
        ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(e[69]), .Q(
        ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(e[70]), .Q(
        ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(e[71]), .Q(
        ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(e[72]), .Q(
        ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(e[73]), .Q(
        ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(e[74]), .Q(
        ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(e[75]), .Q(
        ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(e[76]), .Q(
        ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(e[77]), .Q(
        ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(e[78]), .Q(
        ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(e[79]), .Q(
        ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(e[80]), .Q(
        ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(e[81]), .Q(
        ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(e[82]), .Q(
        ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(e[83]), .Q(
        ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(e[84]), .Q(
        ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(e[85]), .Q(
        ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(e[86]), .Q(
        ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(e[87]), .Q(
        ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(e[88]), .Q(
        ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(e[89]), .Q(
        ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(e[90]), .Q(
        ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(e[91]), .Q(
        ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(e[92]), .Q(
        ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(e[93]), .Q(
        ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(e[94]), .Q(
        ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(e[95]), .Q(
        ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(e[96]), .Q(
        ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(e[97]), .Q(
        ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(e[98]), .Q(
        ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(e[99]), .Q(
        ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(e[100]), 
        .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(e[101]), 
        .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(e[102]), 
        .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(e[103]), 
        .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(e[104]), 
        .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(e[105]), 
        .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(e[106]), 
        .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(e[107]), 
        .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(e[108]), 
        .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(e[109]), 
        .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(e[110]), 
        .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(e[111]), 
        .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(e[112]), 
        .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(e[113]), 
        .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(e[114]), 
        .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(e[115]), 
        .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(e[116]), 
        .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(e[117]), 
        .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(e[118]), 
        .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(e[119]), 
        .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(e[120]), 
        .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(e[121]), 
        .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(e[122]), 
        .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(e[123]), 
        .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(e[124]), 
        .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(e[125]), 
        .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(e[126]), 
        .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(e[127]), 
        .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(e[128]), 
        .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(e[129]), 
        .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(e[130]), 
        .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(e[131]), 
        .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(e[132]), 
        .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(e[133]), 
        .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(e[134]), 
        .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(e[135]), 
        .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(e[136]), 
        .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(e[137]), 
        .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(e[138]), 
        .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(e[139]), 
        .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(e[140]), 
        .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(e[141]), 
        .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(e[142]), 
        .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(e[143]), 
        .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(e[144]), 
        .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(e[145]), 
        .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(e[146]), 
        .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(e[147]), 
        .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(e[148]), 
        .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(e[149]), 
        .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(e[150]), 
        .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(e[151]), 
        .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(e[152]), 
        .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(e[153]), 
        .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(e[154]), 
        .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(e[155]), 
        .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(e[156]), 
        .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(e[157]), 
        .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(e[158]), 
        .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(e[159]), 
        .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(e[160]), 
        .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(e[161]), 
        .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(e[162]), 
        .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(e[163]), 
        .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(e[164]), 
        .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(e[165]), 
        .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(e[166]), 
        .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(e[167]), 
        .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(e[168]), 
        .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(e[169]), 
        .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(e[170]), 
        .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(e[171]), 
        .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(e[172]), 
        .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(e[173]), 
        .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(e[174]), 
        .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(e[175]), 
        .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(e[176]), 
        .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(e[177]), 
        .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(e[178]), 
        .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(e[179]), 
        .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(e[180]), 
        .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(e[181]), 
        .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(e[182]), 
        .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(e[183]), 
        .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(e[184]), 
        .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(e[185]), 
        .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(e[186]), 
        .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(e[187]), 
        .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(e[188]), 
        .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(e[189]), 
        .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(e[190]), 
        .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(e[191]), 
        .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(e[192]), 
        .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(e[193]), 
        .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(e[194]), 
        .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(e[195]), 
        .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(e[196]), 
        .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(e[197]), 
        .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(e[198]), 
        .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(e[199]), 
        .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(e[200]), 
        .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(e[201]), 
        .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(e[202]), 
        .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(e[203]), 
        .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(e[204]), 
        .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(e[205]), 
        .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(e[206]), 
        .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(e[207]), 
        .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(e[208]), 
        .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(e[209]), 
        .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(e[210]), 
        .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(e[211]), 
        .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(e[212]), 
        .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(e[213]), 
        .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(e[214]), 
        .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(e[215]), 
        .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(e[216]), 
        .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(e[217]), 
        .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(e[218]), 
        .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(e[219]), 
        .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(e[220]), 
        .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(e[221]), 
        .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(e[222]), 
        .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(e[223]), 
        .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(e[224]), 
        .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(e[225]), 
        .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(e[226]), 
        .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(e[227]), 
        .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(e[228]), 
        .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(e[229]), 
        .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(e[230]), 
        .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(e[231]), 
        .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(e[232]), 
        .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(e[233]), 
        .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(e[234]), 
        .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(e[235]), 
        .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(e[236]), 
        .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(e[237]), 
        .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(e[238]), 
        .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(e[239]), 
        .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(e[240]), 
        .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(e[241]), 
        .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(e[242]), 
        .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(e[243]), 
        .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(e[244]), 
        .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(e[245]), 
        .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(e[246]), 
        .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(e[247]), 
        .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(e[248]), 
        .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(e[249]), 
        .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(e[250]), 
        .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(e[251]), 
        .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(e[252]), 
        .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(e[253]), 
        .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(e[254]), 
        .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(e[255]), 
        .Q(ein[255]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(creg_next[0]), .CLK(clk), .RST(rst), .I(m[0]), .Q(
        c[0]) );
  DFF \creg_reg[1]  ( .D(creg_next[1]), .CLK(clk), .RST(rst), .I(m[1]), .Q(
        c[1]) );
  DFF \creg_reg[2]  ( .D(creg_next[2]), .CLK(clk), .RST(rst), .I(m[2]), .Q(
        c[2]) );
  DFF \creg_reg[3]  ( .D(creg_next[3]), .CLK(clk), .RST(rst), .I(m[3]), .Q(
        c[3]) );
  DFF \creg_reg[4]  ( .D(creg_next[4]), .CLK(clk), .RST(rst), .I(m[4]), .Q(
        c[4]) );
  DFF \creg_reg[5]  ( .D(creg_next[5]), .CLK(clk), .RST(rst), .I(m[5]), .Q(
        c[5]) );
  DFF \creg_reg[6]  ( .D(creg_next[6]), .CLK(clk), .RST(rst), .I(m[6]), .Q(
        c[6]) );
  DFF \creg_reg[7]  ( .D(creg_next[7]), .CLK(clk), .RST(rst), .I(m[7]), .Q(
        c[7]) );
  DFF \creg_reg[8]  ( .D(creg_next[8]), .CLK(clk), .RST(rst), .I(m[8]), .Q(
        c[8]) );
  DFF \creg_reg[9]  ( .D(creg_next[9]), .CLK(clk), .RST(rst), .I(m[9]), .Q(
        c[9]) );
  DFF \creg_reg[10]  ( .D(creg_next[10]), .CLK(clk), .RST(rst), .I(m[10]), .Q(
        c[10]) );
  DFF \creg_reg[11]  ( .D(creg_next[11]), .CLK(clk), .RST(rst), .I(m[11]), .Q(
        c[11]) );
  DFF \creg_reg[12]  ( .D(creg_next[12]), .CLK(clk), .RST(rst), .I(m[12]), .Q(
        c[12]) );
  DFF \creg_reg[13]  ( .D(creg_next[13]), .CLK(clk), .RST(rst), .I(m[13]), .Q(
        c[13]) );
  DFF \creg_reg[14]  ( .D(creg_next[14]), .CLK(clk), .RST(rst), .I(m[14]), .Q(
        c[14]) );
  DFF \creg_reg[15]  ( .D(creg_next[15]), .CLK(clk), .RST(rst), .I(m[15]), .Q(
        c[15]) );
  DFF \creg_reg[16]  ( .D(creg_next[16]), .CLK(clk), .RST(rst), .I(m[16]), .Q(
        c[16]) );
  DFF \creg_reg[17]  ( .D(creg_next[17]), .CLK(clk), .RST(rst), .I(m[17]), .Q(
        c[17]) );
  DFF \creg_reg[18]  ( .D(creg_next[18]), .CLK(clk), .RST(rst), .I(m[18]), .Q(
        c[18]) );
  DFF \creg_reg[19]  ( .D(creg_next[19]), .CLK(clk), .RST(rst), .I(m[19]), .Q(
        c[19]) );
  DFF \creg_reg[20]  ( .D(creg_next[20]), .CLK(clk), .RST(rst), .I(m[20]), .Q(
        c[20]) );
  DFF \creg_reg[21]  ( .D(creg_next[21]), .CLK(clk), .RST(rst), .I(m[21]), .Q(
        c[21]) );
  DFF \creg_reg[22]  ( .D(creg_next[22]), .CLK(clk), .RST(rst), .I(m[22]), .Q(
        c[22]) );
  DFF \creg_reg[23]  ( .D(creg_next[23]), .CLK(clk), .RST(rst), .I(m[23]), .Q(
        c[23]) );
  DFF \creg_reg[24]  ( .D(creg_next[24]), .CLK(clk), .RST(rst), .I(m[24]), .Q(
        c[24]) );
  DFF \creg_reg[25]  ( .D(creg_next[25]), .CLK(clk), .RST(rst), .I(m[25]), .Q(
        c[25]) );
  DFF \creg_reg[26]  ( .D(creg_next[26]), .CLK(clk), .RST(rst), .I(m[26]), .Q(
        c[26]) );
  DFF \creg_reg[27]  ( .D(creg_next[27]), .CLK(clk), .RST(rst), .I(m[27]), .Q(
        c[27]) );
  DFF \creg_reg[28]  ( .D(creg_next[28]), .CLK(clk), .RST(rst), .I(m[28]), .Q(
        c[28]) );
  DFF \creg_reg[29]  ( .D(creg_next[29]), .CLK(clk), .RST(rst), .I(m[29]), .Q(
        c[29]) );
  DFF \creg_reg[30]  ( .D(creg_next[30]), .CLK(clk), .RST(rst), .I(m[30]), .Q(
        c[30]) );
  DFF \creg_reg[31]  ( .D(creg_next[31]), .CLK(clk), .RST(rst), .I(m[31]), .Q(
        c[31]) );
  DFF \creg_reg[32]  ( .D(creg_next[32]), .CLK(clk), .RST(rst), .I(m[32]), .Q(
        c[32]) );
  DFF \creg_reg[33]  ( .D(creg_next[33]), .CLK(clk), .RST(rst), .I(m[33]), .Q(
        c[33]) );
  DFF \creg_reg[34]  ( .D(creg_next[34]), .CLK(clk), .RST(rst), .I(m[34]), .Q(
        c[34]) );
  DFF \creg_reg[35]  ( .D(creg_next[35]), .CLK(clk), .RST(rst), .I(m[35]), .Q(
        c[35]) );
  DFF \creg_reg[36]  ( .D(creg_next[36]), .CLK(clk), .RST(rst), .I(m[36]), .Q(
        c[36]) );
  DFF \creg_reg[37]  ( .D(creg_next[37]), .CLK(clk), .RST(rst), .I(m[37]), .Q(
        c[37]) );
  DFF \creg_reg[38]  ( .D(creg_next[38]), .CLK(clk), .RST(rst), .I(m[38]), .Q(
        c[38]) );
  DFF \creg_reg[39]  ( .D(creg_next[39]), .CLK(clk), .RST(rst), .I(m[39]), .Q(
        c[39]) );
  DFF \creg_reg[40]  ( .D(creg_next[40]), .CLK(clk), .RST(rst), .I(m[40]), .Q(
        c[40]) );
  DFF \creg_reg[41]  ( .D(creg_next[41]), .CLK(clk), .RST(rst), .I(m[41]), .Q(
        c[41]) );
  DFF \creg_reg[42]  ( .D(creg_next[42]), .CLK(clk), .RST(rst), .I(m[42]), .Q(
        c[42]) );
  DFF \creg_reg[43]  ( .D(creg_next[43]), .CLK(clk), .RST(rst), .I(m[43]), .Q(
        c[43]) );
  DFF \creg_reg[44]  ( .D(creg_next[44]), .CLK(clk), .RST(rst), .I(m[44]), .Q(
        c[44]) );
  DFF \creg_reg[45]  ( .D(creg_next[45]), .CLK(clk), .RST(rst), .I(m[45]), .Q(
        c[45]) );
  DFF \creg_reg[46]  ( .D(creg_next[46]), .CLK(clk), .RST(rst), .I(m[46]), .Q(
        c[46]) );
  DFF \creg_reg[47]  ( .D(creg_next[47]), .CLK(clk), .RST(rst), .I(m[47]), .Q(
        c[47]) );
  DFF \creg_reg[48]  ( .D(creg_next[48]), .CLK(clk), .RST(rst), .I(m[48]), .Q(
        c[48]) );
  DFF \creg_reg[49]  ( .D(creg_next[49]), .CLK(clk), .RST(rst), .I(m[49]), .Q(
        c[49]) );
  DFF \creg_reg[50]  ( .D(creg_next[50]), .CLK(clk), .RST(rst), .I(m[50]), .Q(
        c[50]) );
  DFF \creg_reg[51]  ( .D(creg_next[51]), .CLK(clk), .RST(rst), .I(m[51]), .Q(
        c[51]) );
  DFF \creg_reg[52]  ( .D(creg_next[52]), .CLK(clk), .RST(rst), .I(m[52]), .Q(
        c[52]) );
  DFF \creg_reg[53]  ( .D(creg_next[53]), .CLK(clk), .RST(rst), .I(m[53]), .Q(
        c[53]) );
  DFF \creg_reg[54]  ( .D(creg_next[54]), .CLK(clk), .RST(rst), .I(m[54]), .Q(
        c[54]) );
  DFF \creg_reg[55]  ( .D(creg_next[55]), .CLK(clk), .RST(rst), .I(m[55]), .Q(
        c[55]) );
  DFF \creg_reg[56]  ( .D(creg_next[56]), .CLK(clk), .RST(rst), .I(m[56]), .Q(
        c[56]) );
  DFF \creg_reg[57]  ( .D(creg_next[57]), .CLK(clk), .RST(rst), .I(m[57]), .Q(
        c[57]) );
  DFF \creg_reg[58]  ( .D(creg_next[58]), .CLK(clk), .RST(rst), .I(m[58]), .Q(
        c[58]) );
  DFF \creg_reg[59]  ( .D(creg_next[59]), .CLK(clk), .RST(rst), .I(m[59]), .Q(
        c[59]) );
  DFF \creg_reg[60]  ( .D(creg_next[60]), .CLK(clk), .RST(rst), .I(m[60]), .Q(
        c[60]) );
  DFF \creg_reg[61]  ( .D(creg_next[61]), .CLK(clk), .RST(rst), .I(m[61]), .Q(
        c[61]) );
  DFF \creg_reg[62]  ( .D(creg_next[62]), .CLK(clk), .RST(rst), .I(m[62]), .Q(
        c[62]) );
  DFF \creg_reg[63]  ( .D(creg_next[63]), .CLK(clk), .RST(rst), .I(m[63]), .Q(
        c[63]) );
  DFF \creg_reg[64]  ( .D(creg_next[64]), .CLK(clk), .RST(rst), .I(m[64]), .Q(
        c[64]) );
  DFF \creg_reg[65]  ( .D(creg_next[65]), .CLK(clk), .RST(rst), .I(m[65]), .Q(
        c[65]) );
  DFF \creg_reg[66]  ( .D(creg_next[66]), .CLK(clk), .RST(rst), .I(m[66]), .Q(
        c[66]) );
  DFF \creg_reg[67]  ( .D(creg_next[67]), .CLK(clk), .RST(rst), .I(m[67]), .Q(
        c[67]) );
  DFF \creg_reg[68]  ( .D(creg_next[68]), .CLK(clk), .RST(rst), .I(m[68]), .Q(
        c[68]) );
  DFF \creg_reg[69]  ( .D(creg_next[69]), .CLK(clk), .RST(rst), .I(m[69]), .Q(
        c[69]) );
  DFF \creg_reg[70]  ( .D(creg_next[70]), .CLK(clk), .RST(rst), .I(m[70]), .Q(
        c[70]) );
  DFF \creg_reg[71]  ( .D(creg_next[71]), .CLK(clk), .RST(rst), .I(m[71]), .Q(
        c[71]) );
  DFF \creg_reg[72]  ( .D(creg_next[72]), .CLK(clk), .RST(rst), .I(m[72]), .Q(
        c[72]) );
  DFF \creg_reg[73]  ( .D(creg_next[73]), .CLK(clk), .RST(rst), .I(m[73]), .Q(
        c[73]) );
  DFF \creg_reg[74]  ( .D(creg_next[74]), .CLK(clk), .RST(rst), .I(m[74]), .Q(
        c[74]) );
  DFF \creg_reg[75]  ( .D(creg_next[75]), .CLK(clk), .RST(rst), .I(m[75]), .Q(
        c[75]) );
  DFF \creg_reg[76]  ( .D(creg_next[76]), .CLK(clk), .RST(rst), .I(m[76]), .Q(
        c[76]) );
  DFF \creg_reg[77]  ( .D(creg_next[77]), .CLK(clk), .RST(rst), .I(m[77]), .Q(
        c[77]) );
  DFF \creg_reg[78]  ( .D(creg_next[78]), .CLK(clk), .RST(rst), .I(m[78]), .Q(
        c[78]) );
  DFF \creg_reg[79]  ( .D(creg_next[79]), .CLK(clk), .RST(rst), .I(m[79]), .Q(
        c[79]) );
  DFF \creg_reg[80]  ( .D(creg_next[80]), .CLK(clk), .RST(rst), .I(m[80]), .Q(
        c[80]) );
  DFF \creg_reg[81]  ( .D(creg_next[81]), .CLK(clk), .RST(rst), .I(m[81]), .Q(
        c[81]) );
  DFF \creg_reg[82]  ( .D(creg_next[82]), .CLK(clk), .RST(rst), .I(m[82]), .Q(
        c[82]) );
  DFF \creg_reg[83]  ( .D(creg_next[83]), .CLK(clk), .RST(rst), .I(m[83]), .Q(
        c[83]) );
  DFF \creg_reg[84]  ( .D(creg_next[84]), .CLK(clk), .RST(rst), .I(m[84]), .Q(
        c[84]) );
  DFF \creg_reg[85]  ( .D(creg_next[85]), .CLK(clk), .RST(rst), .I(m[85]), .Q(
        c[85]) );
  DFF \creg_reg[86]  ( .D(creg_next[86]), .CLK(clk), .RST(rst), .I(m[86]), .Q(
        c[86]) );
  DFF \creg_reg[87]  ( .D(creg_next[87]), .CLK(clk), .RST(rst), .I(m[87]), .Q(
        c[87]) );
  DFF \creg_reg[88]  ( .D(creg_next[88]), .CLK(clk), .RST(rst), .I(m[88]), .Q(
        c[88]) );
  DFF \creg_reg[89]  ( .D(creg_next[89]), .CLK(clk), .RST(rst), .I(m[89]), .Q(
        c[89]) );
  DFF \creg_reg[90]  ( .D(creg_next[90]), .CLK(clk), .RST(rst), .I(m[90]), .Q(
        c[90]) );
  DFF \creg_reg[91]  ( .D(creg_next[91]), .CLK(clk), .RST(rst), .I(m[91]), .Q(
        c[91]) );
  DFF \creg_reg[92]  ( .D(creg_next[92]), .CLK(clk), .RST(rst), .I(m[92]), .Q(
        c[92]) );
  DFF \creg_reg[93]  ( .D(creg_next[93]), .CLK(clk), .RST(rst), .I(m[93]), .Q(
        c[93]) );
  DFF \creg_reg[94]  ( .D(creg_next[94]), .CLK(clk), .RST(rst), .I(m[94]), .Q(
        c[94]) );
  DFF \creg_reg[95]  ( .D(creg_next[95]), .CLK(clk), .RST(rst), .I(m[95]), .Q(
        c[95]) );
  DFF \creg_reg[96]  ( .D(creg_next[96]), .CLK(clk), .RST(rst), .I(m[96]), .Q(
        c[96]) );
  DFF \creg_reg[97]  ( .D(creg_next[97]), .CLK(clk), .RST(rst), .I(m[97]), .Q(
        c[97]) );
  DFF \creg_reg[98]  ( .D(creg_next[98]), .CLK(clk), .RST(rst), .I(m[98]), .Q(
        c[98]) );
  DFF \creg_reg[99]  ( .D(creg_next[99]), .CLK(clk), .RST(rst), .I(m[99]), .Q(
        c[99]) );
  DFF \creg_reg[100]  ( .D(creg_next[100]), .CLK(clk), .RST(rst), .I(m[100]), 
        .Q(c[100]) );
  DFF \creg_reg[101]  ( .D(creg_next[101]), .CLK(clk), .RST(rst), .I(m[101]), 
        .Q(c[101]) );
  DFF \creg_reg[102]  ( .D(creg_next[102]), .CLK(clk), .RST(rst), .I(m[102]), 
        .Q(c[102]) );
  DFF \creg_reg[103]  ( .D(creg_next[103]), .CLK(clk), .RST(rst), .I(m[103]), 
        .Q(c[103]) );
  DFF \creg_reg[104]  ( .D(creg_next[104]), .CLK(clk), .RST(rst), .I(m[104]), 
        .Q(c[104]) );
  DFF \creg_reg[105]  ( .D(creg_next[105]), .CLK(clk), .RST(rst), .I(m[105]), 
        .Q(c[105]) );
  DFF \creg_reg[106]  ( .D(creg_next[106]), .CLK(clk), .RST(rst), .I(m[106]), 
        .Q(c[106]) );
  DFF \creg_reg[107]  ( .D(creg_next[107]), .CLK(clk), .RST(rst), .I(m[107]), 
        .Q(c[107]) );
  DFF \creg_reg[108]  ( .D(creg_next[108]), .CLK(clk), .RST(rst), .I(m[108]), 
        .Q(c[108]) );
  DFF \creg_reg[109]  ( .D(creg_next[109]), .CLK(clk), .RST(rst), .I(m[109]), 
        .Q(c[109]) );
  DFF \creg_reg[110]  ( .D(creg_next[110]), .CLK(clk), .RST(rst), .I(m[110]), 
        .Q(c[110]) );
  DFF \creg_reg[111]  ( .D(creg_next[111]), .CLK(clk), .RST(rst), .I(m[111]), 
        .Q(c[111]) );
  DFF \creg_reg[112]  ( .D(creg_next[112]), .CLK(clk), .RST(rst), .I(m[112]), 
        .Q(c[112]) );
  DFF \creg_reg[113]  ( .D(creg_next[113]), .CLK(clk), .RST(rst), .I(m[113]), 
        .Q(c[113]) );
  DFF \creg_reg[114]  ( .D(creg_next[114]), .CLK(clk), .RST(rst), .I(m[114]), 
        .Q(c[114]) );
  DFF \creg_reg[115]  ( .D(creg_next[115]), .CLK(clk), .RST(rst), .I(m[115]), 
        .Q(c[115]) );
  DFF \creg_reg[116]  ( .D(creg_next[116]), .CLK(clk), .RST(rst), .I(m[116]), 
        .Q(c[116]) );
  DFF \creg_reg[117]  ( .D(creg_next[117]), .CLK(clk), .RST(rst), .I(m[117]), 
        .Q(c[117]) );
  DFF \creg_reg[118]  ( .D(creg_next[118]), .CLK(clk), .RST(rst), .I(m[118]), 
        .Q(c[118]) );
  DFF \creg_reg[119]  ( .D(creg_next[119]), .CLK(clk), .RST(rst), .I(m[119]), 
        .Q(c[119]) );
  DFF \creg_reg[120]  ( .D(creg_next[120]), .CLK(clk), .RST(rst), .I(m[120]), 
        .Q(c[120]) );
  DFF \creg_reg[121]  ( .D(creg_next[121]), .CLK(clk), .RST(rst), .I(m[121]), 
        .Q(c[121]) );
  DFF \creg_reg[122]  ( .D(creg_next[122]), .CLK(clk), .RST(rst), .I(m[122]), 
        .Q(c[122]) );
  DFF \creg_reg[123]  ( .D(creg_next[123]), .CLK(clk), .RST(rst), .I(m[123]), 
        .Q(c[123]) );
  DFF \creg_reg[124]  ( .D(creg_next[124]), .CLK(clk), .RST(rst), .I(m[124]), 
        .Q(c[124]) );
  DFF \creg_reg[125]  ( .D(creg_next[125]), .CLK(clk), .RST(rst), .I(m[125]), 
        .Q(c[125]) );
  DFF \creg_reg[126]  ( .D(creg_next[126]), .CLK(clk), .RST(rst), .I(m[126]), 
        .Q(c[126]) );
  DFF \creg_reg[127]  ( .D(creg_next[127]), .CLK(clk), .RST(rst), .I(m[127]), 
        .Q(c[127]) );
  DFF \creg_reg[128]  ( .D(creg_next[128]), .CLK(clk), .RST(rst), .I(m[128]), 
        .Q(c[128]) );
  DFF \creg_reg[129]  ( .D(creg_next[129]), .CLK(clk), .RST(rst), .I(m[129]), 
        .Q(c[129]) );
  DFF \creg_reg[130]  ( .D(creg_next[130]), .CLK(clk), .RST(rst), .I(m[130]), 
        .Q(c[130]) );
  DFF \creg_reg[131]  ( .D(creg_next[131]), .CLK(clk), .RST(rst), .I(m[131]), 
        .Q(c[131]) );
  DFF \creg_reg[132]  ( .D(creg_next[132]), .CLK(clk), .RST(rst), .I(m[132]), 
        .Q(c[132]) );
  DFF \creg_reg[133]  ( .D(creg_next[133]), .CLK(clk), .RST(rst), .I(m[133]), 
        .Q(c[133]) );
  DFF \creg_reg[134]  ( .D(creg_next[134]), .CLK(clk), .RST(rst), .I(m[134]), 
        .Q(c[134]) );
  DFF \creg_reg[135]  ( .D(creg_next[135]), .CLK(clk), .RST(rst), .I(m[135]), 
        .Q(c[135]) );
  DFF \creg_reg[136]  ( .D(creg_next[136]), .CLK(clk), .RST(rst), .I(m[136]), 
        .Q(c[136]) );
  DFF \creg_reg[137]  ( .D(creg_next[137]), .CLK(clk), .RST(rst), .I(m[137]), 
        .Q(c[137]) );
  DFF \creg_reg[138]  ( .D(creg_next[138]), .CLK(clk), .RST(rst), .I(m[138]), 
        .Q(c[138]) );
  DFF \creg_reg[139]  ( .D(creg_next[139]), .CLK(clk), .RST(rst), .I(m[139]), 
        .Q(c[139]) );
  DFF \creg_reg[140]  ( .D(creg_next[140]), .CLK(clk), .RST(rst), .I(m[140]), 
        .Q(c[140]) );
  DFF \creg_reg[141]  ( .D(creg_next[141]), .CLK(clk), .RST(rst), .I(m[141]), 
        .Q(c[141]) );
  DFF \creg_reg[142]  ( .D(creg_next[142]), .CLK(clk), .RST(rst), .I(m[142]), 
        .Q(c[142]) );
  DFF \creg_reg[143]  ( .D(creg_next[143]), .CLK(clk), .RST(rst), .I(m[143]), 
        .Q(c[143]) );
  DFF \creg_reg[144]  ( .D(creg_next[144]), .CLK(clk), .RST(rst), .I(m[144]), 
        .Q(c[144]) );
  DFF \creg_reg[145]  ( .D(creg_next[145]), .CLK(clk), .RST(rst), .I(m[145]), 
        .Q(c[145]) );
  DFF \creg_reg[146]  ( .D(creg_next[146]), .CLK(clk), .RST(rst), .I(m[146]), 
        .Q(c[146]) );
  DFF \creg_reg[147]  ( .D(creg_next[147]), .CLK(clk), .RST(rst), .I(m[147]), 
        .Q(c[147]) );
  DFF \creg_reg[148]  ( .D(creg_next[148]), .CLK(clk), .RST(rst), .I(m[148]), 
        .Q(c[148]) );
  DFF \creg_reg[149]  ( .D(creg_next[149]), .CLK(clk), .RST(rst), .I(m[149]), 
        .Q(c[149]) );
  DFF \creg_reg[150]  ( .D(creg_next[150]), .CLK(clk), .RST(rst), .I(m[150]), 
        .Q(c[150]) );
  DFF \creg_reg[151]  ( .D(creg_next[151]), .CLK(clk), .RST(rst), .I(m[151]), 
        .Q(c[151]) );
  DFF \creg_reg[152]  ( .D(creg_next[152]), .CLK(clk), .RST(rst), .I(m[152]), 
        .Q(c[152]) );
  DFF \creg_reg[153]  ( .D(creg_next[153]), .CLK(clk), .RST(rst), .I(m[153]), 
        .Q(c[153]) );
  DFF \creg_reg[154]  ( .D(creg_next[154]), .CLK(clk), .RST(rst), .I(m[154]), 
        .Q(c[154]) );
  DFF \creg_reg[155]  ( .D(creg_next[155]), .CLK(clk), .RST(rst), .I(m[155]), 
        .Q(c[155]) );
  DFF \creg_reg[156]  ( .D(creg_next[156]), .CLK(clk), .RST(rst), .I(m[156]), 
        .Q(c[156]) );
  DFF \creg_reg[157]  ( .D(creg_next[157]), .CLK(clk), .RST(rst), .I(m[157]), 
        .Q(c[157]) );
  DFF \creg_reg[158]  ( .D(creg_next[158]), .CLK(clk), .RST(rst), .I(m[158]), 
        .Q(c[158]) );
  DFF \creg_reg[159]  ( .D(creg_next[159]), .CLK(clk), .RST(rst), .I(m[159]), 
        .Q(c[159]) );
  DFF \creg_reg[160]  ( .D(creg_next[160]), .CLK(clk), .RST(rst), .I(m[160]), 
        .Q(c[160]) );
  DFF \creg_reg[161]  ( .D(creg_next[161]), .CLK(clk), .RST(rst), .I(m[161]), 
        .Q(c[161]) );
  DFF \creg_reg[162]  ( .D(creg_next[162]), .CLK(clk), .RST(rst), .I(m[162]), 
        .Q(c[162]) );
  DFF \creg_reg[163]  ( .D(creg_next[163]), .CLK(clk), .RST(rst), .I(m[163]), 
        .Q(c[163]) );
  DFF \creg_reg[164]  ( .D(creg_next[164]), .CLK(clk), .RST(rst), .I(m[164]), 
        .Q(c[164]) );
  DFF \creg_reg[165]  ( .D(creg_next[165]), .CLK(clk), .RST(rst), .I(m[165]), 
        .Q(c[165]) );
  DFF \creg_reg[166]  ( .D(creg_next[166]), .CLK(clk), .RST(rst), .I(m[166]), 
        .Q(c[166]) );
  DFF \creg_reg[167]  ( .D(creg_next[167]), .CLK(clk), .RST(rst), .I(m[167]), 
        .Q(c[167]) );
  DFF \creg_reg[168]  ( .D(creg_next[168]), .CLK(clk), .RST(rst), .I(m[168]), 
        .Q(c[168]) );
  DFF \creg_reg[169]  ( .D(creg_next[169]), .CLK(clk), .RST(rst), .I(m[169]), 
        .Q(c[169]) );
  DFF \creg_reg[170]  ( .D(creg_next[170]), .CLK(clk), .RST(rst), .I(m[170]), 
        .Q(c[170]) );
  DFF \creg_reg[171]  ( .D(creg_next[171]), .CLK(clk), .RST(rst), .I(m[171]), 
        .Q(c[171]) );
  DFF \creg_reg[172]  ( .D(creg_next[172]), .CLK(clk), .RST(rst), .I(m[172]), 
        .Q(c[172]) );
  DFF \creg_reg[173]  ( .D(creg_next[173]), .CLK(clk), .RST(rst), .I(m[173]), 
        .Q(c[173]) );
  DFF \creg_reg[174]  ( .D(creg_next[174]), .CLK(clk), .RST(rst), .I(m[174]), 
        .Q(c[174]) );
  DFF \creg_reg[175]  ( .D(creg_next[175]), .CLK(clk), .RST(rst), .I(m[175]), 
        .Q(c[175]) );
  DFF \creg_reg[176]  ( .D(creg_next[176]), .CLK(clk), .RST(rst), .I(m[176]), 
        .Q(c[176]) );
  DFF \creg_reg[177]  ( .D(creg_next[177]), .CLK(clk), .RST(rst), .I(m[177]), 
        .Q(c[177]) );
  DFF \creg_reg[178]  ( .D(creg_next[178]), .CLK(clk), .RST(rst), .I(m[178]), 
        .Q(c[178]) );
  DFF \creg_reg[179]  ( .D(creg_next[179]), .CLK(clk), .RST(rst), .I(m[179]), 
        .Q(c[179]) );
  DFF \creg_reg[180]  ( .D(creg_next[180]), .CLK(clk), .RST(rst), .I(m[180]), 
        .Q(c[180]) );
  DFF \creg_reg[181]  ( .D(creg_next[181]), .CLK(clk), .RST(rst), .I(m[181]), 
        .Q(c[181]) );
  DFF \creg_reg[182]  ( .D(creg_next[182]), .CLK(clk), .RST(rst), .I(m[182]), 
        .Q(c[182]) );
  DFF \creg_reg[183]  ( .D(creg_next[183]), .CLK(clk), .RST(rst), .I(m[183]), 
        .Q(c[183]) );
  DFF \creg_reg[184]  ( .D(creg_next[184]), .CLK(clk), .RST(rst), .I(m[184]), 
        .Q(c[184]) );
  DFF \creg_reg[185]  ( .D(creg_next[185]), .CLK(clk), .RST(rst), .I(m[185]), 
        .Q(c[185]) );
  DFF \creg_reg[186]  ( .D(creg_next[186]), .CLK(clk), .RST(rst), .I(m[186]), 
        .Q(c[186]) );
  DFF \creg_reg[187]  ( .D(creg_next[187]), .CLK(clk), .RST(rst), .I(m[187]), 
        .Q(c[187]) );
  DFF \creg_reg[188]  ( .D(creg_next[188]), .CLK(clk), .RST(rst), .I(m[188]), 
        .Q(c[188]) );
  DFF \creg_reg[189]  ( .D(creg_next[189]), .CLK(clk), .RST(rst), .I(m[189]), 
        .Q(c[189]) );
  DFF \creg_reg[190]  ( .D(creg_next[190]), .CLK(clk), .RST(rst), .I(m[190]), 
        .Q(c[190]) );
  DFF \creg_reg[191]  ( .D(creg_next[191]), .CLK(clk), .RST(rst), .I(m[191]), 
        .Q(c[191]) );
  DFF \creg_reg[192]  ( .D(creg_next[192]), .CLK(clk), .RST(rst), .I(m[192]), 
        .Q(c[192]) );
  DFF \creg_reg[193]  ( .D(creg_next[193]), .CLK(clk), .RST(rst), .I(m[193]), 
        .Q(c[193]) );
  DFF \creg_reg[194]  ( .D(creg_next[194]), .CLK(clk), .RST(rst), .I(m[194]), 
        .Q(c[194]) );
  DFF \creg_reg[195]  ( .D(creg_next[195]), .CLK(clk), .RST(rst), .I(m[195]), 
        .Q(c[195]) );
  DFF \creg_reg[196]  ( .D(creg_next[196]), .CLK(clk), .RST(rst), .I(m[196]), 
        .Q(c[196]) );
  DFF \creg_reg[197]  ( .D(creg_next[197]), .CLK(clk), .RST(rst), .I(m[197]), 
        .Q(c[197]) );
  DFF \creg_reg[198]  ( .D(creg_next[198]), .CLK(clk), .RST(rst), .I(m[198]), 
        .Q(c[198]) );
  DFF \creg_reg[199]  ( .D(creg_next[199]), .CLK(clk), .RST(rst), .I(m[199]), 
        .Q(c[199]) );
  DFF \creg_reg[200]  ( .D(creg_next[200]), .CLK(clk), .RST(rst), .I(m[200]), 
        .Q(c[200]) );
  DFF \creg_reg[201]  ( .D(creg_next[201]), .CLK(clk), .RST(rst), .I(m[201]), 
        .Q(c[201]) );
  DFF \creg_reg[202]  ( .D(creg_next[202]), .CLK(clk), .RST(rst), .I(m[202]), 
        .Q(c[202]) );
  DFF \creg_reg[203]  ( .D(creg_next[203]), .CLK(clk), .RST(rst), .I(m[203]), 
        .Q(c[203]) );
  DFF \creg_reg[204]  ( .D(creg_next[204]), .CLK(clk), .RST(rst), .I(m[204]), 
        .Q(c[204]) );
  DFF \creg_reg[205]  ( .D(creg_next[205]), .CLK(clk), .RST(rst), .I(m[205]), 
        .Q(c[205]) );
  DFF \creg_reg[206]  ( .D(creg_next[206]), .CLK(clk), .RST(rst), .I(m[206]), 
        .Q(c[206]) );
  DFF \creg_reg[207]  ( .D(creg_next[207]), .CLK(clk), .RST(rst), .I(m[207]), 
        .Q(c[207]) );
  DFF \creg_reg[208]  ( .D(creg_next[208]), .CLK(clk), .RST(rst), .I(m[208]), 
        .Q(c[208]) );
  DFF \creg_reg[209]  ( .D(creg_next[209]), .CLK(clk), .RST(rst), .I(m[209]), 
        .Q(c[209]) );
  DFF \creg_reg[210]  ( .D(creg_next[210]), .CLK(clk), .RST(rst), .I(m[210]), 
        .Q(c[210]) );
  DFF \creg_reg[211]  ( .D(creg_next[211]), .CLK(clk), .RST(rst), .I(m[211]), 
        .Q(c[211]) );
  DFF \creg_reg[212]  ( .D(creg_next[212]), .CLK(clk), .RST(rst), .I(m[212]), 
        .Q(c[212]) );
  DFF \creg_reg[213]  ( .D(creg_next[213]), .CLK(clk), .RST(rst), .I(m[213]), 
        .Q(c[213]) );
  DFF \creg_reg[214]  ( .D(creg_next[214]), .CLK(clk), .RST(rst), .I(m[214]), 
        .Q(c[214]) );
  DFF \creg_reg[215]  ( .D(creg_next[215]), .CLK(clk), .RST(rst), .I(m[215]), 
        .Q(c[215]) );
  DFF \creg_reg[216]  ( .D(creg_next[216]), .CLK(clk), .RST(rst), .I(m[216]), 
        .Q(c[216]) );
  DFF \creg_reg[217]  ( .D(creg_next[217]), .CLK(clk), .RST(rst), .I(m[217]), 
        .Q(c[217]) );
  DFF \creg_reg[218]  ( .D(creg_next[218]), .CLK(clk), .RST(rst), .I(m[218]), 
        .Q(c[218]) );
  DFF \creg_reg[219]  ( .D(creg_next[219]), .CLK(clk), .RST(rst), .I(m[219]), 
        .Q(c[219]) );
  DFF \creg_reg[220]  ( .D(creg_next[220]), .CLK(clk), .RST(rst), .I(m[220]), 
        .Q(c[220]) );
  DFF \creg_reg[221]  ( .D(creg_next[221]), .CLK(clk), .RST(rst), .I(m[221]), 
        .Q(c[221]) );
  DFF \creg_reg[222]  ( .D(creg_next[222]), .CLK(clk), .RST(rst), .I(m[222]), 
        .Q(c[222]) );
  DFF \creg_reg[223]  ( .D(creg_next[223]), .CLK(clk), .RST(rst), .I(m[223]), 
        .Q(c[223]) );
  DFF \creg_reg[224]  ( .D(creg_next[224]), .CLK(clk), .RST(rst), .I(m[224]), 
        .Q(c[224]) );
  DFF \creg_reg[225]  ( .D(creg_next[225]), .CLK(clk), .RST(rst), .I(m[225]), 
        .Q(c[225]) );
  DFF \creg_reg[226]  ( .D(creg_next[226]), .CLK(clk), .RST(rst), .I(m[226]), 
        .Q(c[226]) );
  DFF \creg_reg[227]  ( .D(creg_next[227]), .CLK(clk), .RST(rst), .I(m[227]), 
        .Q(c[227]) );
  DFF \creg_reg[228]  ( .D(creg_next[228]), .CLK(clk), .RST(rst), .I(m[228]), 
        .Q(c[228]) );
  DFF \creg_reg[229]  ( .D(creg_next[229]), .CLK(clk), .RST(rst), .I(m[229]), 
        .Q(c[229]) );
  DFF \creg_reg[230]  ( .D(creg_next[230]), .CLK(clk), .RST(rst), .I(m[230]), 
        .Q(c[230]) );
  DFF \creg_reg[231]  ( .D(creg_next[231]), .CLK(clk), .RST(rst), .I(m[231]), 
        .Q(c[231]) );
  DFF \creg_reg[232]  ( .D(creg_next[232]), .CLK(clk), .RST(rst), .I(m[232]), 
        .Q(c[232]) );
  DFF \creg_reg[233]  ( .D(creg_next[233]), .CLK(clk), .RST(rst), .I(m[233]), 
        .Q(c[233]) );
  DFF \creg_reg[234]  ( .D(creg_next[234]), .CLK(clk), .RST(rst), .I(m[234]), 
        .Q(c[234]) );
  DFF \creg_reg[235]  ( .D(creg_next[235]), .CLK(clk), .RST(rst), .I(m[235]), 
        .Q(c[235]) );
  DFF \creg_reg[236]  ( .D(creg_next[236]), .CLK(clk), .RST(rst), .I(m[236]), 
        .Q(c[236]) );
  DFF \creg_reg[237]  ( .D(creg_next[237]), .CLK(clk), .RST(rst), .I(m[237]), 
        .Q(c[237]) );
  DFF \creg_reg[238]  ( .D(creg_next[238]), .CLK(clk), .RST(rst), .I(m[238]), 
        .Q(c[238]) );
  DFF \creg_reg[239]  ( .D(creg_next[239]), .CLK(clk), .RST(rst), .I(m[239]), 
        .Q(c[239]) );
  DFF \creg_reg[240]  ( .D(creg_next[240]), .CLK(clk), .RST(rst), .I(m[240]), 
        .Q(c[240]) );
  DFF \creg_reg[241]  ( .D(creg_next[241]), .CLK(clk), .RST(rst), .I(m[241]), 
        .Q(c[241]) );
  DFF \creg_reg[242]  ( .D(creg_next[242]), .CLK(clk), .RST(rst), .I(m[242]), 
        .Q(c[242]) );
  DFF \creg_reg[243]  ( .D(creg_next[243]), .CLK(clk), .RST(rst), .I(m[243]), 
        .Q(c[243]) );
  DFF \creg_reg[244]  ( .D(creg_next[244]), .CLK(clk), .RST(rst), .I(m[244]), 
        .Q(c[244]) );
  DFF \creg_reg[245]  ( .D(creg_next[245]), .CLK(clk), .RST(rst), .I(m[245]), 
        .Q(c[245]) );
  DFF \creg_reg[246]  ( .D(creg_next[246]), .CLK(clk), .RST(rst), .I(m[246]), 
        .Q(c[246]) );
  DFF \creg_reg[247]  ( .D(creg_next[247]), .CLK(clk), .RST(rst), .I(m[247]), 
        .Q(c[247]) );
  DFF \creg_reg[248]  ( .D(creg_next[248]), .CLK(clk), .RST(rst), .I(m[248]), 
        .Q(c[248]) );
  DFF \creg_reg[249]  ( .D(creg_next[249]), .CLK(clk), .RST(rst), .I(m[249]), 
        .Q(c[249]) );
  DFF \creg_reg[250]  ( .D(creg_next[250]), .CLK(clk), .RST(rst), .I(m[250]), 
        .Q(c[250]) );
  DFF \creg_reg[251]  ( .D(creg_next[251]), .CLK(clk), .RST(rst), .I(m[251]), 
        .Q(c[251]) );
  DFF \creg_reg[252]  ( .D(creg_next[252]), .CLK(clk), .RST(rst), .I(m[252]), 
        .Q(c[252]) );
  DFF \creg_reg[253]  ( .D(creg_next[253]), .CLK(clk), .RST(rst), .I(m[253]), 
        .Q(c[253]) );
  DFF \creg_reg[254]  ( .D(creg_next[254]), .CLK(clk), .RST(rst), .I(m[254]), 
        .Q(c[254]) );
  DFF \creg_reg[255]  ( .D(creg_next[255]), .CLK(clk), .RST(rst), .I(m[255]), 
        .Q(c[255]) );
  XOR U268 ( .A(start_in[255]), .B(mul_pow), .Z(n8) );
  NANDN U269 ( .A(first_one), .B(n265), .Z(n6) );
  NAND U270 ( .A(n266), .B(ein[255]), .Z(n265) );
  AND U271 ( .A(mul_pow), .B(start_in[255]), .Z(n266) );
  NAND U272 ( .A(n267), .B(n268), .Z(_0_net_) );
  NANDN U273 ( .A(mul_pow), .B(first_one), .Z(n268) );
  NAND U274 ( .A(first_one), .B(ein[255]), .Z(n267) );
endmodule

