
module hamming_N16000_CC128 ( clk, rst, x, y, o );
  input [124:0] x;
  input [124:0] y;
  output [13:0] o;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825;
  wire   [13:0] oglobal;

  DFF \oglobal_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(oglobal[13]) );
  DFF \oglobal_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(oglobal[12]) );
  DFF \oglobal_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(oglobal[11]) );
  DFF \oglobal_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(oglobal[10]) );
  DFF \oglobal_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(oglobal[9]) );
  DFF \oglobal_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(oglobal[8]) );
  DFF \oglobal_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(oglobal[7]) );
  DFF \oglobal_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(oglobal[6]) );
  DFF \oglobal_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(oglobal[5]) );
  DFF \oglobal_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(oglobal[4]) );
  DFF \oglobal_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(oglobal[3]) );
  DFF \oglobal_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(oglobal[2]) );
  DFF \oglobal_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(oglobal[1]) );
  DFF \oglobal_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(oglobal[0]) );
  XNOR U128 ( .A(n482), .B(oglobal[0]), .Z(n483) );
  NAND U129 ( .A(n642), .B(n643), .Z(n1) );
  XOR U130 ( .A(n642), .B(n643), .Z(n2) );
  NANDN U131 ( .A(n641), .B(n2), .Z(n3) );
  NAND U132 ( .A(n1), .B(n3), .Z(n712) );
  NAND U133 ( .A(n467), .B(n468), .Z(n4) );
  XOR U134 ( .A(n467), .B(n468), .Z(n5) );
  NANDN U135 ( .A(n466), .B(n5), .Z(n6) );
  NAND U136 ( .A(n4), .B(n6), .Z(n575) );
  NAND U137 ( .A(n651), .B(n653), .Z(n7) );
  XOR U138 ( .A(n651), .B(n653), .Z(n8) );
  NAND U139 ( .A(n8), .B(n652), .Z(n9) );
  NAND U140 ( .A(n7), .B(n9), .Z(n722) );
  NAND U141 ( .A(n570), .B(n572), .Z(n10) );
  XOR U142 ( .A(n570), .B(n572), .Z(n11) );
  NAND U143 ( .A(n11), .B(n571), .Z(n12) );
  NAND U144 ( .A(n10), .B(n12), .Z(n725) );
  NAND U145 ( .A(n426), .B(n427), .Z(n13) );
  XOR U146 ( .A(n426), .B(n427), .Z(n14) );
  NANDN U147 ( .A(n425), .B(n14), .Z(n15) );
  NAND U148 ( .A(n13), .B(n15), .Z(n551) );
  NAND U149 ( .A(n535), .B(n536), .Z(n16) );
  XOR U150 ( .A(n535), .B(n536), .Z(n17) );
  NANDN U151 ( .A(n534), .B(n17), .Z(n18) );
  NAND U152 ( .A(n16), .B(n18), .Z(n736) );
  XOR U153 ( .A(n611), .B(n610), .Z(n19) );
  XNOR U154 ( .A(n613), .B(n19), .Z(n661) );
  NAND U155 ( .A(n732), .B(n733), .Z(n20) );
  XOR U156 ( .A(n732), .B(n733), .Z(n21) );
  NANDN U157 ( .A(n731), .B(n21), .Z(n22) );
  NAND U158 ( .A(n20), .B(n22), .Z(n760) );
  NAND U159 ( .A(n375), .B(n376), .Z(n23) );
  XOR U160 ( .A(n375), .B(n376), .Z(n24) );
  NANDN U161 ( .A(n374), .B(n24), .Z(n25) );
  NAND U162 ( .A(n23), .B(n25), .Z(n567) );
  XNOR U163 ( .A(n247), .B(n246), .Z(n248) );
  XOR U164 ( .A(n517), .B(n515), .Z(n26) );
  NANDN U165 ( .A(n516), .B(n26), .Z(n27) );
  NAND U166 ( .A(n517), .B(n515), .Z(n28) );
  AND U167 ( .A(n27), .B(n28), .Z(n537) );
  NAND U168 ( .A(n632), .B(n633), .Z(n29) );
  XOR U169 ( .A(n632), .B(n633), .Z(n30) );
  NANDN U170 ( .A(n631), .B(n30), .Z(n31) );
  NAND U171 ( .A(n29), .B(n31), .Z(n692) );
  NAND U172 ( .A(n607), .B(n608), .Z(n32) );
  XOR U173 ( .A(n607), .B(n608), .Z(n33) );
  NANDN U174 ( .A(n606), .B(n33), .Z(n34) );
  NAND U175 ( .A(n32), .B(n34), .Z(n715) );
  NAND U176 ( .A(n648), .B(n649), .Z(n35) );
  XOR U177 ( .A(n648), .B(n649), .Z(n36) );
  NANDN U178 ( .A(n647), .B(n36), .Z(n37) );
  NAND U179 ( .A(n35), .B(n37), .Z(n713) );
  XOR U180 ( .A(n658), .B(n656), .Z(n38) );
  NANDN U181 ( .A(n657), .B(n38), .Z(n39) );
  NAND U182 ( .A(n658), .B(n656), .Z(n40) );
  AND U183 ( .A(n39), .B(n40), .Z(n686) );
  NAND U184 ( .A(n725), .B(n726), .Z(n41) );
  XOR U185 ( .A(n725), .B(n726), .Z(n42) );
  NANDN U186 ( .A(n724), .B(n42), .Z(n43) );
  NAND U187 ( .A(n41), .B(n43), .Z(n762) );
  XOR U188 ( .A(n671), .B(n670), .Z(n44) );
  XNOR U189 ( .A(n672), .B(n44), .Z(n673) );
  XOR U190 ( .A(n730), .B(n728), .Z(n45) );
  NANDN U191 ( .A(n729), .B(n45), .Z(n46) );
  NAND U192 ( .A(n730), .B(n728), .Z(n47) );
  AND U193 ( .A(n46), .B(n47), .Z(n761) );
  XOR U194 ( .A(n660), .B(n661), .Z(n48) );
  XNOR U195 ( .A(n659), .B(n48), .Z(n568) );
  XNOR U196 ( .A(n524), .B(n525), .Z(n49) );
  XNOR U197 ( .A(n523), .B(n49), .Z(n527) );
  XNOR U198 ( .A(n477), .B(n476), .Z(n478) );
  XNOR U199 ( .A(n471), .B(n470), .Z(n472) );
  NAND U200 ( .A(n639), .B(n640), .Z(n50) );
  XOR U201 ( .A(n639), .B(n640), .Z(n51) );
  NANDN U202 ( .A(n638), .B(n51), .Z(n52) );
  NAND U203 ( .A(n50), .B(n52), .Z(n694) );
  NAND U204 ( .A(n604), .B(n605), .Z(n53) );
  XOR U205 ( .A(n604), .B(n605), .Z(n54) );
  NANDN U206 ( .A(n603), .B(n54), .Z(n55) );
  NAND U207 ( .A(n53), .B(n55), .Z(n716) );
  NAND U208 ( .A(n645), .B(n646), .Z(n56) );
  XOR U209 ( .A(n645), .B(n646), .Z(n57) );
  NANDN U210 ( .A(n644), .B(n57), .Z(n58) );
  NAND U211 ( .A(n56), .B(n58), .Z(n714) );
  NAND U212 ( .A(n537), .B(n539), .Z(n59) );
  XOR U213 ( .A(n537), .B(n539), .Z(n60) );
  NAND U214 ( .A(n60), .B(n538), .Z(n61) );
  NAND U215 ( .A(n59), .B(n61), .Z(n738) );
  NAND U216 ( .A(n660), .B(n661), .Z(n62) );
  XOR U217 ( .A(n660), .B(n661), .Z(n63) );
  NANDN U218 ( .A(n659), .B(n63), .Z(n64) );
  NAND U219 ( .A(n62), .B(n64), .Z(n685) );
  NAND U220 ( .A(n691), .B(n693), .Z(n65) );
  XOR U221 ( .A(n691), .B(n693), .Z(n66) );
  NAND U222 ( .A(n66), .B(n692), .Z(n67) );
  NAND U223 ( .A(n65), .B(n67), .Z(n766) );
  XOR U224 ( .A(n535), .B(n534), .Z(n68) );
  XNOR U225 ( .A(n536), .B(n68), .Z(n554) );
  XNOR U226 ( .A(n754), .B(n753), .Z(n755) );
  NAND U227 ( .A(n524), .B(n525), .Z(n69) );
  XOR U228 ( .A(n524), .B(n525), .Z(n70) );
  NANDN U229 ( .A(n523), .B(n70), .Z(n71) );
  NAND U230 ( .A(n69), .B(n71), .Z(n563) );
  NAND U231 ( .A(n566), .B(n568), .Z(n72) );
  XOR U232 ( .A(n566), .B(n568), .Z(n73) );
  NAND U233 ( .A(n73), .B(n567), .Z(n74) );
  NAND U234 ( .A(n72), .B(n74), .Z(n675) );
  NANDN U235 ( .A(n680), .B(n683), .Z(n75) );
  OR U236 ( .A(n683), .B(n682), .Z(n76) );
  NANDN U237 ( .A(n681), .B(n76), .Z(n77) );
  NAND U238 ( .A(n75), .B(n77), .Z(n750) );
  XOR U239 ( .A(oglobal[4]), .B(n786), .Z(n78) );
  NAND U240 ( .A(n78), .B(n785), .Z(n79) );
  NAND U241 ( .A(oglobal[4]), .B(n786), .Z(n80) );
  AND U242 ( .A(n79), .B(n80), .Z(n809) );
  XOR U243 ( .A(n423), .B(n422), .Z(n81) );
  XNOR U244 ( .A(n424), .B(n81), .Z(n528) );
  XNOR U245 ( .A(n336), .B(n335), .Z(n337) );
  XNOR U246 ( .A(n253), .B(n252), .Z(n254) );
  XNOR U247 ( .A(n500), .B(n499), .Z(n501) );
  XNOR U248 ( .A(n488), .B(n487), .Z(n489) );
  XNOR U249 ( .A(n601), .B(n602), .Z(n82) );
  XNOR U250 ( .A(n600), .B(n82), .Z(n583) );
  NAND U251 ( .A(n513), .B(n514), .Z(n83) );
  XOR U252 ( .A(n513), .B(n514), .Z(n84) );
  NANDN U253 ( .A(n512), .B(n84), .Z(n85) );
  NAND U254 ( .A(n83), .B(n85), .Z(n538) );
  NAND U255 ( .A(n544), .B(n545), .Z(n86) );
  XOR U256 ( .A(n544), .B(n545), .Z(n87) );
  NAND U257 ( .A(n87), .B(n543), .Z(n88) );
  NAND U258 ( .A(n86), .B(n88), .Z(n706) );
  XNOR U259 ( .A(n368), .B(n367), .Z(n369) );
  XNOR U260 ( .A(n460), .B(n459), .Z(n461) );
  XNOR U261 ( .A(n774), .B(n773), .Z(n767) );
  NAND U262 ( .A(n722), .B(n723), .Z(n89) );
  XOR U263 ( .A(n722), .B(n723), .Z(n90) );
  NANDN U264 ( .A(n721), .B(n90), .Z(n91) );
  NAND U265 ( .A(n89), .B(n91), .Z(n763) );
  XOR U266 ( .A(n619), .B(n618), .Z(n660) );
  XOR U267 ( .A(n728), .B(n729), .Z(n92) );
  XNOR U268 ( .A(n730), .B(n92), .Z(n682) );
  XNOR U269 ( .A(n656), .B(n657), .Z(n93) );
  XNOR U270 ( .A(n658), .B(n93), .Z(n566) );
  NAND U271 ( .A(n564), .B(n565), .Z(n94) );
  XOR U272 ( .A(n564), .B(n565), .Z(n95) );
  NANDN U273 ( .A(n563), .B(n95), .Z(n96) );
  NAND U274 ( .A(n94), .B(n96), .Z(n677) );
  NAND U275 ( .A(n671), .B(n672), .Z(n97) );
  XOR U276 ( .A(n671), .B(n672), .Z(n98) );
  NANDN U277 ( .A(n670), .B(n98), .Z(n99) );
  NAND U278 ( .A(n97), .B(n99), .Z(n751) );
  XNOR U279 ( .A(n797), .B(n796), .Z(n801) );
  NAND U280 ( .A(n528), .B(n529), .Z(n100) );
  XOR U281 ( .A(n528), .B(n529), .Z(n101) );
  NANDN U282 ( .A(n527), .B(n101), .Z(n102) );
  NAND U283 ( .A(n100), .B(n102), .Z(n531) );
  XOR U284 ( .A(n809), .B(n808), .Z(n103) );
  NANDN U285 ( .A(oglobal[5]), .B(n103), .Z(n104) );
  NAND U286 ( .A(n809), .B(n808), .Z(n105) );
  AND U287 ( .A(n104), .B(n105), .Z(n818) );
  XNOR U288 ( .A(n259), .B(n258), .Z(n260) );
  XNOR U289 ( .A(n362), .B(n361), .Z(n363) );
  XNOR U290 ( .A(n494), .B(n493), .Z(n495) );
  XOR U291 ( .A(n581), .B(n582), .Z(n106) );
  XNOR U292 ( .A(n583), .B(n106), .Z(n539) );
  NAND U293 ( .A(n181), .B(n182), .Z(n107) );
  XOR U294 ( .A(n181), .B(n182), .Z(n108) );
  NANDN U295 ( .A(n180), .B(n108), .Z(n109) );
  NAND U296 ( .A(n107), .B(n109), .Z(n589) );
  NAND U297 ( .A(n266), .B(n267), .Z(n110) );
  XOR U298 ( .A(n266), .B(n267), .Z(n111) );
  NANDN U299 ( .A(n265), .B(n111), .Z(n112) );
  NAND U300 ( .A(n110), .B(n112), .Z(n617) );
  NAND U301 ( .A(n636), .B(n637), .Z(n113) );
  XOR U302 ( .A(n636), .B(n637), .Z(n114) );
  NANDN U303 ( .A(n635), .B(n114), .Z(n115) );
  NAND U304 ( .A(n113), .B(n115), .Z(n695) );
  NAND U305 ( .A(n623), .B(n624), .Z(n116) );
  XOR U306 ( .A(n623), .B(n624), .Z(n117) );
  NANDN U307 ( .A(n622), .B(n117), .Z(n118) );
  NAND U308 ( .A(n116), .B(n118), .Z(n691) );
  NAND U309 ( .A(n541), .B(n542), .Z(n119) );
  XOR U310 ( .A(n541), .B(n542), .Z(n120) );
  NANDN U311 ( .A(n540), .B(n120), .Z(n121) );
  NAND U312 ( .A(n119), .B(n121), .Z(n708) );
  NAND U313 ( .A(n548), .B(n549), .Z(n122) );
  XOR U314 ( .A(n548), .B(n549), .Z(n123) );
  NANDN U315 ( .A(n547), .B(n123), .Z(n124) );
  NAND U316 ( .A(n122), .B(n124), .Z(n701) );
  NAND U317 ( .A(n601), .B(n602), .Z(n125) );
  XOR U318 ( .A(n601), .B(n602), .Z(n126) );
  NANDN U319 ( .A(n600), .B(n126), .Z(n127) );
  NAND U320 ( .A(n125), .B(n127), .Z(n718) );
  XNOR U321 ( .A(n356), .B(n355), .Z(n357) );
  NAND U322 ( .A(n315), .B(n316), .Z(n128) );
  XOR U323 ( .A(n315), .B(n316), .Z(n129) );
  NANDN U324 ( .A(n314), .B(n129), .Z(n130) );
  NAND U325 ( .A(n128), .B(n130), .Z(n571) );
  XOR U326 ( .A(n632), .B(n631), .Z(n131) );
  XNOR U327 ( .A(n633), .B(n131), .Z(n651) );
  NANDN U328 ( .A(n519), .B(n522), .Z(n132) );
  OR U329 ( .A(n522), .B(n521), .Z(n133) );
  NANDN U330 ( .A(n520), .B(n133), .Z(n134) );
  NAND U331 ( .A(n132), .B(n134), .Z(n557) );
  NAND U332 ( .A(n423), .B(n424), .Z(n135) );
  XOR U333 ( .A(n423), .B(n424), .Z(n136) );
  NANDN U334 ( .A(n422), .B(n136), .Z(n137) );
  NAND U335 ( .A(n135), .B(n137), .Z(n552) );
  NAND U336 ( .A(n712), .B(n714), .Z(n138) );
  XOR U337 ( .A(n712), .B(n714), .Z(n139) );
  NAND U338 ( .A(n139), .B(n713), .Z(n140) );
  NAND U339 ( .A(n138), .B(n140), .Z(n772) );
  XOR U340 ( .A(n515), .B(n516), .Z(n141) );
  XNOR U341 ( .A(n517), .B(n141), .Z(n427) );
  XNOR U342 ( .A(n507), .B(n506), .Z(n142) );
  XNOR U343 ( .A(n509), .B(n142), .Z(n375) );
  NAND U344 ( .A(n762), .B(n764), .Z(n143) );
  XOR U345 ( .A(n762), .B(n764), .Z(n144) );
  NAND U346 ( .A(n144), .B(n763), .Z(n145) );
  NAND U347 ( .A(n143), .B(n145), .Z(n788) );
  XOR U348 ( .A(n467), .B(n466), .Z(n146) );
  XNOR U349 ( .A(n468), .B(n146), .Z(n525) );
  XNOR U350 ( .A(n756), .B(n755), .Z(n744) );
  NAND U351 ( .A(n759), .B(n761), .Z(n147) );
  XOR U352 ( .A(n759), .B(n761), .Z(n148) );
  NAND U353 ( .A(n148), .B(n760), .Z(n149) );
  NAND U354 ( .A(n147), .B(n149), .Z(n795) );
  NAND U355 ( .A(n532), .B(n533), .Z(n150) );
  XOR U356 ( .A(n532), .B(n533), .Z(n151) );
  NANDN U357 ( .A(n531), .B(n151), .Z(n152) );
  NAND U358 ( .A(n150), .B(n152), .Z(n665) );
  NAND U359 ( .A(n751), .B(n752), .Z(n153) );
  XOR U360 ( .A(n751), .B(n752), .Z(n154) );
  NANDN U361 ( .A(n750), .B(n154), .Z(n155) );
  NAND U362 ( .A(n153), .B(n155), .Z(n804) );
  XOR U363 ( .A(oglobal[6]), .B(n818), .Z(n156) );
  NANDN U364 ( .A(n819), .B(n156), .Z(n157) );
  NAND U365 ( .A(oglobal[6]), .B(n818), .Z(n158) );
  AND U366 ( .A(n157), .B(n158), .Z(n820) );
  NAND U367 ( .A(n825), .B(oglobal[12]), .Z(n159) );
  XNOR U368 ( .A(oglobal[13]), .B(n159), .Z(o[13]) );
  XOR U369 ( .A(x[11]), .B(y[11]), .Z(n370) );
  XOR U370 ( .A(x[15]), .B(y[15]), .Z(n367) );
  XNOR U371 ( .A(x[13]), .B(y[13]), .Z(n368) );
  XOR U372 ( .A(n370), .B(n369), .Z(n175) );
  XOR U373 ( .A(x[17]), .B(y[17]), .Z(n358) );
  XOR U374 ( .A(x[21]), .B(y[21]), .Z(n355) );
  XNOR U375 ( .A(x[19]), .B(y[19]), .Z(n356) );
  XOR U376 ( .A(n358), .B(n357), .Z(n177) );
  XOR U377 ( .A(x[5]), .B(y[5]), .Z(n332) );
  XOR U378 ( .A(x[9]), .B(y[9]), .Z(n330) );
  XOR U379 ( .A(x[7]), .B(y[7]), .Z(n329) );
  XOR U380 ( .A(n330), .B(n329), .Z(n331) );
  XNOR U381 ( .A(n332), .B(n331), .Z(n174) );
  XOR U382 ( .A(n177), .B(n174), .Z(n160) );
  XOR U383 ( .A(n175), .B(n160), .Z(n522) );
  XOR U384 ( .A(x[77]), .B(y[77]), .Z(n261) );
  XOR U385 ( .A(x[81]), .B(y[81]), .Z(n258) );
  XNOR U386 ( .A(x[79]), .B(y[79]), .Z(n259) );
  XOR U387 ( .A(n261), .B(n260), .Z(n184) );
  XOR U388 ( .A(x[83]), .B(y[83]), .Z(n412) );
  XOR U389 ( .A(x[85]), .B(y[85]), .Z(n410) );
  XOR U390 ( .A(x[87]), .B(y[87]), .Z(n409) );
  XOR U391 ( .A(n410), .B(n409), .Z(n411) );
  XOR U392 ( .A(n412), .B(n411), .Z(n186) );
  XOR U393 ( .A(x[115]), .B(y[115]), .Z(n484) );
  XNOR U394 ( .A(x[119]), .B(y[119]), .Z(n482) );
  XNOR U395 ( .A(n484), .B(n483), .Z(n183) );
  XOR U396 ( .A(n186), .B(n183), .Z(n161) );
  XOR U397 ( .A(n184), .B(n161), .Z(n291) );
  XOR U398 ( .A(x[107]), .B(y[107]), .Z(n338) );
  XOR U399 ( .A(x[111]), .B(y[111]), .Z(n335) );
  XNOR U400 ( .A(x[109]), .B(y[109]), .Z(n336) );
  XNOR U401 ( .A(n338), .B(n337), .Z(n290) );
  XOR U402 ( .A(x[101]), .B(y[101]), .Z(n364) );
  XOR U403 ( .A(x[105]), .B(y[105]), .Z(n361) );
  XNOR U404 ( .A(x[103]), .B(y[103]), .Z(n362) );
  XNOR U405 ( .A(n364), .B(n363), .Z(n289) );
  XOR U406 ( .A(n290), .B(n289), .Z(n292) );
  XOR U407 ( .A(n291), .B(n292), .Z(n521) );
  IV U408 ( .A(n521), .Z(n519) );
  XOR U409 ( .A(x[53]), .B(y[53]), .Z(n406) );
  XOR U410 ( .A(x[57]), .B(y[57]), .Z(n404) );
  XOR U411 ( .A(x[55]), .B(y[55]), .Z(n403) );
  XOR U412 ( .A(n404), .B(n403), .Z(n405) );
  XNOR U413 ( .A(n406), .B(n405), .Z(n514) );
  XOR U414 ( .A(x[41]), .B(y[41]), .Z(n387) );
  XOR U415 ( .A(x[45]), .B(y[45]), .Z(n385) );
  XOR U416 ( .A(x[43]), .B(y[43]), .Z(n384) );
  XOR U417 ( .A(n385), .B(n384), .Z(n386) );
  XNOR U418 ( .A(n387), .B(n386), .Z(n513) );
  XOR U419 ( .A(x[47]), .B(y[47]), .Z(n418) );
  XOR U420 ( .A(x[51]), .B(y[51]), .Z(n416) );
  XOR U421 ( .A(x[49]), .B(y[49]), .Z(n415) );
  XOR U422 ( .A(n416), .B(n415), .Z(n417) );
  XOR U423 ( .A(n418), .B(n417), .Z(n512) );
  XOR U424 ( .A(n513), .B(n512), .Z(n162) );
  XOR U425 ( .A(n514), .B(n162), .Z(n520) );
  XOR U426 ( .A(n519), .B(n520), .Z(n163) );
  XNOR U427 ( .A(n522), .B(n163), .Z(n529) );
  XOR U428 ( .A(x[60]), .B(y[60]), .Z(n211) );
  XOR U429 ( .A(x[58]), .B(y[58]), .Z(n208) );
  XOR U430 ( .A(x[56]), .B(y[56]), .Z(n209) );
  XOR U431 ( .A(n208), .B(n209), .Z(n210) );
  XOR U432 ( .A(n211), .B(n210), .Z(n345) );
  XOR U433 ( .A(x[66]), .B(y[66]), .Z(n431) );
  XOR U434 ( .A(x[64]), .B(y[64]), .Z(n429) );
  XOR U435 ( .A(x[62]), .B(y[62]), .Z(n428) );
  XOR U436 ( .A(n429), .B(n428), .Z(n430) );
  XNOR U437 ( .A(n431), .B(n430), .Z(n343) );
  XOR U438 ( .A(x[54]), .B(y[54]), .Z(n223) );
  XOR U439 ( .A(x[52]), .B(y[52]), .Z(n220) );
  XOR U440 ( .A(x[50]), .B(y[50]), .Z(n221) );
  XOR U441 ( .A(n220), .B(n221), .Z(n222) );
  XOR U442 ( .A(n223), .B(n222), .Z(n344) );
  XOR U443 ( .A(n343), .B(n344), .Z(n164) );
  XOR U444 ( .A(n345), .B(n164), .Z(n422) );
  XOR U445 ( .A(x[82]), .B(y[82]), .Z(n236) );
  XOR U446 ( .A(x[118]), .B(y[118]), .Z(n233) );
  XOR U447 ( .A(x[80]), .B(y[80]), .Z(n234) );
  XOR U448 ( .A(n233), .B(n234), .Z(n235) );
  XNOR U449 ( .A(n236), .B(n235), .Z(n349) );
  XOR U450 ( .A(x[98]), .B(y[98]), .Z(n277) );
  XOR U451 ( .A(x[110]), .B(y[110]), .Z(n274) );
  XOR U452 ( .A(x[96]), .B(y[96]), .Z(n275) );
  XOR U453 ( .A(n274), .B(n275), .Z(n276) );
  XOR U454 ( .A(n277), .B(n276), .Z(n450) );
  XOR U455 ( .A(x[106]), .B(y[106]), .Z(n448) );
  XOR U456 ( .A(x[104]), .B(y[104]), .Z(n447) );
  XOR U457 ( .A(n448), .B(n447), .Z(n449) );
  XOR U458 ( .A(n450), .B(n449), .Z(n352) );
  XOR U459 ( .A(x[90]), .B(y[90]), .Z(n456) );
  XOR U460 ( .A(x[114]), .B(y[114]), .Z(n454) );
  XOR U461 ( .A(x[88]), .B(y[88]), .Z(n453) );
  XOR U462 ( .A(n454), .B(n453), .Z(n455) );
  XNOR U463 ( .A(n456), .B(n455), .Z(n350) );
  XOR U464 ( .A(n352), .B(n350), .Z(n165) );
  XOR U465 ( .A(n349), .B(n165), .Z(n424) );
  XOR U466 ( .A(x[74]), .B(y[74]), .Z(n443) );
  XOR U467 ( .A(x[122]), .B(y[122]), .Z(n441) );
  XOR U468 ( .A(x[72]), .B(y[72]), .Z(n440) );
  XOR U469 ( .A(n441), .B(n440), .Z(n442) );
  XNOR U470 ( .A(n443), .B(n442), .Z(n283) );
  XOR U471 ( .A(x[70]), .B(y[70]), .Z(n437) );
  XOR U472 ( .A(x[124]), .B(y[124]), .Z(n435) );
  XOR U473 ( .A(x[68]), .B(y[68]), .Z(n434) );
  XOR U474 ( .A(n435), .B(n434), .Z(n436) );
  XOR U475 ( .A(n437), .B(n436), .Z(n286) );
  XOR U476 ( .A(x[78]), .B(y[78]), .Z(n230) );
  XOR U477 ( .A(x[120]), .B(y[120]), .Z(n227) );
  XOR U478 ( .A(x[76]), .B(y[76]), .Z(n228) );
  XOR U479 ( .A(n227), .B(n228), .Z(n229) );
  XNOR U480 ( .A(n230), .B(n229), .Z(n284) );
  XOR U481 ( .A(n286), .B(n284), .Z(n166) );
  XOR U482 ( .A(n283), .B(n166), .Z(n423) );
  XOR U483 ( .A(x[94]), .B(y[94]), .Z(n462) );
  XOR U484 ( .A(x[112]), .B(y[112]), .Z(n459) );
  XNOR U485 ( .A(x[92]), .B(y[92]), .Z(n460) );
  XNOR U486 ( .A(n462), .B(n461), .Z(n466) );
  XOR U487 ( .A(x[86]), .B(y[86]), .Z(n242) );
  XOR U488 ( .A(x[116]), .B(y[116]), .Z(n239) );
  XOR U489 ( .A(x[84]), .B(y[84]), .Z(n240) );
  XOR U490 ( .A(n239), .B(n240), .Z(n241) );
  XOR U491 ( .A(n242), .B(n241), .Z(n468) );
  XOR U492 ( .A(x[102]), .B(y[102]), .Z(n271) );
  XOR U493 ( .A(x[108]), .B(y[108]), .Z(n268) );
  XOR U494 ( .A(x[100]), .B(y[100]), .Z(n269) );
  XOR U495 ( .A(n268), .B(n269), .Z(n270) );
  XOR U496 ( .A(n271), .B(n270), .Z(n467) );
  XOR U497 ( .A(x[36]), .B(y[36]), .Z(n502) );
  XOR U498 ( .A(x[34]), .B(y[34]), .Z(n499) );
  XNOR U499 ( .A(x[32]), .B(y[32]), .Z(n500) );
  XOR U500 ( .A(n502), .B(n501), .Z(n316) );
  XOR U501 ( .A(x[42]), .B(y[42]), .Z(n490) );
  XOR U502 ( .A(x[40]), .B(y[40]), .Z(n487) );
  XNOR U503 ( .A(x[38]), .B(y[38]), .Z(n488) );
  XNOR U504 ( .A(n490), .B(n489), .Z(n314) );
  XOR U505 ( .A(x[48]), .B(y[48]), .Z(n217) );
  XOR U506 ( .A(x[46]), .B(y[46]), .Z(n214) );
  XOR U507 ( .A(x[44]), .B(y[44]), .Z(n215) );
  XOR U508 ( .A(n214), .B(n215), .Z(n216) );
  XOR U509 ( .A(n217), .B(n216), .Z(n315) );
  XOR U510 ( .A(n314), .B(n315), .Z(n167) );
  XOR U511 ( .A(n316), .B(n167), .Z(n376) );
  XOR U512 ( .A(x[6]), .B(y[6]), .Z(n192) );
  XOR U513 ( .A(x[4]), .B(y[4]), .Z(n189) );
  XOR U514 ( .A(x[2]), .B(y[2]), .Z(n190) );
  XOR U515 ( .A(n189), .B(n190), .Z(n191) );
  XNOR U516 ( .A(n192), .B(n191), .Z(n506) );
  XOR U517 ( .A(x[0]), .B(y[0]), .Z(n326) );
  XOR U518 ( .A(x[3]), .B(y[3]), .Z(n324) );
  XOR U519 ( .A(x[1]), .B(y[1]), .Z(n323) );
  XOR U520 ( .A(n324), .B(n323), .Z(n325) );
  XOR U521 ( .A(n326), .B(n325), .Z(n509) );
  XOR U522 ( .A(x[12]), .B(y[12]), .Z(n204) );
  XOR U523 ( .A(x[10]), .B(y[10]), .Z(n201) );
  XOR U524 ( .A(x[8]), .B(y[8]), .Z(n202) );
  XOR U525 ( .A(n201), .B(n202), .Z(n203) );
  XOR U526 ( .A(n204), .B(n203), .Z(n507) );
  XOR U527 ( .A(x[18]), .B(y[18]), .Z(n479) );
  XOR U528 ( .A(x[16]), .B(y[16]), .Z(n476) );
  XNOR U529 ( .A(x[14]), .B(y[14]), .Z(n477) );
  XOR U530 ( .A(n479), .B(n478), .Z(n319) );
  XOR U531 ( .A(x[24]), .B(y[24]), .Z(n473) );
  XOR U532 ( .A(x[22]), .B(y[22]), .Z(n470) );
  XNOR U533 ( .A(x[20]), .B(y[20]), .Z(n471) );
  XNOR U534 ( .A(n473), .B(n472), .Z(n317) );
  XOR U535 ( .A(x[30]), .B(y[30]), .Z(n496) );
  XOR U536 ( .A(x[28]), .B(y[28]), .Z(n493) );
  XNOR U537 ( .A(x[26]), .B(y[26]), .Z(n494) );
  XOR U538 ( .A(n496), .B(n495), .Z(n318) );
  XOR U539 ( .A(n317), .B(n318), .Z(n168) );
  XNOR U540 ( .A(n319), .B(n168), .Z(n374) );
  XOR U541 ( .A(n375), .B(n374), .Z(n169) );
  XOR U542 ( .A(n376), .B(n169), .Z(n524) );
  XOR U543 ( .A(x[35]), .B(y[35]), .Z(n399) );
  XOR U544 ( .A(x[39]), .B(y[39]), .Z(n397) );
  XOR U545 ( .A(x[37]), .B(y[37]), .Z(n396) );
  XOR U546 ( .A(n397), .B(n396), .Z(n398) );
  XOR U547 ( .A(n399), .B(n398), .Z(n517) );
  XOR U548 ( .A(x[23]), .B(y[23]), .Z(n298) );
  XOR U549 ( .A(x[27]), .B(y[27]), .Z(n296) );
  XOR U550 ( .A(x[25]), .B(y[25]), .Z(n295) );
  XOR U551 ( .A(n296), .B(n295), .Z(n297) );
  XNOR U552 ( .A(n298), .B(n297), .Z(n516) );
  XOR U553 ( .A(x[29]), .B(y[29]), .Z(n304) );
  XOR U554 ( .A(x[33]), .B(y[33]), .Z(n302) );
  XOR U555 ( .A(x[31]), .B(y[31]), .Z(n301) );
  XOR U556 ( .A(n302), .B(n301), .Z(n303) );
  XOR U557 ( .A(n304), .B(n303), .Z(n515) );
  XOR U558 ( .A(x[71]), .B(y[71]), .Z(n381) );
  XOR U559 ( .A(x[75]), .B(y[75]), .Z(n379) );
  XOR U560 ( .A(x[73]), .B(y[73]), .Z(n378) );
  XOR U561 ( .A(n379), .B(n378), .Z(n380) );
  XOR U562 ( .A(n381), .B(n380), .Z(n182) );
  XOR U563 ( .A(x[59]), .B(y[59]), .Z(n255) );
  XOR U564 ( .A(x[63]), .B(y[63]), .Z(n252) );
  XNOR U565 ( .A(x[61]), .B(y[61]), .Z(n253) );
  XNOR U566 ( .A(n255), .B(n254), .Z(n180) );
  XOR U567 ( .A(x[65]), .B(y[65]), .Z(n249) );
  XOR U568 ( .A(x[69]), .B(y[69]), .Z(n246) );
  XNOR U569 ( .A(x[67]), .B(y[67]), .Z(n247) );
  XOR U570 ( .A(n249), .B(n248), .Z(n181) );
  XOR U571 ( .A(n180), .B(n181), .Z(n170) );
  XOR U572 ( .A(n182), .B(n170), .Z(n425) );
  XOR U573 ( .A(x[95]), .B(y[95]), .Z(n310) );
  XOR U574 ( .A(x[97]), .B(y[97]), .Z(n308) );
  XOR U575 ( .A(x[99]), .B(y[99]), .Z(n307) );
  XOR U576 ( .A(n308), .B(n307), .Z(n309) );
  XNOR U577 ( .A(n310), .B(n309), .Z(n267) );
  XOR U578 ( .A(x[89]), .B(y[89]), .Z(n393) );
  XOR U579 ( .A(x[91]), .B(y[91]), .Z(n391) );
  XOR U580 ( .A(x[93]), .B(y[93]), .Z(n390) );
  XOR U581 ( .A(n391), .B(n390), .Z(n392) );
  XNOR U582 ( .A(n393), .B(n392), .Z(n266) );
  XOR U583 ( .A(x[123]), .B(y[123]), .Z(n281) );
  XOR U584 ( .A(x[121]), .B(y[121]), .Z(n280) );
  XOR U585 ( .A(n281), .B(n280), .Z(n198) );
  XOR U586 ( .A(x[113]), .B(y[113]), .Z(n195) );
  XOR U587 ( .A(x[117]), .B(y[117]), .Z(n196) );
  XOR U588 ( .A(n195), .B(n196), .Z(n197) );
  XOR U589 ( .A(n198), .B(n197), .Z(n265) );
  XOR U590 ( .A(n266), .B(n265), .Z(n171) );
  XOR U591 ( .A(n267), .B(n171), .Z(n426) );
  XOR U592 ( .A(n425), .B(n426), .Z(n172) );
  XOR U593 ( .A(n427), .B(n172), .Z(n523) );
  XOR U594 ( .A(n528), .B(n527), .Z(n173) );
  XNOR U595 ( .A(n529), .B(n173), .Z(o[0]) );
  NANDN U596 ( .A(n175), .B(n174), .Z(n179) );
  ANDN U597 ( .B(n175), .A(n174), .Z(n176) );
  OR U598 ( .A(n177), .B(n176), .Z(n178) );
  AND U599 ( .A(n179), .B(n178), .Z(n591) );
  NANDN U600 ( .A(n184), .B(n183), .Z(n188) );
  ANDN U601 ( .B(n184), .A(n183), .Z(n185) );
  OR U602 ( .A(n186), .B(n185), .Z(n187) );
  AND U603 ( .A(n188), .B(n187), .Z(n588) );
  XOR U604 ( .A(n589), .B(n588), .Z(n590) );
  XOR U605 ( .A(n591), .B(n590), .Z(n659) );
  NAND U606 ( .A(n190), .B(n189), .Z(n194) );
  NAND U607 ( .A(n192), .B(n191), .Z(n193) );
  NAND U608 ( .A(n194), .B(n193), .Z(n549) );
  NAND U609 ( .A(n196), .B(n195), .Z(n200) );
  NAND U610 ( .A(n198), .B(n197), .Z(n199) );
  NAND U611 ( .A(n200), .B(n199), .Z(n548) );
  NAND U612 ( .A(n202), .B(n201), .Z(n206) );
  NAND U613 ( .A(n204), .B(n203), .Z(n205) );
  AND U614 ( .A(n206), .B(n205), .Z(n547) );
  XOR U615 ( .A(n548), .B(n547), .Z(n207) );
  XNOR U616 ( .A(n549), .B(n207), .Z(n610) );
  NAND U617 ( .A(n209), .B(n208), .Z(n213) );
  NAND U618 ( .A(n211), .B(n210), .Z(n212) );
  NAND U619 ( .A(n213), .B(n212), .Z(n603) );
  NAND U620 ( .A(n215), .B(n214), .Z(n219) );
  NAND U621 ( .A(n217), .B(n216), .Z(n218) );
  AND U622 ( .A(n219), .B(n218), .Z(n605) );
  NAND U623 ( .A(n221), .B(n220), .Z(n225) );
  NAND U624 ( .A(n223), .B(n222), .Z(n224) );
  AND U625 ( .A(n225), .B(n224), .Z(n604) );
  XNOR U626 ( .A(n605), .B(n604), .Z(n226) );
  XOR U627 ( .A(n603), .B(n226), .Z(n613) );
  NAND U628 ( .A(n228), .B(n227), .Z(n232) );
  NAND U629 ( .A(n230), .B(n229), .Z(n231) );
  NAND U630 ( .A(n232), .B(n231), .Z(n640) );
  NAND U631 ( .A(n234), .B(n233), .Z(n238) );
  NAND U632 ( .A(n236), .B(n235), .Z(n237) );
  NAND U633 ( .A(n238), .B(n237), .Z(n639) );
  NAND U634 ( .A(n240), .B(n239), .Z(n244) );
  NAND U635 ( .A(n242), .B(n241), .Z(n243) );
  AND U636 ( .A(n244), .B(n243), .Z(n638) );
  XOR U637 ( .A(n639), .B(n638), .Z(n245) );
  XOR U638 ( .A(n640), .B(n245), .Z(n611) );
  NANDN U639 ( .A(n247), .B(n246), .Z(n251) );
  NAND U640 ( .A(n249), .B(n248), .Z(n250) );
  NAND U641 ( .A(n251), .B(n250), .Z(n646) );
  NANDN U642 ( .A(n253), .B(n252), .Z(n257) );
  NAND U643 ( .A(n255), .B(n254), .Z(n256) );
  NAND U644 ( .A(n257), .B(n256), .Z(n645) );
  NANDN U645 ( .A(n259), .B(n258), .Z(n263) );
  NAND U646 ( .A(n261), .B(n260), .Z(n262) );
  AND U647 ( .A(n263), .B(n262), .Z(n644) );
  XOR U648 ( .A(n645), .B(n644), .Z(n264) );
  XNOR U649 ( .A(n646), .B(n264), .Z(n618) );
  NAND U650 ( .A(n269), .B(n268), .Z(n273) );
  NAND U651 ( .A(n271), .B(n270), .Z(n272) );
  NAND U652 ( .A(n273), .B(n272), .Z(n545) );
  NAND U653 ( .A(n275), .B(n274), .Z(n279) );
  NAND U654 ( .A(n277), .B(n276), .Z(n278) );
  NAND U655 ( .A(n279), .B(n278), .Z(n543) );
  AND U656 ( .A(n281), .B(n280), .Z(n546) );
  XOR U657 ( .A(oglobal[1]), .B(n546), .Z(n544) );
  XOR U658 ( .A(n543), .B(n544), .Z(n282) );
  XOR U659 ( .A(n545), .B(n282), .Z(n616) );
  XOR U660 ( .A(n617), .B(n616), .Z(n619) );
  NAND U661 ( .A(n284), .B(n283), .Z(n288) );
  NOR U662 ( .A(n284), .B(n283), .Z(n285) );
  OR U663 ( .A(n286), .B(n285), .Z(n287) );
  AND U664 ( .A(n288), .B(n287), .Z(n652) );
  NAND U665 ( .A(n290), .B(n289), .Z(n294) );
  NAND U666 ( .A(n292), .B(n291), .Z(n293) );
  AND U667 ( .A(n294), .B(n293), .Z(n653) );
  NAND U668 ( .A(n296), .B(n295), .Z(n300) );
  NAND U669 ( .A(n298), .B(n297), .Z(n299) );
  AND U670 ( .A(n300), .B(n299), .Z(n631) );
  NAND U671 ( .A(n302), .B(n301), .Z(n306) );
  NAND U672 ( .A(n304), .B(n303), .Z(n305) );
  NAND U673 ( .A(n306), .B(n305), .Z(n633) );
  NAND U674 ( .A(n308), .B(n307), .Z(n312) );
  NAND U675 ( .A(n310), .B(n309), .Z(n311) );
  NAND U676 ( .A(n312), .B(n311), .Z(n632) );
  XOR U677 ( .A(n653), .B(n651), .Z(n313) );
  XOR U678 ( .A(n652), .B(n313), .Z(n658) );
  NANDN U679 ( .A(n318), .B(n317), .Z(n322) );
  ANDN U680 ( .B(n318), .A(n317), .Z(n320) );
  OR U681 ( .A(n320), .B(n319), .Z(n321) );
  AND U682 ( .A(n322), .B(n321), .Z(n572) );
  NAND U683 ( .A(n324), .B(n323), .Z(n328) );
  NAND U684 ( .A(n326), .B(n325), .Z(n327) );
  AND U685 ( .A(n328), .B(n327), .Z(n540) );
  NAND U686 ( .A(n330), .B(n329), .Z(n334) );
  NAND U687 ( .A(n332), .B(n331), .Z(n333) );
  NAND U688 ( .A(n334), .B(n333), .Z(n542) );
  NANDN U689 ( .A(n336), .B(n335), .Z(n340) );
  NAND U690 ( .A(n338), .B(n337), .Z(n339) );
  NAND U691 ( .A(n340), .B(n339), .Z(n541) );
  XNOR U692 ( .A(n542), .B(n541), .Z(n341) );
  XOR U693 ( .A(n540), .B(n341), .Z(n570) );
  XOR U694 ( .A(n572), .B(n570), .Z(n342) );
  XOR U695 ( .A(n571), .B(n342), .Z(n656) );
  NANDN U696 ( .A(n344), .B(n343), .Z(n348) );
  ANDN U697 ( .B(n344), .A(n343), .Z(n346) );
  OR U698 ( .A(n346), .B(n345), .Z(n347) );
  AND U699 ( .A(n348), .B(n347), .Z(n595) );
  NAND U700 ( .A(n350), .B(n349), .Z(n354) );
  NOR U701 ( .A(n350), .B(n349), .Z(n351) );
  OR U702 ( .A(n352), .B(n351), .Z(n353) );
  AND U703 ( .A(n354), .B(n353), .Z(n594) );
  XOR U704 ( .A(n595), .B(n594), .Z(n597) );
  NANDN U705 ( .A(n356), .B(n355), .Z(n360) );
  NAND U706 ( .A(n358), .B(n357), .Z(n359) );
  NAND U707 ( .A(n360), .B(n359), .Z(n649) );
  NANDN U708 ( .A(n362), .B(n361), .Z(n366) );
  NAND U709 ( .A(n364), .B(n363), .Z(n365) );
  NAND U710 ( .A(n366), .B(n365), .Z(n648) );
  NANDN U711 ( .A(n368), .B(n367), .Z(n372) );
  NAND U712 ( .A(n370), .B(n369), .Z(n371) );
  AND U713 ( .A(n372), .B(n371), .Z(n647) );
  XOR U714 ( .A(n648), .B(n647), .Z(n373) );
  XOR U715 ( .A(n649), .B(n373), .Z(n596) );
  XOR U716 ( .A(n597), .B(n596), .Z(n657) );
  XOR U717 ( .A(n566), .B(n567), .Z(n377) );
  XOR U718 ( .A(n568), .B(n377), .Z(n532) );
  NAND U719 ( .A(n379), .B(n378), .Z(n383) );
  NAND U720 ( .A(n381), .B(n380), .Z(n382) );
  NAND U721 ( .A(n383), .B(n382), .Z(n534) );
  NAND U722 ( .A(n385), .B(n384), .Z(n389) );
  NAND U723 ( .A(n387), .B(n386), .Z(n388) );
  NAND U724 ( .A(n389), .B(n388), .Z(n627) );
  NAND U725 ( .A(n391), .B(n390), .Z(n395) );
  NAND U726 ( .A(n393), .B(n392), .Z(n394) );
  NAND U727 ( .A(n395), .B(n394), .Z(n626) );
  NAND U728 ( .A(n397), .B(n396), .Z(n401) );
  NAND U729 ( .A(n399), .B(n398), .Z(n400) );
  AND U730 ( .A(n401), .B(n400), .Z(n625) );
  XOR U731 ( .A(n626), .B(n625), .Z(n402) );
  XOR U732 ( .A(n627), .B(n402), .Z(n536) );
  NAND U733 ( .A(n404), .B(n403), .Z(n408) );
  NAND U734 ( .A(n406), .B(n405), .Z(n407) );
  NAND U735 ( .A(n408), .B(n407), .Z(n624) );
  NAND U736 ( .A(n410), .B(n409), .Z(n414) );
  NAND U737 ( .A(n412), .B(n411), .Z(n413) );
  NAND U738 ( .A(n414), .B(n413), .Z(n623) );
  NAND U739 ( .A(n416), .B(n415), .Z(n420) );
  NAND U740 ( .A(n418), .B(n417), .Z(n419) );
  AND U741 ( .A(n420), .B(n419), .Z(n622) );
  XOR U742 ( .A(n623), .B(n622), .Z(n421) );
  XOR U743 ( .A(n624), .B(n421), .Z(n535) );
  XOR U744 ( .A(n552), .B(n551), .Z(n553) );
  XOR U745 ( .A(n554), .B(n553), .Z(n564) );
  NAND U746 ( .A(n429), .B(n428), .Z(n433) );
  NAND U747 ( .A(n431), .B(n430), .Z(n432) );
  NAND U748 ( .A(n433), .B(n432), .Z(n637) );
  NAND U749 ( .A(n435), .B(n434), .Z(n439) );
  NAND U750 ( .A(n437), .B(n436), .Z(n438) );
  NAND U751 ( .A(n439), .B(n438), .Z(n636) );
  NAND U752 ( .A(n441), .B(n440), .Z(n445) );
  NAND U753 ( .A(n443), .B(n442), .Z(n444) );
  AND U754 ( .A(n445), .B(n444), .Z(n635) );
  XOR U755 ( .A(n636), .B(n635), .Z(n446) );
  XNOR U756 ( .A(n637), .B(n446), .Z(n576) );
  NAND U757 ( .A(n448), .B(n447), .Z(n452) );
  NAND U758 ( .A(n450), .B(n449), .Z(n451) );
  NAND U759 ( .A(n452), .B(n451), .Z(n643) );
  NAND U760 ( .A(n454), .B(n453), .Z(n458) );
  NAND U761 ( .A(n456), .B(n455), .Z(n457) );
  NAND U762 ( .A(n458), .B(n457), .Z(n642) );
  NANDN U763 ( .A(n460), .B(n459), .Z(n464) );
  NAND U764 ( .A(n462), .B(n461), .Z(n463) );
  AND U765 ( .A(n464), .B(n463), .Z(n641) );
  XOR U766 ( .A(n642), .B(n641), .Z(n465) );
  XOR U767 ( .A(n643), .B(n465), .Z(n574) );
  IV U768 ( .A(n574), .Z(n573) );
  XOR U769 ( .A(n573), .B(n575), .Z(n469) );
  XNOR U770 ( .A(n576), .B(n469), .Z(n560) );
  NANDN U771 ( .A(n471), .B(n470), .Z(n475) );
  NAND U772 ( .A(n473), .B(n472), .Z(n474) );
  NAND U773 ( .A(n475), .B(n474), .Z(n600) );
  NANDN U774 ( .A(n477), .B(n476), .Z(n481) );
  NAND U775 ( .A(n479), .B(n478), .Z(n480) );
  AND U776 ( .A(n481), .B(n480), .Z(n602) );
  NANDN U777 ( .A(n482), .B(oglobal[0]), .Z(n486) );
  NAND U778 ( .A(n484), .B(n483), .Z(n485) );
  AND U779 ( .A(n486), .B(n485), .Z(n601) );
  NANDN U780 ( .A(n488), .B(n487), .Z(n492) );
  NAND U781 ( .A(n490), .B(n489), .Z(n491) );
  NAND U782 ( .A(n492), .B(n491), .Z(n606) );
  NANDN U783 ( .A(n494), .B(n493), .Z(n498) );
  NAND U784 ( .A(n496), .B(n495), .Z(n497) );
  AND U785 ( .A(n498), .B(n497), .Z(n608) );
  NANDN U786 ( .A(n500), .B(n499), .Z(n504) );
  NAND U787 ( .A(n502), .B(n501), .Z(n503) );
  AND U788 ( .A(n504), .B(n503), .Z(n607) );
  XNOR U789 ( .A(n608), .B(n607), .Z(n505) );
  XOR U790 ( .A(n606), .B(n505), .Z(n580) );
  IV U791 ( .A(n580), .Z(n582) );
  NANDN U792 ( .A(n507), .B(n506), .Z(n511) );
  ANDN U793 ( .B(n507), .A(n506), .Z(n508) );
  OR U794 ( .A(n509), .B(n508), .Z(n510) );
  AND U795 ( .A(n511), .B(n510), .Z(n581) );
  XNOR U796 ( .A(n538), .B(n537), .Z(n518) );
  XNOR U797 ( .A(n539), .B(n518), .Z(n558) );
  XOR U798 ( .A(n558), .B(n557), .Z(n559) );
  XOR U799 ( .A(n560), .B(n559), .Z(n565) );
  XNOR U800 ( .A(n565), .B(n563), .Z(n526) );
  XOR U801 ( .A(n564), .B(n526), .Z(n533) );
  XNOR U802 ( .A(n533), .B(n531), .Z(n530) );
  XNOR U803 ( .A(n532), .B(n530), .Z(o[1]) );
  AND U804 ( .A(n546), .B(oglobal[1]), .Z(n700) );
  XOR U805 ( .A(oglobal[2]), .B(n700), .Z(n702) );
  XNOR U806 ( .A(n702), .B(n701), .Z(n705) );
  XNOR U807 ( .A(n706), .B(n705), .Z(n707) );
  XOR U808 ( .A(n708), .B(n707), .Z(n735) );
  XOR U809 ( .A(n738), .B(n735), .Z(n550) );
  XOR U810 ( .A(n736), .B(n550), .Z(n670) );
  OR U811 ( .A(n552), .B(n551), .Z(n556) );
  NAND U812 ( .A(n554), .B(n553), .Z(n555) );
  NAND U813 ( .A(n556), .B(n555), .Z(n672) );
  NAND U814 ( .A(n558), .B(n557), .Z(n562) );
  NAND U815 ( .A(n560), .B(n559), .Z(n561) );
  NAND U816 ( .A(n562), .B(n561), .Z(n671) );
  IV U817 ( .A(n673), .Z(n674) );
  XNOR U818 ( .A(n677), .B(n675), .Z(n569) );
  XOR U819 ( .A(n674), .B(n569), .Z(n667) );
  OR U820 ( .A(n575), .B(n573), .Z(n579) );
  ANDN U821 ( .B(n575), .A(n574), .Z(n577) );
  OR U822 ( .A(n577), .B(n576), .Z(n578) );
  AND U823 ( .A(n579), .B(n578), .Z(n726) );
  NANDN U824 ( .A(n580), .B(n581), .Z(n586) );
  NOR U825 ( .A(n582), .B(n581), .Z(n584) );
  NANDN U826 ( .A(n584), .B(n583), .Z(n585) );
  AND U827 ( .A(n586), .B(n585), .Z(n724) );
  XNOR U828 ( .A(n726), .B(n724), .Z(n587) );
  XOR U829 ( .A(n725), .B(n587), .Z(n683) );
  OR U830 ( .A(n589), .B(n588), .Z(n593) );
  NANDN U831 ( .A(n591), .B(n590), .Z(n592) );
  NAND U832 ( .A(n593), .B(n592), .Z(n733) );
  OR U833 ( .A(n595), .B(n594), .Z(n599) );
  NAND U834 ( .A(n597), .B(n596), .Z(n598) );
  NAND U835 ( .A(n599), .B(n598), .Z(n732) );
  XOR U836 ( .A(n716), .B(n715), .Z(n717) );
  XNOR U837 ( .A(n718), .B(n717), .Z(n731) );
  XOR U838 ( .A(n732), .B(n731), .Z(n609) );
  XOR U839 ( .A(n733), .B(n609), .Z(n730) );
  NANDN U840 ( .A(n611), .B(n610), .Z(n615) );
  ANDN U841 ( .B(n611), .A(n610), .Z(n612) );
  OR U842 ( .A(n613), .B(n612), .Z(n614) );
  AND U843 ( .A(n615), .B(n614), .Z(n729) );
  NANDN U844 ( .A(n617), .B(n616), .Z(n621) );
  NANDN U845 ( .A(n619), .B(n618), .Z(n620) );
  NAND U846 ( .A(n621), .B(n620), .Z(n728) );
  IV U847 ( .A(n682), .Z(n680) );
  NANDN U848 ( .A(n626), .B(n625), .Z(n630) );
  ANDN U849 ( .B(n626), .A(n625), .Z(n628) );
  OR U850 ( .A(n628), .B(n627), .Z(n629) );
  AND U851 ( .A(n630), .B(n629), .Z(n693) );
  XNOR U852 ( .A(n693), .B(n692), .Z(n634) );
  XOR U853 ( .A(n691), .B(n634), .Z(n696) );
  XOR U854 ( .A(n695), .B(n694), .Z(n697) );
  XNOR U855 ( .A(n696), .B(n697), .Z(n723) );
  XNOR U856 ( .A(n714), .B(n713), .Z(n650) );
  XOR U857 ( .A(n712), .B(n650), .Z(n721) );
  XOR U858 ( .A(n721), .B(n722), .Z(n654) );
  XOR U859 ( .A(n723), .B(n654), .Z(n681) );
  XOR U860 ( .A(n680), .B(n681), .Z(n655) );
  XOR U861 ( .A(n683), .B(n655), .Z(n688) );
  XOR U862 ( .A(n686), .B(n685), .Z(n687) );
  XOR U863 ( .A(n688), .B(n687), .Z(n664) );
  IV U864 ( .A(n664), .Z(n663) );
  XOR U865 ( .A(n667), .B(n663), .Z(n662) );
  XNOR U866 ( .A(n665), .B(n662), .Z(o[2]) );
  OR U867 ( .A(n665), .B(n663), .Z(n669) );
  ANDN U868 ( .B(n665), .A(n664), .Z(n666) );
  OR U869 ( .A(n667), .B(n666), .Z(n668) );
  AND U870 ( .A(n669), .B(n668), .Z(n745) );
  OR U871 ( .A(n675), .B(n673), .Z(n679) );
  ANDN U872 ( .B(n675), .A(n674), .Z(n676) );
  OR U873 ( .A(n677), .B(n676), .Z(n678) );
  AND U874 ( .A(n679), .B(n678), .Z(n752) );
  XOR U875 ( .A(n752), .B(n750), .Z(n684) );
  XNOR U876 ( .A(n751), .B(n684), .Z(n747) );
  OR U877 ( .A(n686), .B(n685), .Z(n690) );
  NAND U878 ( .A(n688), .B(n687), .Z(n689) );
  AND U879 ( .A(n690), .B(n689), .Z(n756) );
  OR U880 ( .A(n695), .B(n694), .Z(n699) );
  NAND U881 ( .A(n697), .B(n696), .Z(n698) );
  NAND U882 ( .A(n699), .B(n698), .Z(n765) );
  XNOR U883 ( .A(n766), .B(n765), .Z(n768) );
  AND U884 ( .A(oglobal[2]), .B(n700), .Z(n704) );
  NAND U885 ( .A(n702), .B(n701), .Z(n703) );
  NANDN U886 ( .A(n704), .B(n703), .Z(n779) );
  NANDN U887 ( .A(n706), .B(n705), .Z(n710) );
  NANDN U888 ( .A(n708), .B(n707), .Z(n709) );
  NAND U889 ( .A(n710), .B(n709), .Z(n778) );
  IV U890 ( .A(n778), .Z(n777) );
  XOR U891 ( .A(n779), .B(n777), .Z(n711) );
  XNOR U892 ( .A(oglobal[3]), .B(n711), .Z(n773) );
  OR U893 ( .A(n716), .B(n715), .Z(n720) );
  NANDN U894 ( .A(n718), .B(n717), .Z(n719) );
  AND U895 ( .A(n720), .B(n719), .Z(n771) );
  XOR U896 ( .A(n772), .B(n771), .Z(n774) );
  XNOR U897 ( .A(n768), .B(n767), .Z(n764) );
  XNOR U898 ( .A(n763), .B(n762), .Z(n727) );
  XOR U899 ( .A(n764), .B(n727), .Z(n754) );
  IV U900 ( .A(n735), .Z(n734) );
  OR U901 ( .A(n736), .B(n734), .Z(n740) );
  ANDN U902 ( .B(n736), .A(n735), .Z(n737) );
  OR U903 ( .A(n738), .B(n737), .Z(n739) );
  AND U904 ( .A(n740), .B(n739), .Z(n759) );
  XOR U905 ( .A(n760), .B(n759), .Z(n741) );
  XNOR U906 ( .A(n761), .B(n741), .Z(n753) );
  IV U907 ( .A(n744), .Z(n743) );
  XOR U908 ( .A(n747), .B(n743), .Z(n742) );
  XNOR U909 ( .A(n745), .B(n742), .Z(o[3]) );
  OR U910 ( .A(n745), .B(n743), .Z(n749) );
  ANDN U911 ( .B(n745), .A(n744), .Z(n746) );
  OR U912 ( .A(n747), .B(n746), .Z(n748) );
  AND U913 ( .A(n749), .B(n748), .Z(n802) );
  NANDN U914 ( .A(n754), .B(n753), .Z(n758) );
  NANDN U915 ( .A(n756), .B(n755), .Z(n757) );
  NAND U916 ( .A(n758), .B(n757), .Z(n796) );
  NANDN U917 ( .A(n766), .B(n765), .Z(n770) );
  NAND U918 ( .A(n768), .B(n767), .Z(n769) );
  NAND U919 ( .A(n770), .B(n769), .Z(n787) );
  XNOR U920 ( .A(n788), .B(n787), .Z(n790) );
  NANDN U921 ( .A(n772), .B(n771), .Z(n776) );
  NANDN U922 ( .A(n774), .B(n773), .Z(n775) );
  AND U923 ( .A(n776), .B(n775), .Z(n786) );
  OR U924 ( .A(oglobal[3]), .B(n777), .Z(n782) );
  ANDN U925 ( .B(oglobal[3]), .A(n778), .Z(n780) );
  OR U926 ( .A(n780), .B(n779), .Z(n781) );
  AND U927 ( .A(n782), .B(n781), .Z(n785) );
  XNOR U928 ( .A(oglobal[4]), .B(n785), .Z(n783) );
  XOR U929 ( .A(n786), .B(n783), .Z(n789) );
  XNOR U930 ( .A(n790), .B(n789), .Z(n794) );
  XOR U931 ( .A(n795), .B(n794), .Z(n797) );
  IV U932 ( .A(n801), .Z(n800) );
  XOR U933 ( .A(n804), .B(n800), .Z(n784) );
  XNOR U934 ( .A(n802), .B(n784), .Z(o[4]) );
  NANDN U935 ( .A(n788), .B(n787), .Z(n792) );
  NAND U936 ( .A(n790), .B(n789), .Z(n791) );
  NAND U937 ( .A(n792), .B(n791), .Z(n808) );
  XOR U938 ( .A(oglobal[5]), .B(n808), .Z(n793) );
  XOR U939 ( .A(n809), .B(n793), .Z(n811) );
  IV U940 ( .A(n811), .Z(n810) );
  NANDN U941 ( .A(n795), .B(n794), .Z(n799) );
  NANDN U942 ( .A(n797), .B(n796), .Z(n798) );
  AND U943 ( .A(n799), .B(n798), .Z(n814) );
  OR U944 ( .A(n802), .B(n800), .Z(n806) );
  ANDN U945 ( .B(n802), .A(n801), .Z(n803) );
  OR U946 ( .A(n804), .B(n803), .Z(n805) );
  AND U947 ( .A(n806), .B(n805), .Z(n812) );
  XNOR U948 ( .A(n814), .B(n812), .Z(n807) );
  XOR U949 ( .A(n810), .B(n807), .Z(o[5]) );
  OR U950 ( .A(n812), .B(n810), .Z(n816) );
  ANDN U951 ( .B(n812), .A(n811), .Z(n813) );
  OR U952 ( .A(n814), .B(n813), .Z(n815) );
  AND U953 ( .A(n816), .B(n815), .Z(n819) );
  XOR U954 ( .A(n818), .B(n819), .Z(n817) );
  XNOR U955 ( .A(oglobal[6]), .B(n817), .Z(o[6]) );
  XNOR U956 ( .A(n820), .B(oglobal[7]), .Z(o[7]) );
  ANDN U957 ( .B(oglobal[7]), .A(n820), .Z(n821) );
  XOR U958 ( .A(n821), .B(oglobal[8]), .Z(o[8]) );
  AND U959 ( .A(n821), .B(oglobal[8]), .Z(n822) );
  XOR U960 ( .A(n822), .B(oglobal[9]), .Z(o[9]) );
  AND U961 ( .A(n822), .B(oglobal[9]), .Z(n823) );
  XOR U962 ( .A(n823), .B(oglobal[10]), .Z(o[10]) );
  AND U963 ( .A(n823), .B(oglobal[10]), .Z(n824) );
  XOR U964 ( .A(n824), .B(oglobal[11]), .Z(o[11]) );
  AND U965 ( .A(n824), .B(oglobal[11]), .Z(n825) );
  XOR U966 ( .A(oglobal[12]), .B(n825), .Z(o[12]) );
endmodule

