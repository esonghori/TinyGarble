
module MUX_N512_3 ( A, B, S, O );
  input [511:0] A;
  input [511:0] B;
  output [511:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[511]), .B(n109), .Z(O[511]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[511]), .B(A[511]), .Z(n110) );
  XOR U166 ( .A(A[510]), .B(n111), .Z(O[510]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[510]), .B(A[510]), .Z(n112) );
  XOR U169 ( .A(A[50]), .B(n113), .Z(O[50]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[50]), .B(A[50]), .Z(n114) );
  XOR U172 ( .A(A[509]), .B(n115), .Z(O[509]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[509]), .B(A[509]), .Z(n116) );
  XOR U175 ( .A(A[508]), .B(n117), .Z(O[508]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[508]), .B(A[508]), .Z(n118) );
  XOR U178 ( .A(A[507]), .B(n119), .Z(O[507]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[507]), .B(A[507]), .Z(n120) );
  XOR U181 ( .A(A[506]), .B(n121), .Z(O[506]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[506]), .B(A[506]), .Z(n122) );
  XOR U184 ( .A(A[505]), .B(n123), .Z(O[505]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[505]), .B(A[505]), .Z(n124) );
  XOR U187 ( .A(A[504]), .B(n125), .Z(O[504]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[504]), .B(A[504]), .Z(n126) );
  XOR U190 ( .A(A[503]), .B(n127), .Z(O[503]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[503]), .B(A[503]), .Z(n128) );
  XOR U193 ( .A(A[502]), .B(n129), .Z(O[502]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[502]), .B(A[502]), .Z(n130) );
  XOR U196 ( .A(A[501]), .B(n131), .Z(O[501]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[501]), .B(A[501]), .Z(n132) );
  XOR U199 ( .A(A[500]), .B(n133), .Z(O[500]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[500]), .B(A[500]), .Z(n134) );
  XOR U202 ( .A(A[4]), .B(n135), .Z(O[4]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[4]), .B(A[4]), .Z(n136) );
  XOR U205 ( .A(A[49]), .B(n137), .Z(O[49]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[49]), .B(A[49]), .Z(n138) );
  XOR U208 ( .A(A[499]), .B(n139), .Z(O[499]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[499]), .B(A[499]), .Z(n140) );
  XOR U211 ( .A(A[498]), .B(n141), .Z(O[498]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[498]), .B(A[498]), .Z(n142) );
  XOR U214 ( .A(A[497]), .B(n143), .Z(O[497]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[497]), .B(A[497]), .Z(n144) );
  XOR U217 ( .A(A[496]), .B(n145), .Z(O[496]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[496]), .B(A[496]), .Z(n146) );
  XOR U220 ( .A(A[495]), .B(n147), .Z(O[495]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[495]), .B(A[495]), .Z(n148) );
  XOR U223 ( .A(A[494]), .B(n149), .Z(O[494]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[494]), .B(A[494]), .Z(n150) );
  XOR U226 ( .A(A[493]), .B(n151), .Z(O[493]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[493]), .B(A[493]), .Z(n152) );
  XOR U229 ( .A(A[492]), .B(n153), .Z(O[492]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[492]), .B(A[492]), .Z(n154) );
  XOR U232 ( .A(A[491]), .B(n155), .Z(O[491]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[491]), .B(A[491]), .Z(n156) );
  XOR U235 ( .A(A[490]), .B(n157), .Z(O[490]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[490]), .B(A[490]), .Z(n158) );
  XOR U238 ( .A(A[48]), .B(n159), .Z(O[48]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[48]), .B(A[48]), .Z(n160) );
  XOR U241 ( .A(A[489]), .B(n161), .Z(O[489]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[489]), .B(A[489]), .Z(n162) );
  XOR U244 ( .A(A[488]), .B(n163), .Z(O[488]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[488]), .B(A[488]), .Z(n164) );
  XOR U247 ( .A(A[487]), .B(n165), .Z(O[487]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[487]), .B(A[487]), .Z(n166) );
  XOR U250 ( .A(A[486]), .B(n167), .Z(O[486]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[486]), .B(A[486]), .Z(n168) );
  XOR U253 ( .A(A[485]), .B(n169), .Z(O[485]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[485]), .B(A[485]), .Z(n170) );
  XOR U256 ( .A(A[484]), .B(n171), .Z(O[484]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[484]), .B(A[484]), .Z(n172) );
  XOR U259 ( .A(A[483]), .B(n173), .Z(O[483]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[483]), .B(A[483]), .Z(n174) );
  XOR U262 ( .A(A[482]), .B(n175), .Z(O[482]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[482]), .B(A[482]), .Z(n176) );
  XOR U265 ( .A(A[481]), .B(n177), .Z(O[481]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[481]), .B(A[481]), .Z(n178) );
  XOR U268 ( .A(A[480]), .B(n179), .Z(O[480]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[480]), .B(A[480]), .Z(n180) );
  XOR U271 ( .A(A[47]), .B(n181), .Z(O[47]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[47]), .B(A[47]), .Z(n182) );
  XOR U274 ( .A(A[479]), .B(n183), .Z(O[479]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[479]), .B(A[479]), .Z(n184) );
  XOR U277 ( .A(A[478]), .B(n185), .Z(O[478]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[478]), .B(A[478]), .Z(n186) );
  XOR U280 ( .A(A[477]), .B(n187), .Z(O[477]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[477]), .B(A[477]), .Z(n188) );
  XOR U283 ( .A(A[476]), .B(n189), .Z(O[476]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[476]), .B(A[476]), .Z(n190) );
  XOR U286 ( .A(A[475]), .B(n191), .Z(O[475]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[475]), .B(A[475]), .Z(n192) );
  XOR U289 ( .A(A[474]), .B(n193), .Z(O[474]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[474]), .B(A[474]), .Z(n194) );
  XOR U292 ( .A(A[473]), .B(n195), .Z(O[473]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[473]), .B(A[473]), .Z(n196) );
  XOR U295 ( .A(A[472]), .B(n197), .Z(O[472]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[472]), .B(A[472]), .Z(n198) );
  XOR U298 ( .A(A[471]), .B(n199), .Z(O[471]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[471]), .B(A[471]), .Z(n200) );
  XOR U301 ( .A(A[470]), .B(n201), .Z(O[470]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[470]), .B(A[470]), .Z(n202) );
  XOR U304 ( .A(A[46]), .B(n203), .Z(O[46]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[46]), .B(A[46]), .Z(n204) );
  XOR U307 ( .A(A[469]), .B(n205), .Z(O[469]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[469]), .B(A[469]), .Z(n206) );
  XOR U310 ( .A(A[468]), .B(n207), .Z(O[468]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[468]), .B(A[468]), .Z(n208) );
  XOR U313 ( .A(A[467]), .B(n209), .Z(O[467]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[467]), .B(A[467]), .Z(n210) );
  XOR U316 ( .A(A[466]), .B(n211), .Z(O[466]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[466]), .B(A[466]), .Z(n212) );
  XOR U319 ( .A(A[465]), .B(n213), .Z(O[465]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[465]), .B(A[465]), .Z(n214) );
  XOR U322 ( .A(A[464]), .B(n215), .Z(O[464]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[464]), .B(A[464]), .Z(n216) );
  XOR U325 ( .A(A[463]), .B(n217), .Z(O[463]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[463]), .B(A[463]), .Z(n218) );
  XOR U328 ( .A(A[462]), .B(n219), .Z(O[462]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[462]), .B(A[462]), .Z(n220) );
  XOR U331 ( .A(A[461]), .B(n221), .Z(O[461]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[461]), .B(A[461]), .Z(n222) );
  XOR U334 ( .A(A[460]), .B(n223), .Z(O[460]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[460]), .B(A[460]), .Z(n224) );
  XOR U337 ( .A(A[45]), .B(n225), .Z(O[45]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[45]), .B(A[45]), .Z(n226) );
  XOR U340 ( .A(A[459]), .B(n227), .Z(O[459]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[459]), .B(A[459]), .Z(n228) );
  XOR U343 ( .A(A[458]), .B(n229), .Z(O[458]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[458]), .B(A[458]), .Z(n230) );
  XOR U346 ( .A(A[457]), .B(n231), .Z(O[457]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[457]), .B(A[457]), .Z(n232) );
  XOR U349 ( .A(A[456]), .B(n233), .Z(O[456]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[456]), .B(A[456]), .Z(n234) );
  XOR U352 ( .A(A[455]), .B(n235), .Z(O[455]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[455]), .B(A[455]), .Z(n236) );
  XOR U355 ( .A(A[454]), .B(n237), .Z(O[454]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[454]), .B(A[454]), .Z(n238) );
  XOR U358 ( .A(A[453]), .B(n239), .Z(O[453]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[453]), .B(A[453]), .Z(n240) );
  XOR U361 ( .A(A[452]), .B(n241), .Z(O[452]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[452]), .B(A[452]), .Z(n242) );
  XOR U364 ( .A(A[451]), .B(n243), .Z(O[451]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[451]), .B(A[451]), .Z(n244) );
  XOR U367 ( .A(A[450]), .B(n245), .Z(O[450]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[450]), .B(A[450]), .Z(n246) );
  XOR U370 ( .A(A[44]), .B(n247), .Z(O[44]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[44]), .B(A[44]), .Z(n248) );
  XOR U373 ( .A(A[449]), .B(n249), .Z(O[449]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[449]), .B(A[449]), .Z(n250) );
  XOR U376 ( .A(A[448]), .B(n251), .Z(O[448]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[448]), .B(A[448]), .Z(n252) );
  XOR U379 ( .A(A[447]), .B(n253), .Z(O[447]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[447]), .B(A[447]), .Z(n254) );
  XOR U382 ( .A(A[446]), .B(n255), .Z(O[446]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[446]), .B(A[446]), .Z(n256) );
  XOR U385 ( .A(A[445]), .B(n257), .Z(O[445]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[445]), .B(A[445]), .Z(n258) );
  XOR U388 ( .A(A[444]), .B(n259), .Z(O[444]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[444]), .B(A[444]), .Z(n260) );
  XOR U391 ( .A(A[443]), .B(n261), .Z(O[443]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[443]), .B(A[443]), .Z(n262) );
  XOR U394 ( .A(A[442]), .B(n263), .Z(O[442]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[442]), .B(A[442]), .Z(n264) );
  XOR U397 ( .A(A[441]), .B(n265), .Z(O[441]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[441]), .B(A[441]), .Z(n266) );
  XOR U400 ( .A(A[440]), .B(n267), .Z(O[440]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[440]), .B(A[440]), .Z(n268) );
  XOR U403 ( .A(A[43]), .B(n269), .Z(O[43]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[43]), .B(A[43]), .Z(n270) );
  XOR U406 ( .A(A[439]), .B(n271), .Z(O[439]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[439]), .B(A[439]), .Z(n272) );
  XOR U409 ( .A(A[438]), .B(n273), .Z(O[438]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[438]), .B(A[438]), .Z(n274) );
  XOR U412 ( .A(A[437]), .B(n275), .Z(O[437]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[437]), .B(A[437]), .Z(n276) );
  XOR U415 ( .A(A[436]), .B(n277), .Z(O[436]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[436]), .B(A[436]), .Z(n278) );
  XOR U418 ( .A(A[435]), .B(n279), .Z(O[435]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[435]), .B(A[435]), .Z(n280) );
  XOR U421 ( .A(A[434]), .B(n281), .Z(O[434]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[434]), .B(A[434]), .Z(n282) );
  XOR U424 ( .A(A[433]), .B(n283), .Z(O[433]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[433]), .B(A[433]), .Z(n284) );
  XOR U427 ( .A(A[432]), .B(n285), .Z(O[432]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[432]), .B(A[432]), .Z(n286) );
  XOR U430 ( .A(A[431]), .B(n287), .Z(O[431]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[431]), .B(A[431]), .Z(n288) );
  XOR U433 ( .A(A[430]), .B(n289), .Z(O[430]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[430]), .B(A[430]), .Z(n290) );
  XOR U436 ( .A(A[42]), .B(n291), .Z(O[42]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[42]), .B(A[42]), .Z(n292) );
  XOR U439 ( .A(A[429]), .B(n293), .Z(O[429]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[429]), .B(A[429]), .Z(n294) );
  XOR U442 ( .A(A[428]), .B(n295), .Z(O[428]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[428]), .B(A[428]), .Z(n296) );
  XOR U445 ( .A(A[427]), .B(n297), .Z(O[427]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[427]), .B(A[427]), .Z(n298) );
  XOR U448 ( .A(A[426]), .B(n299), .Z(O[426]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[426]), .B(A[426]), .Z(n300) );
  XOR U451 ( .A(A[425]), .B(n301), .Z(O[425]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[425]), .B(A[425]), .Z(n302) );
  XOR U454 ( .A(A[424]), .B(n303), .Z(O[424]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[424]), .B(A[424]), .Z(n304) );
  XOR U457 ( .A(A[423]), .B(n305), .Z(O[423]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[423]), .B(A[423]), .Z(n306) );
  XOR U460 ( .A(A[422]), .B(n307), .Z(O[422]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[422]), .B(A[422]), .Z(n308) );
  XOR U463 ( .A(A[421]), .B(n309), .Z(O[421]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[421]), .B(A[421]), .Z(n310) );
  XOR U466 ( .A(A[420]), .B(n311), .Z(O[420]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[420]), .B(A[420]), .Z(n312) );
  XOR U469 ( .A(A[41]), .B(n313), .Z(O[41]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[41]), .B(A[41]), .Z(n314) );
  XOR U472 ( .A(A[419]), .B(n315), .Z(O[419]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[419]), .B(A[419]), .Z(n316) );
  XOR U475 ( .A(A[418]), .B(n317), .Z(O[418]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[418]), .B(A[418]), .Z(n318) );
  XOR U478 ( .A(A[417]), .B(n319), .Z(O[417]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[417]), .B(A[417]), .Z(n320) );
  XOR U481 ( .A(A[416]), .B(n321), .Z(O[416]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[416]), .B(A[416]), .Z(n322) );
  XOR U484 ( .A(A[415]), .B(n323), .Z(O[415]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[415]), .B(A[415]), .Z(n324) );
  XOR U487 ( .A(A[414]), .B(n325), .Z(O[414]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[414]), .B(A[414]), .Z(n326) );
  XOR U490 ( .A(A[413]), .B(n327), .Z(O[413]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[413]), .B(A[413]), .Z(n328) );
  XOR U493 ( .A(A[412]), .B(n329), .Z(O[412]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[412]), .B(A[412]), .Z(n330) );
  XOR U496 ( .A(A[411]), .B(n331), .Z(O[411]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[411]), .B(A[411]), .Z(n332) );
  XOR U499 ( .A(A[410]), .B(n333), .Z(O[410]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[410]), .B(A[410]), .Z(n334) );
  XOR U502 ( .A(A[40]), .B(n335), .Z(O[40]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[40]), .B(A[40]), .Z(n336) );
  XOR U505 ( .A(A[409]), .B(n337), .Z(O[409]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[409]), .B(A[409]), .Z(n338) );
  XOR U508 ( .A(A[408]), .B(n339), .Z(O[408]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[408]), .B(A[408]), .Z(n340) );
  XOR U511 ( .A(A[407]), .B(n341), .Z(O[407]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[407]), .B(A[407]), .Z(n342) );
  XOR U514 ( .A(A[406]), .B(n343), .Z(O[406]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[406]), .B(A[406]), .Z(n344) );
  XOR U517 ( .A(A[405]), .B(n345), .Z(O[405]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[405]), .B(A[405]), .Z(n346) );
  XOR U520 ( .A(A[404]), .B(n347), .Z(O[404]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[404]), .B(A[404]), .Z(n348) );
  XOR U523 ( .A(A[403]), .B(n349), .Z(O[403]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[403]), .B(A[403]), .Z(n350) );
  XOR U526 ( .A(A[402]), .B(n351), .Z(O[402]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[402]), .B(A[402]), .Z(n352) );
  XOR U529 ( .A(A[401]), .B(n353), .Z(O[401]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[401]), .B(A[401]), .Z(n354) );
  XOR U532 ( .A(A[400]), .B(n355), .Z(O[400]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[400]), .B(A[400]), .Z(n356) );
  XOR U535 ( .A(A[3]), .B(n357), .Z(O[3]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[3]), .B(A[3]), .Z(n358) );
  XOR U538 ( .A(A[39]), .B(n359), .Z(O[39]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[39]), .B(A[39]), .Z(n360) );
  XOR U541 ( .A(A[399]), .B(n361), .Z(O[399]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[399]), .B(A[399]), .Z(n362) );
  XOR U544 ( .A(A[398]), .B(n363), .Z(O[398]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[398]), .B(A[398]), .Z(n364) );
  XOR U547 ( .A(A[397]), .B(n365), .Z(O[397]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[397]), .B(A[397]), .Z(n366) );
  XOR U550 ( .A(A[396]), .B(n367), .Z(O[396]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[396]), .B(A[396]), .Z(n368) );
  XOR U553 ( .A(A[395]), .B(n369), .Z(O[395]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[395]), .B(A[395]), .Z(n370) );
  XOR U556 ( .A(A[394]), .B(n371), .Z(O[394]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[394]), .B(A[394]), .Z(n372) );
  XOR U559 ( .A(A[393]), .B(n373), .Z(O[393]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[393]), .B(A[393]), .Z(n374) );
  XOR U562 ( .A(A[392]), .B(n375), .Z(O[392]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[392]), .B(A[392]), .Z(n376) );
  XOR U565 ( .A(A[391]), .B(n377), .Z(O[391]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[391]), .B(A[391]), .Z(n378) );
  XOR U568 ( .A(A[390]), .B(n379), .Z(O[390]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[390]), .B(A[390]), .Z(n380) );
  XOR U571 ( .A(A[38]), .B(n381), .Z(O[38]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[38]), .B(A[38]), .Z(n382) );
  XOR U574 ( .A(A[389]), .B(n383), .Z(O[389]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[389]), .B(A[389]), .Z(n384) );
  XOR U577 ( .A(A[388]), .B(n385), .Z(O[388]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[388]), .B(A[388]), .Z(n386) );
  XOR U580 ( .A(A[387]), .B(n387), .Z(O[387]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[387]), .B(A[387]), .Z(n388) );
  XOR U583 ( .A(A[386]), .B(n389), .Z(O[386]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[386]), .B(A[386]), .Z(n390) );
  XOR U586 ( .A(A[385]), .B(n391), .Z(O[385]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[385]), .B(A[385]), .Z(n392) );
  XOR U589 ( .A(A[384]), .B(n393), .Z(O[384]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[384]), .B(A[384]), .Z(n394) );
  XOR U592 ( .A(A[383]), .B(n395), .Z(O[383]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[383]), .B(A[383]), .Z(n396) );
  XOR U595 ( .A(A[382]), .B(n397), .Z(O[382]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[382]), .B(A[382]), .Z(n398) );
  XOR U598 ( .A(A[381]), .B(n399), .Z(O[381]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[381]), .B(A[381]), .Z(n400) );
  XOR U601 ( .A(A[380]), .B(n401), .Z(O[380]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[380]), .B(A[380]), .Z(n402) );
  XOR U604 ( .A(A[37]), .B(n403), .Z(O[37]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[37]), .B(A[37]), .Z(n404) );
  XOR U607 ( .A(A[379]), .B(n405), .Z(O[379]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[379]), .B(A[379]), .Z(n406) );
  XOR U610 ( .A(A[378]), .B(n407), .Z(O[378]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[378]), .B(A[378]), .Z(n408) );
  XOR U613 ( .A(A[377]), .B(n409), .Z(O[377]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[377]), .B(A[377]), .Z(n410) );
  XOR U616 ( .A(A[376]), .B(n411), .Z(O[376]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[376]), .B(A[376]), .Z(n412) );
  XOR U619 ( .A(A[375]), .B(n413), .Z(O[375]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[375]), .B(A[375]), .Z(n414) );
  XOR U622 ( .A(A[374]), .B(n415), .Z(O[374]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[374]), .B(A[374]), .Z(n416) );
  XOR U625 ( .A(A[373]), .B(n417), .Z(O[373]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[373]), .B(A[373]), .Z(n418) );
  XOR U628 ( .A(A[372]), .B(n419), .Z(O[372]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[372]), .B(A[372]), .Z(n420) );
  XOR U631 ( .A(A[371]), .B(n421), .Z(O[371]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[371]), .B(A[371]), .Z(n422) );
  XOR U634 ( .A(A[370]), .B(n423), .Z(O[370]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[370]), .B(A[370]), .Z(n424) );
  XOR U637 ( .A(A[36]), .B(n425), .Z(O[36]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[36]), .B(A[36]), .Z(n426) );
  XOR U640 ( .A(A[369]), .B(n427), .Z(O[369]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[369]), .B(A[369]), .Z(n428) );
  XOR U643 ( .A(A[368]), .B(n429), .Z(O[368]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[368]), .B(A[368]), .Z(n430) );
  XOR U646 ( .A(A[367]), .B(n431), .Z(O[367]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[367]), .B(A[367]), .Z(n432) );
  XOR U649 ( .A(A[366]), .B(n433), .Z(O[366]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[366]), .B(A[366]), .Z(n434) );
  XOR U652 ( .A(A[365]), .B(n435), .Z(O[365]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[365]), .B(A[365]), .Z(n436) );
  XOR U655 ( .A(A[364]), .B(n437), .Z(O[364]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[364]), .B(A[364]), .Z(n438) );
  XOR U658 ( .A(A[363]), .B(n439), .Z(O[363]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[363]), .B(A[363]), .Z(n440) );
  XOR U661 ( .A(A[362]), .B(n441), .Z(O[362]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[362]), .B(A[362]), .Z(n442) );
  XOR U664 ( .A(A[361]), .B(n443), .Z(O[361]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[361]), .B(A[361]), .Z(n444) );
  XOR U667 ( .A(A[360]), .B(n445), .Z(O[360]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[360]), .B(A[360]), .Z(n446) );
  XOR U670 ( .A(A[35]), .B(n447), .Z(O[35]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[35]), .B(A[35]), .Z(n448) );
  XOR U673 ( .A(A[359]), .B(n449), .Z(O[359]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[359]), .B(A[359]), .Z(n450) );
  XOR U676 ( .A(A[358]), .B(n451), .Z(O[358]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[358]), .B(A[358]), .Z(n452) );
  XOR U679 ( .A(A[357]), .B(n453), .Z(O[357]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[357]), .B(A[357]), .Z(n454) );
  XOR U682 ( .A(A[356]), .B(n455), .Z(O[356]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[356]), .B(A[356]), .Z(n456) );
  XOR U685 ( .A(A[355]), .B(n457), .Z(O[355]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[355]), .B(A[355]), .Z(n458) );
  XOR U688 ( .A(A[354]), .B(n459), .Z(O[354]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[354]), .B(A[354]), .Z(n460) );
  XOR U691 ( .A(A[353]), .B(n461), .Z(O[353]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[353]), .B(A[353]), .Z(n462) );
  XOR U694 ( .A(A[352]), .B(n463), .Z(O[352]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[352]), .B(A[352]), .Z(n464) );
  XOR U697 ( .A(A[351]), .B(n465), .Z(O[351]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[351]), .B(A[351]), .Z(n466) );
  XOR U700 ( .A(A[350]), .B(n467), .Z(O[350]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[350]), .B(A[350]), .Z(n468) );
  XOR U703 ( .A(A[34]), .B(n469), .Z(O[34]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[34]), .B(A[34]), .Z(n470) );
  XOR U706 ( .A(A[349]), .B(n471), .Z(O[349]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[349]), .B(A[349]), .Z(n472) );
  XOR U709 ( .A(A[348]), .B(n473), .Z(O[348]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[348]), .B(A[348]), .Z(n474) );
  XOR U712 ( .A(A[347]), .B(n475), .Z(O[347]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[347]), .B(A[347]), .Z(n476) );
  XOR U715 ( .A(A[346]), .B(n477), .Z(O[346]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[346]), .B(A[346]), .Z(n478) );
  XOR U718 ( .A(A[345]), .B(n479), .Z(O[345]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[345]), .B(A[345]), .Z(n480) );
  XOR U721 ( .A(A[344]), .B(n481), .Z(O[344]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[344]), .B(A[344]), .Z(n482) );
  XOR U724 ( .A(A[343]), .B(n483), .Z(O[343]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[343]), .B(A[343]), .Z(n484) );
  XOR U727 ( .A(A[342]), .B(n485), .Z(O[342]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[342]), .B(A[342]), .Z(n486) );
  XOR U730 ( .A(A[341]), .B(n487), .Z(O[341]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[341]), .B(A[341]), .Z(n488) );
  XOR U733 ( .A(A[340]), .B(n489), .Z(O[340]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[340]), .B(A[340]), .Z(n490) );
  XOR U736 ( .A(A[33]), .B(n491), .Z(O[33]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[33]), .B(A[33]), .Z(n492) );
  XOR U739 ( .A(A[339]), .B(n493), .Z(O[339]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[339]), .B(A[339]), .Z(n494) );
  XOR U742 ( .A(A[338]), .B(n495), .Z(O[338]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[338]), .B(A[338]), .Z(n496) );
  XOR U745 ( .A(A[337]), .B(n497), .Z(O[337]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[337]), .B(A[337]), .Z(n498) );
  XOR U748 ( .A(A[336]), .B(n499), .Z(O[336]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[336]), .B(A[336]), .Z(n500) );
  XOR U751 ( .A(A[335]), .B(n501), .Z(O[335]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[335]), .B(A[335]), .Z(n502) );
  XOR U754 ( .A(A[334]), .B(n503), .Z(O[334]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[334]), .B(A[334]), .Z(n504) );
  XOR U757 ( .A(A[333]), .B(n505), .Z(O[333]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[333]), .B(A[333]), .Z(n506) );
  XOR U760 ( .A(A[332]), .B(n507), .Z(O[332]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[332]), .B(A[332]), .Z(n508) );
  XOR U763 ( .A(A[331]), .B(n509), .Z(O[331]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[331]), .B(A[331]), .Z(n510) );
  XOR U766 ( .A(A[330]), .B(n511), .Z(O[330]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[330]), .B(A[330]), .Z(n512) );
  XOR U769 ( .A(A[32]), .B(n513), .Z(O[32]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[32]), .B(A[32]), .Z(n514) );
  XOR U772 ( .A(A[329]), .B(n515), .Z(O[329]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[329]), .B(A[329]), .Z(n516) );
  XOR U775 ( .A(A[328]), .B(n517), .Z(O[328]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[328]), .B(A[328]), .Z(n518) );
  XOR U778 ( .A(A[327]), .B(n519), .Z(O[327]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[327]), .B(A[327]), .Z(n520) );
  XOR U781 ( .A(A[326]), .B(n521), .Z(O[326]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[326]), .B(A[326]), .Z(n522) );
  XOR U784 ( .A(A[325]), .B(n523), .Z(O[325]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[325]), .B(A[325]), .Z(n524) );
  XOR U787 ( .A(A[324]), .B(n525), .Z(O[324]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[324]), .B(A[324]), .Z(n526) );
  XOR U790 ( .A(A[323]), .B(n527), .Z(O[323]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[323]), .B(A[323]), .Z(n528) );
  XOR U793 ( .A(A[322]), .B(n529), .Z(O[322]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[322]), .B(A[322]), .Z(n530) );
  XOR U796 ( .A(A[321]), .B(n531), .Z(O[321]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[321]), .B(A[321]), .Z(n532) );
  XOR U799 ( .A(A[320]), .B(n533), .Z(O[320]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[320]), .B(A[320]), .Z(n534) );
  XOR U802 ( .A(A[31]), .B(n535), .Z(O[31]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[31]), .B(A[31]), .Z(n536) );
  XOR U805 ( .A(A[319]), .B(n537), .Z(O[319]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[319]), .B(A[319]), .Z(n538) );
  XOR U808 ( .A(A[318]), .B(n539), .Z(O[318]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[318]), .B(A[318]), .Z(n540) );
  XOR U811 ( .A(A[317]), .B(n541), .Z(O[317]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[317]), .B(A[317]), .Z(n542) );
  XOR U814 ( .A(A[316]), .B(n543), .Z(O[316]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[316]), .B(A[316]), .Z(n544) );
  XOR U817 ( .A(A[315]), .B(n545), .Z(O[315]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[315]), .B(A[315]), .Z(n546) );
  XOR U820 ( .A(A[314]), .B(n547), .Z(O[314]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[314]), .B(A[314]), .Z(n548) );
  XOR U823 ( .A(A[313]), .B(n549), .Z(O[313]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[313]), .B(A[313]), .Z(n550) );
  XOR U826 ( .A(A[312]), .B(n551), .Z(O[312]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[312]), .B(A[312]), .Z(n552) );
  XOR U829 ( .A(A[311]), .B(n553), .Z(O[311]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[311]), .B(A[311]), .Z(n554) );
  XOR U832 ( .A(A[310]), .B(n555), .Z(O[310]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[310]), .B(A[310]), .Z(n556) );
  XOR U835 ( .A(A[30]), .B(n557), .Z(O[30]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[30]), .B(A[30]), .Z(n558) );
  XOR U838 ( .A(A[309]), .B(n559), .Z(O[309]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[309]), .B(A[309]), .Z(n560) );
  XOR U841 ( .A(A[308]), .B(n561), .Z(O[308]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[308]), .B(A[308]), .Z(n562) );
  XOR U844 ( .A(A[307]), .B(n563), .Z(O[307]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[307]), .B(A[307]), .Z(n564) );
  XOR U847 ( .A(A[306]), .B(n565), .Z(O[306]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[306]), .B(A[306]), .Z(n566) );
  XOR U850 ( .A(A[305]), .B(n567), .Z(O[305]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[305]), .B(A[305]), .Z(n568) );
  XOR U853 ( .A(A[304]), .B(n569), .Z(O[304]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[304]), .B(A[304]), .Z(n570) );
  XOR U856 ( .A(A[303]), .B(n571), .Z(O[303]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[303]), .B(A[303]), .Z(n572) );
  XOR U859 ( .A(A[302]), .B(n573), .Z(O[302]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[302]), .B(A[302]), .Z(n574) );
  XOR U862 ( .A(A[301]), .B(n575), .Z(O[301]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[301]), .B(A[301]), .Z(n576) );
  XOR U865 ( .A(A[300]), .B(n577), .Z(O[300]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[300]), .B(A[300]), .Z(n578) );
  XOR U868 ( .A(A[2]), .B(n579), .Z(O[2]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[2]), .B(A[2]), .Z(n580) );
  XOR U871 ( .A(A[29]), .B(n581), .Z(O[29]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[29]), .B(A[29]), .Z(n582) );
  XOR U874 ( .A(A[299]), .B(n583), .Z(O[299]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[299]), .B(A[299]), .Z(n584) );
  XOR U877 ( .A(A[298]), .B(n585), .Z(O[298]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[298]), .B(A[298]), .Z(n586) );
  XOR U880 ( .A(A[297]), .B(n587), .Z(O[297]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[297]), .B(A[297]), .Z(n588) );
  XOR U883 ( .A(A[296]), .B(n589), .Z(O[296]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[296]), .B(A[296]), .Z(n590) );
  XOR U886 ( .A(A[295]), .B(n591), .Z(O[295]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[295]), .B(A[295]), .Z(n592) );
  XOR U889 ( .A(A[294]), .B(n593), .Z(O[294]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[294]), .B(A[294]), .Z(n594) );
  XOR U892 ( .A(A[293]), .B(n595), .Z(O[293]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[293]), .B(A[293]), .Z(n596) );
  XOR U895 ( .A(A[292]), .B(n597), .Z(O[292]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[292]), .B(A[292]), .Z(n598) );
  XOR U898 ( .A(A[291]), .B(n599), .Z(O[291]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[291]), .B(A[291]), .Z(n600) );
  XOR U901 ( .A(A[290]), .B(n601), .Z(O[290]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[290]), .B(A[290]), .Z(n602) );
  XOR U904 ( .A(A[28]), .B(n603), .Z(O[28]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[28]), .B(A[28]), .Z(n604) );
  XOR U907 ( .A(A[289]), .B(n605), .Z(O[289]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[289]), .B(A[289]), .Z(n606) );
  XOR U910 ( .A(A[288]), .B(n607), .Z(O[288]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[288]), .B(A[288]), .Z(n608) );
  XOR U913 ( .A(A[287]), .B(n609), .Z(O[287]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[287]), .B(A[287]), .Z(n610) );
  XOR U916 ( .A(A[286]), .B(n611), .Z(O[286]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[286]), .B(A[286]), .Z(n612) );
  XOR U919 ( .A(A[285]), .B(n613), .Z(O[285]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[285]), .B(A[285]), .Z(n614) );
  XOR U922 ( .A(A[284]), .B(n615), .Z(O[284]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[284]), .B(A[284]), .Z(n616) );
  XOR U925 ( .A(A[283]), .B(n617), .Z(O[283]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[283]), .B(A[283]), .Z(n618) );
  XOR U928 ( .A(A[282]), .B(n619), .Z(O[282]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[282]), .B(A[282]), .Z(n620) );
  XOR U931 ( .A(A[281]), .B(n621), .Z(O[281]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[281]), .B(A[281]), .Z(n622) );
  XOR U934 ( .A(A[280]), .B(n623), .Z(O[280]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[280]), .B(A[280]), .Z(n624) );
  XOR U937 ( .A(A[27]), .B(n625), .Z(O[27]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[27]), .B(A[27]), .Z(n626) );
  XOR U940 ( .A(A[279]), .B(n627), .Z(O[279]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[279]), .B(A[279]), .Z(n628) );
  XOR U943 ( .A(A[278]), .B(n629), .Z(O[278]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[278]), .B(A[278]), .Z(n630) );
  XOR U946 ( .A(A[277]), .B(n631), .Z(O[277]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[277]), .B(A[277]), .Z(n632) );
  XOR U949 ( .A(A[276]), .B(n633), .Z(O[276]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[276]), .B(A[276]), .Z(n634) );
  XOR U952 ( .A(A[275]), .B(n635), .Z(O[275]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[275]), .B(A[275]), .Z(n636) );
  XOR U955 ( .A(A[274]), .B(n637), .Z(O[274]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[274]), .B(A[274]), .Z(n638) );
  XOR U958 ( .A(A[273]), .B(n639), .Z(O[273]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[273]), .B(A[273]), .Z(n640) );
  XOR U961 ( .A(A[272]), .B(n641), .Z(O[272]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[272]), .B(A[272]), .Z(n642) );
  XOR U964 ( .A(A[271]), .B(n643), .Z(O[271]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[271]), .B(A[271]), .Z(n644) );
  XOR U967 ( .A(A[270]), .B(n645), .Z(O[270]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[270]), .B(A[270]), .Z(n646) );
  XOR U970 ( .A(A[26]), .B(n647), .Z(O[26]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[26]), .B(A[26]), .Z(n648) );
  XOR U973 ( .A(A[269]), .B(n649), .Z(O[269]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[269]), .B(A[269]), .Z(n650) );
  XOR U976 ( .A(A[268]), .B(n651), .Z(O[268]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[268]), .B(A[268]), .Z(n652) );
  XOR U979 ( .A(A[267]), .B(n653), .Z(O[267]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[267]), .B(A[267]), .Z(n654) );
  XOR U982 ( .A(A[266]), .B(n655), .Z(O[266]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[266]), .B(A[266]), .Z(n656) );
  XOR U985 ( .A(A[265]), .B(n657), .Z(O[265]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[265]), .B(A[265]), .Z(n658) );
  XOR U988 ( .A(A[264]), .B(n659), .Z(O[264]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[264]), .B(A[264]), .Z(n660) );
  XOR U991 ( .A(A[263]), .B(n661), .Z(O[263]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[263]), .B(A[263]), .Z(n662) );
  XOR U994 ( .A(A[262]), .B(n663), .Z(O[262]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[262]), .B(A[262]), .Z(n664) );
  XOR U997 ( .A(A[261]), .B(n665), .Z(O[261]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[261]), .B(A[261]), .Z(n666) );
  XOR U1000 ( .A(A[260]), .B(n667), .Z(O[260]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[260]), .B(A[260]), .Z(n668) );
  XOR U1003 ( .A(A[25]), .B(n669), .Z(O[25]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[25]), .B(A[25]), .Z(n670) );
  XOR U1006 ( .A(A[259]), .B(n671), .Z(O[259]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[259]), .B(A[259]), .Z(n672) );
  XOR U1009 ( .A(A[258]), .B(n673), .Z(O[258]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[258]), .B(A[258]), .Z(n674) );
  XOR U1012 ( .A(A[257]), .B(n675), .Z(O[257]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[257]), .B(A[257]), .Z(n676) );
  XOR U1015 ( .A(A[256]), .B(n677), .Z(O[256]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[256]), .B(A[256]), .Z(n678) );
  XOR U1018 ( .A(A[255]), .B(n679), .Z(O[255]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[255]), .B(A[255]), .Z(n680) );
  XOR U1021 ( .A(A[254]), .B(n681), .Z(O[254]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[254]), .B(A[254]), .Z(n682) );
  XOR U1024 ( .A(A[253]), .B(n683), .Z(O[253]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[253]), .B(A[253]), .Z(n684) );
  XOR U1027 ( .A(A[252]), .B(n685), .Z(O[252]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[252]), .B(A[252]), .Z(n686) );
  XOR U1030 ( .A(A[251]), .B(n687), .Z(O[251]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[251]), .B(A[251]), .Z(n688) );
  XOR U1033 ( .A(A[250]), .B(n689), .Z(O[250]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[250]), .B(A[250]), .Z(n690) );
  XOR U1036 ( .A(A[24]), .B(n691), .Z(O[24]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[24]), .B(A[24]), .Z(n692) );
  XOR U1039 ( .A(A[249]), .B(n693), .Z(O[249]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[249]), .B(A[249]), .Z(n694) );
  XOR U1042 ( .A(A[248]), .B(n695), .Z(O[248]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[248]), .B(A[248]), .Z(n696) );
  XOR U1045 ( .A(A[247]), .B(n697), .Z(O[247]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[247]), .B(A[247]), .Z(n698) );
  XOR U1048 ( .A(A[246]), .B(n699), .Z(O[246]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[246]), .B(A[246]), .Z(n700) );
  XOR U1051 ( .A(A[245]), .B(n701), .Z(O[245]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[245]), .B(A[245]), .Z(n702) );
  XOR U1054 ( .A(A[244]), .B(n703), .Z(O[244]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[244]), .B(A[244]), .Z(n704) );
  XOR U1057 ( .A(A[243]), .B(n705), .Z(O[243]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[243]), .B(A[243]), .Z(n706) );
  XOR U1060 ( .A(A[242]), .B(n707), .Z(O[242]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[242]), .B(A[242]), .Z(n708) );
  XOR U1063 ( .A(A[241]), .B(n709), .Z(O[241]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[241]), .B(A[241]), .Z(n710) );
  XOR U1066 ( .A(A[240]), .B(n711), .Z(O[240]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[240]), .B(A[240]), .Z(n712) );
  XOR U1069 ( .A(A[23]), .B(n713), .Z(O[23]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[23]), .B(A[23]), .Z(n714) );
  XOR U1072 ( .A(A[239]), .B(n715), .Z(O[239]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[239]), .B(A[239]), .Z(n716) );
  XOR U1075 ( .A(A[238]), .B(n717), .Z(O[238]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[238]), .B(A[238]), .Z(n718) );
  XOR U1078 ( .A(A[237]), .B(n719), .Z(O[237]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[237]), .B(A[237]), .Z(n720) );
  XOR U1081 ( .A(A[236]), .B(n721), .Z(O[236]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[236]), .B(A[236]), .Z(n722) );
  XOR U1084 ( .A(A[235]), .B(n723), .Z(O[235]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[235]), .B(A[235]), .Z(n724) );
  XOR U1087 ( .A(A[234]), .B(n725), .Z(O[234]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[234]), .B(A[234]), .Z(n726) );
  XOR U1090 ( .A(A[233]), .B(n727), .Z(O[233]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[233]), .B(A[233]), .Z(n728) );
  XOR U1093 ( .A(A[232]), .B(n729), .Z(O[232]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[232]), .B(A[232]), .Z(n730) );
  XOR U1096 ( .A(A[231]), .B(n731), .Z(O[231]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[231]), .B(A[231]), .Z(n732) );
  XOR U1099 ( .A(A[230]), .B(n733), .Z(O[230]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[230]), .B(A[230]), .Z(n734) );
  XOR U1102 ( .A(A[22]), .B(n735), .Z(O[22]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[22]), .B(A[22]), .Z(n736) );
  XOR U1105 ( .A(A[229]), .B(n737), .Z(O[229]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[229]), .B(A[229]), .Z(n738) );
  XOR U1108 ( .A(A[228]), .B(n739), .Z(O[228]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[228]), .B(A[228]), .Z(n740) );
  XOR U1111 ( .A(A[227]), .B(n741), .Z(O[227]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[227]), .B(A[227]), .Z(n742) );
  XOR U1114 ( .A(A[226]), .B(n743), .Z(O[226]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[226]), .B(A[226]), .Z(n744) );
  XOR U1117 ( .A(A[225]), .B(n745), .Z(O[225]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[225]), .B(A[225]), .Z(n746) );
  XOR U1120 ( .A(A[224]), .B(n747), .Z(O[224]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[224]), .B(A[224]), .Z(n748) );
  XOR U1123 ( .A(A[223]), .B(n749), .Z(O[223]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[223]), .B(A[223]), .Z(n750) );
  XOR U1126 ( .A(A[222]), .B(n751), .Z(O[222]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[222]), .B(A[222]), .Z(n752) );
  XOR U1129 ( .A(A[221]), .B(n753), .Z(O[221]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[221]), .B(A[221]), .Z(n754) );
  XOR U1132 ( .A(A[220]), .B(n755), .Z(O[220]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[220]), .B(A[220]), .Z(n756) );
  XOR U1135 ( .A(A[21]), .B(n757), .Z(O[21]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[21]), .B(A[21]), .Z(n758) );
  XOR U1138 ( .A(A[219]), .B(n759), .Z(O[219]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[219]), .B(A[219]), .Z(n760) );
  XOR U1141 ( .A(A[218]), .B(n761), .Z(O[218]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[218]), .B(A[218]), .Z(n762) );
  XOR U1144 ( .A(A[217]), .B(n763), .Z(O[217]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[217]), .B(A[217]), .Z(n764) );
  XOR U1147 ( .A(A[216]), .B(n765), .Z(O[216]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[216]), .B(A[216]), .Z(n766) );
  XOR U1150 ( .A(A[215]), .B(n767), .Z(O[215]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[215]), .B(A[215]), .Z(n768) );
  XOR U1153 ( .A(A[214]), .B(n769), .Z(O[214]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[214]), .B(A[214]), .Z(n770) );
  XOR U1156 ( .A(A[213]), .B(n771), .Z(O[213]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[213]), .B(A[213]), .Z(n772) );
  XOR U1159 ( .A(A[212]), .B(n773), .Z(O[212]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[212]), .B(A[212]), .Z(n774) );
  XOR U1162 ( .A(A[211]), .B(n775), .Z(O[211]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[211]), .B(A[211]), .Z(n776) );
  XOR U1165 ( .A(A[210]), .B(n777), .Z(O[210]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[210]), .B(A[210]), .Z(n778) );
  XOR U1168 ( .A(A[20]), .B(n779), .Z(O[20]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[20]), .B(A[20]), .Z(n780) );
  XOR U1171 ( .A(A[209]), .B(n781), .Z(O[209]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[209]), .B(A[209]), .Z(n782) );
  XOR U1174 ( .A(A[208]), .B(n783), .Z(O[208]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[208]), .B(A[208]), .Z(n784) );
  XOR U1177 ( .A(A[207]), .B(n785), .Z(O[207]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[207]), .B(A[207]), .Z(n786) );
  XOR U1180 ( .A(A[206]), .B(n787), .Z(O[206]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[206]), .B(A[206]), .Z(n788) );
  XOR U1183 ( .A(A[205]), .B(n789), .Z(O[205]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[205]), .B(A[205]), .Z(n790) );
  XOR U1186 ( .A(A[204]), .B(n791), .Z(O[204]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[204]), .B(A[204]), .Z(n792) );
  XOR U1189 ( .A(A[203]), .B(n793), .Z(O[203]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[203]), .B(A[203]), .Z(n794) );
  XOR U1192 ( .A(A[202]), .B(n795), .Z(O[202]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[202]), .B(A[202]), .Z(n796) );
  XOR U1195 ( .A(A[201]), .B(n797), .Z(O[201]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[201]), .B(A[201]), .Z(n798) );
  XOR U1198 ( .A(A[200]), .B(n799), .Z(O[200]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[200]), .B(A[200]), .Z(n800) );
  XOR U1201 ( .A(A[1]), .B(n801), .Z(O[1]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[1]), .B(A[1]), .Z(n802) );
  XOR U1204 ( .A(A[19]), .B(n803), .Z(O[19]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[19]), .B(A[19]), .Z(n804) );
  XOR U1207 ( .A(A[199]), .B(n805), .Z(O[199]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[199]), .B(A[199]), .Z(n806) );
  XOR U1210 ( .A(A[198]), .B(n807), .Z(O[198]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[198]), .B(A[198]), .Z(n808) );
  XOR U1213 ( .A(A[197]), .B(n809), .Z(O[197]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[197]), .B(A[197]), .Z(n810) );
  XOR U1216 ( .A(A[196]), .B(n811), .Z(O[196]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[196]), .B(A[196]), .Z(n812) );
  XOR U1219 ( .A(A[195]), .B(n813), .Z(O[195]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[195]), .B(A[195]), .Z(n814) );
  XOR U1222 ( .A(A[194]), .B(n815), .Z(O[194]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[194]), .B(A[194]), .Z(n816) );
  XOR U1225 ( .A(A[193]), .B(n817), .Z(O[193]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[193]), .B(A[193]), .Z(n818) );
  XOR U1228 ( .A(A[192]), .B(n819), .Z(O[192]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[192]), .B(A[192]), .Z(n820) );
  XOR U1231 ( .A(A[191]), .B(n821), .Z(O[191]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[191]), .B(A[191]), .Z(n822) );
  XOR U1234 ( .A(A[190]), .B(n823), .Z(O[190]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[190]), .B(A[190]), .Z(n824) );
  XOR U1237 ( .A(A[18]), .B(n825), .Z(O[18]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[18]), .B(A[18]), .Z(n826) );
  XOR U1240 ( .A(A[189]), .B(n827), .Z(O[189]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[189]), .B(A[189]), .Z(n828) );
  XOR U1243 ( .A(A[188]), .B(n829), .Z(O[188]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[188]), .B(A[188]), .Z(n830) );
  XOR U1246 ( .A(A[187]), .B(n831), .Z(O[187]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[187]), .B(A[187]), .Z(n832) );
  XOR U1249 ( .A(A[186]), .B(n833), .Z(O[186]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[186]), .B(A[186]), .Z(n834) );
  XOR U1252 ( .A(A[185]), .B(n835), .Z(O[185]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[185]), .B(A[185]), .Z(n836) );
  XOR U1255 ( .A(A[184]), .B(n837), .Z(O[184]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[184]), .B(A[184]), .Z(n838) );
  XOR U1258 ( .A(A[183]), .B(n839), .Z(O[183]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[183]), .B(A[183]), .Z(n840) );
  XOR U1261 ( .A(A[182]), .B(n841), .Z(O[182]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[182]), .B(A[182]), .Z(n842) );
  XOR U1264 ( .A(A[181]), .B(n843), .Z(O[181]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[181]), .B(A[181]), .Z(n844) );
  XOR U1267 ( .A(A[180]), .B(n845), .Z(O[180]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[180]), .B(A[180]), .Z(n846) );
  XOR U1270 ( .A(A[17]), .B(n847), .Z(O[17]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[17]), .B(A[17]), .Z(n848) );
  XOR U1273 ( .A(A[179]), .B(n849), .Z(O[179]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[179]), .B(A[179]), .Z(n850) );
  XOR U1276 ( .A(A[178]), .B(n851), .Z(O[178]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[178]), .B(A[178]), .Z(n852) );
  XOR U1279 ( .A(A[177]), .B(n853), .Z(O[177]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[177]), .B(A[177]), .Z(n854) );
  XOR U1282 ( .A(A[176]), .B(n855), .Z(O[176]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[176]), .B(A[176]), .Z(n856) );
  XOR U1285 ( .A(A[175]), .B(n857), .Z(O[175]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[175]), .B(A[175]), .Z(n858) );
  XOR U1288 ( .A(A[174]), .B(n859), .Z(O[174]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[174]), .B(A[174]), .Z(n860) );
  XOR U1291 ( .A(A[173]), .B(n861), .Z(O[173]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[173]), .B(A[173]), .Z(n862) );
  XOR U1294 ( .A(A[172]), .B(n863), .Z(O[172]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[172]), .B(A[172]), .Z(n864) );
  XOR U1297 ( .A(A[171]), .B(n865), .Z(O[171]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[171]), .B(A[171]), .Z(n866) );
  XOR U1300 ( .A(A[170]), .B(n867), .Z(O[170]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[170]), .B(A[170]), .Z(n868) );
  XOR U1303 ( .A(A[16]), .B(n869), .Z(O[16]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[16]), .B(A[16]), .Z(n870) );
  XOR U1306 ( .A(A[169]), .B(n871), .Z(O[169]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[169]), .B(A[169]), .Z(n872) );
  XOR U1309 ( .A(A[168]), .B(n873), .Z(O[168]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[168]), .B(A[168]), .Z(n874) );
  XOR U1312 ( .A(A[167]), .B(n875), .Z(O[167]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[167]), .B(A[167]), .Z(n876) );
  XOR U1315 ( .A(A[166]), .B(n877), .Z(O[166]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[166]), .B(A[166]), .Z(n878) );
  XOR U1318 ( .A(A[165]), .B(n879), .Z(O[165]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[165]), .B(A[165]), .Z(n880) );
  XOR U1321 ( .A(A[164]), .B(n881), .Z(O[164]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[164]), .B(A[164]), .Z(n882) );
  XOR U1324 ( .A(A[163]), .B(n883), .Z(O[163]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[163]), .B(A[163]), .Z(n884) );
  XOR U1327 ( .A(A[162]), .B(n885), .Z(O[162]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[162]), .B(A[162]), .Z(n886) );
  XOR U1330 ( .A(A[161]), .B(n887), .Z(O[161]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[161]), .B(A[161]), .Z(n888) );
  XOR U1333 ( .A(A[160]), .B(n889), .Z(O[160]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[160]), .B(A[160]), .Z(n890) );
  XOR U1336 ( .A(A[15]), .B(n891), .Z(O[15]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[15]), .B(A[15]), .Z(n892) );
  XOR U1339 ( .A(A[159]), .B(n893), .Z(O[159]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[159]), .B(A[159]), .Z(n894) );
  XOR U1342 ( .A(A[158]), .B(n895), .Z(O[158]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[158]), .B(A[158]), .Z(n896) );
  XOR U1345 ( .A(A[157]), .B(n897), .Z(O[157]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[157]), .B(A[157]), .Z(n898) );
  XOR U1348 ( .A(A[156]), .B(n899), .Z(O[156]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[156]), .B(A[156]), .Z(n900) );
  XOR U1351 ( .A(A[155]), .B(n901), .Z(O[155]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[155]), .B(A[155]), .Z(n902) );
  XOR U1354 ( .A(A[154]), .B(n903), .Z(O[154]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[154]), .B(A[154]), .Z(n904) );
  XOR U1357 ( .A(A[153]), .B(n905), .Z(O[153]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[153]), .B(A[153]), .Z(n906) );
  XOR U1360 ( .A(A[152]), .B(n907), .Z(O[152]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[152]), .B(A[152]), .Z(n908) );
  XOR U1363 ( .A(A[151]), .B(n909), .Z(O[151]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[151]), .B(A[151]), .Z(n910) );
  XOR U1366 ( .A(A[150]), .B(n911), .Z(O[150]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[150]), .B(A[150]), .Z(n912) );
  XOR U1369 ( .A(A[14]), .B(n913), .Z(O[14]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[14]), .B(A[14]), .Z(n914) );
  XOR U1372 ( .A(A[149]), .B(n915), .Z(O[149]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[149]), .B(A[149]), .Z(n916) );
  XOR U1375 ( .A(A[148]), .B(n917), .Z(O[148]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[148]), .B(A[148]), .Z(n918) );
  XOR U1378 ( .A(A[147]), .B(n919), .Z(O[147]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[147]), .B(A[147]), .Z(n920) );
  XOR U1381 ( .A(A[146]), .B(n921), .Z(O[146]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[146]), .B(A[146]), .Z(n922) );
  XOR U1384 ( .A(A[145]), .B(n923), .Z(O[145]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[145]), .B(A[145]), .Z(n924) );
  XOR U1387 ( .A(A[144]), .B(n925), .Z(O[144]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[144]), .B(A[144]), .Z(n926) );
  XOR U1390 ( .A(A[143]), .B(n927), .Z(O[143]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[143]), .B(A[143]), .Z(n928) );
  XOR U1393 ( .A(A[142]), .B(n929), .Z(O[142]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[142]), .B(A[142]), .Z(n930) );
  XOR U1396 ( .A(A[141]), .B(n931), .Z(O[141]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[141]), .B(A[141]), .Z(n932) );
  XOR U1399 ( .A(A[140]), .B(n933), .Z(O[140]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[140]), .B(A[140]), .Z(n934) );
  XOR U1402 ( .A(A[13]), .B(n935), .Z(O[13]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[13]), .B(A[13]), .Z(n936) );
  XOR U1405 ( .A(A[139]), .B(n937), .Z(O[139]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[139]), .B(A[139]), .Z(n938) );
  XOR U1408 ( .A(A[138]), .B(n939), .Z(O[138]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[138]), .B(A[138]), .Z(n940) );
  XOR U1411 ( .A(A[137]), .B(n941), .Z(O[137]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[137]), .B(A[137]), .Z(n942) );
  XOR U1414 ( .A(A[136]), .B(n943), .Z(O[136]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[136]), .B(A[136]), .Z(n944) );
  XOR U1417 ( .A(A[135]), .B(n945), .Z(O[135]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[135]), .B(A[135]), .Z(n946) );
  XOR U1420 ( .A(A[134]), .B(n947), .Z(O[134]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[134]), .B(A[134]), .Z(n948) );
  XOR U1423 ( .A(A[133]), .B(n949), .Z(O[133]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[133]), .B(A[133]), .Z(n950) );
  XOR U1426 ( .A(A[132]), .B(n951), .Z(O[132]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[132]), .B(A[132]), .Z(n952) );
  XOR U1429 ( .A(A[131]), .B(n953), .Z(O[131]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[131]), .B(A[131]), .Z(n954) );
  XOR U1432 ( .A(A[130]), .B(n955), .Z(O[130]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[130]), .B(A[130]), .Z(n956) );
  XOR U1435 ( .A(A[12]), .B(n957), .Z(O[12]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[12]), .B(A[12]), .Z(n958) );
  XOR U1438 ( .A(A[129]), .B(n959), .Z(O[129]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[129]), .B(A[129]), .Z(n960) );
  XOR U1441 ( .A(A[128]), .B(n961), .Z(O[128]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[128]), .B(A[128]), .Z(n962) );
  XOR U1444 ( .A(A[127]), .B(n963), .Z(O[127]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[127]), .B(A[127]), .Z(n964) );
  XOR U1447 ( .A(A[126]), .B(n965), .Z(O[126]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[126]), .B(A[126]), .Z(n966) );
  XOR U1450 ( .A(A[125]), .B(n967), .Z(O[125]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[125]), .B(A[125]), .Z(n968) );
  XOR U1453 ( .A(A[124]), .B(n969), .Z(O[124]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[124]), .B(A[124]), .Z(n970) );
  XOR U1456 ( .A(A[123]), .B(n971), .Z(O[123]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[123]), .B(A[123]), .Z(n972) );
  XOR U1459 ( .A(A[122]), .B(n973), .Z(O[122]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[122]), .B(A[122]), .Z(n974) );
  XOR U1462 ( .A(A[121]), .B(n975), .Z(O[121]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[121]), .B(A[121]), .Z(n976) );
  XOR U1465 ( .A(A[120]), .B(n977), .Z(O[120]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[120]), .B(A[120]), .Z(n978) );
  XOR U1468 ( .A(A[11]), .B(n979), .Z(O[11]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[11]), .B(A[11]), .Z(n980) );
  XOR U1471 ( .A(A[119]), .B(n981), .Z(O[119]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[119]), .B(A[119]), .Z(n982) );
  XOR U1474 ( .A(A[118]), .B(n983), .Z(O[118]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[118]), .B(A[118]), .Z(n984) );
  XOR U1477 ( .A(A[117]), .B(n985), .Z(O[117]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[117]), .B(A[117]), .Z(n986) );
  XOR U1480 ( .A(A[116]), .B(n987), .Z(O[116]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[116]), .B(A[116]), .Z(n988) );
  XOR U1483 ( .A(A[115]), .B(n989), .Z(O[115]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[115]), .B(A[115]), .Z(n990) );
  XOR U1486 ( .A(A[114]), .B(n991), .Z(O[114]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[114]), .B(A[114]), .Z(n992) );
  XOR U1489 ( .A(A[113]), .B(n993), .Z(O[113]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[113]), .B(A[113]), .Z(n994) );
  XOR U1492 ( .A(A[112]), .B(n995), .Z(O[112]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[112]), .B(A[112]), .Z(n996) );
  XOR U1495 ( .A(A[111]), .B(n997), .Z(O[111]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[111]), .B(A[111]), .Z(n998) );
  XOR U1498 ( .A(A[110]), .B(n999), .Z(O[110]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[110]), .B(A[110]), .Z(n1000) );
  XOR U1501 ( .A(A[10]), .B(n1001), .Z(O[10]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[10]), .B(A[10]), .Z(n1002) );
  XOR U1504 ( .A(A[109]), .B(n1003), .Z(O[109]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[109]), .B(A[109]), .Z(n1004) );
  XOR U1507 ( .A(A[108]), .B(n1005), .Z(O[108]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[108]), .B(A[108]), .Z(n1006) );
  XOR U1510 ( .A(A[107]), .B(n1007), .Z(O[107]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[107]), .B(A[107]), .Z(n1008) );
  XOR U1513 ( .A(A[106]), .B(n1009), .Z(O[106]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[106]), .B(A[106]), .Z(n1010) );
  XOR U1516 ( .A(A[105]), .B(n1011), .Z(O[105]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[105]), .B(A[105]), .Z(n1012) );
  XOR U1519 ( .A(A[104]), .B(n1013), .Z(O[104]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[104]), .B(A[104]), .Z(n1014) );
  XOR U1522 ( .A(A[103]), .B(n1015), .Z(O[103]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[103]), .B(A[103]), .Z(n1016) );
  XOR U1525 ( .A(A[102]), .B(n1017), .Z(O[102]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[102]), .B(A[102]), .Z(n1018) );
  XOR U1528 ( .A(A[101]), .B(n1019), .Z(O[101]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[101]), .B(A[101]), .Z(n1020) );
  XOR U1531 ( .A(A[100]), .B(n1021), .Z(O[100]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[100]), .B(A[100]), .Z(n1022) );
  XOR U1534 ( .A(A[0]), .B(n1023), .Z(O[0]) );
  AND U1535 ( .A(S), .B(n1024), .Z(n1023) );
  XOR U1536 ( .A(B[0]), .B(A[0]), .Z(n1024) );
endmodule


module MUX_N514_3 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_2580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module FA_11063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_11064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  ANDN U1 ( .B(CI), .A(S), .Z(CO) );
  XOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_11065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_11575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module ADD_N514_1_0 ( A, B, CI, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  input CI;
  output CO;

  wire   [513:1] C;

  FA_2580 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(1'b0), .B(B[0]), .CI(1'b0), .S(
        S[0]) );
  FA_11575 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), 
        .S(S[1]), .CO(C[2]) );
  FA_11574 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), 
        .S(S[2]), .CO(C[3]) );
  FA_11573 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), 
        .S(S[3]), .CO(C[4]) );
  FA_11572 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), 
        .S(S[4]), .CO(C[5]) );
  FA_11571 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), 
        .S(S[5]), .CO(C[6]) );
  FA_11570 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), 
        .S(S[6]), .CO(C[7]) );
  FA_11569 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), 
        .S(S[7]), .CO(C[8]) );
  FA_11568 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), 
        .S(S[8]), .CO(C[9]) );
  FA_11567 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), 
        .S(S[9]), .CO(C[10]) );
  FA_11566 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_11565 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_11564 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_11563 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_11562 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_11561 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_11560 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_11559 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_11558 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_11557 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_11556 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_11555 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_11554 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_11553 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_11552 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_11551 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_11550 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_11549 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_11548 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_11547 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_11546 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_11545 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_11544 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_11543 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_11542 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_11541 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_11540 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_11539 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_11538 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_11537 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_11536 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_11535 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_11534 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_11533 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_11532 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_11531 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_11530 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_11529 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_11528 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_11527 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_11526 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_11525 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_11524 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_11523 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_11522 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_11521 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_11520 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_11519 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_11518 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_11517 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_11516 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_11515 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_11514 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_11513 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_11512 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_11511 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_11510 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_11509 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_11508 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_11507 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_11506 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_11505 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_11504 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_11503 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_11502 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_11501 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_11500 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_11499 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_11498 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_11497 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_11496 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_11495 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_11494 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_11493 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_11492 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_11491 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_11490 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_11489 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_11488 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_11487 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_11486 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_11485 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_11484 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_11483 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_11482 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_11481 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_11480 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_11479 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_11478 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_11477 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_11476 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_11475 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_11474 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_11473 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_11472 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_11471 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_11470 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_11469 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_11468 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_11467 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_11466 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_11465 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_11464 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_11463 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_11462 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_11461 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_11460 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_11459 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_11458 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_11457 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_11456 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_11455 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_11454 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_11453 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_11452 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_11451 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_11450 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_11449 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_11448 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_11447 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_11446 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_11445 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_11444 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_11443 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_11442 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_11441 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_11440 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_11439 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_11438 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_11437 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_11436 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_11435 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_11434 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_11433 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_11432 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_11431 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_11430 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_11429 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_11428 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_11427 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_11426 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_11425 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_11424 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_11423 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_11422 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_11421 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_11420 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_11419 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_11418 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_11417 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_11416 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_11415 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_11414 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_11413 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_11412 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_11411 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_11410 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_11409 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_11408 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_11407 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_11406 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_11405 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_11404 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_11403 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_11402 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_11401 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_11400 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_11399 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_11398 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_11397 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_11396 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_11395 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_11394 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_11393 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_11392 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_11391 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_11390 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_11389 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_11388 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_11387 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_11386 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_11385 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_11384 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_11383 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_11382 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_11381 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_11380 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_11379 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_11378 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_11377 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_11376 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_11375 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_11374 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_11373 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_11372 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_11371 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_11370 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_11369 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_11368 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_11367 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_11366 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_11365 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_11364 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_11363 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_11362 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_11361 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_11360 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_11359 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_11358 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_11357 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_11356 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_11355 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_11354 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_11353 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_11352 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_11351 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_11350 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_11349 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_11348 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_11347 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_11346 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_11345 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_11344 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_11343 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_11342 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_11341 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_11340 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_11339 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_11338 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_11337 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_11336 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_11335 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_11334 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_11333 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_11332 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_11331 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_11330 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_11329 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_11328 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_11327 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_11326 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_11325 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_11324 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_11323 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_11322 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_11321 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_11320 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_11319 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_11318 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_11317 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_11316 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_11315 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_11314 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_11313 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_11312 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_11311 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_11310 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_11309 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_11308 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_11307 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_11306 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_11305 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_11304 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_11303 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_11302 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_11301 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_11300 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_11299 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_11298 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_11297 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_11296 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_11295 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_11294 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_11293 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_11292 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_11291 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_11290 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_11289 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_11288 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_11287 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_11286 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_11285 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_11284 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_11283 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_11282 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_11281 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_11280 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_11279 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_11278 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_11277 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_11276 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_11275 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_11274 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_11273 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_11272 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_11271 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_11270 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_11269 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_11268 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_11267 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_11266 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_11265 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_11264 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_11263 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_11262 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_11261 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_11260 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_11259 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_11258 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_11257 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_11256 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_11255 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_11254 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_11253 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_11252 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_11251 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_11250 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_11249 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_11248 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_11247 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_11246 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_11245 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_11244 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_11243 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_11242 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_11241 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_11240 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_11239 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_11238 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_11237 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_11236 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_11235 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_11234 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_11233 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_11232 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_11231 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_11230 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_11229 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_11228 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_11227 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_11226 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_11225 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_11224 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_11223 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_11222 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_11221 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_11220 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_11219 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_11218 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_11217 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_11216 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_11215 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_11214 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_11213 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_11212 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_11211 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_11210 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_11209 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_11208 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_11207 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_11206 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_11205 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_11204 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_11203 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_11202 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_11201 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_11200 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_11199 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_11198 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_11197 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_11196 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_11195 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_11194 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_11193 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_11192 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_11191 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_11190 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_11189 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_11188 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_11187 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_11186 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_11185 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_11184 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_11183 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_11182 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_11181 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_11180 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_11179 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_11178 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_11177 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_11176 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_11175 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_11174 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_11173 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_11172 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_11171 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_11170 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_11169 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_11168 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_11167 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_11166 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_11165 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_11164 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_11163 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_11162 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_11161 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_11160 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_11159 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_11158 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_11157 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_11156 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_11155 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_11154 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_11153 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_11152 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_11151 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_11150 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_11149 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_11148 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_11147 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_11146 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_11145 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_11144 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_11143 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_11142 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_11141 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_11140 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_11139 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_11138 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_11137 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_11136 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_11135 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_11134 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_11133 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_11132 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_11131 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_11130 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_11129 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_11128 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_11127 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_11126 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_11125 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_11124 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_11123 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_11122 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_11121 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_11120 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_11119 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_11118 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_11117 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_11116 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_11115 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_11114 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_11113 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_11112 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_11111 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_11110 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_11109 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_11108 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_11107 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_11106 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_11105 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_11104 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_11103 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_11102 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_11101 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_11100 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_11099 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_11098 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_11097 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_11096 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_11095 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_11094 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_11093 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_11092 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_11091 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_11090 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_11089 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_11088 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_11087 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_11086 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_11085 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_11084 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_11083 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_11082 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_11081 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_11080 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_11079 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_11078 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_11077 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_11076 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_11075 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_11074 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_11073 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_11072 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_11071 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_11070 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_11069 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_11068 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_11067 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_11066 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_11065 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_11064 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b0), .CI(C[512]), .S(S[512]), .CO(C[513]) );
  FA_11063 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b0), .CI(C[513]), .S(S[513]) );
endmodule


module FA_10549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_10550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_10551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_11062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N514_2 ( A, B, O );
  input [513:0] A;
  input [513:0] B;
  output O;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514;
  wire   [513:1] C;

  FA_11062 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n514), .CI(1'b1), 
        .CO(C[1]) );
  FA_11061 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n513), .CI(C[1]), 
        .CO(C[2]) );
  FA_11060 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n512), .CI(C[2]), 
        .CO(C[3]) );
  FA_11059 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n511), .CI(C[3]), 
        .CO(C[4]) );
  FA_11058 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n510), .CI(C[4]), 
        .CO(C[5]) );
  FA_11057 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n509), .CI(C[5]), 
        .CO(C[6]) );
  FA_11056 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n508), .CI(C[6]), 
        .CO(C[7]) );
  FA_11055 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n507), .CI(C[7]), 
        .CO(C[8]) );
  FA_11054 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n506), .CI(C[8]), 
        .CO(C[9]) );
  FA_11053 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n505), .CI(C[9]), 
        .CO(C[10]) );
  FA_11052 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n504), .CI(C[10]), 
        .CO(C[11]) );
  FA_11051 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n503), .CI(C[11]), 
        .CO(C[12]) );
  FA_11050 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n502), .CI(C[12]), 
        .CO(C[13]) );
  FA_11049 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n501), .CI(C[13]), 
        .CO(C[14]) );
  FA_11048 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n500), .CI(C[14]), 
        .CO(C[15]) );
  FA_11047 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n499), .CI(C[15]), 
        .CO(C[16]) );
  FA_11046 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n498), .CI(C[16]), 
        .CO(C[17]) );
  FA_11045 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n497), .CI(C[17]), 
        .CO(C[18]) );
  FA_11044 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n496), .CI(C[18]), 
        .CO(C[19]) );
  FA_11043 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n495), .CI(C[19]), 
        .CO(C[20]) );
  FA_11042 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n494), .CI(C[20]), 
        .CO(C[21]) );
  FA_11041 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n493), .CI(C[21]), 
        .CO(C[22]) );
  FA_11040 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n492), .CI(C[22]), 
        .CO(C[23]) );
  FA_11039 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n491), .CI(C[23]), 
        .CO(C[24]) );
  FA_11038 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n490), .CI(C[24]), 
        .CO(C[25]) );
  FA_11037 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n489), .CI(C[25]), 
        .CO(C[26]) );
  FA_11036 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n488), .CI(C[26]), 
        .CO(C[27]) );
  FA_11035 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n487), .CI(C[27]), 
        .CO(C[28]) );
  FA_11034 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n486), .CI(C[28]), 
        .CO(C[29]) );
  FA_11033 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n485), .CI(C[29]), 
        .CO(C[30]) );
  FA_11032 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n484), .CI(C[30]), 
        .CO(C[31]) );
  FA_11031 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n483), .CI(C[31]), 
        .CO(C[32]) );
  FA_11030 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n482), .CI(C[32]), 
        .CO(C[33]) );
  FA_11029 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n481), .CI(C[33]), 
        .CO(C[34]) );
  FA_11028 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n480), .CI(C[34]), 
        .CO(C[35]) );
  FA_11027 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n479), .CI(C[35]), 
        .CO(C[36]) );
  FA_11026 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n478), .CI(C[36]), 
        .CO(C[37]) );
  FA_11025 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n477), .CI(C[37]), 
        .CO(C[38]) );
  FA_11024 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n476), .CI(C[38]), 
        .CO(C[39]) );
  FA_11023 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n475), .CI(C[39]), 
        .CO(C[40]) );
  FA_11022 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n474), .CI(C[40]), 
        .CO(C[41]) );
  FA_11021 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n473), .CI(C[41]), 
        .CO(C[42]) );
  FA_11020 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n472), .CI(C[42]), 
        .CO(C[43]) );
  FA_11019 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n471), .CI(C[43]), 
        .CO(C[44]) );
  FA_11018 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n470), .CI(C[44]), 
        .CO(C[45]) );
  FA_11017 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n469), .CI(C[45]), 
        .CO(C[46]) );
  FA_11016 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n468), .CI(C[46]), 
        .CO(C[47]) );
  FA_11015 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n467), .CI(C[47]), 
        .CO(C[48]) );
  FA_11014 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n466), .CI(C[48]), 
        .CO(C[49]) );
  FA_11013 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n465), .CI(C[49]), 
        .CO(C[50]) );
  FA_11012 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n464), .CI(C[50]), 
        .CO(C[51]) );
  FA_11011 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n463), .CI(C[51]), 
        .CO(C[52]) );
  FA_11010 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n462), .CI(C[52]), 
        .CO(C[53]) );
  FA_11009 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n461), .CI(C[53]), 
        .CO(C[54]) );
  FA_11008 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n460), .CI(C[54]), 
        .CO(C[55]) );
  FA_11007 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n459), .CI(C[55]), 
        .CO(C[56]) );
  FA_11006 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n458), .CI(C[56]), 
        .CO(C[57]) );
  FA_11005 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n457), .CI(C[57]), 
        .CO(C[58]) );
  FA_11004 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n456), .CI(C[58]), 
        .CO(C[59]) );
  FA_11003 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n455), .CI(C[59]), 
        .CO(C[60]) );
  FA_11002 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n454), .CI(C[60]), 
        .CO(C[61]) );
  FA_11001 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n453), .CI(C[61]), 
        .CO(C[62]) );
  FA_11000 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n452), .CI(C[62]), 
        .CO(C[63]) );
  FA_10999 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n451), .CI(C[63]), 
        .CO(C[64]) );
  FA_10998 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n450), .CI(C[64]), 
        .CO(C[65]) );
  FA_10997 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n449), .CI(C[65]), 
        .CO(C[66]) );
  FA_10996 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n448), .CI(C[66]), 
        .CO(C[67]) );
  FA_10995 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n447), .CI(C[67]), 
        .CO(C[68]) );
  FA_10994 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n446), .CI(C[68]), 
        .CO(C[69]) );
  FA_10993 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n445), .CI(C[69]), 
        .CO(C[70]) );
  FA_10992 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n444), .CI(C[70]), 
        .CO(C[71]) );
  FA_10991 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n443), .CI(C[71]), 
        .CO(C[72]) );
  FA_10990 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n442), .CI(C[72]), 
        .CO(C[73]) );
  FA_10989 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n441), .CI(C[73]), 
        .CO(C[74]) );
  FA_10988 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n440), .CI(C[74]), 
        .CO(C[75]) );
  FA_10987 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n439), .CI(C[75]), 
        .CO(C[76]) );
  FA_10986 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n438), .CI(C[76]), 
        .CO(C[77]) );
  FA_10985 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n437), .CI(C[77]), 
        .CO(C[78]) );
  FA_10984 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n436), .CI(C[78]), 
        .CO(C[79]) );
  FA_10983 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n435), .CI(C[79]), 
        .CO(C[80]) );
  FA_10982 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n434), .CI(C[80]), 
        .CO(C[81]) );
  FA_10981 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n433), .CI(C[81]), 
        .CO(C[82]) );
  FA_10980 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n432), .CI(C[82]), 
        .CO(C[83]) );
  FA_10979 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n431), .CI(C[83]), 
        .CO(C[84]) );
  FA_10978 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n430), .CI(C[84]), 
        .CO(C[85]) );
  FA_10977 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n429), .CI(C[85]), 
        .CO(C[86]) );
  FA_10976 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n428), .CI(C[86]), 
        .CO(C[87]) );
  FA_10975 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n427), .CI(C[87]), 
        .CO(C[88]) );
  FA_10974 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n426), .CI(C[88]), 
        .CO(C[89]) );
  FA_10973 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n425), .CI(C[89]), 
        .CO(C[90]) );
  FA_10972 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n424), .CI(C[90]), 
        .CO(C[91]) );
  FA_10971 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n423), .CI(C[91]), 
        .CO(C[92]) );
  FA_10970 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n422), .CI(C[92]), 
        .CO(C[93]) );
  FA_10969 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n421), .CI(C[93]), 
        .CO(C[94]) );
  FA_10968 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n420), .CI(C[94]), 
        .CO(C[95]) );
  FA_10967 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n419), .CI(C[95]), 
        .CO(C[96]) );
  FA_10966 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n418), .CI(C[96]), 
        .CO(C[97]) );
  FA_10965 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n417), .CI(C[97]), 
        .CO(C[98]) );
  FA_10964 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n416), .CI(C[98]), 
        .CO(C[99]) );
  FA_10963 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n415), .CI(C[99]), 
        .CO(C[100]) );
  FA_10962 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n414), .CI(
        C[100]), .CO(C[101]) );
  FA_10961 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n413), .CI(
        C[101]), .CO(C[102]) );
  FA_10960 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n412), .CI(
        C[102]), .CO(C[103]) );
  FA_10959 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n411), .CI(
        C[103]), .CO(C[104]) );
  FA_10958 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n410), .CI(
        C[104]), .CO(C[105]) );
  FA_10957 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n409), .CI(
        C[105]), .CO(C[106]) );
  FA_10956 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n408), .CI(
        C[106]), .CO(C[107]) );
  FA_10955 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n407), .CI(
        C[107]), .CO(C[108]) );
  FA_10954 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n406), .CI(
        C[108]), .CO(C[109]) );
  FA_10953 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n405), .CI(
        C[109]), .CO(C[110]) );
  FA_10952 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n404), .CI(
        C[110]), .CO(C[111]) );
  FA_10951 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n403), .CI(
        C[111]), .CO(C[112]) );
  FA_10950 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n402), .CI(
        C[112]), .CO(C[113]) );
  FA_10949 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n401), .CI(
        C[113]), .CO(C[114]) );
  FA_10948 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n400), .CI(
        C[114]), .CO(C[115]) );
  FA_10947 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n399), .CI(
        C[115]), .CO(C[116]) );
  FA_10946 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n398), .CI(
        C[116]), .CO(C[117]) );
  FA_10945 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n397), .CI(
        C[117]), .CO(C[118]) );
  FA_10944 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n396), .CI(
        C[118]), .CO(C[119]) );
  FA_10943 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n395), .CI(
        C[119]), .CO(C[120]) );
  FA_10942 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n394), .CI(
        C[120]), .CO(C[121]) );
  FA_10941 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n393), .CI(
        C[121]), .CO(C[122]) );
  FA_10940 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n392), .CI(
        C[122]), .CO(C[123]) );
  FA_10939 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n391), .CI(
        C[123]), .CO(C[124]) );
  FA_10938 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n390), .CI(
        C[124]), .CO(C[125]) );
  FA_10937 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n389), .CI(
        C[125]), .CO(C[126]) );
  FA_10936 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n388), .CI(
        C[126]), .CO(C[127]) );
  FA_10935 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n387), .CI(
        C[127]), .CO(C[128]) );
  FA_10934 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n386), .CI(
        C[128]), .CO(C[129]) );
  FA_10933 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n385), .CI(
        C[129]), .CO(C[130]) );
  FA_10932 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n384), .CI(
        C[130]), .CO(C[131]) );
  FA_10931 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n383), .CI(
        C[131]), .CO(C[132]) );
  FA_10930 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n382), .CI(
        C[132]), .CO(C[133]) );
  FA_10929 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n381), .CI(
        C[133]), .CO(C[134]) );
  FA_10928 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n380), .CI(
        C[134]), .CO(C[135]) );
  FA_10927 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n379), .CI(
        C[135]), .CO(C[136]) );
  FA_10926 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n378), .CI(
        C[136]), .CO(C[137]) );
  FA_10925 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n377), .CI(
        C[137]), .CO(C[138]) );
  FA_10924 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n376), .CI(
        C[138]), .CO(C[139]) );
  FA_10923 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n375), .CI(
        C[139]), .CO(C[140]) );
  FA_10922 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n374), .CI(
        C[140]), .CO(C[141]) );
  FA_10921 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n373), .CI(
        C[141]), .CO(C[142]) );
  FA_10920 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n372), .CI(
        C[142]), .CO(C[143]) );
  FA_10919 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n371), .CI(
        C[143]), .CO(C[144]) );
  FA_10918 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n370), .CI(
        C[144]), .CO(C[145]) );
  FA_10917 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n369), .CI(
        C[145]), .CO(C[146]) );
  FA_10916 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n368), .CI(
        C[146]), .CO(C[147]) );
  FA_10915 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n367), .CI(
        C[147]), .CO(C[148]) );
  FA_10914 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n366), .CI(
        C[148]), .CO(C[149]) );
  FA_10913 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n365), .CI(
        C[149]), .CO(C[150]) );
  FA_10912 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n364), .CI(
        C[150]), .CO(C[151]) );
  FA_10911 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n363), .CI(
        C[151]), .CO(C[152]) );
  FA_10910 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n362), .CI(
        C[152]), .CO(C[153]) );
  FA_10909 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n361), .CI(
        C[153]), .CO(C[154]) );
  FA_10908 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n360), .CI(
        C[154]), .CO(C[155]) );
  FA_10907 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n359), .CI(
        C[155]), .CO(C[156]) );
  FA_10906 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n358), .CI(
        C[156]), .CO(C[157]) );
  FA_10905 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n357), .CI(
        C[157]), .CO(C[158]) );
  FA_10904 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n356), .CI(
        C[158]), .CO(C[159]) );
  FA_10903 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n355), .CI(
        C[159]), .CO(C[160]) );
  FA_10902 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n354), .CI(
        C[160]), .CO(C[161]) );
  FA_10901 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n353), .CI(
        C[161]), .CO(C[162]) );
  FA_10900 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n352), .CI(
        C[162]), .CO(C[163]) );
  FA_10899 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n351), .CI(
        C[163]), .CO(C[164]) );
  FA_10898 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n350), .CI(
        C[164]), .CO(C[165]) );
  FA_10897 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n349), .CI(
        C[165]), .CO(C[166]) );
  FA_10896 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n348), .CI(
        C[166]), .CO(C[167]) );
  FA_10895 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n347), .CI(
        C[167]), .CO(C[168]) );
  FA_10894 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n346), .CI(
        C[168]), .CO(C[169]) );
  FA_10893 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n345), .CI(
        C[169]), .CO(C[170]) );
  FA_10892 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n344), .CI(
        C[170]), .CO(C[171]) );
  FA_10891 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n343), .CI(
        C[171]), .CO(C[172]) );
  FA_10890 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n342), .CI(
        C[172]), .CO(C[173]) );
  FA_10889 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n341), .CI(
        C[173]), .CO(C[174]) );
  FA_10888 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n340), .CI(
        C[174]), .CO(C[175]) );
  FA_10887 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n339), .CI(
        C[175]), .CO(C[176]) );
  FA_10886 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n338), .CI(
        C[176]), .CO(C[177]) );
  FA_10885 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n337), .CI(
        C[177]), .CO(C[178]) );
  FA_10884 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n336), .CI(
        C[178]), .CO(C[179]) );
  FA_10883 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n335), .CI(
        C[179]), .CO(C[180]) );
  FA_10882 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n334), .CI(
        C[180]), .CO(C[181]) );
  FA_10881 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n333), .CI(
        C[181]), .CO(C[182]) );
  FA_10880 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n332), .CI(
        C[182]), .CO(C[183]) );
  FA_10879 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n331), .CI(
        C[183]), .CO(C[184]) );
  FA_10878 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n330), .CI(
        C[184]), .CO(C[185]) );
  FA_10877 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n329), .CI(
        C[185]), .CO(C[186]) );
  FA_10876 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n328), .CI(
        C[186]), .CO(C[187]) );
  FA_10875 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n327), .CI(
        C[187]), .CO(C[188]) );
  FA_10874 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n326), .CI(
        C[188]), .CO(C[189]) );
  FA_10873 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n325), .CI(
        C[189]), .CO(C[190]) );
  FA_10872 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n324), .CI(
        C[190]), .CO(C[191]) );
  FA_10871 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n323), .CI(
        C[191]), .CO(C[192]) );
  FA_10870 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n322), .CI(
        C[192]), .CO(C[193]) );
  FA_10869 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n321), .CI(
        C[193]), .CO(C[194]) );
  FA_10868 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n320), .CI(
        C[194]), .CO(C[195]) );
  FA_10867 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n319), .CI(
        C[195]), .CO(C[196]) );
  FA_10866 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n318), .CI(
        C[196]), .CO(C[197]) );
  FA_10865 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n317), .CI(
        C[197]), .CO(C[198]) );
  FA_10864 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n316), .CI(
        C[198]), .CO(C[199]) );
  FA_10863 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n315), .CI(
        C[199]), .CO(C[200]) );
  FA_10862 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n314), .CI(
        C[200]), .CO(C[201]) );
  FA_10861 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n313), .CI(
        C[201]), .CO(C[202]) );
  FA_10860 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n312), .CI(
        C[202]), .CO(C[203]) );
  FA_10859 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n311), .CI(
        C[203]), .CO(C[204]) );
  FA_10858 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n310), .CI(
        C[204]), .CO(C[205]) );
  FA_10857 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n309), .CI(
        C[205]), .CO(C[206]) );
  FA_10856 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n308), .CI(
        C[206]), .CO(C[207]) );
  FA_10855 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n307), .CI(
        C[207]), .CO(C[208]) );
  FA_10854 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n306), .CI(
        C[208]), .CO(C[209]) );
  FA_10853 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n305), .CI(
        C[209]), .CO(C[210]) );
  FA_10852 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n304), .CI(
        C[210]), .CO(C[211]) );
  FA_10851 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n303), .CI(
        C[211]), .CO(C[212]) );
  FA_10850 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n302), .CI(
        C[212]), .CO(C[213]) );
  FA_10849 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n301), .CI(
        C[213]), .CO(C[214]) );
  FA_10848 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n300), .CI(
        C[214]), .CO(C[215]) );
  FA_10847 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n299), .CI(
        C[215]), .CO(C[216]) );
  FA_10846 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n298), .CI(
        C[216]), .CO(C[217]) );
  FA_10845 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n297), .CI(
        C[217]), .CO(C[218]) );
  FA_10844 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n296), .CI(
        C[218]), .CO(C[219]) );
  FA_10843 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n295), .CI(
        C[219]), .CO(C[220]) );
  FA_10842 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n294), .CI(
        C[220]), .CO(C[221]) );
  FA_10841 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n293), .CI(
        C[221]), .CO(C[222]) );
  FA_10840 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n292), .CI(
        C[222]), .CO(C[223]) );
  FA_10839 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n291), .CI(
        C[223]), .CO(C[224]) );
  FA_10838 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n290), .CI(
        C[224]), .CO(C[225]) );
  FA_10837 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n289), .CI(
        C[225]), .CO(C[226]) );
  FA_10836 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n288), .CI(
        C[226]), .CO(C[227]) );
  FA_10835 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n287), .CI(
        C[227]), .CO(C[228]) );
  FA_10834 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n286), .CI(
        C[228]), .CO(C[229]) );
  FA_10833 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n285), .CI(
        C[229]), .CO(C[230]) );
  FA_10832 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n284), .CI(
        C[230]), .CO(C[231]) );
  FA_10831 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n283), .CI(
        C[231]), .CO(C[232]) );
  FA_10830 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n282), .CI(
        C[232]), .CO(C[233]) );
  FA_10829 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n281), .CI(
        C[233]), .CO(C[234]) );
  FA_10828 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n280), .CI(
        C[234]), .CO(C[235]) );
  FA_10827 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n279), .CI(
        C[235]), .CO(C[236]) );
  FA_10826 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n278), .CI(
        C[236]), .CO(C[237]) );
  FA_10825 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n277), .CI(
        C[237]), .CO(C[238]) );
  FA_10824 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n276), .CI(
        C[238]), .CO(C[239]) );
  FA_10823 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n275), .CI(
        C[239]), .CO(C[240]) );
  FA_10822 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n274), .CI(
        C[240]), .CO(C[241]) );
  FA_10821 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n273), .CI(
        C[241]), .CO(C[242]) );
  FA_10820 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n272), .CI(
        C[242]), .CO(C[243]) );
  FA_10819 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n271), .CI(
        C[243]), .CO(C[244]) );
  FA_10818 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n270), .CI(
        C[244]), .CO(C[245]) );
  FA_10817 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n269), .CI(
        C[245]), .CO(C[246]) );
  FA_10816 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n268), .CI(
        C[246]), .CO(C[247]) );
  FA_10815 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n267), .CI(
        C[247]), .CO(C[248]) );
  FA_10814 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n266), .CI(
        C[248]), .CO(C[249]) );
  FA_10813 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n265), .CI(
        C[249]), .CO(C[250]) );
  FA_10812 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n264), .CI(
        C[250]), .CO(C[251]) );
  FA_10811 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n263), .CI(
        C[251]), .CO(C[252]) );
  FA_10810 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n262), .CI(
        C[252]), .CO(C[253]) );
  FA_10809 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n261), .CI(
        C[253]), .CO(C[254]) );
  FA_10808 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n260), .CI(
        C[254]), .CO(C[255]) );
  FA_10807 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n259), .CI(
        C[255]), .CO(C[256]) );
  FA_10806 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n258), .CI(
        C[256]), .CO(C[257]) );
  FA_10805 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n257), .CI(
        C[257]), .CO(C[258]) );
  FA_10804 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n256), .CI(
        C[258]), .CO(C[259]) );
  FA_10803 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n255), .CI(
        C[259]), .CO(C[260]) );
  FA_10802 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n254), .CI(
        C[260]), .CO(C[261]) );
  FA_10801 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n253), .CI(
        C[261]), .CO(C[262]) );
  FA_10800 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n252), .CI(
        C[262]), .CO(C[263]) );
  FA_10799 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n251), .CI(
        C[263]), .CO(C[264]) );
  FA_10798 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n250), .CI(
        C[264]), .CO(C[265]) );
  FA_10797 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n249), .CI(
        C[265]), .CO(C[266]) );
  FA_10796 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n248), .CI(
        C[266]), .CO(C[267]) );
  FA_10795 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n247), .CI(
        C[267]), .CO(C[268]) );
  FA_10794 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n246), .CI(
        C[268]), .CO(C[269]) );
  FA_10793 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n245), .CI(
        C[269]), .CO(C[270]) );
  FA_10792 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n244), .CI(
        C[270]), .CO(C[271]) );
  FA_10791 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n243), .CI(
        C[271]), .CO(C[272]) );
  FA_10790 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n242), .CI(
        C[272]), .CO(C[273]) );
  FA_10789 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n241), .CI(
        C[273]), .CO(C[274]) );
  FA_10788 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n240), .CI(
        C[274]), .CO(C[275]) );
  FA_10787 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n239), .CI(
        C[275]), .CO(C[276]) );
  FA_10786 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n238), .CI(
        C[276]), .CO(C[277]) );
  FA_10785 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n237), .CI(
        C[277]), .CO(C[278]) );
  FA_10784 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n236), .CI(
        C[278]), .CO(C[279]) );
  FA_10783 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n235), .CI(
        C[279]), .CO(C[280]) );
  FA_10782 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n234), .CI(
        C[280]), .CO(C[281]) );
  FA_10781 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n233), .CI(
        C[281]), .CO(C[282]) );
  FA_10780 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n232), .CI(
        C[282]), .CO(C[283]) );
  FA_10779 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n231), .CI(
        C[283]), .CO(C[284]) );
  FA_10778 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n230), .CI(
        C[284]), .CO(C[285]) );
  FA_10777 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n229), .CI(
        C[285]), .CO(C[286]) );
  FA_10776 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n228), .CI(
        C[286]), .CO(C[287]) );
  FA_10775 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n227), .CI(
        C[287]), .CO(C[288]) );
  FA_10774 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n226), .CI(
        C[288]), .CO(C[289]) );
  FA_10773 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n225), .CI(
        C[289]), .CO(C[290]) );
  FA_10772 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n224), .CI(
        C[290]), .CO(C[291]) );
  FA_10771 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n223), .CI(
        C[291]), .CO(C[292]) );
  FA_10770 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n222), .CI(
        C[292]), .CO(C[293]) );
  FA_10769 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n221), .CI(
        C[293]), .CO(C[294]) );
  FA_10768 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n220), .CI(
        C[294]), .CO(C[295]) );
  FA_10767 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n219), .CI(
        C[295]), .CO(C[296]) );
  FA_10766 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n218), .CI(
        C[296]), .CO(C[297]) );
  FA_10765 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n217), .CI(
        C[297]), .CO(C[298]) );
  FA_10764 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n216), .CI(
        C[298]), .CO(C[299]) );
  FA_10763 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n215), .CI(
        C[299]), .CO(C[300]) );
  FA_10762 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n214), .CI(
        C[300]), .CO(C[301]) );
  FA_10761 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n213), .CI(
        C[301]), .CO(C[302]) );
  FA_10760 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n212), .CI(
        C[302]), .CO(C[303]) );
  FA_10759 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n211), .CI(
        C[303]), .CO(C[304]) );
  FA_10758 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n210), .CI(
        C[304]), .CO(C[305]) );
  FA_10757 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n209), .CI(
        C[305]), .CO(C[306]) );
  FA_10756 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n208), .CI(
        C[306]), .CO(C[307]) );
  FA_10755 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n207), .CI(
        C[307]), .CO(C[308]) );
  FA_10754 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n206), .CI(
        C[308]), .CO(C[309]) );
  FA_10753 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n205), .CI(
        C[309]), .CO(C[310]) );
  FA_10752 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n204), .CI(
        C[310]), .CO(C[311]) );
  FA_10751 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n203), .CI(
        C[311]), .CO(C[312]) );
  FA_10750 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n202), .CI(
        C[312]), .CO(C[313]) );
  FA_10749 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n201), .CI(
        C[313]), .CO(C[314]) );
  FA_10748 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n200), .CI(
        C[314]), .CO(C[315]) );
  FA_10747 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n199), .CI(
        C[315]), .CO(C[316]) );
  FA_10746 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n198), .CI(
        C[316]), .CO(C[317]) );
  FA_10745 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n197), .CI(
        C[317]), .CO(C[318]) );
  FA_10744 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n196), .CI(
        C[318]), .CO(C[319]) );
  FA_10743 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n195), .CI(
        C[319]), .CO(C[320]) );
  FA_10742 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n194), .CI(
        C[320]), .CO(C[321]) );
  FA_10741 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n193), .CI(
        C[321]), .CO(C[322]) );
  FA_10740 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n192), .CI(
        C[322]), .CO(C[323]) );
  FA_10739 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n191), .CI(
        C[323]), .CO(C[324]) );
  FA_10738 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n190), .CI(
        C[324]), .CO(C[325]) );
  FA_10737 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n189), .CI(
        C[325]), .CO(C[326]) );
  FA_10736 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n188), .CI(
        C[326]), .CO(C[327]) );
  FA_10735 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n187), .CI(
        C[327]), .CO(C[328]) );
  FA_10734 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n186), .CI(
        C[328]), .CO(C[329]) );
  FA_10733 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n185), .CI(
        C[329]), .CO(C[330]) );
  FA_10732 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n184), .CI(
        C[330]), .CO(C[331]) );
  FA_10731 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n183), .CI(
        C[331]), .CO(C[332]) );
  FA_10730 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n182), .CI(
        C[332]), .CO(C[333]) );
  FA_10729 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n181), .CI(
        C[333]), .CO(C[334]) );
  FA_10728 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n180), .CI(
        C[334]), .CO(C[335]) );
  FA_10727 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n179), .CI(
        C[335]), .CO(C[336]) );
  FA_10726 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n178), .CI(
        C[336]), .CO(C[337]) );
  FA_10725 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n177), .CI(
        C[337]), .CO(C[338]) );
  FA_10724 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n176), .CI(
        C[338]), .CO(C[339]) );
  FA_10723 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n175), .CI(
        C[339]), .CO(C[340]) );
  FA_10722 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n174), .CI(
        C[340]), .CO(C[341]) );
  FA_10721 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n173), .CI(
        C[341]), .CO(C[342]) );
  FA_10720 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n172), .CI(
        C[342]), .CO(C[343]) );
  FA_10719 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n171), .CI(
        C[343]), .CO(C[344]) );
  FA_10718 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n170), .CI(
        C[344]), .CO(C[345]) );
  FA_10717 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n169), .CI(
        C[345]), .CO(C[346]) );
  FA_10716 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n168), .CI(
        C[346]), .CO(C[347]) );
  FA_10715 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n167), .CI(
        C[347]), .CO(C[348]) );
  FA_10714 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n166), .CI(
        C[348]), .CO(C[349]) );
  FA_10713 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n165), .CI(
        C[349]), .CO(C[350]) );
  FA_10712 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n164), .CI(
        C[350]), .CO(C[351]) );
  FA_10711 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n163), .CI(
        C[351]), .CO(C[352]) );
  FA_10710 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n162), .CI(
        C[352]), .CO(C[353]) );
  FA_10709 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n161), .CI(
        C[353]), .CO(C[354]) );
  FA_10708 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n160), .CI(
        C[354]), .CO(C[355]) );
  FA_10707 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n159), .CI(
        C[355]), .CO(C[356]) );
  FA_10706 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n158), .CI(
        C[356]), .CO(C[357]) );
  FA_10705 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n157), .CI(
        C[357]), .CO(C[358]) );
  FA_10704 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n156), .CI(
        C[358]), .CO(C[359]) );
  FA_10703 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n155), .CI(
        C[359]), .CO(C[360]) );
  FA_10702 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n154), .CI(
        C[360]), .CO(C[361]) );
  FA_10701 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n153), .CI(
        C[361]), .CO(C[362]) );
  FA_10700 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n152), .CI(
        C[362]), .CO(C[363]) );
  FA_10699 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n151), .CI(
        C[363]), .CO(C[364]) );
  FA_10698 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n150), .CI(
        C[364]), .CO(C[365]) );
  FA_10697 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n149), .CI(
        C[365]), .CO(C[366]) );
  FA_10696 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n148), .CI(
        C[366]), .CO(C[367]) );
  FA_10695 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n147), .CI(
        C[367]), .CO(C[368]) );
  FA_10694 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n146), .CI(
        C[368]), .CO(C[369]) );
  FA_10693 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n145), .CI(
        C[369]), .CO(C[370]) );
  FA_10692 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n144), .CI(
        C[370]), .CO(C[371]) );
  FA_10691 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n143), .CI(
        C[371]), .CO(C[372]) );
  FA_10690 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n142), .CI(
        C[372]), .CO(C[373]) );
  FA_10689 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n141), .CI(
        C[373]), .CO(C[374]) );
  FA_10688 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n140), .CI(
        C[374]), .CO(C[375]) );
  FA_10687 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n139), .CI(
        C[375]), .CO(C[376]) );
  FA_10686 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n138), .CI(
        C[376]), .CO(C[377]) );
  FA_10685 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n137), .CI(
        C[377]), .CO(C[378]) );
  FA_10684 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n136), .CI(
        C[378]), .CO(C[379]) );
  FA_10683 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n135), .CI(
        C[379]), .CO(C[380]) );
  FA_10682 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n134), .CI(
        C[380]), .CO(C[381]) );
  FA_10681 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n133), .CI(
        C[381]), .CO(C[382]) );
  FA_10680 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n132), .CI(
        C[382]), .CO(C[383]) );
  FA_10679 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n131), .CI(
        C[383]), .CO(C[384]) );
  FA_10678 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n130), .CI(
        C[384]), .CO(C[385]) );
  FA_10677 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n129), .CI(
        C[385]), .CO(C[386]) );
  FA_10676 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n128), .CI(
        C[386]), .CO(C[387]) );
  FA_10675 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n127), .CI(
        C[387]), .CO(C[388]) );
  FA_10674 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n126), .CI(
        C[388]), .CO(C[389]) );
  FA_10673 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n125), .CI(
        C[389]), .CO(C[390]) );
  FA_10672 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n124), .CI(
        C[390]), .CO(C[391]) );
  FA_10671 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n123), .CI(
        C[391]), .CO(C[392]) );
  FA_10670 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n122), .CI(
        C[392]), .CO(C[393]) );
  FA_10669 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n121), .CI(
        C[393]), .CO(C[394]) );
  FA_10668 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n120), .CI(
        C[394]), .CO(C[395]) );
  FA_10667 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n119), .CI(
        C[395]), .CO(C[396]) );
  FA_10666 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n118), .CI(
        C[396]), .CO(C[397]) );
  FA_10665 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n117), .CI(
        C[397]), .CO(C[398]) );
  FA_10664 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n116), .CI(
        C[398]), .CO(C[399]) );
  FA_10663 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n115), .CI(
        C[399]), .CO(C[400]) );
  FA_10662 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n114), .CI(
        C[400]), .CO(C[401]) );
  FA_10661 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n113), .CI(
        C[401]), .CO(C[402]) );
  FA_10660 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n112), .CI(
        C[402]), .CO(C[403]) );
  FA_10659 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n111), .CI(
        C[403]), .CO(C[404]) );
  FA_10658 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n110), .CI(
        C[404]), .CO(C[405]) );
  FA_10657 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n109), .CI(
        C[405]), .CO(C[406]) );
  FA_10656 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n108), .CI(
        C[406]), .CO(C[407]) );
  FA_10655 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n107), .CI(
        C[407]), .CO(C[408]) );
  FA_10654 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n106), .CI(
        C[408]), .CO(C[409]) );
  FA_10653 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n105), .CI(
        C[409]), .CO(C[410]) );
  FA_10652 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n104), .CI(
        C[410]), .CO(C[411]) );
  FA_10651 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n103), .CI(
        C[411]), .CO(C[412]) );
  FA_10650 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n102), .CI(
        C[412]), .CO(C[413]) );
  FA_10649 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n101), .CI(
        C[413]), .CO(C[414]) );
  FA_10648 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n100), .CI(
        C[414]), .CO(C[415]) );
  FA_10647 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n99), .CI(C[415]), .CO(C[416]) );
  FA_10646 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n98), .CI(C[416]), .CO(C[417]) );
  FA_10645 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n97), .CI(C[417]), .CO(C[418]) );
  FA_10644 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n96), .CI(C[418]), .CO(C[419]) );
  FA_10643 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n95), .CI(C[419]), .CO(C[420]) );
  FA_10642 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n94), .CI(C[420]), .CO(C[421]) );
  FA_10641 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n93), .CI(C[421]), .CO(C[422]) );
  FA_10640 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n92), .CI(C[422]), .CO(C[423]) );
  FA_10639 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n91), .CI(C[423]), .CO(C[424]) );
  FA_10638 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n90), .CI(C[424]), .CO(C[425]) );
  FA_10637 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n89), .CI(C[425]), .CO(C[426]) );
  FA_10636 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n88), .CI(C[426]), .CO(C[427]) );
  FA_10635 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n87), .CI(C[427]), .CO(C[428]) );
  FA_10634 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n86), .CI(C[428]), .CO(C[429]) );
  FA_10633 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n85), .CI(C[429]), .CO(C[430]) );
  FA_10632 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n84), .CI(C[430]), .CO(C[431]) );
  FA_10631 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n83), .CI(C[431]), .CO(C[432]) );
  FA_10630 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n82), .CI(C[432]), .CO(C[433]) );
  FA_10629 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n81), .CI(C[433]), .CO(C[434]) );
  FA_10628 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n80), .CI(C[434]), .CO(C[435]) );
  FA_10627 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n79), .CI(C[435]), .CO(C[436]) );
  FA_10626 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n78), .CI(C[436]), .CO(C[437]) );
  FA_10625 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n77), .CI(C[437]), .CO(C[438]) );
  FA_10624 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n76), .CI(C[438]), .CO(C[439]) );
  FA_10623 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n75), .CI(C[439]), .CO(C[440]) );
  FA_10622 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n74), .CI(C[440]), .CO(C[441]) );
  FA_10621 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n73), .CI(C[441]), .CO(C[442]) );
  FA_10620 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n72), .CI(C[442]), .CO(C[443]) );
  FA_10619 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n71), .CI(C[443]), .CO(C[444]) );
  FA_10618 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n70), .CI(C[444]), .CO(C[445]) );
  FA_10617 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n69), .CI(C[445]), .CO(C[446]) );
  FA_10616 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n68), .CI(C[446]), .CO(C[447]) );
  FA_10615 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n67), .CI(C[447]), .CO(C[448]) );
  FA_10614 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n66), .CI(C[448]), .CO(C[449]) );
  FA_10613 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n65), .CI(C[449]), .CO(C[450]) );
  FA_10612 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n64), .CI(C[450]), .CO(C[451]) );
  FA_10611 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n63), .CI(C[451]), .CO(C[452]) );
  FA_10610 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n62), .CI(C[452]), .CO(C[453]) );
  FA_10609 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n61), .CI(C[453]), .CO(C[454]) );
  FA_10608 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n60), .CI(C[454]), .CO(C[455]) );
  FA_10607 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n59), .CI(C[455]), .CO(C[456]) );
  FA_10606 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n58), .CI(C[456]), .CO(C[457]) );
  FA_10605 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n57), .CI(C[457]), .CO(C[458]) );
  FA_10604 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n56), .CI(C[458]), .CO(C[459]) );
  FA_10603 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n55), .CI(C[459]), .CO(C[460]) );
  FA_10602 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n54), .CI(C[460]), .CO(C[461]) );
  FA_10601 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n53), .CI(C[461]), .CO(C[462]) );
  FA_10600 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n52), .CI(C[462]), .CO(C[463]) );
  FA_10599 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n51), .CI(C[463]), .CO(C[464]) );
  FA_10598 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n50), .CI(C[464]), .CO(C[465]) );
  FA_10597 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n49), .CI(C[465]), .CO(C[466]) );
  FA_10596 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n48), .CI(C[466]), .CO(C[467]) );
  FA_10595 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n47), .CI(C[467]), .CO(C[468]) );
  FA_10594 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n46), .CI(C[468]), .CO(C[469]) );
  FA_10593 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n45), .CI(C[469]), .CO(C[470]) );
  FA_10592 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n44), .CI(C[470]), .CO(C[471]) );
  FA_10591 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n43), .CI(C[471]), .CO(C[472]) );
  FA_10590 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n42), .CI(C[472]), .CO(C[473]) );
  FA_10589 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n41), .CI(C[473]), .CO(C[474]) );
  FA_10588 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n40), .CI(C[474]), .CO(C[475]) );
  FA_10587 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n39), .CI(C[475]), .CO(C[476]) );
  FA_10586 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n38), .CI(C[476]), .CO(C[477]) );
  FA_10585 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n37), .CI(C[477]), .CO(C[478]) );
  FA_10584 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n36), .CI(C[478]), .CO(C[479]) );
  FA_10583 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n35), .CI(C[479]), .CO(C[480]) );
  FA_10582 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n34), .CI(C[480]), .CO(C[481]) );
  FA_10581 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n33), .CI(C[481]), .CO(C[482]) );
  FA_10580 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n32), .CI(C[482]), .CO(C[483]) );
  FA_10579 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n31), .CI(C[483]), .CO(C[484]) );
  FA_10578 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n30), .CI(C[484]), .CO(C[485]) );
  FA_10577 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n29), .CI(C[485]), .CO(C[486]) );
  FA_10576 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n28), .CI(C[486]), .CO(C[487]) );
  FA_10575 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n27), .CI(C[487]), .CO(C[488]) );
  FA_10574 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n26), .CI(C[488]), .CO(C[489]) );
  FA_10573 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n25), .CI(C[489]), .CO(C[490]) );
  FA_10572 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n24), .CI(C[490]), .CO(C[491]) );
  FA_10571 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n23), .CI(C[491]), .CO(C[492]) );
  FA_10570 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n22), .CI(C[492]), .CO(C[493]) );
  FA_10569 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n21), .CI(C[493]), .CO(C[494]) );
  FA_10568 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n20), .CI(C[494]), .CO(C[495]) );
  FA_10567 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n19), .CI(C[495]), .CO(C[496]) );
  FA_10566 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n18), .CI(C[496]), .CO(C[497]) );
  FA_10565 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n17), .CI(C[497]), .CO(C[498]) );
  FA_10564 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n16), .CI(C[498]), .CO(C[499]) );
  FA_10563 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n15), .CI(C[499]), .CO(C[500]) );
  FA_10562 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n14), .CI(C[500]), .CO(C[501]) );
  FA_10561 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n13), .CI(C[501]), .CO(C[502]) );
  FA_10560 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n12), .CI(C[502]), .CO(C[503]) );
  FA_10559 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n11), .CI(C[503]), .CO(C[504]) );
  FA_10558 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n10), .CI(C[504]), .CO(C[505]) );
  FA_10557 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n9), .CI(C[505]), 
        .CO(C[506]) );
  FA_10556 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n8), .CI(C[506]), 
        .CO(C[507]) );
  FA_10555 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n7), .CI(C[507]), 
        .CO(C[508]) );
  FA_10554 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n6), .CI(C[508]), 
        .CO(C[509]) );
  FA_10553 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n5), .CI(C[509]), 
        .CO(C[510]) );
  FA_10552 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n4), .CI(C[510]), 
        .CO(C[511]) );
  FA_10551 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n3), .CI(C[511]), 
        .CO(C[512]) );
  FA_10550 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .CO(
        C[513]) );
  FA_10549 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b1), .CI(C[513]), .CO(O) );
  IV U2 ( .A(B[415]), .Z(n99) );
  IV U3 ( .A(B[416]), .Z(n98) );
  IV U4 ( .A(B[417]), .Z(n97) );
  IV U5 ( .A(B[418]), .Z(n96) );
  IV U6 ( .A(B[419]), .Z(n95) );
  IV U7 ( .A(B[420]), .Z(n94) );
  IV U8 ( .A(B[421]), .Z(n93) );
  IV U9 ( .A(B[422]), .Z(n92) );
  IV U10 ( .A(B[423]), .Z(n91) );
  IV U11 ( .A(B[424]), .Z(n90) );
  IV U12 ( .A(B[505]), .Z(n9) );
  IV U13 ( .A(B[425]), .Z(n89) );
  IV U14 ( .A(B[426]), .Z(n88) );
  IV U15 ( .A(B[427]), .Z(n87) );
  IV U16 ( .A(B[428]), .Z(n86) );
  IV U17 ( .A(B[429]), .Z(n85) );
  IV U18 ( .A(B[430]), .Z(n84) );
  IV U19 ( .A(B[431]), .Z(n83) );
  IV U20 ( .A(B[432]), .Z(n82) );
  IV U21 ( .A(B[433]), .Z(n81) );
  IV U22 ( .A(B[434]), .Z(n80) );
  IV U23 ( .A(B[506]), .Z(n8) );
  IV U24 ( .A(B[435]), .Z(n79) );
  IV U25 ( .A(B[436]), .Z(n78) );
  IV U26 ( .A(B[437]), .Z(n77) );
  IV U27 ( .A(B[438]), .Z(n76) );
  IV U28 ( .A(B[439]), .Z(n75) );
  IV U29 ( .A(B[440]), .Z(n74) );
  IV U30 ( .A(B[441]), .Z(n73) );
  IV U31 ( .A(B[442]), .Z(n72) );
  IV U32 ( .A(B[443]), .Z(n71) );
  IV U33 ( .A(B[444]), .Z(n70) );
  IV U34 ( .A(B[507]), .Z(n7) );
  IV U35 ( .A(B[445]), .Z(n69) );
  IV U36 ( .A(B[446]), .Z(n68) );
  IV U37 ( .A(B[447]), .Z(n67) );
  IV U38 ( .A(B[448]), .Z(n66) );
  IV U39 ( .A(B[449]), .Z(n65) );
  IV U40 ( .A(B[450]), .Z(n64) );
  IV U41 ( .A(B[451]), .Z(n63) );
  IV U42 ( .A(B[452]), .Z(n62) );
  IV U43 ( .A(B[453]), .Z(n61) );
  IV U44 ( .A(B[454]), .Z(n60) );
  IV U45 ( .A(B[508]), .Z(n6) );
  IV U46 ( .A(B[455]), .Z(n59) );
  IV U47 ( .A(B[456]), .Z(n58) );
  IV U48 ( .A(B[457]), .Z(n57) );
  IV U49 ( .A(B[458]), .Z(n56) );
  IV U50 ( .A(B[459]), .Z(n55) );
  IV U51 ( .A(B[460]), .Z(n54) );
  IV U52 ( .A(B[461]), .Z(n53) );
  IV U53 ( .A(B[462]), .Z(n52) );
  IV U54 ( .A(B[0]), .Z(n514) );
  IV U55 ( .A(B[1]), .Z(n513) );
  IV U56 ( .A(B[2]), .Z(n512) );
  IV U57 ( .A(B[3]), .Z(n511) );
  IV U58 ( .A(B[4]), .Z(n510) );
  IV U59 ( .A(B[463]), .Z(n51) );
  IV U60 ( .A(B[5]), .Z(n509) );
  IV U61 ( .A(B[6]), .Z(n508) );
  IV U62 ( .A(B[7]), .Z(n507) );
  IV U63 ( .A(B[8]), .Z(n506) );
  IV U64 ( .A(B[9]), .Z(n505) );
  IV U65 ( .A(B[10]), .Z(n504) );
  IV U66 ( .A(B[11]), .Z(n503) );
  IV U67 ( .A(B[12]), .Z(n502) );
  IV U68 ( .A(B[13]), .Z(n501) );
  IV U69 ( .A(B[14]), .Z(n500) );
  IV U70 ( .A(B[464]), .Z(n50) );
  IV U71 ( .A(B[509]), .Z(n5) );
  IV U72 ( .A(B[15]), .Z(n499) );
  IV U73 ( .A(B[16]), .Z(n498) );
  IV U74 ( .A(B[17]), .Z(n497) );
  IV U75 ( .A(B[18]), .Z(n496) );
  IV U76 ( .A(B[19]), .Z(n495) );
  IV U77 ( .A(B[20]), .Z(n494) );
  IV U78 ( .A(B[21]), .Z(n493) );
  IV U79 ( .A(B[22]), .Z(n492) );
  IV U80 ( .A(B[23]), .Z(n491) );
  IV U81 ( .A(B[24]), .Z(n490) );
  IV U82 ( .A(B[465]), .Z(n49) );
  IV U83 ( .A(B[25]), .Z(n489) );
  IV U84 ( .A(B[26]), .Z(n488) );
  IV U85 ( .A(B[27]), .Z(n487) );
  IV U86 ( .A(B[28]), .Z(n486) );
  IV U87 ( .A(B[29]), .Z(n485) );
  IV U88 ( .A(B[30]), .Z(n484) );
  IV U89 ( .A(B[31]), .Z(n483) );
  IV U90 ( .A(B[32]), .Z(n482) );
  IV U91 ( .A(B[33]), .Z(n481) );
  IV U92 ( .A(B[34]), .Z(n480) );
  IV U93 ( .A(B[466]), .Z(n48) );
  IV U94 ( .A(B[35]), .Z(n479) );
  IV U95 ( .A(B[36]), .Z(n478) );
  IV U96 ( .A(B[37]), .Z(n477) );
  IV U97 ( .A(B[38]), .Z(n476) );
  IV U98 ( .A(B[39]), .Z(n475) );
  IV U99 ( .A(B[40]), .Z(n474) );
  IV U100 ( .A(B[41]), .Z(n473) );
  IV U101 ( .A(B[42]), .Z(n472) );
  IV U102 ( .A(B[43]), .Z(n471) );
  IV U103 ( .A(B[44]), .Z(n470) );
  IV U104 ( .A(B[467]), .Z(n47) );
  IV U105 ( .A(B[45]), .Z(n469) );
  IV U106 ( .A(B[46]), .Z(n468) );
  IV U107 ( .A(B[47]), .Z(n467) );
  IV U108 ( .A(B[48]), .Z(n466) );
  IV U109 ( .A(B[49]), .Z(n465) );
  IV U110 ( .A(B[50]), .Z(n464) );
  IV U111 ( .A(B[51]), .Z(n463) );
  IV U112 ( .A(B[52]), .Z(n462) );
  IV U113 ( .A(B[53]), .Z(n461) );
  IV U114 ( .A(B[54]), .Z(n460) );
  IV U115 ( .A(B[468]), .Z(n46) );
  IV U116 ( .A(B[55]), .Z(n459) );
  IV U117 ( .A(B[56]), .Z(n458) );
  IV U118 ( .A(B[57]), .Z(n457) );
  IV U119 ( .A(B[58]), .Z(n456) );
  IV U120 ( .A(B[59]), .Z(n455) );
  IV U121 ( .A(B[60]), .Z(n454) );
  IV U122 ( .A(B[61]), .Z(n453) );
  IV U123 ( .A(B[62]), .Z(n452) );
  IV U124 ( .A(B[63]), .Z(n451) );
  IV U125 ( .A(B[64]), .Z(n450) );
  IV U126 ( .A(B[469]), .Z(n45) );
  IV U127 ( .A(B[65]), .Z(n449) );
  IV U128 ( .A(B[66]), .Z(n448) );
  IV U129 ( .A(B[67]), .Z(n447) );
  IV U130 ( .A(B[68]), .Z(n446) );
  IV U131 ( .A(B[69]), .Z(n445) );
  IV U132 ( .A(B[70]), .Z(n444) );
  IV U133 ( .A(B[71]), .Z(n443) );
  IV U134 ( .A(B[72]), .Z(n442) );
  IV U135 ( .A(B[73]), .Z(n441) );
  IV U136 ( .A(B[74]), .Z(n440) );
  IV U137 ( .A(B[470]), .Z(n44) );
  IV U138 ( .A(B[75]), .Z(n439) );
  IV U139 ( .A(B[76]), .Z(n438) );
  IV U140 ( .A(B[77]), .Z(n437) );
  IV U141 ( .A(B[78]), .Z(n436) );
  IV U142 ( .A(B[79]), .Z(n435) );
  IV U143 ( .A(B[80]), .Z(n434) );
  IV U144 ( .A(B[81]), .Z(n433) );
  IV U145 ( .A(B[82]), .Z(n432) );
  IV U146 ( .A(B[83]), .Z(n431) );
  IV U147 ( .A(B[84]), .Z(n430) );
  IV U148 ( .A(B[471]), .Z(n43) );
  IV U149 ( .A(B[85]), .Z(n429) );
  IV U150 ( .A(B[86]), .Z(n428) );
  IV U151 ( .A(B[87]), .Z(n427) );
  IV U152 ( .A(B[88]), .Z(n426) );
  IV U153 ( .A(B[89]), .Z(n425) );
  IV U154 ( .A(B[90]), .Z(n424) );
  IV U155 ( .A(B[91]), .Z(n423) );
  IV U156 ( .A(B[92]), .Z(n422) );
  IV U157 ( .A(B[93]), .Z(n421) );
  IV U158 ( .A(B[94]), .Z(n420) );
  IV U159 ( .A(B[472]), .Z(n42) );
  IV U160 ( .A(B[95]), .Z(n419) );
  IV U161 ( .A(B[96]), .Z(n418) );
  IV U162 ( .A(B[97]), .Z(n417) );
  IV U163 ( .A(B[98]), .Z(n416) );
  IV U164 ( .A(B[99]), .Z(n415) );
  IV U165 ( .A(B[100]), .Z(n414) );
  IV U166 ( .A(B[101]), .Z(n413) );
  IV U167 ( .A(B[102]), .Z(n412) );
  IV U168 ( .A(B[103]), .Z(n411) );
  IV U169 ( .A(B[104]), .Z(n410) );
  IV U170 ( .A(B[473]), .Z(n41) );
  IV U171 ( .A(B[105]), .Z(n409) );
  IV U172 ( .A(B[106]), .Z(n408) );
  IV U173 ( .A(B[107]), .Z(n407) );
  IV U174 ( .A(B[108]), .Z(n406) );
  IV U175 ( .A(B[109]), .Z(n405) );
  IV U176 ( .A(B[110]), .Z(n404) );
  IV U177 ( .A(B[111]), .Z(n403) );
  IV U178 ( .A(B[112]), .Z(n402) );
  IV U179 ( .A(B[113]), .Z(n401) );
  IV U180 ( .A(B[114]), .Z(n400) );
  IV U181 ( .A(B[474]), .Z(n40) );
  IV U182 ( .A(B[510]), .Z(n4) );
  IV U183 ( .A(B[115]), .Z(n399) );
  IV U184 ( .A(B[116]), .Z(n398) );
  IV U185 ( .A(B[117]), .Z(n397) );
  IV U186 ( .A(B[118]), .Z(n396) );
  IV U187 ( .A(B[119]), .Z(n395) );
  IV U188 ( .A(B[120]), .Z(n394) );
  IV U189 ( .A(B[121]), .Z(n393) );
  IV U190 ( .A(B[122]), .Z(n392) );
  IV U191 ( .A(B[123]), .Z(n391) );
  IV U192 ( .A(B[124]), .Z(n390) );
  IV U193 ( .A(B[475]), .Z(n39) );
  IV U194 ( .A(B[125]), .Z(n389) );
  IV U195 ( .A(B[126]), .Z(n388) );
  IV U196 ( .A(B[127]), .Z(n387) );
  IV U197 ( .A(B[128]), .Z(n386) );
  IV U198 ( .A(B[129]), .Z(n385) );
  IV U199 ( .A(B[130]), .Z(n384) );
  IV U200 ( .A(B[131]), .Z(n383) );
  IV U201 ( .A(B[132]), .Z(n382) );
  IV U202 ( .A(B[133]), .Z(n381) );
  IV U203 ( .A(B[134]), .Z(n380) );
  IV U204 ( .A(B[476]), .Z(n38) );
  IV U205 ( .A(B[135]), .Z(n379) );
  IV U206 ( .A(B[136]), .Z(n378) );
  IV U207 ( .A(B[137]), .Z(n377) );
  IV U208 ( .A(B[138]), .Z(n376) );
  IV U209 ( .A(B[139]), .Z(n375) );
  IV U210 ( .A(B[140]), .Z(n374) );
  IV U211 ( .A(B[141]), .Z(n373) );
  IV U212 ( .A(B[142]), .Z(n372) );
  IV U213 ( .A(B[143]), .Z(n371) );
  IV U214 ( .A(B[144]), .Z(n370) );
  IV U215 ( .A(B[477]), .Z(n37) );
  IV U216 ( .A(B[145]), .Z(n369) );
  IV U217 ( .A(B[146]), .Z(n368) );
  IV U218 ( .A(B[147]), .Z(n367) );
  IV U219 ( .A(B[148]), .Z(n366) );
  IV U220 ( .A(B[149]), .Z(n365) );
  IV U221 ( .A(B[150]), .Z(n364) );
  IV U222 ( .A(B[151]), .Z(n363) );
  IV U223 ( .A(B[152]), .Z(n362) );
  IV U224 ( .A(B[153]), .Z(n361) );
  IV U225 ( .A(B[154]), .Z(n360) );
  IV U226 ( .A(B[478]), .Z(n36) );
  IV U227 ( .A(B[155]), .Z(n359) );
  IV U228 ( .A(B[156]), .Z(n358) );
  IV U229 ( .A(B[157]), .Z(n357) );
  IV U230 ( .A(B[158]), .Z(n356) );
  IV U231 ( .A(B[159]), .Z(n355) );
  IV U232 ( .A(B[160]), .Z(n354) );
  IV U233 ( .A(B[161]), .Z(n353) );
  IV U234 ( .A(B[162]), .Z(n352) );
  IV U235 ( .A(B[163]), .Z(n351) );
  IV U236 ( .A(B[164]), .Z(n350) );
  IV U237 ( .A(B[479]), .Z(n35) );
  IV U238 ( .A(B[165]), .Z(n349) );
  IV U239 ( .A(B[166]), .Z(n348) );
  IV U240 ( .A(B[167]), .Z(n347) );
  IV U241 ( .A(B[168]), .Z(n346) );
  IV U242 ( .A(B[169]), .Z(n345) );
  IV U243 ( .A(B[170]), .Z(n344) );
  IV U244 ( .A(B[171]), .Z(n343) );
  IV U245 ( .A(B[172]), .Z(n342) );
  IV U246 ( .A(B[173]), .Z(n341) );
  IV U247 ( .A(B[174]), .Z(n340) );
  IV U248 ( .A(B[480]), .Z(n34) );
  IV U249 ( .A(B[175]), .Z(n339) );
  IV U250 ( .A(B[176]), .Z(n338) );
  IV U251 ( .A(B[177]), .Z(n337) );
  IV U252 ( .A(B[178]), .Z(n336) );
  IV U253 ( .A(B[179]), .Z(n335) );
  IV U254 ( .A(B[180]), .Z(n334) );
  IV U255 ( .A(B[181]), .Z(n333) );
  IV U256 ( .A(B[182]), .Z(n332) );
  IV U257 ( .A(B[183]), .Z(n331) );
  IV U258 ( .A(B[184]), .Z(n330) );
  IV U259 ( .A(B[481]), .Z(n33) );
  IV U260 ( .A(B[185]), .Z(n329) );
  IV U261 ( .A(B[186]), .Z(n328) );
  IV U262 ( .A(B[187]), .Z(n327) );
  IV U263 ( .A(B[188]), .Z(n326) );
  IV U264 ( .A(B[189]), .Z(n325) );
  IV U265 ( .A(B[190]), .Z(n324) );
  IV U266 ( .A(B[191]), .Z(n323) );
  IV U267 ( .A(B[192]), .Z(n322) );
  IV U268 ( .A(B[193]), .Z(n321) );
  IV U269 ( .A(B[194]), .Z(n320) );
  IV U270 ( .A(B[482]), .Z(n32) );
  IV U271 ( .A(B[195]), .Z(n319) );
  IV U272 ( .A(B[196]), .Z(n318) );
  IV U273 ( .A(B[197]), .Z(n317) );
  IV U274 ( .A(B[198]), .Z(n316) );
  IV U275 ( .A(B[199]), .Z(n315) );
  IV U276 ( .A(B[200]), .Z(n314) );
  IV U277 ( .A(B[201]), .Z(n313) );
  IV U278 ( .A(B[202]), .Z(n312) );
  IV U279 ( .A(B[203]), .Z(n311) );
  IV U280 ( .A(B[204]), .Z(n310) );
  IV U281 ( .A(B[483]), .Z(n31) );
  IV U282 ( .A(B[205]), .Z(n309) );
  IV U283 ( .A(B[206]), .Z(n308) );
  IV U284 ( .A(B[207]), .Z(n307) );
  IV U285 ( .A(B[208]), .Z(n306) );
  IV U286 ( .A(B[209]), .Z(n305) );
  IV U287 ( .A(B[210]), .Z(n304) );
  IV U288 ( .A(B[211]), .Z(n303) );
  IV U289 ( .A(B[212]), .Z(n302) );
  IV U290 ( .A(B[213]), .Z(n301) );
  IV U291 ( .A(B[214]), .Z(n300) );
  IV U292 ( .A(B[484]), .Z(n30) );
  IV U293 ( .A(B[511]), .Z(n3) );
  IV U294 ( .A(B[215]), .Z(n299) );
  IV U295 ( .A(B[216]), .Z(n298) );
  IV U296 ( .A(B[217]), .Z(n297) );
  IV U297 ( .A(B[218]), .Z(n296) );
  IV U298 ( .A(B[219]), .Z(n295) );
  IV U299 ( .A(B[220]), .Z(n294) );
  IV U300 ( .A(B[221]), .Z(n293) );
  IV U301 ( .A(B[222]), .Z(n292) );
  IV U302 ( .A(B[223]), .Z(n291) );
  IV U303 ( .A(B[224]), .Z(n290) );
  IV U304 ( .A(B[485]), .Z(n29) );
  IV U305 ( .A(B[225]), .Z(n289) );
  IV U306 ( .A(B[226]), .Z(n288) );
  IV U307 ( .A(B[227]), .Z(n287) );
  IV U308 ( .A(B[228]), .Z(n286) );
  IV U309 ( .A(B[229]), .Z(n285) );
  IV U310 ( .A(B[230]), .Z(n284) );
  IV U311 ( .A(B[231]), .Z(n283) );
  IV U312 ( .A(B[232]), .Z(n282) );
  IV U313 ( .A(B[233]), .Z(n281) );
  IV U314 ( .A(B[234]), .Z(n280) );
  IV U315 ( .A(B[486]), .Z(n28) );
  IV U316 ( .A(B[235]), .Z(n279) );
  IV U317 ( .A(B[236]), .Z(n278) );
  IV U318 ( .A(B[237]), .Z(n277) );
  IV U319 ( .A(B[238]), .Z(n276) );
  IV U320 ( .A(B[239]), .Z(n275) );
  IV U321 ( .A(B[240]), .Z(n274) );
  IV U322 ( .A(B[241]), .Z(n273) );
  IV U323 ( .A(B[242]), .Z(n272) );
  IV U324 ( .A(B[243]), .Z(n271) );
  IV U325 ( .A(B[244]), .Z(n270) );
  IV U326 ( .A(B[487]), .Z(n27) );
  IV U327 ( .A(B[245]), .Z(n269) );
  IV U328 ( .A(B[246]), .Z(n268) );
  IV U329 ( .A(B[247]), .Z(n267) );
  IV U330 ( .A(B[248]), .Z(n266) );
  IV U331 ( .A(B[249]), .Z(n265) );
  IV U332 ( .A(B[250]), .Z(n264) );
  IV U333 ( .A(B[251]), .Z(n263) );
  IV U334 ( .A(B[252]), .Z(n262) );
  IV U335 ( .A(B[253]), .Z(n261) );
  IV U336 ( .A(B[254]), .Z(n260) );
  IV U337 ( .A(B[488]), .Z(n26) );
  IV U338 ( .A(B[255]), .Z(n259) );
  IV U339 ( .A(B[256]), .Z(n258) );
  IV U340 ( .A(B[257]), .Z(n257) );
  IV U341 ( .A(B[258]), .Z(n256) );
  IV U342 ( .A(B[259]), .Z(n255) );
  IV U343 ( .A(B[260]), .Z(n254) );
  IV U344 ( .A(B[261]), .Z(n253) );
  IV U345 ( .A(B[262]), .Z(n252) );
  IV U346 ( .A(B[263]), .Z(n251) );
  IV U347 ( .A(B[264]), .Z(n250) );
  IV U348 ( .A(B[489]), .Z(n25) );
  IV U349 ( .A(B[265]), .Z(n249) );
  IV U350 ( .A(B[266]), .Z(n248) );
  IV U351 ( .A(B[267]), .Z(n247) );
  IV U352 ( .A(B[268]), .Z(n246) );
  IV U353 ( .A(B[269]), .Z(n245) );
  IV U354 ( .A(B[270]), .Z(n244) );
  IV U355 ( .A(B[271]), .Z(n243) );
  IV U356 ( .A(B[272]), .Z(n242) );
  IV U357 ( .A(B[273]), .Z(n241) );
  IV U358 ( .A(B[274]), .Z(n240) );
  IV U359 ( .A(B[490]), .Z(n24) );
  IV U360 ( .A(B[275]), .Z(n239) );
  IV U361 ( .A(B[276]), .Z(n238) );
  IV U362 ( .A(B[277]), .Z(n237) );
  IV U363 ( .A(B[278]), .Z(n236) );
  IV U364 ( .A(B[279]), .Z(n235) );
  IV U365 ( .A(B[280]), .Z(n234) );
  IV U366 ( .A(B[281]), .Z(n233) );
  IV U367 ( .A(B[282]), .Z(n232) );
  IV U368 ( .A(B[283]), .Z(n231) );
  IV U369 ( .A(B[284]), .Z(n230) );
  IV U370 ( .A(B[491]), .Z(n23) );
  IV U371 ( .A(B[285]), .Z(n229) );
  IV U372 ( .A(B[286]), .Z(n228) );
  IV U373 ( .A(B[287]), .Z(n227) );
  IV U374 ( .A(B[288]), .Z(n226) );
  IV U375 ( .A(B[289]), .Z(n225) );
  IV U376 ( .A(B[290]), .Z(n224) );
  IV U377 ( .A(B[291]), .Z(n223) );
  IV U378 ( .A(B[292]), .Z(n222) );
  IV U379 ( .A(B[293]), .Z(n221) );
  IV U380 ( .A(B[294]), .Z(n220) );
  IV U381 ( .A(B[492]), .Z(n22) );
  IV U382 ( .A(B[295]), .Z(n219) );
  IV U383 ( .A(B[296]), .Z(n218) );
  IV U384 ( .A(B[297]), .Z(n217) );
  IV U385 ( .A(B[298]), .Z(n216) );
  IV U386 ( .A(B[299]), .Z(n215) );
  IV U387 ( .A(B[300]), .Z(n214) );
  IV U388 ( .A(B[301]), .Z(n213) );
  IV U389 ( .A(B[302]), .Z(n212) );
  IV U390 ( .A(B[303]), .Z(n211) );
  IV U391 ( .A(B[304]), .Z(n210) );
  IV U392 ( .A(B[493]), .Z(n21) );
  IV U393 ( .A(B[305]), .Z(n209) );
  IV U394 ( .A(B[306]), .Z(n208) );
  IV U395 ( .A(B[307]), .Z(n207) );
  IV U396 ( .A(B[308]), .Z(n206) );
  IV U397 ( .A(B[309]), .Z(n205) );
  IV U398 ( .A(B[310]), .Z(n204) );
  IV U399 ( .A(B[311]), .Z(n203) );
  IV U400 ( .A(B[312]), .Z(n202) );
  IV U401 ( .A(B[313]), .Z(n201) );
  IV U402 ( .A(B[314]), .Z(n200) );
  IV U403 ( .A(B[494]), .Z(n20) );
  IV U404 ( .A(B[315]), .Z(n199) );
  IV U405 ( .A(B[316]), .Z(n198) );
  IV U406 ( .A(B[317]), .Z(n197) );
  IV U407 ( .A(B[318]), .Z(n196) );
  IV U408 ( .A(B[319]), .Z(n195) );
  IV U409 ( .A(B[320]), .Z(n194) );
  IV U410 ( .A(B[321]), .Z(n193) );
  IV U411 ( .A(B[322]), .Z(n192) );
  IV U412 ( .A(B[323]), .Z(n191) );
  IV U413 ( .A(B[324]), .Z(n190) );
  IV U414 ( .A(B[495]), .Z(n19) );
  IV U415 ( .A(B[325]), .Z(n189) );
  IV U416 ( .A(B[326]), .Z(n188) );
  IV U417 ( .A(B[327]), .Z(n187) );
  IV U418 ( .A(B[328]), .Z(n186) );
  IV U419 ( .A(B[329]), .Z(n185) );
  IV U420 ( .A(B[330]), .Z(n184) );
  IV U421 ( .A(B[331]), .Z(n183) );
  IV U422 ( .A(B[332]), .Z(n182) );
  IV U423 ( .A(B[333]), .Z(n181) );
  IV U424 ( .A(B[334]), .Z(n180) );
  IV U425 ( .A(B[496]), .Z(n18) );
  IV U426 ( .A(B[335]), .Z(n179) );
  IV U427 ( .A(B[336]), .Z(n178) );
  IV U428 ( .A(B[337]), .Z(n177) );
  IV U429 ( .A(B[338]), .Z(n176) );
  IV U430 ( .A(B[339]), .Z(n175) );
  IV U431 ( .A(B[340]), .Z(n174) );
  IV U432 ( .A(B[341]), .Z(n173) );
  IV U433 ( .A(B[342]), .Z(n172) );
  IV U434 ( .A(B[343]), .Z(n171) );
  IV U435 ( .A(B[344]), .Z(n170) );
  IV U436 ( .A(B[497]), .Z(n17) );
  IV U437 ( .A(B[345]), .Z(n169) );
  IV U438 ( .A(B[346]), .Z(n168) );
  IV U439 ( .A(B[347]), .Z(n167) );
  IV U440 ( .A(B[348]), .Z(n166) );
  IV U441 ( .A(B[349]), .Z(n165) );
  IV U442 ( .A(B[350]), .Z(n164) );
  IV U443 ( .A(B[351]), .Z(n163) );
  IV U444 ( .A(B[352]), .Z(n162) );
  IV U445 ( .A(B[353]), .Z(n161) );
  IV U446 ( .A(B[354]), .Z(n160) );
  IV U447 ( .A(B[498]), .Z(n16) );
  IV U448 ( .A(B[355]), .Z(n159) );
  IV U449 ( .A(B[356]), .Z(n158) );
  IV U450 ( .A(B[357]), .Z(n157) );
  IV U451 ( .A(B[358]), .Z(n156) );
  IV U452 ( .A(B[359]), .Z(n155) );
  IV U453 ( .A(B[360]), .Z(n154) );
  IV U454 ( .A(B[361]), .Z(n153) );
  IV U455 ( .A(B[362]), .Z(n152) );
  IV U456 ( .A(B[363]), .Z(n151) );
  IV U457 ( .A(B[364]), .Z(n150) );
  IV U458 ( .A(B[499]), .Z(n15) );
  IV U459 ( .A(B[365]), .Z(n149) );
  IV U460 ( .A(B[366]), .Z(n148) );
  IV U461 ( .A(B[367]), .Z(n147) );
  IV U462 ( .A(B[368]), .Z(n146) );
  IV U463 ( .A(B[369]), .Z(n145) );
  IV U464 ( .A(B[370]), .Z(n144) );
  IV U465 ( .A(B[371]), .Z(n143) );
  IV U466 ( .A(B[372]), .Z(n142) );
  IV U467 ( .A(B[373]), .Z(n141) );
  IV U468 ( .A(B[374]), .Z(n140) );
  IV U469 ( .A(B[500]), .Z(n14) );
  IV U470 ( .A(B[375]), .Z(n139) );
  IV U471 ( .A(B[376]), .Z(n138) );
  IV U472 ( .A(B[377]), .Z(n137) );
  IV U473 ( .A(B[378]), .Z(n136) );
  IV U474 ( .A(B[379]), .Z(n135) );
  IV U475 ( .A(B[380]), .Z(n134) );
  IV U476 ( .A(B[381]), .Z(n133) );
  IV U477 ( .A(B[382]), .Z(n132) );
  IV U478 ( .A(B[383]), .Z(n131) );
  IV U479 ( .A(B[384]), .Z(n130) );
  IV U480 ( .A(B[501]), .Z(n13) );
  IV U481 ( .A(B[385]), .Z(n129) );
  IV U482 ( .A(B[386]), .Z(n128) );
  IV U483 ( .A(B[387]), .Z(n127) );
  IV U484 ( .A(B[388]), .Z(n126) );
  IV U485 ( .A(B[389]), .Z(n125) );
  IV U486 ( .A(B[390]), .Z(n124) );
  IV U487 ( .A(B[391]), .Z(n123) );
  IV U488 ( .A(B[392]), .Z(n122) );
  IV U489 ( .A(B[393]), .Z(n121) );
  IV U490 ( .A(B[394]), .Z(n120) );
  IV U491 ( .A(B[502]), .Z(n12) );
  IV U492 ( .A(B[395]), .Z(n119) );
  IV U493 ( .A(B[396]), .Z(n118) );
  IV U494 ( .A(B[397]), .Z(n117) );
  IV U495 ( .A(B[398]), .Z(n116) );
  IV U496 ( .A(B[399]), .Z(n115) );
  IV U497 ( .A(B[400]), .Z(n114) );
  IV U498 ( .A(B[401]), .Z(n113) );
  IV U499 ( .A(B[402]), .Z(n112) );
  IV U500 ( .A(B[403]), .Z(n111) );
  IV U501 ( .A(B[404]), .Z(n110) );
  IV U502 ( .A(B[503]), .Z(n11) );
  IV U503 ( .A(B[405]), .Z(n109) );
  IV U504 ( .A(B[406]), .Z(n108) );
  IV U505 ( .A(B[407]), .Z(n107) );
  IV U506 ( .A(B[408]), .Z(n106) );
  IV U507 ( .A(B[409]), .Z(n105) );
  IV U508 ( .A(B[410]), .Z(n104) );
  IV U509 ( .A(B[411]), .Z(n103) );
  IV U510 ( .A(B[412]), .Z(n102) );
  IV U511 ( .A(B[413]), .Z(n101) );
  IV U512 ( .A(B[414]), .Z(n100) );
  IV U513 ( .A(B[504]), .Z(n10) );
endmodule


module FA_10035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_10036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  NANDN U1 ( .A(CI), .B(S), .Z(CO) );
  XNOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_10037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_10548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N514_2 ( A, B, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  output CO;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514;
  wire   [513:1] C;

  FA_10548 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n514), .CI(1'b1), 
        .S(S[0]), .CO(C[1]) );
  FA_10547 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n513), .CI(C[1]), 
        .S(S[1]), .CO(C[2]) );
  FA_10546 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n512), .CI(C[2]), 
        .S(S[2]), .CO(C[3]) );
  FA_10545 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n511), .CI(C[3]), 
        .S(S[3]), .CO(C[4]) );
  FA_10544 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n510), .CI(C[4]), 
        .S(S[4]), .CO(C[5]) );
  FA_10543 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n509), .CI(C[5]), 
        .S(S[5]), .CO(C[6]) );
  FA_10542 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n508), .CI(C[6]), 
        .S(S[6]), .CO(C[7]) );
  FA_10541 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n507), .CI(C[7]), 
        .S(S[7]), .CO(C[8]) );
  FA_10540 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n506), .CI(C[8]), 
        .S(S[8]), .CO(C[9]) );
  FA_10539 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n505), .CI(C[9]), 
        .S(S[9]), .CO(C[10]) );
  FA_10538 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n504), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_10537 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n503), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_10536 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n502), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_10535 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n501), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_10534 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n500), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_10533 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n499), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_10532 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n498), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_10531 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n497), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_10530 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n496), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_10529 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n495), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_10528 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n494), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_10527 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n493), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_10526 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n492), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_10525 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n491), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_10524 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n490), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_10523 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n489), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_10522 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n488), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_10521 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n487), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_10520 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n486), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_10519 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n485), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_10518 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n484), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_10517 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n483), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_10516 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n482), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_10515 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n481), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_10514 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n480), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_10513 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n479), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_10512 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n478), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_10511 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n477), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_10510 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n476), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_10509 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n475), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_10508 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n474), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_10507 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n473), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_10506 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n472), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_10505 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n471), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_10504 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n470), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_10503 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n469), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_10502 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n468), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_10501 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n467), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_10500 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n466), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_10499 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n465), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_10498 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n464), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_10497 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n463), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_10496 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n462), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_10495 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n461), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_10494 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n460), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_10493 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n459), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_10492 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n458), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_10491 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n457), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_10490 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n456), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_10489 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n455), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_10488 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n454), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_10487 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n453), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_10486 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n452), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_10485 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n451), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_10484 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n450), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_10483 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n449), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_10482 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n448), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_10481 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n447), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_10480 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n446), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_10479 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n445), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_10478 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n444), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_10477 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n443), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_10476 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n442), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_10475 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n441), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_10474 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n440), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_10473 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n439), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_10472 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n438), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_10471 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n437), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_10470 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n436), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_10469 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n435), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_10468 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n434), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_10467 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n433), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_10466 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n432), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_10465 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n431), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_10464 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n430), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_10463 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n429), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_10462 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n428), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_10461 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n427), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_10460 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n426), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_10459 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n425), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_10458 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n424), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_10457 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n423), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_10456 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n422), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_10455 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n421), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_10454 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n420), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_10453 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n419), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_10452 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n418), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_10451 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n417), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_10450 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n416), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_10449 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n415), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_10448 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n414), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_10447 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n413), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_10446 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n412), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_10445 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n411), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_10444 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n410), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_10443 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n409), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_10442 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n408), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_10441 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n407), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_10440 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n406), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_10439 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n405), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_10438 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n404), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_10437 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n403), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_10436 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n402), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_10435 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n401), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_10434 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n400), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_10433 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n399), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_10432 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n398), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_10431 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n397), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_10430 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n396), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_10429 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n395), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_10428 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n394), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_10427 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n393), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_10426 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n392), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_10425 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n391), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_10424 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n390), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_10423 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n389), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_10422 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n388), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_10421 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n387), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_10420 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n386), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_10419 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n385), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_10418 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n384), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_10417 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n383), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_10416 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n382), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_10415 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n381), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_10414 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n380), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_10413 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n379), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_10412 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n378), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_10411 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n377), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_10410 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n376), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_10409 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n375), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_10408 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n374), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_10407 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n373), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_10406 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n372), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_10405 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n371), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_10404 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n370), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_10403 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n369), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_10402 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n368), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_10401 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n367), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_10400 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n366), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_10399 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n365), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_10398 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n364), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_10397 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n363), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_10396 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n362), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_10395 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n361), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_10394 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n360), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_10393 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n359), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_10392 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n358), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_10391 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n357), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_10390 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n356), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_10389 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n355), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_10388 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n354), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_10387 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n353), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_10386 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n352), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_10385 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n351), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_10384 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n350), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_10383 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n349), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_10382 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n348), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_10381 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n347), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_10380 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n346), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_10379 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n345), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_10378 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n344), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_10377 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n343), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_10376 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n342), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_10375 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n341), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_10374 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n340), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_10373 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n339), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_10372 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n338), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_10371 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n337), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_10370 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n336), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_10369 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n335), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_10368 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n334), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_10367 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n333), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_10366 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n332), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_10365 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n331), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_10364 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n330), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_10363 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n329), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_10362 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n328), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_10361 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n327), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_10360 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n326), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_10359 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n325), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_10358 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n324), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_10357 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n323), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_10356 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n322), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_10355 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n321), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_10354 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n320), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_10353 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n319), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_10352 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n318), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_10351 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n317), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_10350 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n316), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_10349 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n315), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_10348 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n314), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_10347 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n313), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_10346 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n312), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_10345 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n311), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_10344 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n310), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_10343 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n309), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_10342 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n308), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_10341 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n307), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_10340 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n306), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_10339 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n305), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_10338 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n304), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_10337 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n303), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_10336 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n302), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_10335 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n301), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_10334 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n300), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_10333 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n299), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_10332 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n298), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_10331 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n297), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_10330 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n296), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_10329 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n295), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_10328 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n294), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_10327 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n293), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_10326 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n292), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_10325 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n291), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_10324 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n290), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_10323 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n289), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_10322 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n288), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_10321 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n287), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_10320 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n286), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_10319 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n285), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_10318 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n284), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_10317 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n283), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_10316 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n282), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_10315 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n281), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_10314 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n280), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_10313 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n279), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_10312 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n278), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_10311 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n277), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_10310 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n276), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_10309 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n275), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_10308 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n274), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_10307 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n273), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_10306 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n272), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_10305 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n271), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_10304 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n270), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_10303 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n269), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_10302 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n268), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_10301 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n267), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_10300 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n266), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_10299 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n265), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_10298 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n264), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_10297 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n263), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_10296 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n262), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_10295 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n261), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_10294 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n260), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_10293 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n259), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_10292 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n258), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_10291 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n257), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_10290 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n256), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_10289 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n255), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_10288 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n254), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_10287 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n253), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_10286 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n252), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_10285 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n251), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_10284 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n250), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_10283 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n249), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_10282 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n248), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_10281 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n247), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_10280 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n246), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_10279 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n245), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_10278 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n244), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_10277 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n243), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_10276 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n242), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_10275 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n241), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_10274 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n240), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_10273 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n239), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_10272 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n238), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_10271 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n237), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_10270 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n236), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_10269 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n235), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_10268 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n234), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_10267 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n233), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_10266 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n232), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_10265 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n231), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_10264 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n230), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_10263 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n229), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_10262 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n228), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_10261 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n227), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_10260 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n226), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_10259 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n225), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_10258 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n224), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_10257 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n223), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_10256 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n222), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_10255 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n221), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_10254 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n220), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_10253 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n219), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_10252 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n218), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_10251 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n217), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_10250 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n216), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_10249 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n215), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_10248 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n214), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_10247 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n213), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_10246 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n212), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_10245 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n211), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_10244 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n210), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_10243 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n209), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_10242 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n208), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_10241 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n207), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_10240 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n206), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_10239 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n205), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_10238 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n204), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_10237 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n203), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_10236 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n202), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_10235 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n201), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_10234 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n200), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_10233 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n199), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_10232 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n198), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_10231 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n197), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_10230 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n196), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_10229 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n195), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_10228 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n194), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_10227 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n193), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_10226 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n192), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_10225 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n191), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_10224 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n190), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_10223 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n189), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_10222 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n188), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_10221 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n187), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_10220 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n186), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_10219 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n185), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_10218 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n184), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_10217 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n183), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_10216 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n182), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_10215 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n181), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_10214 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n180), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_10213 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n179), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_10212 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n178), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_10211 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n177), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_10210 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n176), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_10209 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n175), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_10208 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n174), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_10207 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n173), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_10206 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n172), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_10205 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n171), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_10204 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n170), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_10203 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n169), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_10202 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n168), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_10201 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n167), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_10200 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n166), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_10199 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n165), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_10198 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n164), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_10197 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n163), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_10196 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n162), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_10195 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n161), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_10194 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n160), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_10193 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n159), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_10192 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n158), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_10191 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n157), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_10190 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n156), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_10189 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n155), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_10188 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n154), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_10187 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n153), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_10186 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n152), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_10185 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n151), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_10184 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n150), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_10183 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n149), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_10182 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n148), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_10181 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n147), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_10180 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n146), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_10179 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n145), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_10178 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n144), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_10177 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n143), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_10176 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n142), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_10175 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n141), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_10174 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n140), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_10173 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n139), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_10172 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n138), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_10171 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n137), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_10170 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n136), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_10169 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n135), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_10168 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n134), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_10167 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n133), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_10166 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n132), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_10165 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n131), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_10164 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n130), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_10163 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n129), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_10162 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n128), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_10161 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n127), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_10160 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n126), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_10159 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n125), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_10158 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n124), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_10157 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n123), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_10156 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n122), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_10155 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n121), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_10154 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n120), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_10153 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n119), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_10152 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n118), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_10151 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n117), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_10150 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n116), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_10149 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n115), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_10148 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n114), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_10147 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n113), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_10146 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n112), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_10145 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n111), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_10144 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n110), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_10143 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n109), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_10142 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n108), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_10141 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n107), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_10140 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n106), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_10139 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n105), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_10138 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n104), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_10137 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n103), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_10136 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n102), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_10135 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n101), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_10134 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n100), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_10133 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n99), .CI(C[415]), .S(S[415]), .CO(C[416]) );
  FA_10132 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n98), .CI(C[416]), .S(S[416]), .CO(C[417]) );
  FA_10131 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n97), .CI(C[417]), .S(S[417]), .CO(C[418]) );
  FA_10130 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n96), .CI(C[418]), .S(S[418]), .CO(C[419]) );
  FA_10129 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n95), .CI(C[419]), .S(S[419]), .CO(C[420]) );
  FA_10128 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n94), .CI(C[420]), .S(S[420]), .CO(C[421]) );
  FA_10127 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n93), .CI(C[421]), .S(S[421]), .CO(C[422]) );
  FA_10126 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n92), .CI(C[422]), .S(S[422]), .CO(C[423]) );
  FA_10125 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n91), .CI(C[423]), .S(S[423]), .CO(C[424]) );
  FA_10124 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n90), .CI(C[424]), .S(S[424]), .CO(C[425]) );
  FA_10123 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n89), .CI(C[425]), .S(S[425]), .CO(C[426]) );
  FA_10122 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n88), .CI(C[426]), .S(S[426]), .CO(C[427]) );
  FA_10121 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n87), .CI(C[427]), .S(S[427]), .CO(C[428]) );
  FA_10120 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n86), .CI(C[428]), .S(S[428]), .CO(C[429]) );
  FA_10119 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n85), .CI(C[429]), .S(S[429]), .CO(C[430]) );
  FA_10118 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n84), .CI(C[430]), .S(S[430]), .CO(C[431]) );
  FA_10117 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n83), .CI(C[431]), .S(S[431]), .CO(C[432]) );
  FA_10116 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n82), .CI(C[432]), .S(S[432]), .CO(C[433]) );
  FA_10115 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n81), .CI(C[433]), .S(S[433]), .CO(C[434]) );
  FA_10114 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n80), .CI(C[434]), .S(S[434]), .CO(C[435]) );
  FA_10113 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n79), .CI(C[435]), .S(S[435]), .CO(C[436]) );
  FA_10112 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n78), .CI(C[436]), .S(S[436]), .CO(C[437]) );
  FA_10111 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n77), .CI(C[437]), .S(S[437]), .CO(C[438]) );
  FA_10110 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n76), .CI(C[438]), .S(S[438]), .CO(C[439]) );
  FA_10109 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n75), .CI(C[439]), .S(S[439]), .CO(C[440]) );
  FA_10108 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n74), .CI(C[440]), .S(S[440]), .CO(C[441]) );
  FA_10107 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n73), .CI(C[441]), .S(S[441]), .CO(C[442]) );
  FA_10106 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n72), .CI(C[442]), .S(S[442]), .CO(C[443]) );
  FA_10105 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n71), .CI(C[443]), .S(S[443]), .CO(C[444]) );
  FA_10104 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n70), .CI(C[444]), .S(S[444]), .CO(C[445]) );
  FA_10103 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n69), .CI(C[445]), .S(S[445]), .CO(C[446]) );
  FA_10102 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n68), .CI(C[446]), .S(S[446]), .CO(C[447]) );
  FA_10101 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n67), .CI(C[447]), .S(S[447]), .CO(C[448]) );
  FA_10100 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n66), .CI(C[448]), .S(S[448]), .CO(C[449]) );
  FA_10099 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n65), .CI(C[449]), .S(S[449]), .CO(C[450]) );
  FA_10098 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n64), .CI(C[450]), .S(S[450]), .CO(C[451]) );
  FA_10097 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n63), .CI(C[451]), .S(S[451]), .CO(C[452]) );
  FA_10096 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n62), .CI(C[452]), .S(S[452]), .CO(C[453]) );
  FA_10095 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n61), .CI(C[453]), .S(S[453]), .CO(C[454]) );
  FA_10094 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n60), .CI(C[454]), .S(S[454]), .CO(C[455]) );
  FA_10093 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n59), .CI(C[455]), .S(S[455]), .CO(C[456]) );
  FA_10092 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n58), .CI(C[456]), .S(S[456]), .CO(C[457]) );
  FA_10091 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n57), .CI(C[457]), .S(S[457]), .CO(C[458]) );
  FA_10090 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n56), .CI(C[458]), .S(S[458]), .CO(C[459]) );
  FA_10089 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n55), .CI(C[459]), .S(S[459]), .CO(C[460]) );
  FA_10088 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n54), .CI(C[460]), .S(S[460]), .CO(C[461]) );
  FA_10087 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n53), .CI(C[461]), .S(S[461]), .CO(C[462]) );
  FA_10086 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n52), .CI(C[462]), .S(S[462]), .CO(C[463]) );
  FA_10085 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n51), .CI(C[463]), .S(S[463]), .CO(C[464]) );
  FA_10084 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n50), .CI(C[464]), .S(S[464]), .CO(C[465]) );
  FA_10083 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n49), .CI(C[465]), .S(S[465]), .CO(C[466]) );
  FA_10082 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n48), .CI(C[466]), .S(S[466]), .CO(C[467]) );
  FA_10081 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n47), .CI(C[467]), .S(S[467]), .CO(C[468]) );
  FA_10080 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n46), .CI(C[468]), .S(S[468]), .CO(C[469]) );
  FA_10079 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n45), .CI(C[469]), .S(S[469]), .CO(C[470]) );
  FA_10078 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n44), .CI(C[470]), .S(S[470]), .CO(C[471]) );
  FA_10077 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n43), .CI(C[471]), .S(S[471]), .CO(C[472]) );
  FA_10076 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n42), .CI(C[472]), .S(S[472]), .CO(C[473]) );
  FA_10075 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n41), .CI(C[473]), .S(S[473]), .CO(C[474]) );
  FA_10074 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n40), .CI(C[474]), .S(S[474]), .CO(C[475]) );
  FA_10073 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n39), .CI(C[475]), .S(S[475]), .CO(C[476]) );
  FA_10072 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n38), .CI(C[476]), .S(S[476]), .CO(C[477]) );
  FA_10071 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n37), .CI(C[477]), .S(S[477]), .CO(C[478]) );
  FA_10070 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n36), .CI(C[478]), .S(S[478]), .CO(C[479]) );
  FA_10069 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n35), .CI(C[479]), .S(S[479]), .CO(C[480]) );
  FA_10068 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n34), .CI(C[480]), .S(S[480]), .CO(C[481]) );
  FA_10067 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n33), .CI(C[481]), .S(S[481]), .CO(C[482]) );
  FA_10066 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n32), .CI(C[482]), .S(S[482]), .CO(C[483]) );
  FA_10065 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n31), .CI(C[483]), .S(S[483]), .CO(C[484]) );
  FA_10064 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n30), .CI(C[484]), .S(S[484]), .CO(C[485]) );
  FA_10063 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n29), .CI(C[485]), .S(S[485]), .CO(C[486]) );
  FA_10062 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n28), .CI(C[486]), .S(S[486]), .CO(C[487]) );
  FA_10061 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n27), .CI(C[487]), .S(S[487]), .CO(C[488]) );
  FA_10060 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n26), .CI(C[488]), .S(S[488]), .CO(C[489]) );
  FA_10059 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n25), .CI(C[489]), .S(S[489]), .CO(C[490]) );
  FA_10058 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n24), .CI(C[490]), .S(S[490]), .CO(C[491]) );
  FA_10057 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n23), .CI(C[491]), .S(S[491]), .CO(C[492]) );
  FA_10056 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n22), .CI(C[492]), .S(S[492]), .CO(C[493]) );
  FA_10055 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n21), .CI(C[493]), .S(S[493]), .CO(C[494]) );
  FA_10054 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n20), .CI(C[494]), .S(S[494]), .CO(C[495]) );
  FA_10053 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n19), .CI(C[495]), .S(S[495]), .CO(C[496]) );
  FA_10052 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n18), .CI(C[496]), .S(S[496]), .CO(C[497]) );
  FA_10051 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n17), .CI(C[497]), .S(S[497]), .CO(C[498]) );
  FA_10050 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n16), .CI(C[498]), .S(S[498]), .CO(C[499]) );
  FA_10049 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n15), .CI(C[499]), .S(S[499]), .CO(C[500]) );
  FA_10048 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n14), .CI(C[500]), .S(S[500]), .CO(C[501]) );
  FA_10047 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n13), .CI(C[501]), .S(S[501]), .CO(C[502]) );
  FA_10046 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n12), .CI(C[502]), .S(S[502]), .CO(C[503]) );
  FA_10045 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n11), .CI(C[503]), .S(S[503]), .CO(C[504]) );
  FA_10044 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n10), .CI(C[504]), .S(S[504]), .CO(C[505]) );
  FA_10043 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n9), .CI(C[505]), 
        .S(S[505]), .CO(C[506]) );
  FA_10042 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n8), .CI(C[506]), 
        .S(S[506]), .CO(C[507]) );
  FA_10041 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n7), .CI(C[507]), 
        .S(S[507]), .CO(C[508]) );
  FA_10040 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n6), .CI(C[508]), 
        .S(S[508]), .CO(C[509]) );
  FA_10039 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n5), .CI(C[509]), 
        .S(S[509]), .CO(C[510]) );
  FA_10038 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n4), .CI(C[510]), 
        .S(S[510]), .CO(C[511]) );
  FA_10037 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n3), .CI(C[511]), 
        .S(S[511]), .CO(C[512]) );
  FA_10036 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .S(S[512]), .CO(C[513]) );
  FA_10035 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b1), .CI(C[513]), .S(S[513]) );
  IV U2 ( .A(B[415]), .Z(n99) );
  IV U3 ( .A(B[416]), .Z(n98) );
  IV U4 ( .A(B[417]), .Z(n97) );
  IV U5 ( .A(B[418]), .Z(n96) );
  IV U6 ( .A(B[419]), .Z(n95) );
  IV U7 ( .A(B[420]), .Z(n94) );
  IV U8 ( .A(B[421]), .Z(n93) );
  IV U9 ( .A(B[422]), .Z(n92) );
  IV U10 ( .A(B[423]), .Z(n91) );
  IV U11 ( .A(B[424]), .Z(n90) );
  IV U12 ( .A(B[505]), .Z(n9) );
  IV U13 ( .A(B[425]), .Z(n89) );
  IV U14 ( .A(B[426]), .Z(n88) );
  IV U15 ( .A(B[427]), .Z(n87) );
  IV U16 ( .A(B[428]), .Z(n86) );
  IV U17 ( .A(B[429]), .Z(n85) );
  IV U18 ( .A(B[430]), .Z(n84) );
  IV U19 ( .A(B[431]), .Z(n83) );
  IV U20 ( .A(B[432]), .Z(n82) );
  IV U21 ( .A(B[433]), .Z(n81) );
  IV U22 ( .A(B[434]), .Z(n80) );
  IV U23 ( .A(B[506]), .Z(n8) );
  IV U24 ( .A(B[435]), .Z(n79) );
  IV U25 ( .A(B[436]), .Z(n78) );
  IV U26 ( .A(B[437]), .Z(n77) );
  IV U27 ( .A(B[438]), .Z(n76) );
  IV U28 ( .A(B[439]), .Z(n75) );
  IV U29 ( .A(B[440]), .Z(n74) );
  IV U30 ( .A(B[441]), .Z(n73) );
  IV U31 ( .A(B[442]), .Z(n72) );
  IV U32 ( .A(B[443]), .Z(n71) );
  IV U33 ( .A(B[444]), .Z(n70) );
  IV U34 ( .A(B[507]), .Z(n7) );
  IV U35 ( .A(B[445]), .Z(n69) );
  IV U36 ( .A(B[446]), .Z(n68) );
  IV U37 ( .A(B[447]), .Z(n67) );
  IV U38 ( .A(B[448]), .Z(n66) );
  IV U39 ( .A(B[449]), .Z(n65) );
  IV U40 ( .A(B[450]), .Z(n64) );
  IV U41 ( .A(B[451]), .Z(n63) );
  IV U42 ( .A(B[452]), .Z(n62) );
  IV U43 ( .A(B[453]), .Z(n61) );
  IV U44 ( .A(B[454]), .Z(n60) );
  IV U45 ( .A(B[508]), .Z(n6) );
  IV U46 ( .A(B[455]), .Z(n59) );
  IV U47 ( .A(B[456]), .Z(n58) );
  IV U48 ( .A(B[457]), .Z(n57) );
  IV U49 ( .A(B[458]), .Z(n56) );
  IV U50 ( .A(B[459]), .Z(n55) );
  IV U51 ( .A(B[460]), .Z(n54) );
  IV U52 ( .A(B[461]), .Z(n53) );
  IV U53 ( .A(B[462]), .Z(n52) );
  IV U54 ( .A(B[0]), .Z(n514) );
  IV U55 ( .A(B[1]), .Z(n513) );
  IV U56 ( .A(B[2]), .Z(n512) );
  IV U57 ( .A(B[3]), .Z(n511) );
  IV U58 ( .A(B[4]), .Z(n510) );
  IV U59 ( .A(B[463]), .Z(n51) );
  IV U60 ( .A(B[5]), .Z(n509) );
  IV U61 ( .A(B[6]), .Z(n508) );
  IV U62 ( .A(B[7]), .Z(n507) );
  IV U63 ( .A(B[8]), .Z(n506) );
  IV U64 ( .A(B[9]), .Z(n505) );
  IV U65 ( .A(B[10]), .Z(n504) );
  IV U66 ( .A(B[11]), .Z(n503) );
  IV U67 ( .A(B[12]), .Z(n502) );
  IV U68 ( .A(B[13]), .Z(n501) );
  IV U69 ( .A(B[14]), .Z(n500) );
  IV U70 ( .A(B[464]), .Z(n50) );
  IV U71 ( .A(B[509]), .Z(n5) );
  IV U72 ( .A(B[15]), .Z(n499) );
  IV U73 ( .A(B[16]), .Z(n498) );
  IV U74 ( .A(B[17]), .Z(n497) );
  IV U75 ( .A(B[18]), .Z(n496) );
  IV U76 ( .A(B[19]), .Z(n495) );
  IV U77 ( .A(B[20]), .Z(n494) );
  IV U78 ( .A(B[21]), .Z(n493) );
  IV U79 ( .A(B[22]), .Z(n492) );
  IV U80 ( .A(B[23]), .Z(n491) );
  IV U81 ( .A(B[24]), .Z(n490) );
  IV U82 ( .A(B[465]), .Z(n49) );
  IV U83 ( .A(B[25]), .Z(n489) );
  IV U84 ( .A(B[26]), .Z(n488) );
  IV U85 ( .A(B[27]), .Z(n487) );
  IV U86 ( .A(B[28]), .Z(n486) );
  IV U87 ( .A(B[29]), .Z(n485) );
  IV U88 ( .A(B[30]), .Z(n484) );
  IV U89 ( .A(B[31]), .Z(n483) );
  IV U90 ( .A(B[32]), .Z(n482) );
  IV U91 ( .A(B[33]), .Z(n481) );
  IV U92 ( .A(B[34]), .Z(n480) );
  IV U93 ( .A(B[466]), .Z(n48) );
  IV U94 ( .A(B[35]), .Z(n479) );
  IV U95 ( .A(B[36]), .Z(n478) );
  IV U96 ( .A(B[37]), .Z(n477) );
  IV U97 ( .A(B[38]), .Z(n476) );
  IV U98 ( .A(B[39]), .Z(n475) );
  IV U99 ( .A(B[40]), .Z(n474) );
  IV U100 ( .A(B[41]), .Z(n473) );
  IV U101 ( .A(B[42]), .Z(n472) );
  IV U102 ( .A(B[43]), .Z(n471) );
  IV U103 ( .A(B[44]), .Z(n470) );
  IV U104 ( .A(B[467]), .Z(n47) );
  IV U105 ( .A(B[45]), .Z(n469) );
  IV U106 ( .A(B[46]), .Z(n468) );
  IV U107 ( .A(B[47]), .Z(n467) );
  IV U108 ( .A(B[48]), .Z(n466) );
  IV U109 ( .A(B[49]), .Z(n465) );
  IV U110 ( .A(B[50]), .Z(n464) );
  IV U111 ( .A(B[51]), .Z(n463) );
  IV U112 ( .A(B[52]), .Z(n462) );
  IV U113 ( .A(B[53]), .Z(n461) );
  IV U114 ( .A(B[54]), .Z(n460) );
  IV U115 ( .A(B[468]), .Z(n46) );
  IV U116 ( .A(B[55]), .Z(n459) );
  IV U117 ( .A(B[56]), .Z(n458) );
  IV U118 ( .A(B[57]), .Z(n457) );
  IV U119 ( .A(B[58]), .Z(n456) );
  IV U120 ( .A(B[59]), .Z(n455) );
  IV U121 ( .A(B[60]), .Z(n454) );
  IV U122 ( .A(B[61]), .Z(n453) );
  IV U123 ( .A(B[62]), .Z(n452) );
  IV U124 ( .A(B[63]), .Z(n451) );
  IV U125 ( .A(B[64]), .Z(n450) );
  IV U126 ( .A(B[469]), .Z(n45) );
  IV U127 ( .A(B[65]), .Z(n449) );
  IV U128 ( .A(B[66]), .Z(n448) );
  IV U129 ( .A(B[67]), .Z(n447) );
  IV U130 ( .A(B[68]), .Z(n446) );
  IV U131 ( .A(B[69]), .Z(n445) );
  IV U132 ( .A(B[70]), .Z(n444) );
  IV U133 ( .A(B[71]), .Z(n443) );
  IV U134 ( .A(B[72]), .Z(n442) );
  IV U135 ( .A(B[73]), .Z(n441) );
  IV U136 ( .A(B[74]), .Z(n440) );
  IV U137 ( .A(B[470]), .Z(n44) );
  IV U138 ( .A(B[75]), .Z(n439) );
  IV U139 ( .A(B[76]), .Z(n438) );
  IV U140 ( .A(B[77]), .Z(n437) );
  IV U141 ( .A(B[78]), .Z(n436) );
  IV U142 ( .A(B[79]), .Z(n435) );
  IV U143 ( .A(B[80]), .Z(n434) );
  IV U144 ( .A(B[81]), .Z(n433) );
  IV U145 ( .A(B[82]), .Z(n432) );
  IV U146 ( .A(B[83]), .Z(n431) );
  IV U147 ( .A(B[84]), .Z(n430) );
  IV U148 ( .A(B[471]), .Z(n43) );
  IV U149 ( .A(B[85]), .Z(n429) );
  IV U150 ( .A(B[86]), .Z(n428) );
  IV U151 ( .A(B[87]), .Z(n427) );
  IV U152 ( .A(B[88]), .Z(n426) );
  IV U153 ( .A(B[89]), .Z(n425) );
  IV U154 ( .A(B[90]), .Z(n424) );
  IV U155 ( .A(B[91]), .Z(n423) );
  IV U156 ( .A(B[92]), .Z(n422) );
  IV U157 ( .A(B[93]), .Z(n421) );
  IV U158 ( .A(B[94]), .Z(n420) );
  IV U159 ( .A(B[472]), .Z(n42) );
  IV U160 ( .A(B[95]), .Z(n419) );
  IV U161 ( .A(B[96]), .Z(n418) );
  IV U162 ( .A(B[97]), .Z(n417) );
  IV U163 ( .A(B[98]), .Z(n416) );
  IV U164 ( .A(B[99]), .Z(n415) );
  IV U165 ( .A(B[100]), .Z(n414) );
  IV U166 ( .A(B[101]), .Z(n413) );
  IV U167 ( .A(B[102]), .Z(n412) );
  IV U168 ( .A(B[103]), .Z(n411) );
  IV U169 ( .A(B[104]), .Z(n410) );
  IV U170 ( .A(B[473]), .Z(n41) );
  IV U171 ( .A(B[105]), .Z(n409) );
  IV U172 ( .A(B[106]), .Z(n408) );
  IV U173 ( .A(B[107]), .Z(n407) );
  IV U174 ( .A(B[108]), .Z(n406) );
  IV U175 ( .A(B[109]), .Z(n405) );
  IV U176 ( .A(B[110]), .Z(n404) );
  IV U177 ( .A(B[111]), .Z(n403) );
  IV U178 ( .A(B[112]), .Z(n402) );
  IV U179 ( .A(B[113]), .Z(n401) );
  IV U180 ( .A(B[114]), .Z(n400) );
  IV U181 ( .A(B[474]), .Z(n40) );
  IV U182 ( .A(B[510]), .Z(n4) );
  IV U183 ( .A(B[115]), .Z(n399) );
  IV U184 ( .A(B[116]), .Z(n398) );
  IV U185 ( .A(B[117]), .Z(n397) );
  IV U186 ( .A(B[118]), .Z(n396) );
  IV U187 ( .A(B[119]), .Z(n395) );
  IV U188 ( .A(B[120]), .Z(n394) );
  IV U189 ( .A(B[121]), .Z(n393) );
  IV U190 ( .A(B[122]), .Z(n392) );
  IV U191 ( .A(B[123]), .Z(n391) );
  IV U192 ( .A(B[124]), .Z(n390) );
  IV U193 ( .A(B[475]), .Z(n39) );
  IV U194 ( .A(B[125]), .Z(n389) );
  IV U195 ( .A(B[126]), .Z(n388) );
  IV U196 ( .A(B[127]), .Z(n387) );
  IV U197 ( .A(B[128]), .Z(n386) );
  IV U198 ( .A(B[129]), .Z(n385) );
  IV U199 ( .A(B[130]), .Z(n384) );
  IV U200 ( .A(B[131]), .Z(n383) );
  IV U201 ( .A(B[132]), .Z(n382) );
  IV U202 ( .A(B[133]), .Z(n381) );
  IV U203 ( .A(B[134]), .Z(n380) );
  IV U204 ( .A(B[476]), .Z(n38) );
  IV U205 ( .A(B[135]), .Z(n379) );
  IV U206 ( .A(B[136]), .Z(n378) );
  IV U207 ( .A(B[137]), .Z(n377) );
  IV U208 ( .A(B[138]), .Z(n376) );
  IV U209 ( .A(B[139]), .Z(n375) );
  IV U210 ( .A(B[140]), .Z(n374) );
  IV U211 ( .A(B[141]), .Z(n373) );
  IV U212 ( .A(B[142]), .Z(n372) );
  IV U213 ( .A(B[143]), .Z(n371) );
  IV U214 ( .A(B[144]), .Z(n370) );
  IV U215 ( .A(B[477]), .Z(n37) );
  IV U216 ( .A(B[145]), .Z(n369) );
  IV U217 ( .A(B[146]), .Z(n368) );
  IV U218 ( .A(B[147]), .Z(n367) );
  IV U219 ( .A(B[148]), .Z(n366) );
  IV U220 ( .A(B[149]), .Z(n365) );
  IV U221 ( .A(B[150]), .Z(n364) );
  IV U222 ( .A(B[151]), .Z(n363) );
  IV U223 ( .A(B[152]), .Z(n362) );
  IV U224 ( .A(B[153]), .Z(n361) );
  IV U225 ( .A(B[154]), .Z(n360) );
  IV U226 ( .A(B[478]), .Z(n36) );
  IV U227 ( .A(B[155]), .Z(n359) );
  IV U228 ( .A(B[156]), .Z(n358) );
  IV U229 ( .A(B[157]), .Z(n357) );
  IV U230 ( .A(B[158]), .Z(n356) );
  IV U231 ( .A(B[159]), .Z(n355) );
  IV U232 ( .A(B[160]), .Z(n354) );
  IV U233 ( .A(B[161]), .Z(n353) );
  IV U234 ( .A(B[162]), .Z(n352) );
  IV U235 ( .A(B[163]), .Z(n351) );
  IV U236 ( .A(B[164]), .Z(n350) );
  IV U237 ( .A(B[479]), .Z(n35) );
  IV U238 ( .A(B[165]), .Z(n349) );
  IV U239 ( .A(B[166]), .Z(n348) );
  IV U240 ( .A(B[167]), .Z(n347) );
  IV U241 ( .A(B[168]), .Z(n346) );
  IV U242 ( .A(B[169]), .Z(n345) );
  IV U243 ( .A(B[170]), .Z(n344) );
  IV U244 ( .A(B[171]), .Z(n343) );
  IV U245 ( .A(B[172]), .Z(n342) );
  IV U246 ( .A(B[173]), .Z(n341) );
  IV U247 ( .A(B[174]), .Z(n340) );
  IV U248 ( .A(B[480]), .Z(n34) );
  IV U249 ( .A(B[175]), .Z(n339) );
  IV U250 ( .A(B[176]), .Z(n338) );
  IV U251 ( .A(B[177]), .Z(n337) );
  IV U252 ( .A(B[178]), .Z(n336) );
  IV U253 ( .A(B[179]), .Z(n335) );
  IV U254 ( .A(B[180]), .Z(n334) );
  IV U255 ( .A(B[181]), .Z(n333) );
  IV U256 ( .A(B[182]), .Z(n332) );
  IV U257 ( .A(B[183]), .Z(n331) );
  IV U258 ( .A(B[184]), .Z(n330) );
  IV U259 ( .A(B[481]), .Z(n33) );
  IV U260 ( .A(B[185]), .Z(n329) );
  IV U261 ( .A(B[186]), .Z(n328) );
  IV U262 ( .A(B[187]), .Z(n327) );
  IV U263 ( .A(B[188]), .Z(n326) );
  IV U264 ( .A(B[189]), .Z(n325) );
  IV U265 ( .A(B[190]), .Z(n324) );
  IV U266 ( .A(B[191]), .Z(n323) );
  IV U267 ( .A(B[192]), .Z(n322) );
  IV U268 ( .A(B[193]), .Z(n321) );
  IV U269 ( .A(B[194]), .Z(n320) );
  IV U270 ( .A(B[482]), .Z(n32) );
  IV U271 ( .A(B[195]), .Z(n319) );
  IV U272 ( .A(B[196]), .Z(n318) );
  IV U273 ( .A(B[197]), .Z(n317) );
  IV U274 ( .A(B[198]), .Z(n316) );
  IV U275 ( .A(B[199]), .Z(n315) );
  IV U276 ( .A(B[200]), .Z(n314) );
  IV U277 ( .A(B[201]), .Z(n313) );
  IV U278 ( .A(B[202]), .Z(n312) );
  IV U279 ( .A(B[203]), .Z(n311) );
  IV U280 ( .A(B[204]), .Z(n310) );
  IV U281 ( .A(B[483]), .Z(n31) );
  IV U282 ( .A(B[205]), .Z(n309) );
  IV U283 ( .A(B[206]), .Z(n308) );
  IV U284 ( .A(B[207]), .Z(n307) );
  IV U285 ( .A(B[208]), .Z(n306) );
  IV U286 ( .A(B[209]), .Z(n305) );
  IV U287 ( .A(B[210]), .Z(n304) );
  IV U288 ( .A(B[211]), .Z(n303) );
  IV U289 ( .A(B[212]), .Z(n302) );
  IV U290 ( .A(B[213]), .Z(n301) );
  IV U291 ( .A(B[214]), .Z(n300) );
  IV U292 ( .A(B[484]), .Z(n30) );
  IV U293 ( .A(B[511]), .Z(n3) );
  IV U294 ( .A(B[215]), .Z(n299) );
  IV U295 ( .A(B[216]), .Z(n298) );
  IV U296 ( .A(B[217]), .Z(n297) );
  IV U297 ( .A(B[218]), .Z(n296) );
  IV U298 ( .A(B[219]), .Z(n295) );
  IV U299 ( .A(B[220]), .Z(n294) );
  IV U300 ( .A(B[221]), .Z(n293) );
  IV U301 ( .A(B[222]), .Z(n292) );
  IV U302 ( .A(B[223]), .Z(n291) );
  IV U303 ( .A(B[224]), .Z(n290) );
  IV U304 ( .A(B[485]), .Z(n29) );
  IV U305 ( .A(B[225]), .Z(n289) );
  IV U306 ( .A(B[226]), .Z(n288) );
  IV U307 ( .A(B[227]), .Z(n287) );
  IV U308 ( .A(B[228]), .Z(n286) );
  IV U309 ( .A(B[229]), .Z(n285) );
  IV U310 ( .A(B[230]), .Z(n284) );
  IV U311 ( .A(B[231]), .Z(n283) );
  IV U312 ( .A(B[232]), .Z(n282) );
  IV U313 ( .A(B[233]), .Z(n281) );
  IV U314 ( .A(B[234]), .Z(n280) );
  IV U315 ( .A(B[486]), .Z(n28) );
  IV U316 ( .A(B[235]), .Z(n279) );
  IV U317 ( .A(B[236]), .Z(n278) );
  IV U318 ( .A(B[237]), .Z(n277) );
  IV U319 ( .A(B[238]), .Z(n276) );
  IV U320 ( .A(B[239]), .Z(n275) );
  IV U321 ( .A(B[240]), .Z(n274) );
  IV U322 ( .A(B[241]), .Z(n273) );
  IV U323 ( .A(B[242]), .Z(n272) );
  IV U324 ( .A(B[243]), .Z(n271) );
  IV U325 ( .A(B[244]), .Z(n270) );
  IV U326 ( .A(B[487]), .Z(n27) );
  IV U327 ( .A(B[245]), .Z(n269) );
  IV U328 ( .A(B[246]), .Z(n268) );
  IV U329 ( .A(B[247]), .Z(n267) );
  IV U330 ( .A(B[248]), .Z(n266) );
  IV U331 ( .A(B[249]), .Z(n265) );
  IV U332 ( .A(B[250]), .Z(n264) );
  IV U333 ( .A(B[251]), .Z(n263) );
  IV U334 ( .A(B[252]), .Z(n262) );
  IV U335 ( .A(B[253]), .Z(n261) );
  IV U336 ( .A(B[254]), .Z(n260) );
  IV U337 ( .A(B[488]), .Z(n26) );
  IV U338 ( .A(B[255]), .Z(n259) );
  IV U339 ( .A(B[256]), .Z(n258) );
  IV U340 ( .A(B[257]), .Z(n257) );
  IV U341 ( .A(B[258]), .Z(n256) );
  IV U342 ( .A(B[259]), .Z(n255) );
  IV U343 ( .A(B[260]), .Z(n254) );
  IV U344 ( .A(B[261]), .Z(n253) );
  IV U345 ( .A(B[262]), .Z(n252) );
  IV U346 ( .A(B[263]), .Z(n251) );
  IV U347 ( .A(B[264]), .Z(n250) );
  IV U348 ( .A(B[489]), .Z(n25) );
  IV U349 ( .A(B[265]), .Z(n249) );
  IV U350 ( .A(B[266]), .Z(n248) );
  IV U351 ( .A(B[267]), .Z(n247) );
  IV U352 ( .A(B[268]), .Z(n246) );
  IV U353 ( .A(B[269]), .Z(n245) );
  IV U354 ( .A(B[270]), .Z(n244) );
  IV U355 ( .A(B[271]), .Z(n243) );
  IV U356 ( .A(B[272]), .Z(n242) );
  IV U357 ( .A(B[273]), .Z(n241) );
  IV U358 ( .A(B[274]), .Z(n240) );
  IV U359 ( .A(B[490]), .Z(n24) );
  IV U360 ( .A(B[275]), .Z(n239) );
  IV U361 ( .A(B[276]), .Z(n238) );
  IV U362 ( .A(B[277]), .Z(n237) );
  IV U363 ( .A(B[278]), .Z(n236) );
  IV U364 ( .A(B[279]), .Z(n235) );
  IV U365 ( .A(B[280]), .Z(n234) );
  IV U366 ( .A(B[281]), .Z(n233) );
  IV U367 ( .A(B[282]), .Z(n232) );
  IV U368 ( .A(B[283]), .Z(n231) );
  IV U369 ( .A(B[284]), .Z(n230) );
  IV U370 ( .A(B[491]), .Z(n23) );
  IV U371 ( .A(B[285]), .Z(n229) );
  IV U372 ( .A(B[286]), .Z(n228) );
  IV U373 ( .A(B[287]), .Z(n227) );
  IV U374 ( .A(B[288]), .Z(n226) );
  IV U375 ( .A(B[289]), .Z(n225) );
  IV U376 ( .A(B[290]), .Z(n224) );
  IV U377 ( .A(B[291]), .Z(n223) );
  IV U378 ( .A(B[292]), .Z(n222) );
  IV U379 ( .A(B[293]), .Z(n221) );
  IV U380 ( .A(B[294]), .Z(n220) );
  IV U381 ( .A(B[492]), .Z(n22) );
  IV U382 ( .A(B[295]), .Z(n219) );
  IV U383 ( .A(B[296]), .Z(n218) );
  IV U384 ( .A(B[297]), .Z(n217) );
  IV U385 ( .A(B[298]), .Z(n216) );
  IV U386 ( .A(B[299]), .Z(n215) );
  IV U387 ( .A(B[300]), .Z(n214) );
  IV U388 ( .A(B[301]), .Z(n213) );
  IV U389 ( .A(B[302]), .Z(n212) );
  IV U390 ( .A(B[303]), .Z(n211) );
  IV U391 ( .A(B[304]), .Z(n210) );
  IV U392 ( .A(B[493]), .Z(n21) );
  IV U393 ( .A(B[305]), .Z(n209) );
  IV U394 ( .A(B[306]), .Z(n208) );
  IV U395 ( .A(B[307]), .Z(n207) );
  IV U396 ( .A(B[308]), .Z(n206) );
  IV U397 ( .A(B[309]), .Z(n205) );
  IV U398 ( .A(B[310]), .Z(n204) );
  IV U399 ( .A(B[311]), .Z(n203) );
  IV U400 ( .A(B[312]), .Z(n202) );
  IV U401 ( .A(B[313]), .Z(n201) );
  IV U402 ( .A(B[314]), .Z(n200) );
  IV U403 ( .A(B[494]), .Z(n20) );
  IV U404 ( .A(B[315]), .Z(n199) );
  IV U405 ( .A(B[316]), .Z(n198) );
  IV U406 ( .A(B[317]), .Z(n197) );
  IV U407 ( .A(B[318]), .Z(n196) );
  IV U408 ( .A(B[319]), .Z(n195) );
  IV U409 ( .A(B[320]), .Z(n194) );
  IV U410 ( .A(B[321]), .Z(n193) );
  IV U411 ( .A(B[322]), .Z(n192) );
  IV U412 ( .A(B[323]), .Z(n191) );
  IV U413 ( .A(B[324]), .Z(n190) );
  IV U414 ( .A(B[495]), .Z(n19) );
  IV U415 ( .A(B[325]), .Z(n189) );
  IV U416 ( .A(B[326]), .Z(n188) );
  IV U417 ( .A(B[327]), .Z(n187) );
  IV U418 ( .A(B[328]), .Z(n186) );
  IV U419 ( .A(B[329]), .Z(n185) );
  IV U420 ( .A(B[330]), .Z(n184) );
  IV U421 ( .A(B[331]), .Z(n183) );
  IV U422 ( .A(B[332]), .Z(n182) );
  IV U423 ( .A(B[333]), .Z(n181) );
  IV U424 ( .A(B[334]), .Z(n180) );
  IV U425 ( .A(B[496]), .Z(n18) );
  IV U426 ( .A(B[335]), .Z(n179) );
  IV U427 ( .A(B[336]), .Z(n178) );
  IV U428 ( .A(B[337]), .Z(n177) );
  IV U429 ( .A(B[338]), .Z(n176) );
  IV U430 ( .A(B[339]), .Z(n175) );
  IV U431 ( .A(B[340]), .Z(n174) );
  IV U432 ( .A(B[341]), .Z(n173) );
  IV U433 ( .A(B[342]), .Z(n172) );
  IV U434 ( .A(B[343]), .Z(n171) );
  IV U435 ( .A(B[344]), .Z(n170) );
  IV U436 ( .A(B[497]), .Z(n17) );
  IV U437 ( .A(B[345]), .Z(n169) );
  IV U438 ( .A(B[346]), .Z(n168) );
  IV U439 ( .A(B[347]), .Z(n167) );
  IV U440 ( .A(B[348]), .Z(n166) );
  IV U441 ( .A(B[349]), .Z(n165) );
  IV U442 ( .A(B[350]), .Z(n164) );
  IV U443 ( .A(B[351]), .Z(n163) );
  IV U444 ( .A(B[352]), .Z(n162) );
  IV U445 ( .A(B[353]), .Z(n161) );
  IV U446 ( .A(B[354]), .Z(n160) );
  IV U447 ( .A(B[498]), .Z(n16) );
  IV U448 ( .A(B[355]), .Z(n159) );
  IV U449 ( .A(B[356]), .Z(n158) );
  IV U450 ( .A(B[357]), .Z(n157) );
  IV U451 ( .A(B[358]), .Z(n156) );
  IV U452 ( .A(B[359]), .Z(n155) );
  IV U453 ( .A(B[360]), .Z(n154) );
  IV U454 ( .A(B[361]), .Z(n153) );
  IV U455 ( .A(B[362]), .Z(n152) );
  IV U456 ( .A(B[363]), .Z(n151) );
  IV U457 ( .A(B[364]), .Z(n150) );
  IV U458 ( .A(B[499]), .Z(n15) );
  IV U459 ( .A(B[365]), .Z(n149) );
  IV U460 ( .A(B[366]), .Z(n148) );
  IV U461 ( .A(B[367]), .Z(n147) );
  IV U462 ( .A(B[368]), .Z(n146) );
  IV U463 ( .A(B[369]), .Z(n145) );
  IV U464 ( .A(B[370]), .Z(n144) );
  IV U465 ( .A(B[371]), .Z(n143) );
  IV U466 ( .A(B[372]), .Z(n142) );
  IV U467 ( .A(B[373]), .Z(n141) );
  IV U468 ( .A(B[374]), .Z(n140) );
  IV U469 ( .A(B[500]), .Z(n14) );
  IV U470 ( .A(B[375]), .Z(n139) );
  IV U471 ( .A(B[376]), .Z(n138) );
  IV U472 ( .A(B[377]), .Z(n137) );
  IV U473 ( .A(B[378]), .Z(n136) );
  IV U474 ( .A(B[379]), .Z(n135) );
  IV U475 ( .A(B[380]), .Z(n134) );
  IV U476 ( .A(B[381]), .Z(n133) );
  IV U477 ( .A(B[382]), .Z(n132) );
  IV U478 ( .A(B[383]), .Z(n131) );
  IV U479 ( .A(B[384]), .Z(n130) );
  IV U480 ( .A(B[501]), .Z(n13) );
  IV U481 ( .A(B[385]), .Z(n129) );
  IV U482 ( .A(B[386]), .Z(n128) );
  IV U483 ( .A(B[387]), .Z(n127) );
  IV U484 ( .A(B[388]), .Z(n126) );
  IV U485 ( .A(B[389]), .Z(n125) );
  IV U486 ( .A(B[390]), .Z(n124) );
  IV U487 ( .A(B[391]), .Z(n123) );
  IV U488 ( .A(B[392]), .Z(n122) );
  IV U489 ( .A(B[393]), .Z(n121) );
  IV U490 ( .A(B[394]), .Z(n120) );
  IV U491 ( .A(B[502]), .Z(n12) );
  IV U492 ( .A(B[395]), .Z(n119) );
  IV U493 ( .A(B[396]), .Z(n118) );
  IV U494 ( .A(B[397]), .Z(n117) );
  IV U495 ( .A(B[398]), .Z(n116) );
  IV U496 ( .A(B[399]), .Z(n115) );
  IV U497 ( .A(B[400]), .Z(n114) );
  IV U498 ( .A(B[401]), .Z(n113) );
  IV U499 ( .A(B[402]), .Z(n112) );
  IV U500 ( .A(B[403]), .Z(n111) );
  IV U501 ( .A(B[404]), .Z(n110) );
  IV U502 ( .A(B[503]), .Z(n11) );
  IV U503 ( .A(B[405]), .Z(n109) );
  IV U504 ( .A(B[406]), .Z(n108) );
  IV U505 ( .A(B[407]), .Z(n107) );
  IV U506 ( .A(B[408]), .Z(n106) );
  IV U507 ( .A(B[409]), .Z(n105) );
  IV U508 ( .A(B[410]), .Z(n104) );
  IV U509 ( .A(B[411]), .Z(n103) );
  IV U510 ( .A(B[412]), .Z(n102) );
  IV U511 ( .A(B[413]), .Z(n101) );
  IV U512 ( .A(B[414]), .Z(n100) );
  IV U513 ( .A(B[504]), .Z(n10) );
endmodule


module MUX_N514_7 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N514_8 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_9521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_9522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_9523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_9999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_10034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N514_5 ( A, B, O );
  input [513:0] A;
  input [513:0] B;
  output O;
  wire   n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  wire   [513:1] C;

  FA_10034 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n516), .CI(1'b1), 
        .CO(C[1]) );
  FA_10033 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n517), .CI(C[1]), 
        .CO(C[2]) );
  FA_10032 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n518), .CI(C[2]), 
        .CO(C[3]) );
  FA_10031 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n519), .CI(C[3]), 
        .CO(C[4]) );
  FA_10030 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n520), .CI(C[4]), 
        .CO(C[5]) );
  FA_10029 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n521), .CI(C[5]), 
        .CO(C[6]) );
  FA_10028 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n522), .CI(C[6]), 
        .CO(C[7]) );
  FA_10027 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n523), .CI(C[7]), 
        .CO(C[8]) );
  FA_10026 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n524), .CI(C[8]), 
        .CO(C[9]) );
  FA_10025 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n525), .CI(C[9]), 
        .CO(C[10]) );
  FA_10024 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n526), .CI(C[10]), 
        .CO(C[11]) );
  FA_10023 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n527), .CI(C[11]), 
        .CO(C[12]) );
  FA_10022 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n528), .CI(C[12]), 
        .CO(C[13]) );
  FA_10021 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n529), .CI(C[13]), 
        .CO(C[14]) );
  FA_10020 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n530), .CI(C[14]), 
        .CO(C[15]) );
  FA_10019 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n531), .CI(C[15]), 
        .CO(C[16]) );
  FA_10018 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n532), .CI(C[16]), 
        .CO(C[17]) );
  FA_10017 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n533), .CI(C[17]), 
        .CO(C[18]) );
  FA_10016 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n534), .CI(C[18]), 
        .CO(C[19]) );
  FA_10015 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n535), .CI(C[19]), 
        .CO(C[20]) );
  FA_10014 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n536), .CI(C[20]), 
        .CO(C[21]) );
  FA_10013 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n537), .CI(C[21]), 
        .CO(C[22]) );
  FA_10012 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n538), .CI(C[22]), 
        .CO(C[23]) );
  FA_10011 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n539), .CI(C[23]), 
        .CO(C[24]) );
  FA_10010 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n540), .CI(C[24]), 
        .CO(C[25]) );
  FA_10009 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n541), .CI(C[25]), 
        .CO(C[26]) );
  FA_10008 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n542), .CI(C[26]), 
        .CO(C[27]) );
  FA_10007 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n543), .CI(C[27]), 
        .CO(C[28]) );
  FA_10006 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n544), .CI(C[28]), 
        .CO(C[29]) );
  FA_10005 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n545), .CI(C[29]), 
        .CO(C[30]) );
  FA_10004 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n546), .CI(C[30]), 
        .CO(C[31]) );
  FA_10003 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n547), .CI(C[31]), 
        .CO(C[32]) );
  FA_10002 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n548), .CI(C[32]), 
        .CO(C[33]) );
  FA_10001 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n549), .CI(C[33]), 
        .CO(C[34]) );
  FA_10000 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n550), .CI(C[34]), 
        .CO(C[35]) );
  FA_9999 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n551), .CI(C[35]), 
        .CO(C[36]) );
  FA_9998 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n552), .CI(C[36]), 
        .CO(C[37]) );
  FA_9997 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n553), .CI(C[37]), 
        .CO(C[38]) );
  FA_9996 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n554), .CI(C[38]), 
        .CO(C[39]) );
  FA_9995 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n555), .CI(C[39]), 
        .CO(C[40]) );
  FA_9994 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n556), .CI(C[40]), 
        .CO(C[41]) );
  FA_9993 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n557), .CI(C[41]), 
        .CO(C[42]) );
  FA_9992 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n558), .CI(C[42]), 
        .CO(C[43]) );
  FA_9991 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n559), .CI(C[43]), 
        .CO(C[44]) );
  FA_9990 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n560), .CI(C[44]), 
        .CO(C[45]) );
  FA_9989 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n561), .CI(C[45]), 
        .CO(C[46]) );
  FA_9988 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n562), .CI(C[46]), 
        .CO(C[47]) );
  FA_9987 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n563), .CI(C[47]), 
        .CO(C[48]) );
  FA_9986 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n564), .CI(C[48]), 
        .CO(C[49]) );
  FA_9985 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n565), .CI(C[49]), 
        .CO(C[50]) );
  FA_9984 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n566), .CI(C[50]), 
        .CO(C[51]) );
  FA_9983 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n567), .CI(C[51]), 
        .CO(C[52]) );
  FA_9982 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n568), .CI(C[52]), 
        .CO(C[53]) );
  FA_9981 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n569), .CI(C[53]), 
        .CO(C[54]) );
  FA_9980 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n570), .CI(C[54]), 
        .CO(C[55]) );
  FA_9979 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n571), .CI(C[55]), 
        .CO(C[56]) );
  FA_9978 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n572), .CI(C[56]), 
        .CO(C[57]) );
  FA_9977 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n573), .CI(C[57]), 
        .CO(C[58]) );
  FA_9976 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n574), .CI(C[58]), 
        .CO(C[59]) );
  FA_9975 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n575), .CI(C[59]), 
        .CO(C[60]) );
  FA_9974 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n576), .CI(C[60]), 
        .CO(C[61]) );
  FA_9973 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n577), .CI(C[61]), 
        .CO(C[62]) );
  FA_9972 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n578), .CI(C[62]), 
        .CO(C[63]) );
  FA_9971 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n579), .CI(C[63]), 
        .CO(C[64]) );
  FA_9970 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n580), .CI(C[64]), 
        .CO(C[65]) );
  FA_9969 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n581), .CI(C[65]), 
        .CO(C[66]) );
  FA_9968 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n582), .CI(C[66]), 
        .CO(C[67]) );
  FA_9967 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n583), .CI(C[67]), 
        .CO(C[68]) );
  FA_9966 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n584), .CI(C[68]), 
        .CO(C[69]) );
  FA_9965 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n585), .CI(C[69]), 
        .CO(C[70]) );
  FA_9964 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n586), .CI(C[70]), 
        .CO(C[71]) );
  FA_9963 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n587), .CI(C[71]), 
        .CO(C[72]) );
  FA_9962 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n588), .CI(C[72]), 
        .CO(C[73]) );
  FA_9961 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n589), .CI(C[73]), 
        .CO(C[74]) );
  FA_9960 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n590), .CI(C[74]), 
        .CO(C[75]) );
  FA_9959 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n591), .CI(C[75]), 
        .CO(C[76]) );
  FA_9958 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n592), .CI(C[76]), 
        .CO(C[77]) );
  FA_9957 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n593), .CI(C[77]), 
        .CO(C[78]) );
  FA_9956 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n594), .CI(C[78]), 
        .CO(C[79]) );
  FA_9955 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n595), .CI(C[79]), 
        .CO(C[80]) );
  FA_9954 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n596), .CI(C[80]), 
        .CO(C[81]) );
  FA_9953 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n597), .CI(C[81]), 
        .CO(C[82]) );
  FA_9952 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n598), .CI(C[82]), 
        .CO(C[83]) );
  FA_9951 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n599), .CI(C[83]), 
        .CO(C[84]) );
  FA_9950 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n600), .CI(C[84]), 
        .CO(C[85]) );
  FA_9949 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n601), .CI(C[85]), 
        .CO(C[86]) );
  FA_9948 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n602), .CI(C[86]), 
        .CO(C[87]) );
  FA_9947 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n603), .CI(C[87]), 
        .CO(C[88]) );
  FA_9946 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n604), .CI(C[88]), 
        .CO(C[89]) );
  FA_9945 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n605), .CI(C[89]), 
        .CO(C[90]) );
  FA_9944 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n606), .CI(C[90]), 
        .CO(C[91]) );
  FA_9943 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n607), .CI(C[91]), 
        .CO(C[92]) );
  FA_9942 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n608), .CI(C[92]), 
        .CO(C[93]) );
  FA_9941 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n609), .CI(C[93]), 
        .CO(C[94]) );
  FA_9940 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n610), .CI(C[94]), 
        .CO(C[95]) );
  FA_9939 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n611), .CI(C[95]), 
        .CO(C[96]) );
  FA_9938 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n612), .CI(C[96]), 
        .CO(C[97]) );
  FA_9937 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n613), .CI(C[97]), 
        .CO(C[98]) );
  FA_9936 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n614), .CI(C[98]), 
        .CO(C[99]) );
  FA_9935 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n615), .CI(C[99]), 
        .CO(C[100]) );
  FA_9934 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n616), .CI(C[100]), .CO(C[101]) );
  FA_9933 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n617), .CI(C[101]), .CO(C[102]) );
  FA_9932 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n618), .CI(C[102]), .CO(C[103]) );
  FA_9931 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n619), .CI(C[103]), .CO(C[104]) );
  FA_9930 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n620), .CI(C[104]), .CO(C[105]) );
  FA_9929 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n621), .CI(C[105]), .CO(C[106]) );
  FA_9928 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n622), .CI(C[106]), .CO(C[107]) );
  FA_9927 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n623), .CI(C[107]), .CO(C[108]) );
  FA_9926 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n624), .CI(C[108]), .CO(C[109]) );
  FA_9925 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n625), .CI(C[109]), .CO(C[110]) );
  FA_9924 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n626), .CI(C[110]), .CO(C[111]) );
  FA_9923 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n627), .CI(C[111]), .CO(C[112]) );
  FA_9922 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n628), .CI(C[112]), .CO(C[113]) );
  FA_9921 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n629), .CI(C[113]), .CO(C[114]) );
  FA_9920 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n630), .CI(C[114]), .CO(C[115]) );
  FA_9919 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n631), .CI(C[115]), .CO(C[116]) );
  FA_9918 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n632), .CI(C[116]), .CO(C[117]) );
  FA_9917 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n633), .CI(C[117]), .CO(C[118]) );
  FA_9916 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n634), .CI(C[118]), .CO(C[119]) );
  FA_9915 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n635), .CI(C[119]), .CO(C[120]) );
  FA_9914 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n636), .CI(C[120]), .CO(C[121]) );
  FA_9913 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n637), .CI(C[121]), .CO(C[122]) );
  FA_9912 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n638), .CI(C[122]), .CO(C[123]) );
  FA_9911 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n639), .CI(C[123]), .CO(C[124]) );
  FA_9910 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n640), .CI(C[124]), .CO(C[125]) );
  FA_9909 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n641), .CI(C[125]), .CO(C[126]) );
  FA_9908 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n642), .CI(C[126]), .CO(C[127]) );
  FA_9907 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n643), .CI(C[127]), .CO(C[128]) );
  FA_9906 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n644), .CI(C[128]), .CO(C[129]) );
  FA_9905 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n645), .CI(C[129]), .CO(C[130]) );
  FA_9904 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n646), .CI(C[130]), .CO(C[131]) );
  FA_9903 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n647), .CI(C[131]), .CO(C[132]) );
  FA_9902 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n648), .CI(C[132]), .CO(C[133]) );
  FA_9901 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n649), .CI(C[133]), .CO(C[134]) );
  FA_9900 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n650), .CI(C[134]), .CO(C[135]) );
  FA_9899 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n651), .CI(C[135]), .CO(C[136]) );
  FA_9898 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n652), .CI(C[136]), .CO(C[137]) );
  FA_9897 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n653), .CI(C[137]), .CO(C[138]) );
  FA_9896 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n654), .CI(C[138]), .CO(C[139]) );
  FA_9895 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n655), .CI(C[139]), .CO(C[140]) );
  FA_9894 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n656), .CI(C[140]), .CO(C[141]) );
  FA_9893 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n657), .CI(C[141]), .CO(C[142]) );
  FA_9892 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n658), .CI(C[142]), .CO(C[143]) );
  FA_9891 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n659), .CI(C[143]), .CO(C[144]) );
  FA_9890 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n660), .CI(C[144]), .CO(C[145]) );
  FA_9889 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n661), .CI(C[145]), .CO(C[146]) );
  FA_9888 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n662), .CI(C[146]), .CO(C[147]) );
  FA_9887 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n663), .CI(C[147]), .CO(C[148]) );
  FA_9886 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n664), .CI(C[148]), .CO(C[149]) );
  FA_9885 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n665), .CI(C[149]), .CO(C[150]) );
  FA_9884 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n666), .CI(C[150]), .CO(C[151]) );
  FA_9883 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n667), .CI(C[151]), .CO(C[152]) );
  FA_9882 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n668), .CI(C[152]), .CO(C[153]) );
  FA_9881 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n669), .CI(C[153]), .CO(C[154]) );
  FA_9880 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n670), .CI(C[154]), .CO(C[155]) );
  FA_9879 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n671), .CI(C[155]), .CO(C[156]) );
  FA_9878 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n672), .CI(C[156]), .CO(C[157]) );
  FA_9877 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n673), .CI(C[157]), .CO(C[158]) );
  FA_9876 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n674), .CI(C[158]), .CO(C[159]) );
  FA_9875 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n675), .CI(C[159]), .CO(C[160]) );
  FA_9874 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n676), .CI(C[160]), .CO(C[161]) );
  FA_9873 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n677), .CI(C[161]), .CO(C[162]) );
  FA_9872 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n678), .CI(C[162]), .CO(C[163]) );
  FA_9871 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n679), .CI(C[163]), .CO(C[164]) );
  FA_9870 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n680), .CI(C[164]), .CO(C[165]) );
  FA_9869 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n681), .CI(C[165]), .CO(C[166]) );
  FA_9868 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n682), .CI(C[166]), .CO(C[167]) );
  FA_9867 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n683), .CI(C[167]), .CO(C[168]) );
  FA_9866 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n684), .CI(C[168]), .CO(C[169]) );
  FA_9865 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n685), .CI(C[169]), .CO(C[170]) );
  FA_9864 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n686), .CI(C[170]), .CO(C[171]) );
  FA_9863 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n687), .CI(C[171]), .CO(C[172]) );
  FA_9862 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n688), .CI(C[172]), .CO(C[173]) );
  FA_9861 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n689), .CI(C[173]), .CO(C[174]) );
  FA_9860 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n690), .CI(C[174]), .CO(C[175]) );
  FA_9859 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n691), .CI(C[175]), .CO(C[176]) );
  FA_9858 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n692), .CI(C[176]), .CO(C[177]) );
  FA_9857 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n693), .CI(C[177]), .CO(C[178]) );
  FA_9856 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n694), .CI(C[178]), .CO(C[179]) );
  FA_9855 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n695), .CI(C[179]), .CO(C[180]) );
  FA_9854 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n696), .CI(C[180]), .CO(C[181]) );
  FA_9853 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n697), .CI(C[181]), .CO(C[182]) );
  FA_9852 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n698), .CI(C[182]), .CO(C[183]) );
  FA_9851 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n699), .CI(C[183]), .CO(C[184]) );
  FA_9850 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n700), .CI(C[184]), .CO(C[185]) );
  FA_9849 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n701), .CI(C[185]), .CO(C[186]) );
  FA_9848 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n702), .CI(C[186]), .CO(C[187]) );
  FA_9847 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n703), .CI(C[187]), .CO(C[188]) );
  FA_9846 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n704), .CI(C[188]), .CO(C[189]) );
  FA_9845 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n705), .CI(C[189]), .CO(C[190]) );
  FA_9844 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n706), .CI(C[190]), .CO(C[191]) );
  FA_9843 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n707), .CI(C[191]), .CO(C[192]) );
  FA_9842 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n708), .CI(C[192]), .CO(C[193]) );
  FA_9841 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n709), .CI(C[193]), .CO(C[194]) );
  FA_9840 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n710), .CI(C[194]), .CO(C[195]) );
  FA_9839 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n711), .CI(C[195]), .CO(C[196]) );
  FA_9838 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n712), .CI(C[196]), .CO(C[197]) );
  FA_9837 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n713), .CI(C[197]), .CO(C[198]) );
  FA_9836 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n714), .CI(C[198]), .CO(C[199]) );
  FA_9835 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n715), .CI(C[199]), .CO(C[200]) );
  FA_9834 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n716), .CI(C[200]), .CO(C[201]) );
  FA_9833 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n717), .CI(C[201]), .CO(C[202]) );
  FA_9832 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n718), .CI(C[202]), .CO(C[203]) );
  FA_9831 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n719), .CI(C[203]), .CO(C[204]) );
  FA_9830 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n720), .CI(C[204]), .CO(C[205]) );
  FA_9829 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n721), .CI(C[205]), .CO(C[206]) );
  FA_9828 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n722), .CI(C[206]), .CO(C[207]) );
  FA_9827 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n723), .CI(C[207]), .CO(C[208]) );
  FA_9826 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n724), .CI(C[208]), .CO(C[209]) );
  FA_9825 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n725), .CI(C[209]), .CO(C[210]) );
  FA_9824 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n726), .CI(C[210]), .CO(C[211]) );
  FA_9823 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n727), .CI(C[211]), .CO(C[212]) );
  FA_9822 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n728), .CI(C[212]), .CO(C[213]) );
  FA_9821 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n729), .CI(C[213]), .CO(C[214]) );
  FA_9820 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n730), .CI(C[214]), .CO(C[215]) );
  FA_9819 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n731), .CI(C[215]), .CO(C[216]) );
  FA_9818 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n732), .CI(C[216]), .CO(C[217]) );
  FA_9817 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n733), .CI(C[217]), .CO(C[218]) );
  FA_9816 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n734), .CI(C[218]), .CO(C[219]) );
  FA_9815 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n735), .CI(C[219]), .CO(C[220]) );
  FA_9814 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n736), .CI(C[220]), .CO(C[221]) );
  FA_9813 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n737), .CI(C[221]), .CO(C[222]) );
  FA_9812 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n738), .CI(C[222]), .CO(C[223]) );
  FA_9811 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n739), .CI(C[223]), .CO(C[224]) );
  FA_9810 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n740), .CI(C[224]), .CO(C[225]) );
  FA_9809 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n741), .CI(C[225]), .CO(C[226]) );
  FA_9808 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n742), .CI(C[226]), .CO(C[227]) );
  FA_9807 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n743), .CI(C[227]), .CO(C[228]) );
  FA_9806 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n744), .CI(C[228]), .CO(C[229]) );
  FA_9805 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n745), .CI(C[229]), .CO(C[230]) );
  FA_9804 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n746), .CI(C[230]), .CO(C[231]) );
  FA_9803 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n747), .CI(C[231]), .CO(C[232]) );
  FA_9802 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n748), .CI(C[232]), .CO(C[233]) );
  FA_9801 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n749), .CI(C[233]), .CO(C[234]) );
  FA_9800 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n750), .CI(C[234]), .CO(C[235]) );
  FA_9799 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n751), .CI(C[235]), .CO(C[236]) );
  FA_9798 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n752), .CI(C[236]), .CO(C[237]) );
  FA_9797 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n753), .CI(C[237]), .CO(C[238]) );
  FA_9796 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n754), .CI(C[238]), .CO(C[239]) );
  FA_9795 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n755), .CI(C[239]), .CO(C[240]) );
  FA_9794 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n756), .CI(C[240]), .CO(C[241]) );
  FA_9793 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n757), .CI(C[241]), .CO(C[242]) );
  FA_9792 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n758), .CI(C[242]), .CO(C[243]) );
  FA_9791 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n759), .CI(C[243]), .CO(C[244]) );
  FA_9790 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n760), .CI(C[244]), .CO(C[245]) );
  FA_9789 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n761), .CI(C[245]), .CO(C[246]) );
  FA_9788 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n762), .CI(C[246]), .CO(C[247]) );
  FA_9787 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n763), .CI(C[247]), .CO(C[248]) );
  FA_9786 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n764), .CI(C[248]), .CO(C[249]) );
  FA_9785 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n765), .CI(C[249]), .CO(C[250]) );
  FA_9784 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n766), .CI(C[250]), .CO(C[251]) );
  FA_9783 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n767), .CI(C[251]), .CO(C[252]) );
  FA_9782 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n768), .CI(C[252]), .CO(C[253]) );
  FA_9781 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n769), .CI(C[253]), .CO(C[254]) );
  FA_9780 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n770), .CI(C[254]), .CO(C[255]) );
  FA_9779 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n771), .CI(C[255]), .CO(C[256]) );
  FA_9778 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n772), .CI(C[256]), .CO(C[257]) );
  FA_9777 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n773), .CI(C[257]), .CO(C[258]) );
  FA_9776 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n774), .CI(C[258]), .CO(C[259]) );
  FA_9775 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n775), .CI(C[259]), .CO(C[260]) );
  FA_9774 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n776), .CI(C[260]), .CO(C[261]) );
  FA_9773 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n777), .CI(C[261]), .CO(C[262]) );
  FA_9772 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n778), .CI(C[262]), .CO(C[263]) );
  FA_9771 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n779), .CI(C[263]), .CO(C[264]) );
  FA_9770 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n780), .CI(C[264]), .CO(C[265]) );
  FA_9769 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n781), .CI(C[265]), .CO(C[266]) );
  FA_9768 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n782), .CI(C[266]), .CO(C[267]) );
  FA_9767 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n783), .CI(C[267]), .CO(C[268]) );
  FA_9766 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n784), .CI(C[268]), .CO(C[269]) );
  FA_9765 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n785), .CI(C[269]), .CO(C[270]) );
  FA_9764 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n786), .CI(C[270]), .CO(C[271]) );
  FA_9763 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n787), .CI(C[271]), .CO(C[272]) );
  FA_9762 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n788), .CI(C[272]), .CO(C[273]) );
  FA_9761 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n789), .CI(C[273]), .CO(C[274]) );
  FA_9760 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n790), .CI(C[274]), .CO(C[275]) );
  FA_9759 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n791), .CI(C[275]), .CO(C[276]) );
  FA_9758 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n792), .CI(C[276]), .CO(C[277]) );
  FA_9757 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n793), .CI(C[277]), .CO(C[278]) );
  FA_9756 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n794), .CI(C[278]), .CO(C[279]) );
  FA_9755 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n795), .CI(C[279]), .CO(C[280]) );
  FA_9754 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n796), .CI(C[280]), .CO(C[281]) );
  FA_9753 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n797), .CI(C[281]), .CO(C[282]) );
  FA_9752 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n798), .CI(C[282]), .CO(C[283]) );
  FA_9751 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n799), .CI(C[283]), .CO(C[284]) );
  FA_9750 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n800), .CI(C[284]), .CO(C[285]) );
  FA_9749 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n801), .CI(C[285]), .CO(C[286]) );
  FA_9748 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n802), .CI(C[286]), .CO(C[287]) );
  FA_9747 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n803), .CI(C[287]), .CO(C[288]) );
  FA_9746 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n804), .CI(C[288]), .CO(C[289]) );
  FA_9745 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n805), .CI(C[289]), .CO(C[290]) );
  FA_9744 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n806), .CI(C[290]), .CO(C[291]) );
  FA_9743 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n807), .CI(C[291]), .CO(C[292]) );
  FA_9742 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n808), .CI(C[292]), .CO(C[293]) );
  FA_9741 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n809), .CI(C[293]), .CO(C[294]) );
  FA_9740 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n810), .CI(C[294]), .CO(C[295]) );
  FA_9739 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n811), .CI(C[295]), .CO(C[296]) );
  FA_9738 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n812), .CI(C[296]), .CO(C[297]) );
  FA_9737 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n813), .CI(C[297]), .CO(C[298]) );
  FA_9736 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n814), .CI(C[298]), .CO(C[299]) );
  FA_9735 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n815), .CI(C[299]), .CO(C[300]) );
  FA_9734 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n816), .CI(C[300]), .CO(C[301]) );
  FA_9733 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n817), .CI(C[301]), .CO(C[302]) );
  FA_9732 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n818), .CI(C[302]), .CO(C[303]) );
  FA_9731 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n819), .CI(C[303]), .CO(C[304]) );
  FA_9730 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n820), .CI(C[304]), .CO(C[305]) );
  FA_9729 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n821), .CI(C[305]), .CO(C[306]) );
  FA_9728 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n822), .CI(C[306]), .CO(C[307]) );
  FA_9727 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n823), .CI(C[307]), .CO(C[308]) );
  FA_9726 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n824), .CI(C[308]), .CO(C[309]) );
  FA_9725 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n825), .CI(C[309]), .CO(C[310]) );
  FA_9724 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n826), .CI(C[310]), .CO(C[311]) );
  FA_9723 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n827), .CI(C[311]), .CO(C[312]) );
  FA_9722 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n828), .CI(C[312]), .CO(C[313]) );
  FA_9721 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n829), .CI(C[313]), .CO(C[314]) );
  FA_9720 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n830), .CI(C[314]), .CO(C[315]) );
  FA_9719 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n831), .CI(C[315]), .CO(C[316]) );
  FA_9718 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n832), .CI(C[316]), .CO(C[317]) );
  FA_9717 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n833), .CI(C[317]), .CO(C[318]) );
  FA_9716 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n834), .CI(C[318]), .CO(C[319]) );
  FA_9715 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n835), .CI(C[319]), .CO(C[320]) );
  FA_9714 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n836), .CI(C[320]), .CO(C[321]) );
  FA_9713 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n837), .CI(C[321]), .CO(C[322]) );
  FA_9712 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n838), .CI(C[322]), .CO(C[323]) );
  FA_9711 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n839), .CI(C[323]), .CO(C[324]) );
  FA_9710 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n840), .CI(C[324]), .CO(C[325]) );
  FA_9709 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n841), .CI(C[325]), .CO(C[326]) );
  FA_9708 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n842), .CI(C[326]), .CO(C[327]) );
  FA_9707 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n843), .CI(C[327]), .CO(C[328]) );
  FA_9706 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n844), .CI(C[328]), .CO(C[329]) );
  FA_9705 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n845), .CI(C[329]), .CO(C[330]) );
  FA_9704 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n846), .CI(C[330]), .CO(C[331]) );
  FA_9703 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n847), .CI(C[331]), .CO(C[332]) );
  FA_9702 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n848), .CI(C[332]), .CO(C[333]) );
  FA_9701 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n849), .CI(C[333]), .CO(C[334]) );
  FA_9700 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n850), .CI(C[334]), .CO(C[335]) );
  FA_9699 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n851), .CI(C[335]), .CO(C[336]) );
  FA_9698 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n852), .CI(C[336]), .CO(C[337]) );
  FA_9697 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n853), .CI(C[337]), .CO(C[338]) );
  FA_9696 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n854), .CI(C[338]), .CO(C[339]) );
  FA_9695 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n855), .CI(C[339]), .CO(C[340]) );
  FA_9694 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n856), .CI(C[340]), .CO(C[341]) );
  FA_9693 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n857), .CI(C[341]), .CO(C[342]) );
  FA_9692 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n858), .CI(C[342]), .CO(C[343]) );
  FA_9691 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n859), .CI(C[343]), .CO(C[344]) );
  FA_9690 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n860), .CI(C[344]), .CO(C[345]) );
  FA_9689 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n861), .CI(C[345]), .CO(C[346]) );
  FA_9688 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n862), .CI(C[346]), .CO(C[347]) );
  FA_9687 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n863), .CI(C[347]), .CO(C[348]) );
  FA_9686 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n864), .CI(C[348]), .CO(C[349]) );
  FA_9685 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n865), .CI(C[349]), .CO(C[350]) );
  FA_9684 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n866), .CI(C[350]), .CO(C[351]) );
  FA_9683 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n867), .CI(C[351]), .CO(C[352]) );
  FA_9682 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n868), .CI(C[352]), .CO(C[353]) );
  FA_9681 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n869), .CI(C[353]), .CO(C[354]) );
  FA_9680 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n870), .CI(C[354]), .CO(C[355]) );
  FA_9679 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n871), .CI(C[355]), .CO(C[356]) );
  FA_9678 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n872), .CI(C[356]), .CO(C[357]) );
  FA_9677 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n873), .CI(C[357]), .CO(C[358]) );
  FA_9676 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n874), .CI(C[358]), .CO(C[359]) );
  FA_9675 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n875), .CI(C[359]), .CO(C[360]) );
  FA_9674 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n876), .CI(C[360]), .CO(C[361]) );
  FA_9673 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n877), .CI(C[361]), .CO(C[362]) );
  FA_9672 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n878), .CI(C[362]), .CO(C[363]) );
  FA_9671 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n879), .CI(C[363]), .CO(C[364]) );
  FA_9670 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n880), .CI(C[364]), .CO(C[365]) );
  FA_9669 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n881), .CI(C[365]), .CO(C[366]) );
  FA_9668 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n882), .CI(C[366]), .CO(C[367]) );
  FA_9667 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n883), .CI(C[367]), .CO(C[368]) );
  FA_9666 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n884), .CI(C[368]), .CO(C[369]) );
  FA_9665 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n885), .CI(C[369]), .CO(C[370]) );
  FA_9664 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n886), .CI(C[370]), .CO(C[371]) );
  FA_9663 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n887), .CI(C[371]), .CO(C[372]) );
  FA_9662 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n888), .CI(C[372]), .CO(C[373]) );
  FA_9661 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n889), .CI(C[373]), .CO(C[374]) );
  FA_9660 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n890), .CI(C[374]), .CO(C[375]) );
  FA_9659 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n891), .CI(C[375]), .CO(C[376]) );
  FA_9658 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n892), .CI(C[376]), .CO(C[377]) );
  FA_9657 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n893), .CI(C[377]), .CO(C[378]) );
  FA_9656 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n894), .CI(C[378]), .CO(C[379]) );
  FA_9655 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n895), .CI(C[379]), .CO(C[380]) );
  FA_9654 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n896), .CI(C[380]), .CO(C[381]) );
  FA_9653 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n897), .CI(C[381]), .CO(C[382]) );
  FA_9652 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n898), .CI(C[382]), .CO(C[383]) );
  FA_9651 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n899), .CI(C[383]), .CO(C[384]) );
  FA_9650 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n900), .CI(C[384]), .CO(C[385]) );
  FA_9649 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n901), .CI(C[385]), .CO(C[386]) );
  FA_9648 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n902), .CI(C[386]), .CO(C[387]) );
  FA_9647 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n903), .CI(C[387]), .CO(C[388]) );
  FA_9646 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n904), .CI(C[388]), .CO(C[389]) );
  FA_9645 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n905), .CI(C[389]), .CO(C[390]) );
  FA_9644 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n906), .CI(C[390]), .CO(C[391]) );
  FA_9643 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n907), .CI(C[391]), .CO(C[392]) );
  FA_9642 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n908), .CI(C[392]), .CO(C[393]) );
  FA_9641 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n909), .CI(C[393]), .CO(C[394]) );
  FA_9640 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n910), .CI(C[394]), .CO(C[395]) );
  FA_9639 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n911), .CI(C[395]), .CO(C[396]) );
  FA_9638 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n912), .CI(C[396]), .CO(C[397]) );
  FA_9637 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n913), .CI(C[397]), .CO(C[398]) );
  FA_9636 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n914), .CI(C[398]), .CO(C[399]) );
  FA_9635 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n915), .CI(C[399]), .CO(C[400]) );
  FA_9634 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n916), .CI(C[400]), .CO(C[401]) );
  FA_9633 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n917), .CI(C[401]), .CO(C[402]) );
  FA_9632 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n918), .CI(C[402]), .CO(C[403]) );
  FA_9631 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n919), .CI(C[403]), .CO(C[404]) );
  FA_9630 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n920), .CI(C[404]), .CO(C[405]) );
  FA_9629 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n921), .CI(C[405]), .CO(C[406]) );
  FA_9628 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n922), .CI(C[406]), .CO(C[407]) );
  FA_9627 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n923), .CI(C[407]), .CO(C[408]) );
  FA_9626 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n924), .CI(C[408]), .CO(C[409]) );
  FA_9625 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n925), .CI(C[409]), .CO(C[410]) );
  FA_9624 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n926), .CI(C[410]), .CO(C[411]) );
  FA_9623 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n927), .CI(C[411]), .CO(C[412]) );
  FA_9622 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n928), .CI(C[412]), .CO(C[413]) );
  FA_9621 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n929), .CI(C[413]), .CO(C[414]) );
  FA_9620 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n930), .CI(C[414]), .CO(C[415]) );
  FA_9619 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n931), .CI(C[415]), .CO(C[416]) );
  FA_9618 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n932), .CI(C[416]), .CO(C[417]) );
  FA_9617 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n933), .CI(C[417]), .CO(C[418]) );
  FA_9616 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n934), .CI(C[418]), .CO(C[419]) );
  FA_9615 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n935), .CI(C[419]), .CO(C[420]) );
  FA_9614 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n936), .CI(C[420]), .CO(C[421]) );
  FA_9613 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n937), .CI(C[421]), .CO(C[422]) );
  FA_9612 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n938), .CI(C[422]), .CO(C[423]) );
  FA_9611 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n939), .CI(C[423]), .CO(C[424]) );
  FA_9610 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n940), .CI(C[424]), .CO(C[425]) );
  FA_9609 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n941), .CI(C[425]), .CO(C[426]) );
  FA_9608 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n942), .CI(C[426]), .CO(C[427]) );
  FA_9607 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n943), .CI(C[427]), .CO(C[428]) );
  FA_9606 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n944), .CI(C[428]), .CO(C[429]) );
  FA_9605 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n945), .CI(C[429]), .CO(C[430]) );
  FA_9604 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n946), .CI(C[430]), .CO(C[431]) );
  FA_9603 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n947), .CI(C[431]), .CO(C[432]) );
  FA_9602 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n948), .CI(C[432]), .CO(C[433]) );
  FA_9601 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n949), .CI(C[433]), .CO(C[434]) );
  FA_9600 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n950), .CI(C[434]), .CO(C[435]) );
  FA_9599 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n951), .CI(C[435]), .CO(C[436]) );
  FA_9598 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n952), .CI(C[436]), .CO(C[437]) );
  FA_9597 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n953), .CI(C[437]), .CO(C[438]) );
  FA_9596 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n954), .CI(C[438]), .CO(C[439]) );
  FA_9595 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n955), .CI(C[439]), .CO(C[440]) );
  FA_9594 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n956), .CI(C[440]), .CO(C[441]) );
  FA_9593 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n957), .CI(C[441]), .CO(C[442]) );
  FA_9592 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n958), .CI(C[442]), .CO(C[443]) );
  FA_9591 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n959), .CI(C[443]), .CO(C[444]) );
  FA_9590 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n960), .CI(C[444]), .CO(C[445]) );
  FA_9589 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n961), .CI(C[445]), .CO(C[446]) );
  FA_9588 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n962), .CI(C[446]), .CO(C[447]) );
  FA_9587 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n963), .CI(C[447]), .CO(C[448]) );
  FA_9586 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n964), .CI(C[448]), .CO(C[449]) );
  FA_9585 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n965), .CI(C[449]), .CO(C[450]) );
  FA_9584 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n966), .CI(C[450]), .CO(C[451]) );
  FA_9583 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n967), .CI(C[451]), .CO(C[452]) );
  FA_9582 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n968), .CI(C[452]), .CO(C[453]) );
  FA_9581 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n969), .CI(C[453]), .CO(C[454]) );
  FA_9580 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n970), .CI(C[454]), .CO(C[455]) );
  FA_9579 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n971), .CI(C[455]), .CO(C[456]) );
  FA_9578 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n972), .CI(C[456]), .CO(C[457]) );
  FA_9577 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n973), .CI(C[457]), .CO(C[458]) );
  FA_9576 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n974), .CI(C[458]), .CO(C[459]) );
  FA_9575 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n975), .CI(C[459]), .CO(C[460]) );
  FA_9574 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n976), .CI(C[460]), .CO(C[461]) );
  FA_9573 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n977), .CI(C[461]), .CO(C[462]) );
  FA_9572 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n978), .CI(C[462]), .CO(C[463]) );
  FA_9571 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n979), .CI(C[463]), .CO(C[464]) );
  FA_9570 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n980), .CI(C[464]), .CO(C[465]) );
  FA_9569 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n981), .CI(C[465]), .CO(C[466]) );
  FA_9568 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n982), .CI(C[466]), .CO(C[467]) );
  FA_9567 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n983), .CI(C[467]), .CO(C[468]) );
  FA_9566 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n984), .CI(C[468]), .CO(C[469]) );
  FA_9565 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n985), .CI(C[469]), .CO(C[470]) );
  FA_9564 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n986), .CI(C[470]), .CO(C[471]) );
  FA_9563 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n987), .CI(C[471]), .CO(C[472]) );
  FA_9562 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n988), .CI(C[472]), .CO(C[473]) );
  FA_9561 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n989), .CI(C[473]), .CO(C[474]) );
  FA_9560 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n990), .CI(C[474]), .CO(C[475]) );
  FA_9559 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n991), .CI(C[475]), .CO(C[476]) );
  FA_9558 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n992), .CI(C[476]), .CO(C[477]) );
  FA_9557 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n993), .CI(C[477]), .CO(C[478]) );
  FA_9556 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n994), .CI(C[478]), .CO(C[479]) );
  FA_9555 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n995), .CI(C[479]), .CO(C[480]) );
  FA_9554 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n996), .CI(C[480]), .CO(C[481]) );
  FA_9553 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n997), .CI(C[481]), .CO(C[482]) );
  FA_9552 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n998), .CI(C[482]), .CO(C[483]) );
  FA_9551 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n999), .CI(C[483]), .CO(C[484]) );
  FA_9550 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n1000), .CI(
        C[484]), .CO(C[485]) );
  FA_9549 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n1001), .CI(
        C[485]), .CO(C[486]) );
  FA_9548 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n1002), .CI(
        C[486]), .CO(C[487]) );
  FA_9547 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1003), .CI(
        C[487]), .CO(C[488]) );
  FA_9546 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1004), .CI(
        C[488]), .CO(C[489]) );
  FA_9545 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1005), .CI(
        C[489]), .CO(C[490]) );
  FA_9544 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1006), .CI(
        C[490]), .CO(C[491]) );
  FA_9543 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1007), .CI(
        C[491]), .CO(C[492]) );
  FA_9542 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1008), .CI(
        C[492]), .CO(C[493]) );
  FA_9541 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1009), .CI(
        C[493]), .CO(C[494]) );
  FA_9540 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1010), .CI(
        C[494]), .CO(C[495]) );
  FA_9539 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1011), .CI(
        C[495]), .CO(C[496]) );
  FA_9538 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1012), .CI(
        C[496]), .CO(C[497]) );
  FA_9537 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1013), .CI(
        C[497]), .CO(C[498]) );
  FA_9536 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1014), .CI(
        C[498]), .CO(C[499]) );
  FA_9535 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1015), .CI(
        C[499]), .CO(C[500]) );
  FA_9534 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1016), .CI(
        C[500]), .CO(C[501]) );
  FA_9533 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1017), .CI(
        C[501]), .CO(C[502]) );
  FA_9532 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1018), .CI(
        C[502]), .CO(C[503]) );
  FA_9531 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1019), .CI(
        C[503]), .CO(C[504]) );
  FA_9530 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1020), .CI(
        C[504]), .CO(C[505]) );
  FA_9529 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1021), .CI(
        C[505]), .CO(C[506]) );
  FA_9528 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1022), .CI(
        C[506]), .CO(C[507]) );
  FA_9527 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1023), .CI(
        C[507]), .CO(C[508]) );
  FA_9526 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1024), .CI(
        C[508]), .CO(C[509]) );
  FA_9525 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1025), .CI(
        C[509]), .CO(C[510]) );
  FA_9524 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1026), .CI(
        C[510]), .CO(C[511]) );
  FA_9523 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1027), .CI(
        C[511]), .CO(C[512]) );
  FA_9522 \FA_INST_1[512].FA_  ( .A(1'b0), .B(n1028), .CI(C[512]), .CO(C[513])
         );
  FA_9521 \FA_INST_1[513].FA_  ( .A(1'b0), .B(n1029), .CI(C[513]), .CO(O) );
  IV U2 ( .A(B[415]), .Z(n931) );
  IV U3 ( .A(B[416]), .Z(n932) );
  IV U4 ( .A(B[417]), .Z(n933) );
  IV U5 ( .A(B[418]), .Z(n934) );
  IV U6 ( .A(B[419]), .Z(n935) );
  IV U7 ( .A(B[420]), .Z(n936) );
  IV U8 ( .A(B[421]), .Z(n937) );
  IV U9 ( .A(B[422]), .Z(n938) );
  IV U10 ( .A(B[423]), .Z(n939) );
  IV U11 ( .A(B[424]), .Z(n940) );
  IV U12 ( .A(B[505]), .Z(n1021) );
  IV U13 ( .A(B[425]), .Z(n941) );
  IV U14 ( .A(B[426]), .Z(n942) );
  IV U15 ( .A(B[427]), .Z(n943) );
  IV U16 ( .A(B[428]), .Z(n944) );
  IV U17 ( .A(B[429]), .Z(n945) );
  IV U18 ( .A(B[430]), .Z(n946) );
  IV U19 ( .A(B[431]), .Z(n947) );
  IV U20 ( .A(B[432]), .Z(n948) );
  IV U21 ( .A(B[433]), .Z(n949) );
  IV U22 ( .A(B[434]), .Z(n950) );
  IV U23 ( .A(B[506]), .Z(n1022) );
  IV U24 ( .A(B[435]), .Z(n951) );
  IV U25 ( .A(B[436]), .Z(n952) );
  IV U26 ( .A(B[437]), .Z(n953) );
  IV U27 ( .A(B[438]), .Z(n954) );
  IV U28 ( .A(B[439]), .Z(n955) );
  IV U29 ( .A(B[440]), .Z(n956) );
  IV U30 ( .A(B[441]), .Z(n957) );
  IV U31 ( .A(B[442]), .Z(n958) );
  IV U32 ( .A(B[443]), .Z(n959) );
  IV U33 ( .A(B[444]), .Z(n960) );
  IV U34 ( .A(B[507]), .Z(n1023) );
  IV U35 ( .A(B[445]), .Z(n961) );
  IV U36 ( .A(B[446]), .Z(n962) );
  IV U37 ( .A(B[447]), .Z(n963) );
  IV U38 ( .A(B[448]), .Z(n964) );
  IV U39 ( .A(B[449]), .Z(n965) );
  IV U40 ( .A(B[450]), .Z(n966) );
  IV U41 ( .A(B[451]), .Z(n967) );
  IV U42 ( .A(B[452]), .Z(n968) );
  IV U43 ( .A(B[453]), .Z(n969) );
  IV U44 ( .A(B[454]), .Z(n970) );
  IV U45 ( .A(B[508]), .Z(n1024) );
  IV U46 ( .A(B[455]), .Z(n971) );
  IV U47 ( .A(B[456]), .Z(n972) );
  IV U48 ( .A(B[457]), .Z(n973) );
  IV U49 ( .A(B[458]), .Z(n974) );
  IV U50 ( .A(B[459]), .Z(n975) );
  IV U51 ( .A(B[460]), .Z(n976) );
  IV U52 ( .A(B[461]), .Z(n977) );
  IV U53 ( .A(B[462]), .Z(n978) );
  IV U54 ( .A(B[0]), .Z(n516) );
  IV U55 ( .A(B[1]), .Z(n517) );
  IV U56 ( .A(B[2]), .Z(n518) );
  IV U57 ( .A(B[3]), .Z(n519) );
  IV U58 ( .A(B[4]), .Z(n520) );
  IV U59 ( .A(B[463]), .Z(n979) );
  IV U60 ( .A(B[5]), .Z(n521) );
  IV U61 ( .A(B[6]), .Z(n522) );
  IV U62 ( .A(B[7]), .Z(n523) );
  IV U63 ( .A(B[8]), .Z(n524) );
  IV U64 ( .A(B[9]), .Z(n525) );
  IV U65 ( .A(B[10]), .Z(n526) );
  IV U66 ( .A(B[11]), .Z(n527) );
  IV U67 ( .A(B[12]), .Z(n528) );
  IV U68 ( .A(B[13]), .Z(n529) );
  IV U69 ( .A(B[14]), .Z(n530) );
  IV U70 ( .A(B[464]), .Z(n980) );
  IV U71 ( .A(B[509]), .Z(n1025) );
  IV U72 ( .A(B[15]), .Z(n531) );
  IV U73 ( .A(B[16]), .Z(n532) );
  IV U74 ( .A(B[17]), .Z(n533) );
  IV U75 ( .A(B[18]), .Z(n534) );
  IV U76 ( .A(B[19]), .Z(n535) );
  IV U77 ( .A(B[20]), .Z(n536) );
  IV U78 ( .A(B[21]), .Z(n537) );
  IV U79 ( .A(B[22]), .Z(n538) );
  IV U80 ( .A(B[23]), .Z(n539) );
  IV U81 ( .A(B[24]), .Z(n540) );
  IV U82 ( .A(B[465]), .Z(n981) );
  IV U83 ( .A(B[25]), .Z(n541) );
  IV U84 ( .A(B[26]), .Z(n542) );
  IV U85 ( .A(B[27]), .Z(n543) );
  IV U86 ( .A(B[28]), .Z(n544) );
  IV U87 ( .A(B[29]), .Z(n545) );
  IV U88 ( .A(B[30]), .Z(n546) );
  IV U89 ( .A(B[31]), .Z(n547) );
  IV U90 ( .A(B[32]), .Z(n548) );
  IV U91 ( .A(B[33]), .Z(n549) );
  IV U92 ( .A(B[34]), .Z(n550) );
  IV U93 ( .A(B[466]), .Z(n982) );
  IV U94 ( .A(B[35]), .Z(n551) );
  IV U95 ( .A(B[36]), .Z(n552) );
  IV U96 ( .A(B[37]), .Z(n553) );
  IV U97 ( .A(B[38]), .Z(n554) );
  IV U98 ( .A(B[39]), .Z(n555) );
  IV U99 ( .A(B[40]), .Z(n556) );
  IV U100 ( .A(B[41]), .Z(n557) );
  IV U101 ( .A(B[42]), .Z(n558) );
  IV U102 ( .A(B[43]), .Z(n559) );
  IV U103 ( .A(B[44]), .Z(n560) );
  IV U104 ( .A(B[467]), .Z(n983) );
  IV U105 ( .A(B[45]), .Z(n561) );
  IV U106 ( .A(B[46]), .Z(n562) );
  IV U107 ( .A(B[47]), .Z(n563) );
  IV U108 ( .A(B[48]), .Z(n564) );
  IV U109 ( .A(B[49]), .Z(n565) );
  IV U110 ( .A(B[50]), .Z(n566) );
  IV U111 ( .A(B[51]), .Z(n567) );
  IV U112 ( .A(B[52]), .Z(n568) );
  IV U113 ( .A(B[53]), .Z(n569) );
  IV U114 ( .A(B[54]), .Z(n570) );
  IV U115 ( .A(B[468]), .Z(n984) );
  IV U116 ( .A(B[55]), .Z(n571) );
  IV U117 ( .A(B[56]), .Z(n572) );
  IV U118 ( .A(B[57]), .Z(n573) );
  IV U119 ( .A(B[58]), .Z(n574) );
  IV U120 ( .A(B[59]), .Z(n575) );
  IV U121 ( .A(B[60]), .Z(n576) );
  IV U122 ( .A(B[61]), .Z(n577) );
  IV U123 ( .A(B[62]), .Z(n578) );
  IV U124 ( .A(B[63]), .Z(n579) );
  IV U125 ( .A(B[64]), .Z(n580) );
  IV U126 ( .A(B[469]), .Z(n985) );
  IV U127 ( .A(B[65]), .Z(n581) );
  IV U128 ( .A(B[66]), .Z(n582) );
  IV U129 ( .A(B[67]), .Z(n583) );
  IV U130 ( .A(B[68]), .Z(n584) );
  IV U131 ( .A(B[69]), .Z(n585) );
  IV U132 ( .A(B[70]), .Z(n586) );
  IV U133 ( .A(B[71]), .Z(n587) );
  IV U134 ( .A(B[72]), .Z(n588) );
  IV U135 ( .A(B[73]), .Z(n589) );
  IV U136 ( .A(B[74]), .Z(n590) );
  IV U137 ( .A(B[470]), .Z(n986) );
  IV U138 ( .A(B[75]), .Z(n591) );
  IV U139 ( .A(B[76]), .Z(n592) );
  IV U140 ( .A(B[77]), .Z(n593) );
  IV U141 ( .A(B[78]), .Z(n594) );
  IV U142 ( .A(B[79]), .Z(n595) );
  IV U143 ( .A(B[80]), .Z(n596) );
  IV U144 ( .A(B[81]), .Z(n597) );
  IV U145 ( .A(B[82]), .Z(n598) );
  IV U146 ( .A(B[83]), .Z(n599) );
  IV U147 ( .A(B[84]), .Z(n600) );
  IV U148 ( .A(B[471]), .Z(n987) );
  IV U149 ( .A(B[85]), .Z(n601) );
  IV U150 ( .A(B[86]), .Z(n602) );
  IV U151 ( .A(B[87]), .Z(n603) );
  IV U152 ( .A(B[88]), .Z(n604) );
  IV U153 ( .A(B[89]), .Z(n605) );
  IV U154 ( .A(B[90]), .Z(n606) );
  IV U155 ( .A(B[91]), .Z(n607) );
  IV U156 ( .A(B[92]), .Z(n608) );
  IV U157 ( .A(B[93]), .Z(n609) );
  IV U158 ( .A(B[94]), .Z(n610) );
  IV U159 ( .A(B[472]), .Z(n988) );
  IV U160 ( .A(B[95]), .Z(n611) );
  IV U161 ( .A(B[96]), .Z(n612) );
  IV U162 ( .A(B[97]), .Z(n613) );
  IV U163 ( .A(B[98]), .Z(n614) );
  IV U164 ( .A(B[99]), .Z(n615) );
  IV U165 ( .A(B[100]), .Z(n616) );
  IV U166 ( .A(B[101]), .Z(n617) );
  IV U167 ( .A(B[102]), .Z(n618) );
  IV U168 ( .A(B[103]), .Z(n619) );
  IV U169 ( .A(B[104]), .Z(n620) );
  IV U170 ( .A(B[473]), .Z(n989) );
  IV U171 ( .A(B[105]), .Z(n621) );
  IV U172 ( .A(B[106]), .Z(n622) );
  IV U173 ( .A(B[107]), .Z(n623) );
  IV U174 ( .A(B[108]), .Z(n624) );
  IV U175 ( .A(B[109]), .Z(n625) );
  IV U176 ( .A(B[110]), .Z(n626) );
  IV U177 ( .A(B[111]), .Z(n627) );
  IV U178 ( .A(B[112]), .Z(n628) );
  IV U179 ( .A(B[113]), .Z(n629) );
  IV U180 ( .A(B[114]), .Z(n630) );
  IV U181 ( .A(B[474]), .Z(n990) );
  IV U182 ( .A(B[510]), .Z(n1026) );
  IV U183 ( .A(B[115]), .Z(n631) );
  IV U184 ( .A(B[116]), .Z(n632) );
  IV U185 ( .A(B[117]), .Z(n633) );
  IV U186 ( .A(B[118]), .Z(n634) );
  IV U187 ( .A(B[119]), .Z(n635) );
  IV U188 ( .A(B[120]), .Z(n636) );
  IV U189 ( .A(B[121]), .Z(n637) );
  IV U190 ( .A(B[122]), .Z(n638) );
  IV U191 ( .A(B[123]), .Z(n639) );
  IV U192 ( .A(B[124]), .Z(n640) );
  IV U193 ( .A(B[475]), .Z(n991) );
  IV U194 ( .A(B[125]), .Z(n641) );
  IV U195 ( .A(B[126]), .Z(n642) );
  IV U196 ( .A(B[127]), .Z(n643) );
  IV U197 ( .A(B[128]), .Z(n644) );
  IV U198 ( .A(B[129]), .Z(n645) );
  IV U199 ( .A(B[130]), .Z(n646) );
  IV U200 ( .A(B[131]), .Z(n647) );
  IV U201 ( .A(B[132]), .Z(n648) );
  IV U202 ( .A(B[133]), .Z(n649) );
  IV U203 ( .A(B[134]), .Z(n650) );
  IV U204 ( .A(B[476]), .Z(n992) );
  IV U205 ( .A(B[135]), .Z(n651) );
  IV U206 ( .A(B[136]), .Z(n652) );
  IV U207 ( .A(B[137]), .Z(n653) );
  IV U208 ( .A(B[138]), .Z(n654) );
  IV U209 ( .A(B[139]), .Z(n655) );
  IV U210 ( .A(B[140]), .Z(n656) );
  IV U211 ( .A(B[141]), .Z(n657) );
  IV U212 ( .A(B[142]), .Z(n658) );
  IV U213 ( .A(B[143]), .Z(n659) );
  IV U214 ( .A(B[144]), .Z(n660) );
  IV U215 ( .A(B[477]), .Z(n993) );
  IV U216 ( .A(B[145]), .Z(n661) );
  IV U217 ( .A(B[146]), .Z(n662) );
  IV U218 ( .A(B[147]), .Z(n663) );
  IV U219 ( .A(B[148]), .Z(n664) );
  IV U220 ( .A(B[149]), .Z(n665) );
  IV U221 ( .A(B[150]), .Z(n666) );
  IV U222 ( .A(B[151]), .Z(n667) );
  IV U223 ( .A(B[152]), .Z(n668) );
  IV U224 ( .A(B[153]), .Z(n669) );
  IV U225 ( .A(B[154]), .Z(n670) );
  IV U226 ( .A(B[478]), .Z(n994) );
  IV U227 ( .A(B[155]), .Z(n671) );
  IV U228 ( .A(B[156]), .Z(n672) );
  IV U229 ( .A(B[157]), .Z(n673) );
  IV U230 ( .A(B[158]), .Z(n674) );
  IV U231 ( .A(B[159]), .Z(n675) );
  IV U232 ( .A(B[160]), .Z(n676) );
  IV U233 ( .A(B[161]), .Z(n677) );
  IV U234 ( .A(B[162]), .Z(n678) );
  IV U235 ( .A(B[163]), .Z(n679) );
  IV U236 ( .A(B[164]), .Z(n680) );
  IV U237 ( .A(B[479]), .Z(n995) );
  IV U238 ( .A(B[165]), .Z(n681) );
  IV U239 ( .A(B[166]), .Z(n682) );
  IV U240 ( .A(B[167]), .Z(n683) );
  IV U241 ( .A(B[168]), .Z(n684) );
  IV U242 ( .A(B[169]), .Z(n685) );
  IV U243 ( .A(B[170]), .Z(n686) );
  IV U244 ( .A(B[171]), .Z(n687) );
  IV U245 ( .A(B[172]), .Z(n688) );
  IV U246 ( .A(B[173]), .Z(n689) );
  IV U247 ( .A(B[174]), .Z(n690) );
  IV U248 ( .A(B[480]), .Z(n996) );
  IV U249 ( .A(B[175]), .Z(n691) );
  IV U250 ( .A(B[176]), .Z(n692) );
  IV U251 ( .A(B[177]), .Z(n693) );
  IV U252 ( .A(B[178]), .Z(n694) );
  IV U253 ( .A(B[179]), .Z(n695) );
  IV U254 ( .A(B[180]), .Z(n696) );
  IV U255 ( .A(B[181]), .Z(n697) );
  IV U256 ( .A(B[182]), .Z(n698) );
  IV U257 ( .A(B[183]), .Z(n699) );
  IV U258 ( .A(B[184]), .Z(n700) );
  IV U259 ( .A(B[481]), .Z(n997) );
  IV U260 ( .A(B[185]), .Z(n701) );
  IV U261 ( .A(B[186]), .Z(n702) );
  IV U262 ( .A(B[187]), .Z(n703) );
  IV U263 ( .A(B[188]), .Z(n704) );
  IV U264 ( .A(B[189]), .Z(n705) );
  IV U265 ( .A(B[190]), .Z(n706) );
  IV U266 ( .A(B[191]), .Z(n707) );
  IV U267 ( .A(B[192]), .Z(n708) );
  IV U268 ( .A(B[193]), .Z(n709) );
  IV U269 ( .A(B[194]), .Z(n710) );
  IV U270 ( .A(B[482]), .Z(n998) );
  IV U271 ( .A(B[195]), .Z(n711) );
  IV U272 ( .A(B[196]), .Z(n712) );
  IV U273 ( .A(B[197]), .Z(n713) );
  IV U274 ( .A(B[198]), .Z(n714) );
  IV U275 ( .A(B[199]), .Z(n715) );
  IV U276 ( .A(B[200]), .Z(n716) );
  IV U277 ( .A(B[201]), .Z(n717) );
  IV U278 ( .A(B[202]), .Z(n718) );
  IV U279 ( .A(B[203]), .Z(n719) );
  IV U280 ( .A(B[204]), .Z(n720) );
  IV U281 ( .A(B[483]), .Z(n999) );
  IV U282 ( .A(B[205]), .Z(n721) );
  IV U283 ( .A(B[206]), .Z(n722) );
  IV U284 ( .A(B[207]), .Z(n723) );
  IV U285 ( .A(B[208]), .Z(n724) );
  IV U286 ( .A(B[209]), .Z(n725) );
  IV U287 ( .A(B[210]), .Z(n726) );
  IV U288 ( .A(B[211]), .Z(n727) );
  IV U289 ( .A(B[212]), .Z(n728) );
  IV U290 ( .A(B[213]), .Z(n729) );
  IV U291 ( .A(B[214]), .Z(n730) );
  IV U292 ( .A(B[484]), .Z(n1000) );
  IV U293 ( .A(B[511]), .Z(n1027) );
  IV U294 ( .A(B[215]), .Z(n731) );
  IV U295 ( .A(B[216]), .Z(n732) );
  IV U296 ( .A(B[217]), .Z(n733) );
  IV U297 ( .A(B[218]), .Z(n734) );
  IV U298 ( .A(B[219]), .Z(n735) );
  IV U299 ( .A(B[220]), .Z(n736) );
  IV U300 ( .A(B[221]), .Z(n737) );
  IV U301 ( .A(B[222]), .Z(n738) );
  IV U302 ( .A(B[223]), .Z(n739) );
  IV U303 ( .A(B[224]), .Z(n740) );
  IV U304 ( .A(B[485]), .Z(n1001) );
  IV U305 ( .A(B[225]), .Z(n741) );
  IV U306 ( .A(B[226]), .Z(n742) );
  IV U307 ( .A(B[227]), .Z(n743) );
  IV U308 ( .A(B[228]), .Z(n744) );
  IV U309 ( .A(B[229]), .Z(n745) );
  IV U310 ( .A(B[230]), .Z(n746) );
  IV U311 ( .A(B[231]), .Z(n747) );
  IV U312 ( .A(B[232]), .Z(n748) );
  IV U313 ( .A(B[233]), .Z(n749) );
  IV U314 ( .A(B[234]), .Z(n750) );
  IV U315 ( .A(B[486]), .Z(n1002) );
  IV U316 ( .A(B[235]), .Z(n751) );
  IV U317 ( .A(B[236]), .Z(n752) );
  IV U318 ( .A(B[237]), .Z(n753) );
  IV U319 ( .A(B[238]), .Z(n754) );
  IV U320 ( .A(B[239]), .Z(n755) );
  IV U321 ( .A(B[240]), .Z(n756) );
  IV U322 ( .A(B[241]), .Z(n757) );
  IV U323 ( .A(B[242]), .Z(n758) );
  IV U324 ( .A(B[243]), .Z(n759) );
  IV U325 ( .A(B[244]), .Z(n760) );
  IV U326 ( .A(B[487]), .Z(n1003) );
  IV U327 ( .A(B[245]), .Z(n761) );
  IV U328 ( .A(B[246]), .Z(n762) );
  IV U329 ( .A(B[247]), .Z(n763) );
  IV U330 ( .A(B[248]), .Z(n764) );
  IV U331 ( .A(B[249]), .Z(n765) );
  IV U332 ( .A(B[250]), .Z(n766) );
  IV U333 ( .A(B[251]), .Z(n767) );
  IV U334 ( .A(B[252]), .Z(n768) );
  IV U335 ( .A(B[253]), .Z(n769) );
  IV U336 ( .A(B[254]), .Z(n770) );
  IV U337 ( .A(B[488]), .Z(n1004) );
  IV U338 ( .A(B[255]), .Z(n771) );
  IV U339 ( .A(B[256]), .Z(n772) );
  IV U340 ( .A(B[257]), .Z(n773) );
  IV U341 ( .A(B[258]), .Z(n774) );
  IV U342 ( .A(B[259]), .Z(n775) );
  IV U343 ( .A(B[260]), .Z(n776) );
  IV U344 ( .A(B[261]), .Z(n777) );
  IV U345 ( .A(B[262]), .Z(n778) );
  IV U346 ( .A(B[263]), .Z(n779) );
  IV U347 ( .A(B[264]), .Z(n780) );
  IV U348 ( .A(B[489]), .Z(n1005) );
  IV U349 ( .A(B[265]), .Z(n781) );
  IV U350 ( .A(B[266]), .Z(n782) );
  IV U351 ( .A(B[267]), .Z(n783) );
  IV U352 ( .A(B[268]), .Z(n784) );
  IV U353 ( .A(B[269]), .Z(n785) );
  IV U354 ( .A(B[270]), .Z(n786) );
  IV U355 ( .A(B[271]), .Z(n787) );
  IV U356 ( .A(B[272]), .Z(n788) );
  IV U357 ( .A(B[273]), .Z(n789) );
  IV U358 ( .A(B[274]), .Z(n790) );
  IV U359 ( .A(B[490]), .Z(n1006) );
  IV U360 ( .A(B[275]), .Z(n791) );
  IV U361 ( .A(B[276]), .Z(n792) );
  IV U362 ( .A(B[277]), .Z(n793) );
  IV U363 ( .A(B[278]), .Z(n794) );
  IV U364 ( .A(B[279]), .Z(n795) );
  IV U365 ( .A(B[280]), .Z(n796) );
  IV U366 ( .A(B[281]), .Z(n797) );
  IV U367 ( .A(B[282]), .Z(n798) );
  IV U368 ( .A(B[283]), .Z(n799) );
  IV U369 ( .A(B[284]), .Z(n800) );
  IV U370 ( .A(B[491]), .Z(n1007) );
  IV U371 ( .A(B[285]), .Z(n801) );
  IV U372 ( .A(B[286]), .Z(n802) );
  IV U373 ( .A(B[287]), .Z(n803) );
  IV U374 ( .A(B[288]), .Z(n804) );
  IV U375 ( .A(B[289]), .Z(n805) );
  IV U376 ( .A(B[290]), .Z(n806) );
  IV U377 ( .A(B[291]), .Z(n807) );
  IV U378 ( .A(B[292]), .Z(n808) );
  IV U379 ( .A(B[293]), .Z(n809) );
  IV U380 ( .A(B[294]), .Z(n810) );
  IV U381 ( .A(B[492]), .Z(n1008) );
  IV U382 ( .A(B[295]), .Z(n811) );
  IV U383 ( .A(B[296]), .Z(n812) );
  IV U384 ( .A(B[297]), .Z(n813) );
  IV U385 ( .A(B[298]), .Z(n814) );
  IV U386 ( .A(B[299]), .Z(n815) );
  IV U387 ( .A(B[300]), .Z(n816) );
  IV U388 ( .A(B[301]), .Z(n817) );
  IV U389 ( .A(B[302]), .Z(n818) );
  IV U390 ( .A(B[303]), .Z(n819) );
  IV U391 ( .A(B[304]), .Z(n820) );
  IV U392 ( .A(B[493]), .Z(n1009) );
  IV U393 ( .A(B[305]), .Z(n821) );
  IV U394 ( .A(B[306]), .Z(n822) );
  IV U395 ( .A(B[307]), .Z(n823) );
  IV U396 ( .A(B[308]), .Z(n824) );
  IV U397 ( .A(B[309]), .Z(n825) );
  IV U398 ( .A(B[310]), .Z(n826) );
  IV U399 ( .A(B[311]), .Z(n827) );
  IV U400 ( .A(B[312]), .Z(n828) );
  IV U401 ( .A(B[313]), .Z(n829) );
  IV U402 ( .A(B[314]), .Z(n830) );
  IV U403 ( .A(B[494]), .Z(n1010) );
  IV U404 ( .A(B[512]), .Z(n1028) );
  IV U405 ( .A(B[315]), .Z(n831) );
  IV U406 ( .A(B[316]), .Z(n832) );
  IV U407 ( .A(B[317]), .Z(n833) );
  IV U408 ( .A(B[318]), .Z(n834) );
  IV U409 ( .A(B[319]), .Z(n835) );
  IV U410 ( .A(B[320]), .Z(n836) );
  IV U411 ( .A(B[321]), .Z(n837) );
  IV U412 ( .A(B[322]), .Z(n838) );
  IV U413 ( .A(B[323]), .Z(n839) );
  IV U414 ( .A(B[324]), .Z(n840) );
  IV U415 ( .A(B[495]), .Z(n1011) );
  IV U416 ( .A(B[325]), .Z(n841) );
  IV U417 ( .A(B[326]), .Z(n842) );
  IV U418 ( .A(B[327]), .Z(n843) );
  IV U419 ( .A(B[328]), .Z(n844) );
  IV U420 ( .A(B[329]), .Z(n845) );
  IV U421 ( .A(B[330]), .Z(n846) );
  IV U422 ( .A(B[331]), .Z(n847) );
  IV U423 ( .A(B[332]), .Z(n848) );
  IV U424 ( .A(B[333]), .Z(n849) );
  IV U425 ( .A(B[334]), .Z(n850) );
  IV U426 ( .A(B[496]), .Z(n1012) );
  IV U427 ( .A(B[335]), .Z(n851) );
  IV U428 ( .A(B[336]), .Z(n852) );
  IV U429 ( .A(B[337]), .Z(n853) );
  IV U430 ( .A(B[338]), .Z(n854) );
  IV U431 ( .A(B[339]), .Z(n855) );
  IV U432 ( .A(B[340]), .Z(n856) );
  IV U433 ( .A(B[341]), .Z(n857) );
  IV U434 ( .A(B[342]), .Z(n858) );
  IV U435 ( .A(B[343]), .Z(n859) );
  IV U436 ( .A(B[344]), .Z(n860) );
  IV U437 ( .A(B[497]), .Z(n1013) );
  IV U438 ( .A(B[345]), .Z(n861) );
  IV U439 ( .A(B[346]), .Z(n862) );
  IV U440 ( .A(B[347]), .Z(n863) );
  IV U441 ( .A(B[348]), .Z(n864) );
  IV U442 ( .A(B[349]), .Z(n865) );
  IV U443 ( .A(B[350]), .Z(n866) );
  IV U444 ( .A(B[351]), .Z(n867) );
  IV U445 ( .A(B[352]), .Z(n868) );
  IV U446 ( .A(B[353]), .Z(n869) );
  IV U447 ( .A(B[354]), .Z(n870) );
  IV U448 ( .A(B[498]), .Z(n1014) );
  IV U449 ( .A(B[355]), .Z(n871) );
  IV U450 ( .A(B[356]), .Z(n872) );
  IV U451 ( .A(B[357]), .Z(n873) );
  IV U452 ( .A(B[358]), .Z(n874) );
  IV U453 ( .A(B[359]), .Z(n875) );
  IV U454 ( .A(B[360]), .Z(n876) );
  IV U455 ( .A(B[361]), .Z(n877) );
  IV U456 ( .A(B[362]), .Z(n878) );
  IV U457 ( .A(B[363]), .Z(n879) );
  IV U458 ( .A(B[364]), .Z(n880) );
  IV U459 ( .A(B[499]), .Z(n1015) );
  IV U460 ( .A(B[365]), .Z(n881) );
  IV U461 ( .A(B[366]), .Z(n882) );
  IV U462 ( .A(B[367]), .Z(n883) );
  IV U463 ( .A(B[368]), .Z(n884) );
  IV U464 ( .A(B[369]), .Z(n885) );
  IV U465 ( .A(B[370]), .Z(n886) );
  IV U466 ( .A(B[371]), .Z(n887) );
  IV U467 ( .A(B[372]), .Z(n888) );
  IV U468 ( .A(B[373]), .Z(n889) );
  IV U469 ( .A(B[374]), .Z(n890) );
  IV U470 ( .A(B[500]), .Z(n1016) );
  IV U471 ( .A(B[375]), .Z(n891) );
  IV U472 ( .A(B[376]), .Z(n892) );
  IV U473 ( .A(B[377]), .Z(n893) );
  IV U474 ( .A(B[378]), .Z(n894) );
  IV U475 ( .A(B[379]), .Z(n895) );
  IV U476 ( .A(B[380]), .Z(n896) );
  IV U477 ( .A(B[381]), .Z(n897) );
  IV U478 ( .A(B[382]), .Z(n898) );
  IV U479 ( .A(B[383]), .Z(n899) );
  IV U480 ( .A(B[384]), .Z(n900) );
  IV U481 ( .A(B[501]), .Z(n1017) );
  IV U482 ( .A(B[385]), .Z(n901) );
  IV U483 ( .A(B[386]), .Z(n902) );
  IV U484 ( .A(B[387]), .Z(n903) );
  IV U485 ( .A(B[388]), .Z(n904) );
  IV U486 ( .A(B[389]), .Z(n905) );
  IV U487 ( .A(B[390]), .Z(n906) );
  IV U488 ( .A(B[391]), .Z(n907) );
  IV U489 ( .A(B[392]), .Z(n908) );
  IV U490 ( .A(B[393]), .Z(n909) );
  IV U491 ( .A(B[394]), .Z(n910) );
  IV U492 ( .A(B[502]), .Z(n1018) );
  IV U493 ( .A(B[395]), .Z(n911) );
  IV U494 ( .A(B[396]), .Z(n912) );
  IV U495 ( .A(B[397]), .Z(n913) );
  IV U496 ( .A(B[398]), .Z(n914) );
  IV U497 ( .A(B[399]), .Z(n915) );
  IV U498 ( .A(B[400]), .Z(n916) );
  IV U499 ( .A(B[401]), .Z(n917) );
  IV U500 ( .A(B[402]), .Z(n918) );
  IV U501 ( .A(B[403]), .Z(n919) );
  IV U502 ( .A(B[404]), .Z(n920) );
  IV U503 ( .A(B[503]), .Z(n1019) );
  IV U504 ( .A(B[405]), .Z(n921) );
  IV U505 ( .A(B[406]), .Z(n922) );
  IV U506 ( .A(B[407]), .Z(n923) );
  IV U507 ( .A(B[408]), .Z(n924) );
  IV U508 ( .A(B[409]), .Z(n925) );
  IV U509 ( .A(B[410]), .Z(n926) );
  IV U510 ( .A(B[411]), .Z(n927) );
  IV U511 ( .A(B[412]), .Z(n928) );
  IV U512 ( .A(B[413]), .Z(n929) );
  IV U513 ( .A(B[414]), .Z(n930) );
  IV U514 ( .A(B[504]), .Z(n1020) );
  IV U515 ( .A(B[513]), .Z(n1029) );
endmodule


module FA_9008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_9009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N514_5 ( A, B, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  output CO;
  wire   n2, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  wire   [513:1] C;

  FA_9520 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(
        S[0]), .CO(C[1]) );
  FA_9519 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n514), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_9518 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n515), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_9517 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n516), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_9516 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n517), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_9515 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n518), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_9514 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n519), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_9513 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n520), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_9512 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n521), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_9511 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n522), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_9510 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n523), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_9509 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n524), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_9508 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n525), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_9507 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n526), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_9506 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n527), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_9505 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n528), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_9504 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n529), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_9503 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n530), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_9502 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n531), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_9501 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n532), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_9500 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n533), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_9499 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n534), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_9498 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n535), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_9497 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n536), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_9496 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n537), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_9495 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n538), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_9494 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n539), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_9493 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n540), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_9492 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n541), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_9491 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n542), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_9490 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n543), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_9489 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n544), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_9488 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n545), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_9487 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n546), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_9486 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n547), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_9485 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n548), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_9484 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n549), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_9483 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n550), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_9482 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n551), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_9481 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n552), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_9480 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n553), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_9479 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n554), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_9478 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n555), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_9477 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n556), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_9476 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n557), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_9475 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n558), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_9474 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n559), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_9473 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n560), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_9472 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n561), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_9471 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n562), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_9470 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n563), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_9469 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n564), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_9468 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n565), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_9467 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n566), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_9466 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n567), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_9465 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n568), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_9464 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n569), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_9463 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n570), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_9462 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n571), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_9461 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n572), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_9460 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n573), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_9459 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n574), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_9458 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n575), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_9457 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n576), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_9456 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n577), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_9455 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n578), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_9454 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n579), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_9453 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n580), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_9452 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n581), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_9451 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n582), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_9450 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n583), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_9449 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n584), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_9448 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n585), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_9447 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n586), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_9446 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n587), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_9445 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n588), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_9444 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n589), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_9443 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n590), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_9442 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n591), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_9441 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n592), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_9440 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n593), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_9439 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n594), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_9438 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n595), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_9437 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n596), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_9436 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n597), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_9435 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n598), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_9434 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n599), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_9433 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n600), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_9432 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n601), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_9431 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n602), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_9430 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n603), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_9429 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n604), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_9428 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n605), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_9427 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n606), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_9426 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n607), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_9425 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n608), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_9424 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n609), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_9423 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n610), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_9422 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n611), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_9421 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n612), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_9420 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n613), .CI(C[100]), .S(S[100]), .CO(C[101]) );
  FA_9419 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n614), .CI(C[101]), .S(S[101]), .CO(C[102]) );
  FA_9418 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n615), .CI(C[102]), .S(S[102]), .CO(C[103]) );
  FA_9417 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n616), .CI(C[103]), .S(S[103]), .CO(C[104]) );
  FA_9416 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n617), .CI(C[104]), .S(S[104]), .CO(C[105]) );
  FA_9415 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n618), .CI(C[105]), .S(S[105]), .CO(C[106]) );
  FA_9414 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n619), .CI(C[106]), .S(S[106]), .CO(C[107]) );
  FA_9413 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n620), .CI(C[107]), .S(S[107]), .CO(C[108]) );
  FA_9412 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n621), .CI(C[108]), .S(S[108]), .CO(C[109]) );
  FA_9411 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n622), .CI(C[109]), .S(S[109]), .CO(C[110]) );
  FA_9410 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n623), .CI(C[110]), .S(S[110]), .CO(C[111]) );
  FA_9409 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n624), .CI(C[111]), .S(S[111]), .CO(C[112]) );
  FA_9408 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n625), .CI(C[112]), .S(S[112]), .CO(C[113]) );
  FA_9407 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n626), .CI(C[113]), .S(S[113]), .CO(C[114]) );
  FA_9406 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n627), .CI(C[114]), .S(S[114]), .CO(C[115]) );
  FA_9405 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n628), .CI(C[115]), .S(S[115]), .CO(C[116]) );
  FA_9404 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n629), .CI(C[116]), .S(S[116]), .CO(C[117]) );
  FA_9403 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n630), .CI(C[117]), .S(S[117]), .CO(C[118]) );
  FA_9402 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n631), .CI(C[118]), .S(S[118]), .CO(C[119]) );
  FA_9401 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n632), .CI(C[119]), .S(S[119]), .CO(C[120]) );
  FA_9400 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n633), .CI(C[120]), .S(S[120]), .CO(C[121]) );
  FA_9399 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n634), .CI(C[121]), .S(S[121]), .CO(C[122]) );
  FA_9398 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n635), .CI(C[122]), .S(S[122]), .CO(C[123]) );
  FA_9397 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n636), .CI(C[123]), .S(S[123]), .CO(C[124]) );
  FA_9396 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n637), .CI(C[124]), .S(S[124]), .CO(C[125]) );
  FA_9395 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n638), .CI(C[125]), .S(S[125]), .CO(C[126]) );
  FA_9394 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n639), .CI(C[126]), .S(S[126]), .CO(C[127]) );
  FA_9393 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n640), .CI(C[127]), .S(S[127]), .CO(C[128]) );
  FA_9392 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n641), .CI(C[128]), .S(S[128]), .CO(C[129]) );
  FA_9391 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n642), .CI(C[129]), .S(S[129]), .CO(C[130]) );
  FA_9390 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n643), .CI(C[130]), .S(S[130]), .CO(C[131]) );
  FA_9389 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n644), .CI(C[131]), .S(S[131]), .CO(C[132]) );
  FA_9388 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n645), .CI(C[132]), .S(S[132]), .CO(C[133]) );
  FA_9387 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n646), .CI(C[133]), .S(S[133]), .CO(C[134]) );
  FA_9386 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n647), .CI(C[134]), .S(S[134]), .CO(C[135]) );
  FA_9385 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n648), .CI(C[135]), .S(S[135]), .CO(C[136]) );
  FA_9384 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n649), .CI(C[136]), .S(S[136]), .CO(C[137]) );
  FA_9383 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n650), .CI(C[137]), .S(S[137]), .CO(C[138]) );
  FA_9382 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n651), .CI(C[138]), .S(S[138]), .CO(C[139]) );
  FA_9381 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n652), .CI(C[139]), .S(S[139]), .CO(C[140]) );
  FA_9380 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n653), .CI(C[140]), .S(S[140]), .CO(C[141]) );
  FA_9379 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n654), .CI(C[141]), .S(S[141]), .CO(C[142]) );
  FA_9378 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n655), .CI(C[142]), .S(S[142]), .CO(C[143]) );
  FA_9377 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n656), .CI(C[143]), .S(S[143]), .CO(C[144]) );
  FA_9376 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n657), .CI(C[144]), .S(S[144]), .CO(C[145]) );
  FA_9375 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n658), .CI(C[145]), .S(S[145]), .CO(C[146]) );
  FA_9374 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n659), .CI(C[146]), .S(S[146]), .CO(C[147]) );
  FA_9373 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n660), .CI(C[147]), .S(S[147]), .CO(C[148]) );
  FA_9372 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n661), .CI(C[148]), .S(S[148]), .CO(C[149]) );
  FA_9371 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n662), .CI(C[149]), .S(S[149]), .CO(C[150]) );
  FA_9370 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n663), .CI(C[150]), .S(S[150]), .CO(C[151]) );
  FA_9369 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n664), .CI(C[151]), .S(S[151]), .CO(C[152]) );
  FA_9368 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n665), .CI(C[152]), .S(S[152]), .CO(C[153]) );
  FA_9367 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n666), .CI(C[153]), .S(S[153]), .CO(C[154]) );
  FA_9366 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n667), .CI(C[154]), .S(S[154]), .CO(C[155]) );
  FA_9365 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n668), .CI(C[155]), .S(S[155]), .CO(C[156]) );
  FA_9364 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n669), .CI(C[156]), .S(S[156]), .CO(C[157]) );
  FA_9363 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n670), .CI(C[157]), .S(S[157]), .CO(C[158]) );
  FA_9362 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n671), .CI(C[158]), .S(S[158]), .CO(C[159]) );
  FA_9361 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n672), .CI(C[159]), .S(S[159]), .CO(C[160]) );
  FA_9360 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n673), .CI(C[160]), .S(S[160]), .CO(C[161]) );
  FA_9359 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n674), .CI(C[161]), .S(S[161]), .CO(C[162]) );
  FA_9358 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n675), .CI(C[162]), .S(S[162]), .CO(C[163]) );
  FA_9357 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n676), .CI(C[163]), .S(S[163]), .CO(C[164]) );
  FA_9356 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n677), .CI(C[164]), .S(S[164]), .CO(C[165]) );
  FA_9355 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n678), .CI(C[165]), .S(S[165]), .CO(C[166]) );
  FA_9354 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n679), .CI(C[166]), .S(S[166]), .CO(C[167]) );
  FA_9353 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n680), .CI(C[167]), .S(S[167]), .CO(C[168]) );
  FA_9352 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n681), .CI(C[168]), .S(S[168]), .CO(C[169]) );
  FA_9351 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n682), .CI(C[169]), .S(S[169]), .CO(C[170]) );
  FA_9350 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n683), .CI(C[170]), .S(S[170]), .CO(C[171]) );
  FA_9349 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n684), .CI(C[171]), .S(S[171]), .CO(C[172]) );
  FA_9348 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n685), .CI(C[172]), .S(S[172]), .CO(C[173]) );
  FA_9347 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n686), .CI(C[173]), .S(S[173]), .CO(C[174]) );
  FA_9346 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n687), .CI(C[174]), .S(S[174]), .CO(C[175]) );
  FA_9345 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n688), .CI(C[175]), .S(S[175]), .CO(C[176]) );
  FA_9344 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n689), .CI(C[176]), .S(S[176]), .CO(C[177]) );
  FA_9343 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n690), .CI(C[177]), .S(S[177]), .CO(C[178]) );
  FA_9342 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n691), .CI(C[178]), .S(S[178]), .CO(C[179]) );
  FA_9341 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n692), .CI(C[179]), .S(S[179]), .CO(C[180]) );
  FA_9340 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n693), .CI(C[180]), .S(S[180]), .CO(C[181]) );
  FA_9339 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n694), .CI(C[181]), .S(S[181]), .CO(C[182]) );
  FA_9338 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n695), .CI(C[182]), .S(S[182]), .CO(C[183]) );
  FA_9337 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n696), .CI(C[183]), .S(S[183]), .CO(C[184]) );
  FA_9336 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n697), .CI(C[184]), .S(S[184]), .CO(C[185]) );
  FA_9335 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n698), .CI(C[185]), .S(S[185]), .CO(C[186]) );
  FA_9334 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n699), .CI(C[186]), .S(S[186]), .CO(C[187]) );
  FA_9333 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n700), .CI(C[187]), .S(S[187]), .CO(C[188]) );
  FA_9332 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n701), .CI(C[188]), .S(S[188]), .CO(C[189]) );
  FA_9331 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n702), .CI(C[189]), .S(S[189]), .CO(C[190]) );
  FA_9330 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n703), .CI(C[190]), .S(S[190]), .CO(C[191]) );
  FA_9329 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n704), .CI(C[191]), .S(S[191]), .CO(C[192]) );
  FA_9328 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n705), .CI(C[192]), .S(S[192]), .CO(C[193]) );
  FA_9327 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n706), .CI(C[193]), .S(S[193]), .CO(C[194]) );
  FA_9326 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n707), .CI(C[194]), .S(S[194]), .CO(C[195]) );
  FA_9325 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n708), .CI(C[195]), .S(S[195]), .CO(C[196]) );
  FA_9324 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n709), .CI(C[196]), .S(S[196]), .CO(C[197]) );
  FA_9323 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n710), .CI(C[197]), .S(S[197]), .CO(C[198]) );
  FA_9322 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n711), .CI(C[198]), .S(S[198]), .CO(C[199]) );
  FA_9321 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n712), .CI(C[199]), .S(S[199]), .CO(C[200]) );
  FA_9320 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n713), .CI(C[200]), .S(S[200]), .CO(C[201]) );
  FA_9319 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n714), .CI(C[201]), .S(S[201]), .CO(C[202]) );
  FA_9318 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n715), .CI(C[202]), .S(S[202]), .CO(C[203]) );
  FA_9317 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n716), .CI(C[203]), .S(S[203]), .CO(C[204]) );
  FA_9316 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n717), .CI(C[204]), .S(S[204]), .CO(C[205]) );
  FA_9315 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n718), .CI(C[205]), .S(S[205]), .CO(C[206]) );
  FA_9314 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n719), .CI(C[206]), .S(S[206]), .CO(C[207]) );
  FA_9313 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n720), .CI(C[207]), .S(S[207]), .CO(C[208]) );
  FA_9312 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n721), .CI(C[208]), .S(S[208]), .CO(C[209]) );
  FA_9311 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n722), .CI(C[209]), .S(S[209]), .CO(C[210]) );
  FA_9310 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n723), .CI(C[210]), .S(S[210]), .CO(C[211]) );
  FA_9309 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n724), .CI(C[211]), .S(S[211]), .CO(C[212]) );
  FA_9308 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n725), .CI(C[212]), .S(S[212]), .CO(C[213]) );
  FA_9307 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n726), .CI(C[213]), .S(S[213]), .CO(C[214]) );
  FA_9306 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n727), .CI(C[214]), .S(S[214]), .CO(C[215]) );
  FA_9305 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n728), .CI(C[215]), .S(S[215]), .CO(C[216]) );
  FA_9304 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n729), .CI(C[216]), .S(S[216]), .CO(C[217]) );
  FA_9303 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n730), .CI(C[217]), .S(S[217]), .CO(C[218]) );
  FA_9302 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n731), .CI(C[218]), .S(S[218]), .CO(C[219]) );
  FA_9301 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n732), .CI(C[219]), .S(S[219]), .CO(C[220]) );
  FA_9300 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n733), .CI(C[220]), .S(S[220]), .CO(C[221]) );
  FA_9299 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n734), .CI(C[221]), .S(S[221]), .CO(C[222]) );
  FA_9298 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n735), .CI(C[222]), .S(S[222]), .CO(C[223]) );
  FA_9297 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n736), .CI(C[223]), .S(S[223]), .CO(C[224]) );
  FA_9296 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n737), .CI(C[224]), .S(S[224]), .CO(C[225]) );
  FA_9295 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n738), .CI(C[225]), .S(S[225]), .CO(C[226]) );
  FA_9294 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n739), .CI(C[226]), .S(S[226]), .CO(C[227]) );
  FA_9293 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n740), .CI(C[227]), .S(S[227]), .CO(C[228]) );
  FA_9292 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n741), .CI(C[228]), .S(S[228]), .CO(C[229]) );
  FA_9291 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n742), .CI(C[229]), .S(S[229]), .CO(C[230]) );
  FA_9290 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n743), .CI(C[230]), .S(S[230]), .CO(C[231]) );
  FA_9289 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n744), .CI(C[231]), .S(S[231]), .CO(C[232]) );
  FA_9288 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n745), .CI(C[232]), .S(S[232]), .CO(C[233]) );
  FA_9287 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n746), .CI(C[233]), .S(S[233]), .CO(C[234]) );
  FA_9286 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n747), .CI(C[234]), .S(S[234]), .CO(C[235]) );
  FA_9285 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n748), .CI(C[235]), .S(S[235]), .CO(C[236]) );
  FA_9284 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n749), .CI(C[236]), .S(S[236]), .CO(C[237]) );
  FA_9283 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n750), .CI(C[237]), .S(S[237]), .CO(C[238]) );
  FA_9282 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n751), .CI(C[238]), .S(S[238]), .CO(C[239]) );
  FA_9281 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n752), .CI(C[239]), .S(S[239]), .CO(C[240]) );
  FA_9280 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n753), .CI(C[240]), .S(S[240]), .CO(C[241]) );
  FA_9279 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n754), .CI(C[241]), .S(S[241]), .CO(C[242]) );
  FA_9278 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n755), .CI(C[242]), .S(S[242]), .CO(C[243]) );
  FA_9277 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n756), .CI(C[243]), .S(S[243]), .CO(C[244]) );
  FA_9276 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n757), .CI(C[244]), .S(S[244]), .CO(C[245]) );
  FA_9275 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n758), .CI(C[245]), .S(S[245]), .CO(C[246]) );
  FA_9274 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n759), .CI(C[246]), .S(S[246]), .CO(C[247]) );
  FA_9273 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n760), .CI(C[247]), .S(S[247]), .CO(C[248]) );
  FA_9272 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n761), .CI(C[248]), .S(S[248]), .CO(C[249]) );
  FA_9271 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n762), .CI(C[249]), .S(S[249]), .CO(C[250]) );
  FA_9270 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n763), .CI(C[250]), .S(S[250]), .CO(C[251]) );
  FA_9269 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n764), .CI(C[251]), .S(S[251]), .CO(C[252]) );
  FA_9268 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n765), .CI(C[252]), .S(S[252]), .CO(C[253]) );
  FA_9267 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n766), .CI(C[253]), .S(S[253]), .CO(C[254]) );
  FA_9266 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n767), .CI(C[254]), .S(S[254]), .CO(C[255]) );
  FA_9265 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n768), .CI(C[255]), .S(S[255]), .CO(C[256]) );
  FA_9264 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n769), .CI(C[256]), .S(S[256]), .CO(C[257]) );
  FA_9263 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n770), .CI(C[257]), .S(S[257]), .CO(C[258]) );
  FA_9262 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n771), .CI(C[258]), .S(S[258]), .CO(C[259]) );
  FA_9261 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n772), .CI(C[259]), .S(S[259]), .CO(C[260]) );
  FA_9260 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n773), .CI(C[260]), .S(S[260]), .CO(C[261]) );
  FA_9259 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n774), .CI(C[261]), .S(S[261]), .CO(C[262]) );
  FA_9258 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n775), .CI(C[262]), .S(S[262]), .CO(C[263]) );
  FA_9257 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n776), .CI(C[263]), .S(S[263]), .CO(C[264]) );
  FA_9256 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n777), .CI(C[264]), .S(S[264]), .CO(C[265]) );
  FA_9255 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n778), .CI(C[265]), .S(S[265]), .CO(C[266]) );
  FA_9254 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n779), .CI(C[266]), .S(S[266]), .CO(C[267]) );
  FA_9253 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n780), .CI(C[267]), .S(S[267]), .CO(C[268]) );
  FA_9252 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n781), .CI(C[268]), .S(S[268]), .CO(C[269]) );
  FA_9251 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n782), .CI(C[269]), .S(S[269]), .CO(C[270]) );
  FA_9250 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n783), .CI(C[270]), .S(S[270]), .CO(C[271]) );
  FA_9249 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n784), .CI(C[271]), .S(S[271]), .CO(C[272]) );
  FA_9248 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n785), .CI(C[272]), .S(S[272]), .CO(C[273]) );
  FA_9247 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n786), .CI(C[273]), .S(S[273]), .CO(C[274]) );
  FA_9246 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n787), .CI(C[274]), .S(S[274]), .CO(C[275]) );
  FA_9245 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n788), .CI(C[275]), .S(S[275]), .CO(C[276]) );
  FA_9244 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n789), .CI(C[276]), .S(S[276]), .CO(C[277]) );
  FA_9243 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n790), .CI(C[277]), .S(S[277]), .CO(C[278]) );
  FA_9242 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n791), .CI(C[278]), .S(S[278]), .CO(C[279]) );
  FA_9241 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n792), .CI(C[279]), .S(S[279]), .CO(C[280]) );
  FA_9240 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n793), .CI(C[280]), .S(S[280]), .CO(C[281]) );
  FA_9239 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n794), .CI(C[281]), .S(S[281]), .CO(C[282]) );
  FA_9238 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n795), .CI(C[282]), .S(S[282]), .CO(C[283]) );
  FA_9237 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n796), .CI(C[283]), .S(S[283]), .CO(C[284]) );
  FA_9236 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n797), .CI(C[284]), .S(S[284]), .CO(C[285]) );
  FA_9235 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n798), .CI(C[285]), .S(S[285]), .CO(C[286]) );
  FA_9234 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n799), .CI(C[286]), .S(S[286]), .CO(C[287]) );
  FA_9233 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n800), .CI(C[287]), .S(S[287]), .CO(C[288]) );
  FA_9232 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n801), .CI(C[288]), .S(S[288]), .CO(C[289]) );
  FA_9231 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n802), .CI(C[289]), .S(S[289]), .CO(C[290]) );
  FA_9230 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n803), .CI(C[290]), .S(S[290]), .CO(C[291]) );
  FA_9229 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n804), .CI(C[291]), .S(S[291]), .CO(C[292]) );
  FA_9228 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n805), .CI(C[292]), .S(S[292]), .CO(C[293]) );
  FA_9227 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n806), .CI(C[293]), .S(S[293]), .CO(C[294]) );
  FA_9226 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n807), .CI(C[294]), .S(S[294]), .CO(C[295]) );
  FA_9225 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n808), .CI(C[295]), .S(S[295]), .CO(C[296]) );
  FA_9224 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n809), .CI(C[296]), .S(S[296]), .CO(C[297]) );
  FA_9223 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n810), .CI(C[297]), .S(S[297]), .CO(C[298]) );
  FA_9222 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n811), .CI(C[298]), .S(S[298]), .CO(C[299]) );
  FA_9221 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n812), .CI(C[299]), .S(S[299]), .CO(C[300]) );
  FA_9220 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n813), .CI(C[300]), .S(S[300]), .CO(C[301]) );
  FA_9219 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n814), .CI(C[301]), .S(S[301]), .CO(C[302]) );
  FA_9218 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n815), .CI(C[302]), .S(S[302]), .CO(C[303]) );
  FA_9217 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n816), .CI(C[303]), .S(S[303]), .CO(C[304]) );
  FA_9216 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n817), .CI(C[304]), .S(S[304]), .CO(C[305]) );
  FA_9215 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n818), .CI(C[305]), .S(S[305]), .CO(C[306]) );
  FA_9214 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n819), .CI(C[306]), .S(S[306]), .CO(C[307]) );
  FA_9213 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n820), .CI(C[307]), .S(S[307]), .CO(C[308]) );
  FA_9212 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n821), .CI(C[308]), .S(S[308]), .CO(C[309]) );
  FA_9211 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n822), .CI(C[309]), .S(S[309]), .CO(C[310]) );
  FA_9210 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n823), .CI(C[310]), .S(S[310]), .CO(C[311]) );
  FA_9209 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n824), .CI(C[311]), .S(S[311]), .CO(C[312]) );
  FA_9208 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n825), .CI(C[312]), .S(S[312]), .CO(C[313]) );
  FA_9207 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n826), .CI(C[313]), .S(S[313]), .CO(C[314]) );
  FA_9206 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n827), .CI(C[314]), .S(S[314]), .CO(C[315]) );
  FA_9205 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n828), .CI(C[315]), .S(S[315]), .CO(C[316]) );
  FA_9204 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n829), .CI(C[316]), .S(S[316]), .CO(C[317]) );
  FA_9203 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n830), .CI(C[317]), .S(S[317]), .CO(C[318]) );
  FA_9202 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n831), .CI(C[318]), .S(S[318]), .CO(C[319]) );
  FA_9201 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n832), .CI(C[319]), .S(S[319]), .CO(C[320]) );
  FA_9200 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n833), .CI(C[320]), .S(S[320]), .CO(C[321]) );
  FA_9199 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n834), .CI(C[321]), .S(S[321]), .CO(C[322]) );
  FA_9198 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n835), .CI(C[322]), .S(S[322]), .CO(C[323]) );
  FA_9197 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n836), .CI(C[323]), .S(S[323]), .CO(C[324]) );
  FA_9196 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n837), .CI(C[324]), .S(S[324]), .CO(C[325]) );
  FA_9195 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n838), .CI(C[325]), .S(S[325]), .CO(C[326]) );
  FA_9194 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n839), .CI(C[326]), .S(S[326]), .CO(C[327]) );
  FA_9193 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n840), .CI(C[327]), .S(S[327]), .CO(C[328]) );
  FA_9192 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n841), .CI(C[328]), .S(S[328]), .CO(C[329]) );
  FA_9191 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n842), .CI(C[329]), .S(S[329]), .CO(C[330]) );
  FA_9190 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n843), .CI(C[330]), .S(S[330]), .CO(C[331]) );
  FA_9189 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n844), .CI(C[331]), .S(S[331]), .CO(C[332]) );
  FA_9188 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n845), .CI(C[332]), .S(S[332]), .CO(C[333]) );
  FA_9187 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n846), .CI(C[333]), .S(S[333]), .CO(C[334]) );
  FA_9186 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n847), .CI(C[334]), .S(S[334]), .CO(C[335]) );
  FA_9185 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n848), .CI(C[335]), .S(S[335]), .CO(C[336]) );
  FA_9184 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n849), .CI(C[336]), .S(S[336]), .CO(C[337]) );
  FA_9183 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n850), .CI(C[337]), .S(S[337]), .CO(C[338]) );
  FA_9182 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n851), .CI(C[338]), .S(S[338]), .CO(C[339]) );
  FA_9181 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n852), .CI(C[339]), .S(S[339]), .CO(C[340]) );
  FA_9180 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n853), .CI(C[340]), .S(S[340]), .CO(C[341]) );
  FA_9179 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n854), .CI(C[341]), .S(S[341]), .CO(C[342]) );
  FA_9178 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n855), .CI(C[342]), .S(S[342]), .CO(C[343]) );
  FA_9177 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n856), .CI(C[343]), .S(S[343]), .CO(C[344]) );
  FA_9176 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n857), .CI(C[344]), .S(S[344]), .CO(C[345]) );
  FA_9175 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n858), .CI(C[345]), .S(S[345]), .CO(C[346]) );
  FA_9174 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n859), .CI(C[346]), .S(S[346]), .CO(C[347]) );
  FA_9173 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n860), .CI(C[347]), .S(S[347]), .CO(C[348]) );
  FA_9172 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n861), .CI(C[348]), .S(S[348]), .CO(C[349]) );
  FA_9171 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n862), .CI(C[349]), .S(S[349]), .CO(C[350]) );
  FA_9170 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n863), .CI(C[350]), .S(S[350]), .CO(C[351]) );
  FA_9169 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n864), .CI(C[351]), .S(S[351]), .CO(C[352]) );
  FA_9168 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n865), .CI(C[352]), .S(S[352]), .CO(C[353]) );
  FA_9167 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n866), .CI(C[353]), .S(S[353]), .CO(C[354]) );
  FA_9166 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n867), .CI(C[354]), .S(S[354]), .CO(C[355]) );
  FA_9165 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n868), .CI(C[355]), .S(S[355]), .CO(C[356]) );
  FA_9164 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n869), .CI(C[356]), .S(S[356]), .CO(C[357]) );
  FA_9163 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n870), .CI(C[357]), .S(S[357]), .CO(C[358]) );
  FA_9162 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n871), .CI(C[358]), .S(S[358]), .CO(C[359]) );
  FA_9161 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n872), .CI(C[359]), .S(S[359]), .CO(C[360]) );
  FA_9160 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n873), .CI(C[360]), .S(S[360]), .CO(C[361]) );
  FA_9159 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n874), .CI(C[361]), .S(S[361]), .CO(C[362]) );
  FA_9158 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n875), .CI(C[362]), .S(S[362]), .CO(C[363]) );
  FA_9157 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n876), .CI(C[363]), .S(S[363]), .CO(C[364]) );
  FA_9156 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n877), .CI(C[364]), .S(S[364]), .CO(C[365]) );
  FA_9155 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n878), .CI(C[365]), .S(S[365]), .CO(C[366]) );
  FA_9154 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n879), .CI(C[366]), .S(S[366]), .CO(C[367]) );
  FA_9153 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n880), .CI(C[367]), .S(S[367]), .CO(C[368]) );
  FA_9152 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n881), .CI(C[368]), .S(S[368]), .CO(C[369]) );
  FA_9151 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n882), .CI(C[369]), .S(S[369]), .CO(C[370]) );
  FA_9150 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n883), .CI(C[370]), .S(S[370]), .CO(C[371]) );
  FA_9149 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n884), .CI(C[371]), .S(S[371]), .CO(C[372]) );
  FA_9148 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n885), .CI(C[372]), .S(S[372]), .CO(C[373]) );
  FA_9147 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n886), .CI(C[373]), .S(S[373]), .CO(C[374]) );
  FA_9146 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n887), .CI(C[374]), .S(S[374]), .CO(C[375]) );
  FA_9145 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n888), .CI(C[375]), .S(S[375]), .CO(C[376]) );
  FA_9144 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n889), .CI(C[376]), .S(S[376]), .CO(C[377]) );
  FA_9143 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n890), .CI(C[377]), .S(S[377]), .CO(C[378]) );
  FA_9142 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n891), .CI(C[378]), .S(S[378]), .CO(C[379]) );
  FA_9141 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n892), .CI(C[379]), .S(S[379]), .CO(C[380]) );
  FA_9140 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n893), .CI(C[380]), .S(S[380]), .CO(C[381]) );
  FA_9139 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n894), .CI(C[381]), .S(S[381]), .CO(C[382]) );
  FA_9138 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n895), .CI(C[382]), .S(S[382]), .CO(C[383]) );
  FA_9137 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n896), .CI(C[383]), .S(S[383]), .CO(C[384]) );
  FA_9136 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n897), .CI(C[384]), .S(S[384]), .CO(C[385]) );
  FA_9135 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n898), .CI(C[385]), .S(S[385]), .CO(C[386]) );
  FA_9134 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n899), .CI(C[386]), .S(S[386]), .CO(C[387]) );
  FA_9133 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n900), .CI(C[387]), .S(S[387]), .CO(C[388]) );
  FA_9132 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n901), .CI(C[388]), .S(S[388]), .CO(C[389]) );
  FA_9131 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n902), .CI(C[389]), .S(S[389]), .CO(C[390]) );
  FA_9130 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n903), .CI(C[390]), .S(S[390]), .CO(C[391]) );
  FA_9129 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n904), .CI(C[391]), .S(S[391]), .CO(C[392]) );
  FA_9128 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n905), .CI(C[392]), .S(S[392]), .CO(C[393]) );
  FA_9127 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n906), .CI(C[393]), .S(S[393]), .CO(C[394]) );
  FA_9126 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n907), .CI(C[394]), .S(S[394]), .CO(C[395]) );
  FA_9125 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n908), .CI(C[395]), .S(S[395]), .CO(C[396]) );
  FA_9124 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n909), .CI(C[396]), .S(S[396]), .CO(C[397]) );
  FA_9123 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n910), .CI(C[397]), .S(S[397]), .CO(C[398]) );
  FA_9122 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n911), .CI(C[398]), .S(S[398]), .CO(C[399]) );
  FA_9121 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n912), .CI(C[399]), .S(S[399]), .CO(C[400]) );
  FA_9120 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n913), .CI(C[400]), .S(S[400]), .CO(C[401]) );
  FA_9119 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n914), .CI(C[401]), .S(S[401]), .CO(C[402]) );
  FA_9118 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n915), .CI(C[402]), .S(S[402]), .CO(C[403]) );
  FA_9117 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n916), .CI(C[403]), .S(S[403]), .CO(C[404]) );
  FA_9116 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n917), .CI(C[404]), .S(S[404]), .CO(C[405]) );
  FA_9115 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n918), .CI(C[405]), .S(S[405]), .CO(C[406]) );
  FA_9114 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n919), .CI(C[406]), .S(S[406]), .CO(C[407]) );
  FA_9113 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n920), .CI(C[407]), .S(S[407]), .CO(C[408]) );
  FA_9112 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n921), .CI(C[408]), .S(S[408]), .CO(C[409]) );
  FA_9111 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n922), .CI(C[409]), .S(S[409]), .CO(C[410]) );
  FA_9110 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n923), .CI(C[410]), .S(S[410]), .CO(C[411]) );
  FA_9109 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n924), .CI(C[411]), .S(S[411]), .CO(C[412]) );
  FA_9108 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n925), .CI(C[412]), .S(S[412]), .CO(C[413]) );
  FA_9107 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n926), .CI(C[413]), .S(S[413]), .CO(C[414]) );
  FA_9106 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n927), .CI(C[414]), .S(S[414]), .CO(C[415]) );
  FA_9105 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n928), .CI(C[415]), .S(S[415]), .CO(C[416]) );
  FA_9104 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n929), .CI(C[416]), .S(S[416]), .CO(C[417]) );
  FA_9103 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n930), .CI(C[417]), .S(S[417]), .CO(C[418]) );
  FA_9102 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n931), .CI(C[418]), .S(S[418]), .CO(C[419]) );
  FA_9101 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n932), .CI(C[419]), .S(S[419]), .CO(C[420]) );
  FA_9100 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n933), .CI(C[420]), .S(S[420]), .CO(C[421]) );
  FA_9099 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n934), .CI(C[421]), .S(S[421]), .CO(C[422]) );
  FA_9098 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n935), .CI(C[422]), .S(S[422]), .CO(C[423]) );
  FA_9097 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n936), .CI(C[423]), .S(S[423]), .CO(C[424]) );
  FA_9096 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n937), .CI(C[424]), .S(S[424]), .CO(C[425]) );
  FA_9095 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n938), .CI(C[425]), .S(S[425]), .CO(C[426]) );
  FA_9094 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n939), .CI(C[426]), .S(S[426]), .CO(C[427]) );
  FA_9093 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n940), .CI(C[427]), .S(S[427]), .CO(C[428]) );
  FA_9092 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n941), .CI(C[428]), .S(S[428]), .CO(C[429]) );
  FA_9091 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n942), .CI(C[429]), .S(S[429]), .CO(C[430]) );
  FA_9090 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n943), .CI(C[430]), .S(S[430]), .CO(C[431]) );
  FA_9089 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n944), .CI(C[431]), .S(S[431]), .CO(C[432]) );
  FA_9088 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n945), .CI(C[432]), .S(S[432]), .CO(C[433]) );
  FA_9087 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n946), .CI(C[433]), .S(S[433]), .CO(C[434]) );
  FA_9086 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n947), .CI(C[434]), .S(S[434]), .CO(C[435]) );
  FA_9085 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n948), .CI(C[435]), .S(S[435]), .CO(C[436]) );
  FA_9084 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n949), .CI(C[436]), .S(S[436]), .CO(C[437]) );
  FA_9083 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n950), .CI(C[437]), .S(S[437]), .CO(C[438]) );
  FA_9082 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n951), .CI(C[438]), .S(S[438]), .CO(C[439]) );
  FA_9081 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n952), .CI(C[439]), .S(S[439]), .CO(C[440]) );
  FA_9080 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n953), .CI(C[440]), .S(S[440]), .CO(C[441]) );
  FA_9079 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n954), .CI(C[441]), .S(S[441]), .CO(C[442]) );
  FA_9078 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n955), .CI(C[442]), .S(S[442]), .CO(C[443]) );
  FA_9077 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n956), .CI(C[443]), .S(S[443]), .CO(C[444]) );
  FA_9076 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n957), .CI(C[444]), .S(S[444]), .CO(C[445]) );
  FA_9075 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n958), .CI(C[445]), .S(S[445]), .CO(C[446]) );
  FA_9074 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n959), .CI(C[446]), .S(S[446]), .CO(C[447]) );
  FA_9073 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n960), .CI(C[447]), .S(S[447]), .CO(C[448]) );
  FA_9072 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n961), .CI(C[448]), .S(S[448]), .CO(C[449]) );
  FA_9071 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n962), .CI(C[449]), .S(S[449]), .CO(C[450]) );
  FA_9070 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n963), .CI(C[450]), .S(S[450]), .CO(C[451]) );
  FA_9069 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n964), .CI(C[451]), .S(S[451]), .CO(C[452]) );
  FA_9068 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n965), .CI(C[452]), .S(S[452]), .CO(C[453]) );
  FA_9067 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n966), .CI(C[453]), .S(S[453]), .CO(C[454]) );
  FA_9066 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n967), .CI(C[454]), .S(S[454]), .CO(C[455]) );
  FA_9065 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n968), .CI(C[455]), .S(S[455]), .CO(C[456]) );
  FA_9064 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n969), .CI(C[456]), .S(S[456]), .CO(C[457]) );
  FA_9063 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n970), .CI(C[457]), .S(S[457]), .CO(C[458]) );
  FA_9062 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n971), .CI(C[458]), .S(S[458]), .CO(C[459]) );
  FA_9061 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n972), .CI(C[459]), .S(S[459]), .CO(C[460]) );
  FA_9060 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n973), .CI(C[460]), .S(S[460]), .CO(C[461]) );
  FA_9059 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n974), .CI(C[461]), .S(S[461]), .CO(C[462]) );
  FA_9058 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n975), .CI(C[462]), .S(S[462]), .CO(C[463]) );
  FA_9057 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n976), .CI(C[463]), .S(S[463]), .CO(C[464]) );
  FA_9056 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n977), .CI(C[464]), .S(S[464]), .CO(C[465]) );
  FA_9055 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n978), .CI(C[465]), .S(S[465]), .CO(C[466]) );
  FA_9054 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n979), .CI(C[466]), .S(S[466]), .CO(C[467]) );
  FA_9053 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n980), .CI(C[467]), .S(S[467]), .CO(C[468]) );
  FA_9052 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n981), .CI(C[468]), .S(S[468]), .CO(C[469]) );
  FA_9051 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n982), .CI(C[469]), .S(S[469]), .CO(C[470]) );
  FA_9050 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n983), .CI(C[470]), .S(S[470]), .CO(C[471]) );
  FA_9049 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n984), .CI(C[471]), .S(S[471]), .CO(C[472]) );
  FA_9048 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n985), .CI(C[472]), .S(S[472]), .CO(C[473]) );
  FA_9047 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n986), .CI(C[473]), .S(S[473]), .CO(C[474]) );
  FA_9046 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n987), .CI(C[474]), .S(S[474]), .CO(C[475]) );
  FA_9045 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n988), .CI(C[475]), .S(S[475]), .CO(C[476]) );
  FA_9044 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n989), .CI(C[476]), .S(S[476]), .CO(C[477]) );
  FA_9043 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n990), .CI(C[477]), .S(S[477]), .CO(C[478]) );
  FA_9042 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n991), .CI(C[478]), .S(S[478]), .CO(C[479]) );
  FA_9041 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n992), .CI(C[479]), .S(S[479]), .CO(C[480]) );
  FA_9040 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n993), .CI(C[480]), .S(S[480]), .CO(C[481]) );
  FA_9039 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n994), .CI(C[481]), .S(S[481]), .CO(C[482]) );
  FA_9038 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n995), .CI(C[482]), .S(S[482]), .CO(C[483]) );
  FA_9037 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n996), .CI(C[483]), .S(S[483]), .CO(C[484]) );
  FA_9036 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n997), .CI(C[484]), .S(S[484]), .CO(C[485]) );
  FA_9035 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n998), .CI(C[485]), .S(S[485]), .CO(C[486]) );
  FA_9034 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n999), .CI(C[486]), .S(S[486]), .CO(C[487]) );
  FA_9033 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1000), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_9032 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1001), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_9031 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1002), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_9030 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1003), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_9029 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1004), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_9028 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1005), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_9027 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1006), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_9026 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1007), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_9025 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1008), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_9024 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1009), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_9023 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1010), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_9022 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1011), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_9021 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1012), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_9020 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1013), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_9019 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1014), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_9018 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1015), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_9017 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1016), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_9016 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1017), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_9015 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1018), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_9014 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1019), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_9013 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1020), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_9012 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1021), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_9011 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1022), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_9010 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1023), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_9009 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1024), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_9008 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .S(S[512])
         );
  IV U2 ( .A(B[415]), .Z(n928) );
  IV U3 ( .A(B[416]), .Z(n929) );
  IV U4 ( .A(B[417]), .Z(n930) );
  IV U5 ( .A(B[418]), .Z(n931) );
  IV U6 ( .A(B[419]), .Z(n932) );
  IV U7 ( .A(B[420]), .Z(n933) );
  IV U8 ( .A(B[421]), .Z(n934) );
  IV U9 ( .A(B[422]), .Z(n935) );
  IV U10 ( .A(B[423]), .Z(n936) );
  IV U11 ( .A(B[424]), .Z(n937) );
  IV U12 ( .A(B[505]), .Z(n1018) );
  IV U13 ( .A(B[425]), .Z(n938) );
  IV U14 ( .A(B[426]), .Z(n939) );
  IV U15 ( .A(B[427]), .Z(n940) );
  IV U16 ( .A(B[428]), .Z(n941) );
  IV U17 ( .A(B[429]), .Z(n942) );
  IV U18 ( .A(B[430]), .Z(n943) );
  IV U19 ( .A(B[431]), .Z(n944) );
  IV U20 ( .A(B[432]), .Z(n945) );
  IV U21 ( .A(B[433]), .Z(n946) );
  IV U22 ( .A(B[434]), .Z(n947) );
  IV U23 ( .A(B[506]), .Z(n1019) );
  IV U24 ( .A(B[435]), .Z(n948) );
  IV U25 ( .A(B[436]), .Z(n949) );
  IV U26 ( .A(B[437]), .Z(n950) );
  IV U27 ( .A(B[438]), .Z(n951) );
  IV U28 ( .A(B[439]), .Z(n952) );
  IV U29 ( .A(B[440]), .Z(n953) );
  IV U30 ( .A(B[441]), .Z(n954) );
  IV U31 ( .A(B[442]), .Z(n955) );
  IV U32 ( .A(B[443]), .Z(n956) );
  IV U33 ( .A(B[444]), .Z(n957) );
  IV U34 ( .A(B[507]), .Z(n1020) );
  IV U35 ( .A(B[445]), .Z(n958) );
  IV U36 ( .A(B[446]), .Z(n959) );
  IV U37 ( .A(B[447]), .Z(n960) );
  IV U38 ( .A(B[448]), .Z(n961) );
  IV U39 ( .A(B[449]), .Z(n962) );
  IV U40 ( .A(B[450]), .Z(n963) );
  IV U41 ( .A(B[451]), .Z(n964) );
  IV U42 ( .A(B[452]), .Z(n965) );
  IV U43 ( .A(B[453]), .Z(n966) );
  IV U44 ( .A(B[454]), .Z(n967) );
  IV U45 ( .A(B[508]), .Z(n1021) );
  IV U46 ( .A(B[455]), .Z(n968) );
  IV U47 ( .A(B[456]), .Z(n969) );
  IV U48 ( .A(B[457]), .Z(n970) );
  IV U49 ( .A(B[458]), .Z(n971) );
  IV U50 ( .A(B[459]), .Z(n972) );
  IV U51 ( .A(B[460]), .Z(n973) );
  IV U52 ( .A(B[461]), .Z(n974) );
  IV U53 ( .A(B[462]), .Z(n975) );
  IV U54 ( .A(B[0]), .Z(n2) );
  IV U55 ( .A(B[1]), .Z(n514) );
  IV U56 ( .A(B[2]), .Z(n515) );
  IV U57 ( .A(B[3]), .Z(n516) );
  IV U58 ( .A(B[4]), .Z(n517) );
  IV U59 ( .A(B[463]), .Z(n976) );
  IV U60 ( .A(B[5]), .Z(n518) );
  IV U61 ( .A(B[6]), .Z(n519) );
  IV U62 ( .A(B[7]), .Z(n520) );
  IV U63 ( .A(B[8]), .Z(n521) );
  IV U64 ( .A(B[9]), .Z(n522) );
  IV U65 ( .A(B[10]), .Z(n523) );
  IV U66 ( .A(B[11]), .Z(n524) );
  IV U67 ( .A(B[12]), .Z(n525) );
  IV U68 ( .A(B[13]), .Z(n526) );
  IV U69 ( .A(B[14]), .Z(n527) );
  IV U70 ( .A(B[464]), .Z(n977) );
  IV U71 ( .A(B[509]), .Z(n1022) );
  IV U72 ( .A(B[15]), .Z(n528) );
  IV U73 ( .A(B[16]), .Z(n529) );
  IV U74 ( .A(B[17]), .Z(n530) );
  IV U75 ( .A(B[18]), .Z(n531) );
  IV U76 ( .A(B[19]), .Z(n532) );
  IV U77 ( .A(B[20]), .Z(n533) );
  IV U78 ( .A(B[21]), .Z(n534) );
  IV U79 ( .A(B[22]), .Z(n535) );
  IV U80 ( .A(B[23]), .Z(n536) );
  IV U81 ( .A(B[24]), .Z(n537) );
  IV U82 ( .A(B[465]), .Z(n978) );
  IV U83 ( .A(B[25]), .Z(n538) );
  IV U84 ( .A(B[26]), .Z(n539) );
  IV U85 ( .A(B[27]), .Z(n540) );
  IV U86 ( .A(B[28]), .Z(n541) );
  IV U87 ( .A(B[29]), .Z(n542) );
  IV U88 ( .A(B[30]), .Z(n543) );
  IV U89 ( .A(B[31]), .Z(n544) );
  IV U90 ( .A(B[32]), .Z(n545) );
  IV U91 ( .A(B[33]), .Z(n546) );
  IV U92 ( .A(B[34]), .Z(n547) );
  IV U93 ( .A(B[466]), .Z(n979) );
  IV U94 ( .A(B[35]), .Z(n548) );
  IV U95 ( .A(B[36]), .Z(n549) );
  IV U96 ( .A(B[37]), .Z(n550) );
  IV U97 ( .A(B[38]), .Z(n551) );
  IV U98 ( .A(B[39]), .Z(n552) );
  IV U99 ( .A(B[40]), .Z(n553) );
  IV U100 ( .A(B[41]), .Z(n554) );
  IV U101 ( .A(B[42]), .Z(n555) );
  IV U102 ( .A(B[43]), .Z(n556) );
  IV U103 ( .A(B[44]), .Z(n557) );
  IV U104 ( .A(B[467]), .Z(n980) );
  IV U105 ( .A(B[45]), .Z(n558) );
  IV U106 ( .A(B[46]), .Z(n559) );
  IV U107 ( .A(B[47]), .Z(n560) );
  IV U108 ( .A(B[48]), .Z(n561) );
  IV U109 ( .A(B[49]), .Z(n562) );
  IV U110 ( .A(B[50]), .Z(n563) );
  IV U111 ( .A(B[51]), .Z(n564) );
  IV U112 ( .A(B[52]), .Z(n565) );
  IV U113 ( .A(B[53]), .Z(n566) );
  IV U114 ( .A(B[54]), .Z(n567) );
  IV U115 ( .A(B[468]), .Z(n981) );
  IV U116 ( .A(B[55]), .Z(n568) );
  IV U117 ( .A(B[56]), .Z(n569) );
  IV U118 ( .A(B[57]), .Z(n570) );
  IV U119 ( .A(B[58]), .Z(n571) );
  IV U120 ( .A(B[59]), .Z(n572) );
  IV U121 ( .A(B[60]), .Z(n573) );
  IV U122 ( .A(B[61]), .Z(n574) );
  IV U123 ( .A(B[62]), .Z(n575) );
  IV U124 ( .A(B[63]), .Z(n576) );
  IV U125 ( .A(B[64]), .Z(n577) );
  IV U126 ( .A(B[469]), .Z(n982) );
  IV U127 ( .A(B[65]), .Z(n578) );
  IV U128 ( .A(B[66]), .Z(n579) );
  IV U129 ( .A(B[67]), .Z(n580) );
  IV U130 ( .A(B[68]), .Z(n581) );
  IV U131 ( .A(B[69]), .Z(n582) );
  IV U132 ( .A(B[70]), .Z(n583) );
  IV U133 ( .A(B[71]), .Z(n584) );
  IV U134 ( .A(B[72]), .Z(n585) );
  IV U135 ( .A(B[73]), .Z(n586) );
  IV U136 ( .A(B[74]), .Z(n587) );
  IV U137 ( .A(B[470]), .Z(n983) );
  IV U138 ( .A(B[75]), .Z(n588) );
  IV U139 ( .A(B[76]), .Z(n589) );
  IV U140 ( .A(B[77]), .Z(n590) );
  IV U141 ( .A(B[78]), .Z(n591) );
  IV U142 ( .A(B[79]), .Z(n592) );
  IV U143 ( .A(B[80]), .Z(n593) );
  IV U144 ( .A(B[81]), .Z(n594) );
  IV U145 ( .A(B[82]), .Z(n595) );
  IV U146 ( .A(B[83]), .Z(n596) );
  IV U147 ( .A(B[84]), .Z(n597) );
  IV U148 ( .A(B[471]), .Z(n984) );
  IV U149 ( .A(B[85]), .Z(n598) );
  IV U150 ( .A(B[86]), .Z(n599) );
  IV U151 ( .A(B[87]), .Z(n600) );
  IV U152 ( .A(B[88]), .Z(n601) );
  IV U153 ( .A(B[89]), .Z(n602) );
  IV U154 ( .A(B[90]), .Z(n603) );
  IV U155 ( .A(B[91]), .Z(n604) );
  IV U156 ( .A(B[92]), .Z(n605) );
  IV U157 ( .A(B[93]), .Z(n606) );
  IV U158 ( .A(B[94]), .Z(n607) );
  IV U159 ( .A(B[472]), .Z(n985) );
  IV U160 ( .A(B[95]), .Z(n608) );
  IV U161 ( .A(B[96]), .Z(n609) );
  IV U162 ( .A(B[97]), .Z(n610) );
  IV U163 ( .A(B[98]), .Z(n611) );
  IV U164 ( .A(B[99]), .Z(n612) );
  IV U165 ( .A(B[100]), .Z(n613) );
  IV U166 ( .A(B[101]), .Z(n614) );
  IV U167 ( .A(B[102]), .Z(n615) );
  IV U168 ( .A(B[103]), .Z(n616) );
  IV U169 ( .A(B[104]), .Z(n617) );
  IV U170 ( .A(B[473]), .Z(n986) );
  IV U171 ( .A(B[105]), .Z(n618) );
  IV U172 ( .A(B[106]), .Z(n619) );
  IV U173 ( .A(B[107]), .Z(n620) );
  IV U174 ( .A(B[108]), .Z(n621) );
  IV U175 ( .A(B[109]), .Z(n622) );
  IV U176 ( .A(B[110]), .Z(n623) );
  IV U177 ( .A(B[111]), .Z(n624) );
  IV U178 ( .A(B[112]), .Z(n625) );
  IV U179 ( .A(B[113]), .Z(n626) );
  IV U180 ( .A(B[114]), .Z(n627) );
  IV U181 ( .A(B[474]), .Z(n987) );
  IV U182 ( .A(B[510]), .Z(n1023) );
  IV U183 ( .A(B[115]), .Z(n628) );
  IV U184 ( .A(B[116]), .Z(n629) );
  IV U185 ( .A(B[117]), .Z(n630) );
  IV U186 ( .A(B[118]), .Z(n631) );
  IV U187 ( .A(B[119]), .Z(n632) );
  IV U188 ( .A(B[120]), .Z(n633) );
  IV U189 ( .A(B[121]), .Z(n634) );
  IV U190 ( .A(B[122]), .Z(n635) );
  IV U191 ( .A(B[123]), .Z(n636) );
  IV U192 ( .A(B[124]), .Z(n637) );
  IV U193 ( .A(B[475]), .Z(n988) );
  IV U194 ( .A(B[125]), .Z(n638) );
  IV U195 ( .A(B[126]), .Z(n639) );
  IV U196 ( .A(B[127]), .Z(n640) );
  IV U197 ( .A(B[128]), .Z(n641) );
  IV U198 ( .A(B[129]), .Z(n642) );
  IV U199 ( .A(B[130]), .Z(n643) );
  IV U200 ( .A(B[131]), .Z(n644) );
  IV U201 ( .A(B[132]), .Z(n645) );
  IV U202 ( .A(B[133]), .Z(n646) );
  IV U203 ( .A(B[134]), .Z(n647) );
  IV U204 ( .A(B[476]), .Z(n989) );
  IV U205 ( .A(B[135]), .Z(n648) );
  IV U206 ( .A(B[136]), .Z(n649) );
  IV U207 ( .A(B[137]), .Z(n650) );
  IV U208 ( .A(B[138]), .Z(n651) );
  IV U209 ( .A(B[139]), .Z(n652) );
  IV U210 ( .A(B[140]), .Z(n653) );
  IV U211 ( .A(B[141]), .Z(n654) );
  IV U212 ( .A(B[142]), .Z(n655) );
  IV U213 ( .A(B[143]), .Z(n656) );
  IV U214 ( .A(B[144]), .Z(n657) );
  IV U215 ( .A(B[477]), .Z(n990) );
  IV U216 ( .A(B[145]), .Z(n658) );
  IV U217 ( .A(B[146]), .Z(n659) );
  IV U218 ( .A(B[147]), .Z(n660) );
  IV U219 ( .A(B[148]), .Z(n661) );
  IV U220 ( .A(B[149]), .Z(n662) );
  IV U221 ( .A(B[150]), .Z(n663) );
  IV U222 ( .A(B[151]), .Z(n664) );
  IV U223 ( .A(B[152]), .Z(n665) );
  IV U224 ( .A(B[153]), .Z(n666) );
  IV U225 ( .A(B[154]), .Z(n667) );
  IV U226 ( .A(B[478]), .Z(n991) );
  IV U227 ( .A(B[155]), .Z(n668) );
  IV U228 ( .A(B[156]), .Z(n669) );
  IV U229 ( .A(B[157]), .Z(n670) );
  IV U230 ( .A(B[158]), .Z(n671) );
  IV U231 ( .A(B[159]), .Z(n672) );
  IV U232 ( .A(B[160]), .Z(n673) );
  IV U233 ( .A(B[161]), .Z(n674) );
  IV U234 ( .A(B[162]), .Z(n675) );
  IV U235 ( .A(B[163]), .Z(n676) );
  IV U236 ( .A(B[164]), .Z(n677) );
  IV U237 ( .A(B[479]), .Z(n992) );
  IV U238 ( .A(B[165]), .Z(n678) );
  IV U239 ( .A(B[166]), .Z(n679) );
  IV U240 ( .A(B[167]), .Z(n680) );
  IV U241 ( .A(B[168]), .Z(n681) );
  IV U242 ( .A(B[169]), .Z(n682) );
  IV U243 ( .A(B[170]), .Z(n683) );
  IV U244 ( .A(B[171]), .Z(n684) );
  IV U245 ( .A(B[172]), .Z(n685) );
  IV U246 ( .A(B[173]), .Z(n686) );
  IV U247 ( .A(B[174]), .Z(n687) );
  IV U248 ( .A(B[480]), .Z(n993) );
  IV U249 ( .A(B[175]), .Z(n688) );
  IV U250 ( .A(B[176]), .Z(n689) );
  IV U251 ( .A(B[177]), .Z(n690) );
  IV U252 ( .A(B[178]), .Z(n691) );
  IV U253 ( .A(B[179]), .Z(n692) );
  IV U254 ( .A(B[180]), .Z(n693) );
  IV U255 ( .A(B[181]), .Z(n694) );
  IV U256 ( .A(B[182]), .Z(n695) );
  IV U257 ( .A(B[183]), .Z(n696) );
  IV U258 ( .A(B[184]), .Z(n697) );
  IV U259 ( .A(B[481]), .Z(n994) );
  IV U260 ( .A(B[185]), .Z(n698) );
  IV U261 ( .A(B[186]), .Z(n699) );
  IV U262 ( .A(B[187]), .Z(n700) );
  IV U263 ( .A(B[188]), .Z(n701) );
  IV U264 ( .A(B[189]), .Z(n702) );
  IV U265 ( .A(B[190]), .Z(n703) );
  IV U266 ( .A(B[191]), .Z(n704) );
  IV U267 ( .A(B[192]), .Z(n705) );
  IV U268 ( .A(B[193]), .Z(n706) );
  IV U269 ( .A(B[194]), .Z(n707) );
  IV U270 ( .A(B[482]), .Z(n995) );
  IV U271 ( .A(B[195]), .Z(n708) );
  IV U272 ( .A(B[196]), .Z(n709) );
  IV U273 ( .A(B[197]), .Z(n710) );
  IV U274 ( .A(B[198]), .Z(n711) );
  IV U275 ( .A(B[199]), .Z(n712) );
  IV U276 ( .A(B[200]), .Z(n713) );
  IV U277 ( .A(B[201]), .Z(n714) );
  IV U278 ( .A(B[202]), .Z(n715) );
  IV U279 ( .A(B[203]), .Z(n716) );
  IV U280 ( .A(B[204]), .Z(n717) );
  IV U281 ( .A(B[483]), .Z(n996) );
  IV U282 ( .A(B[205]), .Z(n718) );
  IV U283 ( .A(B[206]), .Z(n719) );
  IV U284 ( .A(B[207]), .Z(n720) );
  IV U285 ( .A(B[208]), .Z(n721) );
  IV U286 ( .A(B[209]), .Z(n722) );
  IV U287 ( .A(B[210]), .Z(n723) );
  IV U288 ( .A(B[211]), .Z(n724) );
  IV U289 ( .A(B[212]), .Z(n725) );
  IV U290 ( .A(B[213]), .Z(n726) );
  IV U291 ( .A(B[214]), .Z(n727) );
  IV U292 ( .A(B[484]), .Z(n997) );
  IV U293 ( .A(B[511]), .Z(n1024) );
  IV U294 ( .A(B[215]), .Z(n728) );
  IV U295 ( .A(B[216]), .Z(n729) );
  IV U296 ( .A(B[217]), .Z(n730) );
  IV U297 ( .A(B[218]), .Z(n731) );
  IV U298 ( .A(B[219]), .Z(n732) );
  IV U299 ( .A(B[220]), .Z(n733) );
  IV U300 ( .A(B[221]), .Z(n734) );
  IV U301 ( .A(B[222]), .Z(n735) );
  IV U302 ( .A(B[223]), .Z(n736) );
  IV U303 ( .A(B[224]), .Z(n737) );
  IV U304 ( .A(B[485]), .Z(n998) );
  IV U305 ( .A(B[225]), .Z(n738) );
  IV U306 ( .A(B[226]), .Z(n739) );
  IV U307 ( .A(B[227]), .Z(n740) );
  IV U308 ( .A(B[228]), .Z(n741) );
  IV U309 ( .A(B[229]), .Z(n742) );
  IV U310 ( .A(B[230]), .Z(n743) );
  IV U311 ( .A(B[231]), .Z(n744) );
  IV U312 ( .A(B[232]), .Z(n745) );
  IV U313 ( .A(B[233]), .Z(n746) );
  IV U314 ( .A(B[234]), .Z(n747) );
  IV U315 ( .A(B[486]), .Z(n999) );
  IV U316 ( .A(B[235]), .Z(n748) );
  IV U317 ( .A(B[236]), .Z(n749) );
  IV U318 ( .A(B[237]), .Z(n750) );
  IV U319 ( .A(B[238]), .Z(n751) );
  IV U320 ( .A(B[239]), .Z(n752) );
  IV U321 ( .A(B[240]), .Z(n753) );
  IV U322 ( .A(B[241]), .Z(n754) );
  IV U323 ( .A(B[242]), .Z(n755) );
  IV U324 ( .A(B[243]), .Z(n756) );
  IV U325 ( .A(B[244]), .Z(n757) );
  IV U326 ( .A(B[487]), .Z(n1000) );
  IV U327 ( .A(B[245]), .Z(n758) );
  IV U328 ( .A(B[246]), .Z(n759) );
  IV U329 ( .A(B[247]), .Z(n760) );
  IV U330 ( .A(B[248]), .Z(n761) );
  IV U331 ( .A(B[249]), .Z(n762) );
  IV U332 ( .A(B[250]), .Z(n763) );
  IV U333 ( .A(B[251]), .Z(n764) );
  IV U334 ( .A(B[252]), .Z(n765) );
  IV U335 ( .A(B[253]), .Z(n766) );
  IV U336 ( .A(B[254]), .Z(n767) );
  IV U337 ( .A(B[488]), .Z(n1001) );
  IV U338 ( .A(B[255]), .Z(n768) );
  IV U339 ( .A(B[256]), .Z(n769) );
  IV U340 ( .A(B[257]), .Z(n770) );
  IV U341 ( .A(B[258]), .Z(n771) );
  IV U342 ( .A(B[259]), .Z(n772) );
  IV U343 ( .A(B[260]), .Z(n773) );
  IV U344 ( .A(B[261]), .Z(n774) );
  IV U345 ( .A(B[262]), .Z(n775) );
  IV U346 ( .A(B[263]), .Z(n776) );
  IV U347 ( .A(B[264]), .Z(n777) );
  IV U348 ( .A(B[489]), .Z(n1002) );
  IV U349 ( .A(B[265]), .Z(n778) );
  IV U350 ( .A(B[266]), .Z(n779) );
  IV U351 ( .A(B[267]), .Z(n780) );
  IV U352 ( .A(B[268]), .Z(n781) );
  IV U353 ( .A(B[269]), .Z(n782) );
  IV U354 ( .A(B[270]), .Z(n783) );
  IV U355 ( .A(B[271]), .Z(n784) );
  IV U356 ( .A(B[272]), .Z(n785) );
  IV U357 ( .A(B[273]), .Z(n786) );
  IV U358 ( .A(B[274]), .Z(n787) );
  IV U359 ( .A(B[490]), .Z(n1003) );
  IV U360 ( .A(B[275]), .Z(n788) );
  IV U361 ( .A(B[276]), .Z(n789) );
  IV U362 ( .A(B[277]), .Z(n790) );
  IV U363 ( .A(B[278]), .Z(n791) );
  IV U364 ( .A(B[279]), .Z(n792) );
  IV U365 ( .A(B[280]), .Z(n793) );
  IV U366 ( .A(B[281]), .Z(n794) );
  IV U367 ( .A(B[282]), .Z(n795) );
  IV U368 ( .A(B[283]), .Z(n796) );
  IV U369 ( .A(B[284]), .Z(n797) );
  IV U370 ( .A(B[491]), .Z(n1004) );
  IV U371 ( .A(B[285]), .Z(n798) );
  IV U372 ( .A(B[286]), .Z(n799) );
  IV U373 ( .A(B[287]), .Z(n800) );
  IV U374 ( .A(B[288]), .Z(n801) );
  IV U375 ( .A(B[289]), .Z(n802) );
  IV U376 ( .A(B[290]), .Z(n803) );
  IV U377 ( .A(B[291]), .Z(n804) );
  IV U378 ( .A(B[292]), .Z(n805) );
  IV U379 ( .A(B[293]), .Z(n806) );
  IV U380 ( .A(B[294]), .Z(n807) );
  IV U381 ( .A(B[492]), .Z(n1005) );
  IV U382 ( .A(B[295]), .Z(n808) );
  IV U383 ( .A(B[296]), .Z(n809) );
  IV U384 ( .A(B[297]), .Z(n810) );
  IV U385 ( .A(B[298]), .Z(n811) );
  IV U386 ( .A(B[299]), .Z(n812) );
  IV U387 ( .A(B[300]), .Z(n813) );
  IV U388 ( .A(B[301]), .Z(n814) );
  IV U389 ( .A(B[302]), .Z(n815) );
  IV U390 ( .A(B[303]), .Z(n816) );
  IV U391 ( .A(B[304]), .Z(n817) );
  IV U392 ( .A(B[493]), .Z(n1006) );
  IV U393 ( .A(B[305]), .Z(n818) );
  IV U394 ( .A(B[306]), .Z(n819) );
  IV U395 ( .A(B[307]), .Z(n820) );
  IV U396 ( .A(B[308]), .Z(n821) );
  IV U397 ( .A(B[309]), .Z(n822) );
  IV U398 ( .A(B[310]), .Z(n823) );
  IV U399 ( .A(B[311]), .Z(n824) );
  IV U400 ( .A(B[312]), .Z(n825) );
  IV U401 ( .A(B[313]), .Z(n826) );
  IV U402 ( .A(B[314]), .Z(n827) );
  IV U403 ( .A(B[494]), .Z(n1007) );
  IV U404 ( .A(B[315]), .Z(n828) );
  IV U405 ( .A(B[316]), .Z(n829) );
  IV U406 ( .A(B[317]), .Z(n830) );
  IV U407 ( .A(B[318]), .Z(n831) );
  IV U408 ( .A(B[319]), .Z(n832) );
  IV U409 ( .A(B[320]), .Z(n833) );
  IV U410 ( .A(B[321]), .Z(n834) );
  IV U411 ( .A(B[322]), .Z(n835) );
  IV U412 ( .A(B[323]), .Z(n836) );
  IV U413 ( .A(B[324]), .Z(n837) );
  IV U414 ( .A(B[495]), .Z(n1008) );
  IV U415 ( .A(B[325]), .Z(n838) );
  IV U416 ( .A(B[326]), .Z(n839) );
  IV U417 ( .A(B[327]), .Z(n840) );
  IV U418 ( .A(B[328]), .Z(n841) );
  IV U419 ( .A(B[329]), .Z(n842) );
  IV U420 ( .A(B[330]), .Z(n843) );
  IV U421 ( .A(B[331]), .Z(n844) );
  IV U422 ( .A(B[332]), .Z(n845) );
  IV U423 ( .A(B[333]), .Z(n846) );
  IV U424 ( .A(B[334]), .Z(n847) );
  IV U425 ( .A(B[496]), .Z(n1009) );
  IV U426 ( .A(B[335]), .Z(n848) );
  IV U427 ( .A(B[336]), .Z(n849) );
  IV U428 ( .A(B[337]), .Z(n850) );
  IV U429 ( .A(B[338]), .Z(n851) );
  IV U430 ( .A(B[339]), .Z(n852) );
  IV U431 ( .A(B[340]), .Z(n853) );
  IV U432 ( .A(B[341]), .Z(n854) );
  IV U433 ( .A(B[342]), .Z(n855) );
  IV U434 ( .A(B[343]), .Z(n856) );
  IV U435 ( .A(B[344]), .Z(n857) );
  IV U436 ( .A(B[497]), .Z(n1010) );
  IV U437 ( .A(B[345]), .Z(n858) );
  IV U438 ( .A(B[346]), .Z(n859) );
  IV U439 ( .A(B[347]), .Z(n860) );
  IV U440 ( .A(B[348]), .Z(n861) );
  IV U441 ( .A(B[349]), .Z(n862) );
  IV U442 ( .A(B[350]), .Z(n863) );
  IV U443 ( .A(B[351]), .Z(n864) );
  IV U444 ( .A(B[352]), .Z(n865) );
  IV U445 ( .A(B[353]), .Z(n866) );
  IV U446 ( .A(B[354]), .Z(n867) );
  IV U447 ( .A(B[498]), .Z(n1011) );
  IV U448 ( .A(B[355]), .Z(n868) );
  IV U449 ( .A(B[356]), .Z(n869) );
  IV U450 ( .A(B[357]), .Z(n870) );
  IV U451 ( .A(B[358]), .Z(n871) );
  IV U452 ( .A(B[359]), .Z(n872) );
  IV U453 ( .A(B[360]), .Z(n873) );
  IV U454 ( .A(B[361]), .Z(n874) );
  IV U455 ( .A(B[362]), .Z(n875) );
  IV U456 ( .A(B[363]), .Z(n876) );
  IV U457 ( .A(B[364]), .Z(n877) );
  IV U458 ( .A(B[499]), .Z(n1012) );
  IV U459 ( .A(B[365]), .Z(n878) );
  IV U460 ( .A(B[366]), .Z(n879) );
  IV U461 ( .A(B[367]), .Z(n880) );
  IV U462 ( .A(B[368]), .Z(n881) );
  IV U463 ( .A(B[369]), .Z(n882) );
  IV U464 ( .A(B[370]), .Z(n883) );
  IV U465 ( .A(B[371]), .Z(n884) );
  IV U466 ( .A(B[372]), .Z(n885) );
  IV U467 ( .A(B[373]), .Z(n886) );
  IV U468 ( .A(B[374]), .Z(n887) );
  IV U469 ( .A(B[500]), .Z(n1013) );
  IV U470 ( .A(B[375]), .Z(n888) );
  IV U471 ( .A(B[376]), .Z(n889) );
  IV U472 ( .A(B[377]), .Z(n890) );
  IV U473 ( .A(B[378]), .Z(n891) );
  IV U474 ( .A(B[379]), .Z(n892) );
  IV U475 ( .A(B[380]), .Z(n893) );
  IV U476 ( .A(B[381]), .Z(n894) );
  IV U477 ( .A(B[382]), .Z(n895) );
  IV U478 ( .A(B[383]), .Z(n896) );
  IV U479 ( .A(B[384]), .Z(n897) );
  IV U480 ( .A(B[501]), .Z(n1014) );
  IV U481 ( .A(B[385]), .Z(n898) );
  IV U482 ( .A(B[386]), .Z(n899) );
  IV U483 ( .A(B[387]), .Z(n900) );
  IV U484 ( .A(B[388]), .Z(n901) );
  IV U485 ( .A(B[389]), .Z(n902) );
  IV U486 ( .A(B[390]), .Z(n903) );
  IV U487 ( .A(B[391]), .Z(n904) );
  IV U488 ( .A(B[392]), .Z(n905) );
  IV U489 ( .A(B[393]), .Z(n906) );
  IV U490 ( .A(B[394]), .Z(n907) );
  IV U491 ( .A(B[502]), .Z(n1015) );
  IV U492 ( .A(B[395]), .Z(n908) );
  IV U493 ( .A(B[396]), .Z(n909) );
  IV U494 ( .A(B[397]), .Z(n910) );
  IV U495 ( .A(B[398]), .Z(n911) );
  IV U496 ( .A(B[399]), .Z(n912) );
  IV U497 ( .A(B[400]), .Z(n913) );
  IV U498 ( .A(B[401]), .Z(n914) );
  IV U499 ( .A(B[402]), .Z(n915) );
  IV U500 ( .A(B[403]), .Z(n916) );
  IV U501 ( .A(B[404]), .Z(n917) );
  IV U502 ( .A(B[503]), .Z(n1016) );
  IV U503 ( .A(B[405]), .Z(n918) );
  IV U504 ( .A(B[406]), .Z(n919) );
  IV U505 ( .A(B[407]), .Z(n920) );
  IV U506 ( .A(B[408]), .Z(n921) );
  IV U507 ( .A(B[409]), .Z(n922) );
  IV U508 ( .A(B[410]), .Z(n923) );
  IV U509 ( .A(B[411]), .Z(n924) );
  IV U510 ( .A(B[412]), .Z(n925) );
  IV U511 ( .A(B[413]), .Z(n926) );
  IV U512 ( .A(B[414]), .Z(n927) );
  IV U513 ( .A(B[504]), .Z(n1017) );
endmodule


module modmult_step_N512_1_0 ( xregN_1, y, n, zin, zout );
  input [511:0] y;
  input [511:0] n;
  input [513:0] zin;
  output [513:0] zout;
  input xregN_1;
  wire   c1, c2, n1;
  wire   [513:0] w1;
  wire   [513:0] w2;
  wire   [513:0] w3;
  wire   [513:0] z2;
  wire   [513:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  MUX_N514_3 MUX_1 ( .A({1'b0, 1'b0, y}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(xregN_1), .O({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, w1[511:0]}) );
  MUX_N514_8 MUX_2 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(c1), .O({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, w2[511:0]}) );
  MUX_N514_7 MUX_3 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(n1), .O({SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, w3[511:0]}) );
  ADD_N514_1_0 ADD_1 ( .A({zin[512:0], 1'b0}), .B({1'b0, 1'b0, w1[511:0]}), 
        .CI(1'b0), .S(z2) );
  COMP_N514_2 COMP_1 ( .A(z2), .B({1'b0, 1'b0, n}), .O(c1) );
  SUB_N514_2 SUB_1 ( .A(z2), .B({1'b0, 1'b0, w2[511:0]}), .S(z3) );
  COMP_N514_5 COMP_2 ( .A({1'b0, 1'b0, n}), .B(z3), .O(c2) );
  SUB_N514_5 SUB_2 ( .A({1'b0, z3[512:0]}), .B({1'b0, 1'b0, w3[511:0]}), .S({
        SYNOPSYS_UNCONNECTED__6, zout[512:0]}) );
  IV U2 ( .A(c2), .Z(n1) );
endmodule


module MUX_N514_4 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N514_5 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module MUX_N514_6 ( A, B, S, O );
  input [513:0] A;
  input [513:0] B;
  output [513:0] O;
  input S;


  ANDN U1 ( .B(A[9]), .A(S), .Z(O[9]) );
  ANDN U2 ( .B(A[99]), .A(S), .Z(O[99]) );
  ANDN U3 ( .B(A[98]), .A(S), .Z(O[98]) );
  ANDN U4 ( .B(A[97]), .A(S), .Z(O[97]) );
  ANDN U5 ( .B(A[96]), .A(S), .Z(O[96]) );
  ANDN U6 ( .B(A[95]), .A(S), .Z(O[95]) );
  ANDN U7 ( .B(A[94]), .A(S), .Z(O[94]) );
  ANDN U8 ( .B(A[93]), .A(S), .Z(O[93]) );
  ANDN U9 ( .B(A[92]), .A(S), .Z(O[92]) );
  ANDN U10 ( .B(A[91]), .A(S), .Z(O[91]) );
  ANDN U11 ( .B(A[90]), .A(S), .Z(O[90]) );
  ANDN U12 ( .B(A[8]), .A(S), .Z(O[8]) );
  ANDN U13 ( .B(A[89]), .A(S), .Z(O[89]) );
  ANDN U14 ( .B(A[88]), .A(S), .Z(O[88]) );
  ANDN U15 ( .B(A[87]), .A(S), .Z(O[87]) );
  ANDN U16 ( .B(A[86]), .A(S), .Z(O[86]) );
  ANDN U17 ( .B(A[85]), .A(S), .Z(O[85]) );
  ANDN U18 ( .B(A[84]), .A(S), .Z(O[84]) );
  ANDN U19 ( .B(A[83]), .A(S), .Z(O[83]) );
  ANDN U20 ( .B(A[82]), .A(S), .Z(O[82]) );
  ANDN U21 ( .B(A[81]), .A(S), .Z(O[81]) );
  ANDN U22 ( .B(A[80]), .A(S), .Z(O[80]) );
  ANDN U23 ( .B(A[7]), .A(S), .Z(O[7]) );
  ANDN U24 ( .B(A[79]), .A(S), .Z(O[79]) );
  ANDN U25 ( .B(A[78]), .A(S), .Z(O[78]) );
  ANDN U26 ( .B(A[77]), .A(S), .Z(O[77]) );
  ANDN U27 ( .B(A[76]), .A(S), .Z(O[76]) );
  ANDN U28 ( .B(A[75]), .A(S), .Z(O[75]) );
  ANDN U29 ( .B(A[74]), .A(S), .Z(O[74]) );
  ANDN U30 ( .B(A[73]), .A(S), .Z(O[73]) );
  ANDN U31 ( .B(A[72]), .A(S), .Z(O[72]) );
  ANDN U32 ( .B(A[71]), .A(S), .Z(O[71]) );
  ANDN U33 ( .B(A[70]), .A(S), .Z(O[70]) );
  ANDN U34 ( .B(A[6]), .A(S), .Z(O[6]) );
  ANDN U35 ( .B(A[69]), .A(S), .Z(O[69]) );
  ANDN U36 ( .B(A[68]), .A(S), .Z(O[68]) );
  ANDN U37 ( .B(A[67]), .A(S), .Z(O[67]) );
  ANDN U38 ( .B(A[66]), .A(S), .Z(O[66]) );
  ANDN U39 ( .B(A[65]), .A(S), .Z(O[65]) );
  ANDN U40 ( .B(A[64]), .A(S), .Z(O[64]) );
  ANDN U41 ( .B(A[63]), .A(S), .Z(O[63]) );
  ANDN U42 ( .B(A[62]), .A(S), .Z(O[62]) );
  ANDN U43 ( .B(A[61]), .A(S), .Z(O[61]) );
  ANDN U44 ( .B(A[60]), .A(S), .Z(O[60]) );
  ANDN U45 ( .B(A[5]), .A(S), .Z(O[5]) );
  ANDN U46 ( .B(A[59]), .A(S), .Z(O[59]) );
  ANDN U47 ( .B(A[58]), .A(S), .Z(O[58]) );
  ANDN U48 ( .B(A[57]), .A(S), .Z(O[57]) );
  ANDN U49 ( .B(A[56]), .A(S), .Z(O[56]) );
  ANDN U50 ( .B(A[55]), .A(S), .Z(O[55]) );
  ANDN U51 ( .B(A[54]), .A(S), .Z(O[54]) );
  ANDN U52 ( .B(A[53]), .A(S), .Z(O[53]) );
  ANDN U53 ( .B(A[52]), .A(S), .Z(O[52]) );
  ANDN U54 ( .B(A[51]), .A(S), .Z(O[51]) );
  ANDN U55 ( .B(A[511]), .A(S), .Z(O[511]) );
  ANDN U56 ( .B(A[510]), .A(S), .Z(O[510]) );
  ANDN U57 ( .B(A[50]), .A(S), .Z(O[50]) );
  ANDN U58 ( .B(A[509]), .A(S), .Z(O[509]) );
  ANDN U59 ( .B(A[508]), .A(S), .Z(O[508]) );
  ANDN U60 ( .B(A[507]), .A(S), .Z(O[507]) );
  ANDN U61 ( .B(A[506]), .A(S), .Z(O[506]) );
  ANDN U62 ( .B(A[505]), .A(S), .Z(O[505]) );
  ANDN U63 ( .B(A[504]), .A(S), .Z(O[504]) );
  ANDN U64 ( .B(A[503]), .A(S), .Z(O[503]) );
  ANDN U65 ( .B(A[502]), .A(S), .Z(O[502]) );
  ANDN U66 ( .B(A[501]), .A(S), .Z(O[501]) );
  ANDN U67 ( .B(A[500]), .A(S), .Z(O[500]) );
  ANDN U68 ( .B(A[4]), .A(S), .Z(O[4]) );
  ANDN U69 ( .B(A[49]), .A(S), .Z(O[49]) );
  ANDN U70 ( .B(A[499]), .A(S), .Z(O[499]) );
  ANDN U71 ( .B(A[498]), .A(S), .Z(O[498]) );
  ANDN U72 ( .B(A[497]), .A(S), .Z(O[497]) );
  ANDN U73 ( .B(A[496]), .A(S), .Z(O[496]) );
  ANDN U74 ( .B(A[495]), .A(S), .Z(O[495]) );
  ANDN U75 ( .B(A[494]), .A(S), .Z(O[494]) );
  ANDN U76 ( .B(A[493]), .A(S), .Z(O[493]) );
  ANDN U77 ( .B(A[492]), .A(S), .Z(O[492]) );
  ANDN U78 ( .B(A[491]), .A(S), .Z(O[491]) );
  ANDN U79 ( .B(A[490]), .A(S), .Z(O[490]) );
  ANDN U80 ( .B(A[48]), .A(S), .Z(O[48]) );
  ANDN U81 ( .B(A[489]), .A(S), .Z(O[489]) );
  ANDN U82 ( .B(A[488]), .A(S), .Z(O[488]) );
  ANDN U83 ( .B(A[487]), .A(S), .Z(O[487]) );
  ANDN U84 ( .B(A[486]), .A(S), .Z(O[486]) );
  ANDN U85 ( .B(A[485]), .A(S), .Z(O[485]) );
  ANDN U86 ( .B(A[484]), .A(S), .Z(O[484]) );
  ANDN U87 ( .B(A[483]), .A(S), .Z(O[483]) );
  ANDN U88 ( .B(A[482]), .A(S), .Z(O[482]) );
  ANDN U89 ( .B(A[481]), .A(S), .Z(O[481]) );
  ANDN U90 ( .B(A[480]), .A(S), .Z(O[480]) );
  ANDN U91 ( .B(A[47]), .A(S), .Z(O[47]) );
  ANDN U92 ( .B(A[479]), .A(S), .Z(O[479]) );
  ANDN U93 ( .B(A[478]), .A(S), .Z(O[478]) );
  ANDN U94 ( .B(A[477]), .A(S), .Z(O[477]) );
  ANDN U95 ( .B(A[476]), .A(S), .Z(O[476]) );
  ANDN U96 ( .B(A[475]), .A(S), .Z(O[475]) );
  ANDN U97 ( .B(A[474]), .A(S), .Z(O[474]) );
  ANDN U98 ( .B(A[473]), .A(S), .Z(O[473]) );
  ANDN U99 ( .B(A[472]), .A(S), .Z(O[472]) );
  ANDN U100 ( .B(A[471]), .A(S), .Z(O[471]) );
  ANDN U101 ( .B(A[470]), .A(S), .Z(O[470]) );
  ANDN U102 ( .B(A[46]), .A(S), .Z(O[46]) );
  ANDN U103 ( .B(A[469]), .A(S), .Z(O[469]) );
  ANDN U104 ( .B(A[468]), .A(S), .Z(O[468]) );
  ANDN U105 ( .B(A[467]), .A(S), .Z(O[467]) );
  ANDN U106 ( .B(A[466]), .A(S), .Z(O[466]) );
  ANDN U107 ( .B(A[465]), .A(S), .Z(O[465]) );
  ANDN U108 ( .B(A[464]), .A(S), .Z(O[464]) );
  ANDN U109 ( .B(A[463]), .A(S), .Z(O[463]) );
  ANDN U110 ( .B(A[462]), .A(S), .Z(O[462]) );
  ANDN U111 ( .B(A[461]), .A(S), .Z(O[461]) );
  ANDN U112 ( .B(A[460]), .A(S), .Z(O[460]) );
  ANDN U113 ( .B(A[45]), .A(S), .Z(O[45]) );
  ANDN U114 ( .B(A[459]), .A(S), .Z(O[459]) );
  ANDN U115 ( .B(A[458]), .A(S), .Z(O[458]) );
  ANDN U116 ( .B(A[457]), .A(S), .Z(O[457]) );
  ANDN U117 ( .B(A[456]), .A(S), .Z(O[456]) );
  ANDN U118 ( .B(A[455]), .A(S), .Z(O[455]) );
  ANDN U119 ( .B(A[454]), .A(S), .Z(O[454]) );
  ANDN U120 ( .B(A[453]), .A(S), .Z(O[453]) );
  ANDN U121 ( .B(A[452]), .A(S), .Z(O[452]) );
  ANDN U122 ( .B(A[451]), .A(S), .Z(O[451]) );
  ANDN U123 ( .B(A[450]), .A(S), .Z(O[450]) );
  ANDN U124 ( .B(A[44]), .A(S), .Z(O[44]) );
  ANDN U125 ( .B(A[449]), .A(S), .Z(O[449]) );
  ANDN U126 ( .B(A[448]), .A(S), .Z(O[448]) );
  ANDN U127 ( .B(A[447]), .A(S), .Z(O[447]) );
  ANDN U128 ( .B(A[446]), .A(S), .Z(O[446]) );
  ANDN U129 ( .B(A[445]), .A(S), .Z(O[445]) );
  ANDN U130 ( .B(A[444]), .A(S), .Z(O[444]) );
  ANDN U131 ( .B(A[443]), .A(S), .Z(O[443]) );
  ANDN U132 ( .B(A[442]), .A(S), .Z(O[442]) );
  ANDN U133 ( .B(A[441]), .A(S), .Z(O[441]) );
  ANDN U134 ( .B(A[440]), .A(S), .Z(O[440]) );
  ANDN U135 ( .B(A[43]), .A(S), .Z(O[43]) );
  ANDN U136 ( .B(A[439]), .A(S), .Z(O[439]) );
  ANDN U137 ( .B(A[438]), .A(S), .Z(O[438]) );
  ANDN U138 ( .B(A[437]), .A(S), .Z(O[437]) );
  ANDN U139 ( .B(A[436]), .A(S), .Z(O[436]) );
  ANDN U140 ( .B(A[435]), .A(S), .Z(O[435]) );
  ANDN U141 ( .B(A[434]), .A(S), .Z(O[434]) );
  ANDN U142 ( .B(A[433]), .A(S), .Z(O[433]) );
  ANDN U143 ( .B(A[432]), .A(S), .Z(O[432]) );
  ANDN U144 ( .B(A[431]), .A(S), .Z(O[431]) );
  ANDN U145 ( .B(A[430]), .A(S), .Z(O[430]) );
  ANDN U146 ( .B(A[42]), .A(S), .Z(O[42]) );
  ANDN U147 ( .B(A[429]), .A(S), .Z(O[429]) );
  ANDN U148 ( .B(A[428]), .A(S), .Z(O[428]) );
  ANDN U149 ( .B(A[427]), .A(S), .Z(O[427]) );
  ANDN U150 ( .B(A[426]), .A(S), .Z(O[426]) );
  ANDN U151 ( .B(A[425]), .A(S), .Z(O[425]) );
  ANDN U152 ( .B(A[424]), .A(S), .Z(O[424]) );
  ANDN U153 ( .B(A[423]), .A(S), .Z(O[423]) );
  ANDN U154 ( .B(A[422]), .A(S), .Z(O[422]) );
  ANDN U155 ( .B(A[421]), .A(S), .Z(O[421]) );
  ANDN U156 ( .B(A[420]), .A(S), .Z(O[420]) );
  ANDN U157 ( .B(A[41]), .A(S), .Z(O[41]) );
  ANDN U158 ( .B(A[419]), .A(S), .Z(O[419]) );
  ANDN U159 ( .B(A[418]), .A(S), .Z(O[418]) );
  ANDN U160 ( .B(A[417]), .A(S), .Z(O[417]) );
  ANDN U161 ( .B(A[416]), .A(S), .Z(O[416]) );
  ANDN U162 ( .B(A[415]), .A(S), .Z(O[415]) );
  ANDN U163 ( .B(A[414]), .A(S), .Z(O[414]) );
  ANDN U164 ( .B(A[413]), .A(S), .Z(O[413]) );
  ANDN U165 ( .B(A[412]), .A(S), .Z(O[412]) );
  ANDN U166 ( .B(A[411]), .A(S), .Z(O[411]) );
  ANDN U167 ( .B(A[410]), .A(S), .Z(O[410]) );
  ANDN U168 ( .B(A[40]), .A(S), .Z(O[40]) );
  ANDN U169 ( .B(A[409]), .A(S), .Z(O[409]) );
  ANDN U170 ( .B(A[408]), .A(S), .Z(O[408]) );
  ANDN U171 ( .B(A[407]), .A(S), .Z(O[407]) );
  ANDN U172 ( .B(A[406]), .A(S), .Z(O[406]) );
  ANDN U173 ( .B(A[405]), .A(S), .Z(O[405]) );
  ANDN U174 ( .B(A[404]), .A(S), .Z(O[404]) );
  ANDN U175 ( .B(A[403]), .A(S), .Z(O[403]) );
  ANDN U176 ( .B(A[402]), .A(S), .Z(O[402]) );
  ANDN U177 ( .B(A[401]), .A(S), .Z(O[401]) );
  ANDN U178 ( .B(A[400]), .A(S), .Z(O[400]) );
  ANDN U179 ( .B(A[3]), .A(S), .Z(O[3]) );
  ANDN U180 ( .B(A[39]), .A(S), .Z(O[39]) );
  ANDN U181 ( .B(A[399]), .A(S), .Z(O[399]) );
  ANDN U182 ( .B(A[398]), .A(S), .Z(O[398]) );
  ANDN U183 ( .B(A[397]), .A(S), .Z(O[397]) );
  ANDN U184 ( .B(A[396]), .A(S), .Z(O[396]) );
  ANDN U185 ( .B(A[395]), .A(S), .Z(O[395]) );
  ANDN U186 ( .B(A[394]), .A(S), .Z(O[394]) );
  ANDN U187 ( .B(A[393]), .A(S), .Z(O[393]) );
  ANDN U188 ( .B(A[392]), .A(S), .Z(O[392]) );
  ANDN U189 ( .B(A[391]), .A(S), .Z(O[391]) );
  ANDN U190 ( .B(A[390]), .A(S), .Z(O[390]) );
  ANDN U191 ( .B(A[38]), .A(S), .Z(O[38]) );
  ANDN U192 ( .B(A[389]), .A(S), .Z(O[389]) );
  ANDN U193 ( .B(A[388]), .A(S), .Z(O[388]) );
  ANDN U194 ( .B(A[387]), .A(S), .Z(O[387]) );
  ANDN U195 ( .B(A[386]), .A(S), .Z(O[386]) );
  ANDN U196 ( .B(A[385]), .A(S), .Z(O[385]) );
  ANDN U197 ( .B(A[384]), .A(S), .Z(O[384]) );
  ANDN U198 ( .B(A[383]), .A(S), .Z(O[383]) );
  ANDN U199 ( .B(A[382]), .A(S), .Z(O[382]) );
  ANDN U200 ( .B(A[381]), .A(S), .Z(O[381]) );
  ANDN U201 ( .B(A[380]), .A(S), .Z(O[380]) );
  ANDN U202 ( .B(A[37]), .A(S), .Z(O[37]) );
  ANDN U203 ( .B(A[379]), .A(S), .Z(O[379]) );
  ANDN U204 ( .B(A[378]), .A(S), .Z(O[378]) );
  ANDN U205 ( .B(A[377]), .A(S), .Z(O[377]) );
  ANDN U206 ( .B(A[376]), .A(S), .Z(O[376]) );
  ANDN U207 ( .B(A[375]), .A(S), .Z(O[375]) );
  ANDN U208 ( .B(A[374]), .A(S), .Z(O[374]) );
  ANDN U209 ( .B(A[373]), .A(S), .Z(O[373]) );
  ANDN U210 ( .B(A[372]), .A(S), .Z(O[372]) );
  ANDN U211 ( .B(A[371]), .A(S), .Z(O[371]) );
  ANDN U212 ( .B(A[370]), .A(S), .Z(O[370]) );
  ANDN U213 ( .B(A[36]), .A(S), .Z(O[36]) );
  ANDN U214 ( .B(A[369]), .A(S), .Z(O[369]) );
  ANDN U215 ( .B(A[368]), .A(S), .Z(O[368]) );
  ANDN U216 ( .B(A[367]), .A(S), .Z(O[367]) );
  ANDN U217 ( .B(A[366]), .A(S), .Z(O[366]) );
  ANDN U218 ( .B(A[365]), .A(S), .Z(O[365]) );
  ANDN U219 ( .B(A[364]), .A(S), .Z(O[364]) );
  ANDN U220 ( .B(A[363]), .A(S), .Z(O[363]) );
  ANDN U221 ( .B(A[362]), .A(S), .Z(O[362]) );
  ANDN U222 ( .B(A[361]), .A(S), .Z(O[361]) );
  ANDN U223 ( .B(A[360]), .A(S), .Z(O[360]) );
  ANDN U224 ( .B(A[35]), .A(S), .Z(O[35]) );
  ANDN U225 ( .B(A[359]), .A(S), .Z(O[359]) );
  ANDN U226 ( .B(A[358]), .A(S), .Z(O[358]) );
  ANDN U227 ( .B(A[357]), .A(S), .Z(O[357]) );
  ANDN U228 ( .B(A[356]), .A(S), .Z(O[356]) );
  ANDN U229 ( .B(A[355]), .A(S), .Z(O[355]) );
  ANDN U230 ( .B(A[354]), .A(S), .Z(O[354]) );
  ANDN U231 ( .B(A[353]), .A(S), .Z(O[353]) );
  ANDN U232 ( .B(A[352]), .A(S), .Z(O[352]) );
  ANDN U233 ( .B(A[351]), .A(S), .Z(O[351]) );
  ANDN U234 ( .B(A[350]), .A(S), .Z(O[350]) );
  ANDN U235 ( .B(A[34]), .A(S), .Z(O[34]) );
  ANDN U236 ( .B(A[349]), .A(S), .Z(O[349]) );
  ANDN U237 ( .B(A[348]), .A(S), .Z(O[348]) );
  ANDN U238 ( .B(A[347]), .A(S), .Z(O[347]) );
  ANDN U239 ( .B(A[346]), .A(S), .Z(O[346]) );
  ANDN U240 ( .B(A[345]), .A(S), .Z(O[345]) );
  ANDN U241 ( .B(A[344]), .A(S), .Z(O[344]) );
  ANDN U242 ( .B(A[343]), .A(S), .Z(O[343]) );
  ANDN U243 ( .B(A[342]), .A(S), .Z(O[342]) );
  ANDN U244 ( .B(A[341]), .A(S), .Z(O[341]) );
  ANDN U245 ( .B(A[340]), .A(S), .Z(O[340]) );
  ANDN U246 ( .B(A[33]), .A(S), .Z(O[33]) );
  ANDN U247 ( .B(A[339]), .A(S), .Z(O[339]) );
  ANDN U248 ( .B(A[338]), .A(S), .Z(O[338]) );
  ANDN U249 ( .B(A[337]), .A(S), .Z(O[337]) );
  ANDN U250 ( .B(A[336]), .A(S), .Z(O[336]) );
  ANDN U251 ( .B(A[335]), .A(S), .Z(O[335]) );
  ANDN U252 ( .B(A[334]), .A(S), .Z(O[334]) );
  ANDN U253 ( .B(A[333]), .A(S), .Z(O[333]) );
  ANDN U254 ( .B(A[332]), .A(S), .Z(O[332]) );
  ANDN U255 ( .B(A[331]), .A(S), .Z(O[331]) );
  ANDN U256 ( .B(A[330]), .A(S), .Z(O[330]) );
  ANDN U257 ( .B(A[32]), .A(S), .Z(O[32]) );
  ANDN U258 ( .B(A[329]), .A(S), .Z(O[329]) );
  ANDN U259 ( .B(A[328]), .A(S), .Z(O[328]) );
  ANDN U260 ( .B(A[327]), .A(S), .Z(O[327]) );
  ANDN U261 ( .B(A[326]), .A(S), .Z(O[326]) );
  ANDN U262 ( .B(A[325]), .A(S), .Z(O[325]) );
  ANDN U263 ( .B(A[324]), .A(S), .Z(O[324]) );
  ANDN U264 ( .B(A[323]), .A(S), .Z(O[323]) );
  ANDN U265 ( .B(A[322]), .A(S), .Z(O[322]) );
  ANDN U266 ( .B(A[321]), .A(S), .Z(O[321]) );
  ANDN U267 ( .B(A[320]), .A(S), .Z(O[320]) );
  ANDN U268 ( .B(A[31]), .A(S), .Z(O[31]) );
  ANDN U269 ( .B(A[319]), .A(S), .Z(O[319]) );
  ANDN U270 ( .B(A[318]), .A(S), .Z(O[318]) );
  ANDN U271 ( .B(A[317]), .A(S), .Z(O[317]) );
  ANDN U272 ( .B(A[316]), .A(S), .Z(O[316]) );
  ANDN U273 ( .B(A[315]), .A(S), .Z(O[315]) );
  ANDN U274 ( .B(A[314]), .A(S), .Z(O[314]) );
  ANDN U275 ( .B(A[313]), .A(S), .Z(O[313]) );
  ANDN U276 ( .B(A[312]), .A(S), .Z(O[312]) );
  ANDN U277 ( .B(A[311]), .A(S), .Z(O[311]) );
  ANDN U278 ( .B(A[310]), .A(S), .Z(O[310]) );
  ANDN U279 ( .B(A[30]), .A(S), .Z(O[30]) );
  ANDN U280 ( .B(A[309]), .A(S), .Z(O[309]) );
  ANDN U281 ( .B(A[308]), .A(S), .Z(O[308]) );
  ANDN U282 ( .B(A[307]), .A(S), .Z(O[307]) );
  ANDN U283 ( .B(A[306]), .A(S), .Z(O[306]) );
  ANDN U284 ( .B(A[305]), .A(S), .Z(O[305]) );
  ANDN U285 ( .B(A[304]), .A(S), .Z(O[304]) );
  ANDN U286 ( .B(A[303]), .A(S), .Z(O[303]) );
  ANDN U287 ( .B(A[302]), .A(S), .Z(O[302]) );
  ANDN U288 ( .B(A[301]), .A(S), .Z(O[301]) );
  ANDN U289 ( .B(A[300]), .A(S), .Z(O[300]) );
  ANDN U290 ( .B(A[2]), .A(S), .Z(O[2]) );
  ANDN U291 ( .B(A[29]), .A(S), .Z(O[29]) );
  ANDN U292 ( .B(A[299]), .A(S), .Z(O[299]) );
  ANDN U293 ( .B(A[298]), .A(S), .Z(O[298]) );
  ANDN U294 ( .B(A[297]), .A(S), .Z(O[297]) );
  ANDN U295 ( .B(A[296]), .A(S), .Z(O[296]) );
  ANDN U296 ( .B(A[295]), .A(S), .Z(O[295]) );
  ANDN U297 ( .B(A[294]), .A(S), .Z(O[294]) );
  ANDN U298 ( .B(A[293]), .A(S), .Z(O[293]) );
  ANDN U299 ( .B(A[292]), .A(S), .Z(O[292]) );
  ANDN U300 ( .B(A[291]), .A(S), .Z(O[291]) );
  ANDN U301 ( .B(A[290]), .A(S), .Z(O[290]) );
  ANDN U302 ( .B(A[28]), .A(S), .Z(O[28]) );
  ANDN U303 ( .B(A[289]), .A(S), .Z(O[289]) );
  ANDN U304 ( .B(A[288]), .A(S), .Z(O[288]) );
  ANDN U305 ( .B(A[287]), .A(S), .Z(O[287]) );
  ANDN U306 ( .B(A[286]), .A(S), .Z(O[286]) );
  ANDN U307 ( .B(A[285]), .A(S), .Z(O[285]) );
  ANDN U308 ( .B(A[284]), .A(S), .Z(O[284]) );
  ANDN U309 ( .B(A[283]), .A(S), .Z(O[283]) );
  ANDN U310 ( .B(A[282]), .A(S), .Z(O[282]) );
  ANDN U311 ( .B(A[281]), .A(S), .Z(O[281]) );
  ANDN U312 ( .B(A[280]), .A(S), .Z(O[280]) );
  ANDN U313 ( .B(A[27]), .A(S), .Z(O[27]) );
  ANDN U314 ( .B(A[279]), .A(S), .Z(O[279]) );
  ANDN U315 ( .B(A[278]), .A(S), .Z(O[278]) );
  ANDN U316 ( .B(A[277]), .A(S), .Z(O[277]) );
  ANDN U317 ( .B(A[276]), .A(S), .Z(O[276]) );
  ANDN U318 ( .B(A[275]), .A(S), .Z(O[275]) );
  ANDN U319 ( .B(A[274]), .A(S), .Z(O[274]) );
  ANDN U320 ( .B(A[273]), .A(S), .Z(O[273]) );
  ANDN U321 ( .B(A[272]), .A(S), .Z(O[272]) );
  ANDN U322 ( .B(A[271]), .A(S), .Z(O[271]) );
  ANDN U323 ( .B(A[270]), .A(S), .Z(O[270]) );
  ANDN U324 ( .B(A[26]), .A(S), .Z(O[26]) );
  ANDN U325 ( .B(A[269]), .A(S), .Z(O[269]) );
  ANDN U326 ( .B(A[268]), .A(S), .Z(O[268]) );
  ANDN U327 ( .B(A[267]), .A(S), .Z(O[267]) );
  ANDN U328 ( .B(A[266]), .A(S), .Z(O[266]) );
  ANDN U329 ( .B(A[265]), .A(S), .Z(O[265]) );
  ANDN U330 ( .B(A[264]), .A(S), .Z(O[264]) );
  ANDN U331 ( .B(A[263]), .A(S), .Z(O[263]) );
  ANDN U332 ( .B(A[262]), .A(S), .Z(O[262]) );
  ANDN U333 ( .B(A[261]), .A(S), .Z(O[261]) );
  ANDN U334 ( .B(A[260]), .A(S), .Z(O[260]) );
  ANDN U335 ( .B(A[25]), .A(S), .Z(O[25]) );
  ANDN U336 ( .B(A[259]), .A(S), .Z(O[259]) );
  ANDN U337 ( .B(A[258]), .A(S), .Z(O[258]) );
  ANDN U338 ( .B(A[257]), .A(S), .Z(O[257]) );
  ANDN U339 ( .B(A[256]), .A(S), .Z(O[256]) );
  ANDN U340 ( .B(A[255]), .A(S), .Z(O[255]) );
  ANDN U341 ( .B(A[254]), .A(S), .Z(O[254]) );
  ANDN U342 ( .B(A[253]), .A(S), .Z(O[253]) );
  ANDN U343 ( .B(A[252]), .A(S), .Z(O[252]) );
  ANDN U344 ( .B(A[251]), .A(S), .Z(O[251]) );
  ANDN U345 ( .B(A[250]), .A(S), .Z(O[250]) );
  ANDN U346 ( .B(A[24]), .A(S), .Z(O[24]) );
  ANDN U347 ( .B(A[249]), .A(S), .Z(O[249]) );
  ANDN U348 ( .B(A[248]), .A(S), .Z(O[248]) );
  ANDN U349 ( .B(A[247]), .A(S), .Z(O[247]) );
  ANDN U350 ( .B(A[246]), .A(S), .Z(O[246]) );
  ANDN U351 ( .B(A[245]), .A(S), .Z(O[245]) );
  ANDN U352 ( .B(A[244]), .A(S), .Z(O[244]) );
  ANDN U353 ( .B(A[243]), .A(S), .Z(O[243]) );
  ANDN U354 ( .B(A[242]), .A(S), .Z(O[242]) );
  ANDN U355 ( .B(A[241]), .A(S), .Z(O[241]) );
  ANDN U356 ( .B(A[240]), .A(S), .Z(O[240]) );
  ANDN U357 ( .B(A[23]), .A(S), .Z(O[23]) );
  ANDN U358 ( .B(A[239]), .A(S), .Z(O[239]) );
  ANDN U359 ( .B(A[238]), .A(S), .Z(O[238]) );
  ANDN U360 ( .B(A[237]), .A(S), .Z(O[237]) );
  ANDN U361 ( .B(A[236]), .A(S), .Z(O[236]) );
  ANDN U362 ( .B(A[235]), .A(S), .Z(O[235]) );
  ANDN U363 ( .B(A[234]), .A(S), .Z(O[234]) );
  ANDN U364 ( .B(A[233]), .A(S), .Z(O[233]) );
  ANDN U365 ( .B(A[232]), .A(S), .Z(O[232]) );
  ANDN U366 ( .B(A[231]), .A(S), .Z(O[231]) );
  ANDN U367 ( .B(A[230]), .A(S), .Z(O[230]) );
  ANDN U368 ( .B(A[22]), .A(S), .Z(O[22]) );
  ANDN U369 ( .B(A[229]), .A(S), .Z(O[229]) );
  ANDN U370 ( .B(A[228]), .A(S), .Z(O[228]) );
  ANDN U371 ( .B(A[227]), .A(S), .Z(O[227]) );
  ANDN U372 ( .B(A[226]), .A(S), .Z(O[226]) );
  ANDN U373 ( .B(A[225]), .A(S), .Z(O[225]) );
  ANDN U374 ( .B(A[224]), .A(S), .Z(O[224]) );
  ANDN U375 ( .B(A[223]), .A(S), .Z(O[223]) );
  ANDN U376 ( .B(A[222]), .A(S), .Z(O[222]) );
  ANDN U377 ( .B(A[221]), .A(S), .Z(O[221]) );
  ANDN U378 ( .B(A[220]), .A(S), .Z(O[220]) );
  ANDN U379 ( .B(A[21]), .A(S), .Z(O[21]) );
  ANDN U380 ( .B(A[219]), .A(S), .Z(O[219]) );
  ANDN U381 ( .B(A[218]), .A(S), .Z(O[218]) );
  ANDN U382 ( .B(A[217]), .A(S), .Z(O[217]) );
  ANDN U383 ( .B(A[216]), .A(S), .Z(O[216]) );
  ANDN U384 ( .B(A[215]), .A(S), .Z(O[215]) );
  ANDN U385 ( .B(A[214]), .A(S), .Z(O[214]) );
  ANDN U386 ( .B(A[213]), .A(S), .Z(O[213]) );
  ANDN U387 ( .B(A[212]), .A(S), .Z(O[212]) );
  ANDN U388 ( .B(A[211]), .A(S), .Z(O[211]) );
  ANDN U389 ( .B(A[210]), .A(S), .Z(O[210]) );
  ANDN U390 ( .B(A[20]), .A(S), .Z(O[20]) );
  ANDN U391 ( .B(A[209]), .A(S), .Z(O[209]) );
  ANDN U392 ( .B(A[208]), .A(S), .Z(O[208]) );
  ANDN U393 ( .B(A[207]), .A(S), .Z(O[207]) );
  ANDN U394 ( .B(A[206]), .A(S), .Z(O[206]) );
  ANDN U395 ( .B(A[205]), .A(S), .Z(O[205]) );
  ANDN U396 ( .B(A[204]), .A(S), .Z(O[204]) );
  ANDN U397 ( .B(A[203]), .A(S), .Z(O[203]) );
  ANDN U398 ( .B(A[202]), .A(S), .Z(O[202]) );
  ANDN U399 ( .B(A[201]), .A(S), .Z(O[201]) );
  ANDN U400 ( .B(A[200]), .A(S), .Z(O[200]) );
  ANDN U401 ( .B(A[1]), .A(S), .Z(O[1]) );
  ANDN U402 ( .B(A[19]), .A(S), .Z(O[19]) );
  ANDN U403 ( .B(A[199]), .A(S), .Z(O[199]) );
  ANDN U404 ( .B(A[198]), .A(S), .Z(O[198]) );
  ANDN U405 ( .B(A[197]), .A(S), .Z(O[197]) );
  ANDN U406 ( .B(A[196]), .A(S), .Z(O[196]) );
  ANDN U407 ( .B(A[195]), .A(S), .Z(O[195]) );
  ANDN U408 ( .B(A[194]), .A(S), .Z(O[194]) );
  ANDN U409 ( .B(A[193]), .A(S), .Z(O[193]) );
  ANDN U410 ( .B(A[192]), .A(S), .Z(O[192]) );
  ANDN U411 ( .B(A[191]), .A(S), .Z(O[191]) );
  ANDN U412 ( .B(A[190]), .A(S), .Z(O[190]) );
  ANDN U413 ( .B(A[18]), .A(S), .Z(O[18]) );
  ANDN U414 ( .B(A[189]), .A(S), .Z(O[189]) );
  ANDN U415 ( .B(A[188]), .A(S), .Z(O[188]) );
  ANDN U416 ( .B(A[187]), .A(S), .Z(O[187]) );
  ANDN U417 ( .B(A[186]), .A(S), .Z(O[186]) );
  ANDN U418 ( .B(A[185]), .A(S), .Z(O[185]) );
  ANDN U419 ( .B(A[184]), .A(S), .Z(O[184]) );
  ANDN U420 ( .B(A[183]), .A(S), .Z(O[183]) );
  ANDN U421 ( .B(A[182]), .A(S), .Z(O[182]) );
  ANDN U422 ( .B(A[181]), .A(S), .Z(O[181]) );
  ANDN U423 ( .B(A[180]), .A(S), .Z(O[180]) );
  ANDN U424 ( .B(A[17]), .A(S), .Z(O[17]) );
  ANDN U425 ( .B(A[179]), .A(S), .Z(O[179]) );
  ANDN U426 ( .B(A[178]), .A(S), .Z(O[178]) );
  ANDN U427 ( .B(A[177]), .A(S), .Z(O[177]) );
  ANDN U428 ( .B(A[176]), .A(S), .Z(O[176]) );
  ANDN U429 ( .B(A[175]), .A(S), .Z(O[175]) );
  ANDN U430 ( .B(A[174]), .A(S), .Z(O[174]) );
  ANDN U431 ( .B(A[173]), .A(S), .Z(O[173]) );
  ANDN U432 ( .B(A[172]), .A(S), .Z(O[172]) );
  ANDN U433 ( .B(A[171]), .A(S), .Z(O[171]) );
  ANDN U434 ( .B(A[170]), .A(S), .Z(O[170]) );
  ANDN U435 ( .B(A[16]), .A(S), .Z(O[16]) );
  ANDN U436 ( .B(A[169]), .A(S), .Z(O[169]) );
  ANDN U437 ( .B(A[168]), .A(S), .Z(O[168]) );
  ANDN U438 ( .B(A[167]), .A(S), .Z(O[167]) );
  ANDN U439 ( .B(A[166]), .A(S), .Z(O[166]) );
  ANDN U440 ( .B(A[165]), .A(S), .Z(O[165]) );
  ANDN U441 ( .B(A[164]), .A(S), .Z(O[164]) );
  ANDN U442 ( .B(A[163]), .A(S), .Z(O[163]) );
  ANDN U443 ( .B(A[162]), .A(S), .Z(O[162]) );
  ANDN U444 ( .B(A[161]), .A(S), .Z(O[161]) );
  ANDN U445 ( .B(A[160]), .A(S), .Z(O[160]) );
  ANDN U446 ( .B(A[15]), .A(S), .Z(O[15]) );
  ANDN U447 ( .B(A[159]), .A(S), .Z(O[159]) );
  ANDN U448 ( .B(A[158]), .A(S), .Z(O[158]) );
  ANDN U449 ( .B(A[157]), .A(S), .Z(O[157]) );
  ANDN U450 ( .B(A[156]), .A(S), .Z(O[156]) );
  ANDN U451 ( .B(A[155]), .A(S), .Z(O[155]) );
  ANDN U452 ( .B(A[154]), .A(S), .Z(O[154]) );
  ANDN U453 ( .B(A[153]), .A(S), .Z(O[153]) );
  ANDN U454 ( .B(A[152]), .A(S), .Z(O[152]) );
  ANDN U455 ( .B(A[151]), .A(S), .Z(O[151]) );
  ANDN U456 ( .B(A[150]), .A(S), .Z(O[150]) );
  ANDN U457 ( .B(A[14]), .A(S), .Z(O[14]) );
  ANDN U458 ( .B(A[149]), .A(S), .Z(O[149]) );
  ANDN U459 ( .B(A[148]), .A(S), .Z(O[148]) );
  ANDN U460 ( .B(A[147]), .A(S), .Z(O[147]) );
  ANDN U461 ( .B(A[146]), .A(S), .Z(O[146]) );
  ANDN U462 ( .B(A[145]), .A(S), .Z(O[145]) );
  ANDN U463 ( .B(A[144]), .A(S), .Z(O[144]) );
  ANDN U464 ( .B(A[143]), .A(S), .Z(O[143]) );
  ANDN U465 ( .B(A[142]), .A(S), .Z(O[142]) );
  ANDN U466 ( .B(A[141]), .A(S), .Z(O[141]) );
  ANDN U467 ( .B(A[140]), .A(S), .Z(O[140]) );
  ANDN U468 ( .B(A[13]), .A(S), .Z(O[13]) );
  ANDN U469 ( .B(A[139]), .A(S), .Z(O[139]) );
  ANDN U470 ( .B(A[138]), .A(S), .Z(O[138]) );
  ANDN U471 ( .B(A[137]), .A(S), .Z(O[137]) );
  ANDN U472 ( .B(A[136]), .A(S), .Z(O[136]) );
  ANDN U473 ( .B(A[135]), .A(S), .Z(O[135]) );
  ANDN U474 ( .B(A[134]), .A(S), .Z(O[134]) );
  ANDN U475 ( .B(A[133]), .A(S), .Z(O[133]) );
  ANDN U476 ( .B(A[132]), .A(S), .Z(O[132]) );
  ANDN U477 ( .B(A[131]), .A(S), .Z(O[131]) );
  ANDN U478 ( .B(A[130]), .A(S), .Z(O[130]) );
  ANDN U479 ( .B(A[12]), .A(S), .Z(O[12]) );
  ANDN U480 ( .B(A[129]), .A(S), .Z(O[129]) );
  ANDN U481 ( .B(A[128]), .A(S), .Z(O[128]) );
  ANDN U482 ( .B(A[127]), .A(S), .Z(O[127]) );
  ANDN U483 ( .B(A[126]), .A(S), .Z(O[126]) );
  ANDN U484 ( .B(A[125]), .A(S), .Z(O[125]) );
  ANDN U485 ( .B(A[124]), .A(S), .Z(O[124]) );
  ANDN U486 ( .B(A[123]), .A(S), .Z(O[123]) );
  ANDN U487 ( .B(A[122]), .A(S), .Z(O[122]) );
  ANDN U488 ( .B(A[121]), .A(S), .Z(O[121]) );
  ANDN U489 ( .B(A[120]), .A(S), .Z(O[120]) );
  ANDN U490 ( .B(A[11]), .A(S), .Z(O[11]) );
  ANDN U491 ( .B(A[119]), .A(S), .Z(O[119]) );
  ANDN U492 ( .B(A[118]), .A(S), .Z(O[118]) );
  ANDN U493 ( .B(A[117]), .A(S), .Z(O[117]) );
  ANDN U494 ( .B(A[116]), .A(S), .Z(O[116]) );
  ANDN U495 ( .B(A[115]), .A(S), .Z(O[115]) );
  ANDN U496 ( .B(A[114]), .A(S), .Z(O[114]) );
  ANDN U497 ( .B(A[113]), .A(S), .Z(O[113]) );
  ANDN U498 ( .B(A[112]), .A(S), .Z(O[112]) );
  ANDN U499 ( .B(A[111]), .A(S), .Z(O[111]) );
  ANDN U500 ( .B(A[110]), .A(S), .Z(O[110]) );
  ANDN U501 ( .B(A[10]), .A(S), .Z(O[10]) );
  ANDN U502 ( .B(A[109]), .A(S), .Z(O[109]) );
  ANDN U503 ( .B(A[108]), .A(S), .Z(O[108]) );
  ANDN U504 ( .B(A[107]), .A(S), .Z(O[107]) );
  ANDN U505 ( .B(A[106]), .A(S), .Z(O[106]) );
  ANDN U506 ( .B(A[105]), .A(S), .Z(O[105]) );
  ANDN U507 ( .B(A[104]), .A(S), .Z(O[104]) );
  ANDN U508 ( .B(A[103]), .A(S), .Z(O[103]) );
  ANDN U509 ( .B(A[102]), .A(S), .Z(O[102]) );
  ANDN U510 ( .B(A[101]), .A(S), .Z(O[101]) );
  ANDN U511 ( .B(A[100]), .A(S), .Z(O[100]) );
  ANDN U512 ( .B(A[0]), .A(S), .Z(O[0]) );
endmodule


module FA_8493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_8494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  ANDN U1 ( .B(CI), .A(S), .Z(CO) );
  XOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_8495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_8999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_9005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XOR U1 ( .A(B), .B(A), .Z(S) );
  AND U2 ( .A(A), .B(B), .Z(CO) );
endmodule


module FA_9006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N514_1_1 ( A, B, CI, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  input CI;
  output CO;

  wire   [513:1] C;

  FA_9006 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(1'b0), .B(B[0]), .CI(1'b0), .S(
        S[0]) );
  FA_9005 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(B[1]), .CI(1'b0), .S(
        S[1]), .CO(C[2]) );
  FA_9004 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_9003 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_9002 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_9001 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_9000 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_8999 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_8998 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_8997 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_8996 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_8995 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_8994 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_8993 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_8992 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_8991 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_8990 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_8989 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_8988 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_8987 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_8986 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_8985 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_8984 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_8983 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_8982 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_8981 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_8980 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_8979 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_8978 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_8977 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_8976 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_8975 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_8974 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_8973 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_8972 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_8971 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_8970 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_8969 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_8968 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_8967 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_8966 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_8965 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_8964 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_8963 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_8962 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_8961 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_8960 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_8959 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_8958 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_8957 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_8956 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_8955 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_8954 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_8953 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_8952 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_8951 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_8950 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_8949 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_8948 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_8947 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_8946 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_8945 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_8944 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_8943 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_8942 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_8941 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_8940 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_8939 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_8938 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_8937 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_8936 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_8935 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_8934 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_8933 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_8932 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_8931 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_8930 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_8929 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_8928 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_8927 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_8926 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_8925 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_8924 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_8923 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_8922 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_8921 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_8920 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_8919 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_8918 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_8917 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_8916 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_8915 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_8914 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_8913 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_8912 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_8911 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_8910 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_8909 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_8908 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_8907 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_8906 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(B[100]), .CI(
        C[100]), .S(S[100]), .CO(C[101]) );
  FA_8905 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(B[101]), .CI(
        C[101]), .S(S[101]), .CO(C[102]) );
  FA_8904 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(B[102]), .CI(
        C[102]), .S(S[102]), .CO(C[103]) );
  FA_8903 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(B[103]), .CI(
        C[103]), .S(S[103]), .CO(C[104]) );
  FA_8902 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(B[104]), .CI(
        C[104]), .S(S[104]), .CO(C[105]) );
  FA_8901 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(B[105]), .CI(
        C[105]), .S(S[105]), .CO(C[106]) );
  FA_8900 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(B[106]), .CI(
        C[106]), .S(S[106]), .CO(C[107]) );
  FA_8899 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(B[107]), .CI(
        C[107]), .S(S[107]), .CO(C[108]) );
  FA_8898 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(B[108]), .CI(
        C[108]), .S(S[108]), .CO(C[109]) );
  FA_8897 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(B[109]), .CI(
        C[109]), .S(S[109]), .CO(C[110]) );
  FA_8896 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(B[110]), .CI(
        C[110]), .S(S[110]), .CO(C[111]) );
  FA_8895 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(B[111]), .CI(
        C[111]), .S(S[111]), .CO(C[112]) );
  FA_8894 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(B[112]), .CI(
        C[112]), .S(S[112]), .CO(C[113]) );
  FA_8893 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(B[113]), .CI(
        C[113]), .S(S[113]), .CO(C[114]) );
  FA_8892 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(B[114]), .CI(
        C[114]), .S(S[114]), .CO(C[115]) );
  FA_8891 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(B[115]), .CI(
        C[115]), .S(S[115]), .CO(C[116]) );
  FA_8890 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(B[116]), .CI(
        C[116]), .S(S[116]), .CO(C[117]) );
  FA_8889 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(B[117]), .CI(
        C[117]), .S(S[117]), .CO(C[118]) );
  FA_8888 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(B[118]), .CI(
        C[118]), .S(S[118]), .CO(C[119]) );
  FA_8887 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(B[119]), .CI(
        C[119]), .S(S[119]), .CO(C[120]) );
  FA_8886 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(B[120]), .CI(
        C[120]), .S(S[120]), .CO(C[121]) );
  FA_8885 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(B[121]), .CI(
        C[121]), .S(S[121]), .CO(C[122]) );
  FA_8884 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(B[122]), .CI(
        C[122]), .S(S[122]), .CO(C[123]) );
  FA_8883 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(B[123]), .CI(
        C[123]), .S(S[123]), .CO(C[124]) );
  FA_8882 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(B[124]), .CI(
        C[124]), .S(S[124]), .CO(C[125]) );
  FA_8881 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(B[125]), .CI(
        C[125]), .S(S[125]), .CO(C[126]) );
  FA_8880 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(B[126]), .CI(
        C[126]), .S(S[126]), .CO(C[127]) );
  FA_8879 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(B[127]), .CI(
        C[127]), .S(S[127]), .CO(C[128]) );
  FA_8878 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(B[128]), .CI(
        C[128]), .S(S[128]), .CO(C[129]) );
  FA_8877 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(B[129]), .CI(
        C[129]), .S(S[129]), .CO(C[130]) );
  FA_8876 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(B[130]), .CI(
        C[130]), .S(S[130]), .CO(C[131]) );
  FA_8875 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(B[131]), .CI(
        C[131]), .S(S[131]), .CO(C[132]) );
  FA_8874 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(B[132]), .CI(
        C[132]), .S(S[132]), .CO(C[133]) );
  FA_8873 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(B[133]), .CI(
        C[133]), .S(S[133]), .CO(C[134]) );
  FA_8872 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(B[134]), .CI(
        C[134]), .S(S[134]), .CO(C[135]) );
  FA_8871 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(B[135]), .CI(
        C[135]), .S(S[135]), .CO(C[136]) );
  FA_8870 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(B[136]), .CI(
        C[136]), .S(S[136]), .CO(C[137]) );
  FA_8869 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(B[137]), .CI(
        C[137]), .S(S[137]), .CO(C[138]) );
  FA_8868 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(B[138]), .CI(
        C[138]), .S(S[138]), .CO(C[139]) );
  FA_8867 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(B[139]), .CI(
        C[139]), .S(S[139]), .CO(C[140]) );
  FA_8866 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(B[140]), .CI(
        C[140]), .S(S[140]), .CO(C[141]) );
  FA_8865 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(B[141]), .CI(
        C[141]), .S(S[141]), .CO(C[142]) );
  FA_8864 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(B[142]), .CI(
        C[142]), .S(S[142]), .CO(C[143]) );
  FA_8863 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(B[143]), .CI(
        C[143]), .S(S[143]), .CO(C[144]) );
  FA_8862 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(B[144]), .CI(
        C[144]), .S(S[144]), .CO(C[145]) );
  FA_8861 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(B[145]), .CI(
        C[145]), .S(S[145]), .CO(C[146]) );
  FA_8860 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(B[146]), .CI(
        C[146]), .S(S[146]), .CO(C[147]) );
  FA_8859 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(B[147]), .CI(
        C[147]), .S(S[147]), .CO(C[148]) );
  FA_8858 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(B[148]), .CI(
        C[148]), .S(S[148]), .CO(C[149]) );
  FA_8857 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(B[149]), .CI(
        C[149]), .S(S[149]), .CO(C[150]) );
  FA_8856 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(B[150]), .CI(
        C[150]), .S(S[150]), .CO(C[151]) );
  FA_8855 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(B[151]), .CI(
        C[151]), .S(S[151]), .CO(C[152]) );
  FA_8854 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(B[152]), .CI(
        C[152]), .S(S[152]), .CO(C[153]) );
  FA_8853 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(B[153]), .CI(
        C[153]), .S(S[153]), .CO(C[154]) );
  FA_8852 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(B[154]), .CI(
        C[154]), .S(S[154]), .CO(C[155]) );
  FA_8851 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(B[155]), .CI(
        C[155]), .S(S[155]), .CO(C[156]) );
  FA_8850 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(B[156]), .CI(
        C[156]), .S(S[156]), .CO(C[157]) );
  FA_8849 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(B[157]), .CI(
        C[157]), .S(S[157]), .CO(C[158]) );
  FA_8848 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(B[158]), .CI(
        C[158]), .S(S[158]), .CO(C[159]) );
  FA_8847 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(B[159]), .CI(
        C[159]), .S(S[159]), .CO(C[160]) );
  FA_8846 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(B[160]), .CI(
        C[160]), .S(S[160]), .CO(C[161]) );
  FA_8845 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(B[161]), .CI(
        C[161]), .S(S[161]), .CO(C[162]) );
  FA_8844 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(B[162]), .CI(
        C[162]), .S(S[162]), .CO(C[163]) );
  FA_8843 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(B[163]), .CI(
        C[163]), .S(S[163]), .CO(C[164]) );
  FA_8842 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(B[164]), .CI(
        C[164]), .S(S[164]), .CO(C[165]) );
  FA_8841 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(B[165]), .CI(
        C[165]), .S(S[165]), .CO(C[166]) );
  FA_8840 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(B[166]), .CI(
        C[166]), .S(S[166]), .CO(C[167]) );
  FA_8839 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(B[167]), .CI(
        C[167]), .S(S[167]), .CO(C[168]) );
  FA_8838 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(B[168]), .CI(
        C[168]), .S(S[168]), .CO(C[169]) );
  FA_8837 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(B[169]), .CI(
        C[169]), .S(S[169]), .CO(C[170]) );
  FA_8836 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(B[170]), .CI(
        C[170]), .S(S[170]), .CO(C[171]) );
  FA_8835 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(B[171]), .CI(
        C[171]), .S(S[171]), .CO(C[172]) );
  FA_8834 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(B[172]), .CI(
        C[172]), .S(S[172]), .CO(C[173]) );
  FA_8833 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(B[173]), .CI(
        C[173]), .S(S[173]), .CO(C[174]) );
  FA_8832 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(B[174]), .CI(
        C[174]), .S(S[174]), .CO(C[175]) );
  FA_8831 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(B[175]), .CI(
        C[175]), .S(S[175]), .CO(C[176]) );
  FA_8830 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(B[176]), .CI(
        C[176]), .S(S[176]), .CO(C[177]) );
  FA_8829 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(B[177]), .CI(
        C[177]), .S(S[177]), .CO(C[178]) );
  FA_8828 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(B[178]), .CI(
        C[178]), .S(S[178]), .CO(C[179]) );
  FA_8827 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(B[179]), .CI(
        C[179]), .S(S[179]), .CO(C[180]) );
  FA_8826 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(B[180]), .CI(
        C[180]), .S(S[180]), .CO(C[181]) );
  FA_8825 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(B[181]), .CI(
        C[181]), .S(S[181]), .CO(C[182]) );
  FA_8824 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(B[182]), .CI(
        C[182]), .S(S[182]), .CO(C[183]) );
  FA_8823 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(B[183]), .CI(
        C[183]), .S(S[183]), .CO(C[184]) );
  FA_8822 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(B[184]), .CI(
        C[184]), .S(S[184]), .CO(C[185]) );
  FA_8821 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(B[185]), .CI(
        C[185]), .S(S[185]), .CO(C[186]) );
  FA_8820 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(B[186]), .CI(
        C[186]), .S(S[186]), .CO(C[187]) );
  FA_8819 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(B[187]), .CI(
        C[187]), .S(S[187]), .CO(C[188]) );
  FA_8818 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(B[188]), .CI(
        C[188]), .S(S[188]), .CO(C[189]) );
  FA_8817 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(B[189]), .CI(
        C[189]), .S(S[189]), .CO(C[190]) );
  FA_8816 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(B[190]), .CI(
        C[190]), .S(S[190]), .CO(C[191]) );
  FA_8815 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(B[191]), .CI(
        C[191]), .S(S[191]), .CO(C[192]) );
  FA_8814 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(B[192]), .CI(
        C[192]), .S(S[192]), .CO(C[193]) );
  FA_8813 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(B[193]), .CI(
        C[193]), .S(S[193]), .CO(C[194]) );
  FA_8812 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(B[194]), .CI(
        C[194]), .S(S[194]), .CO(C[195]) );
  FA_8811 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(B[195]), .CI(
        C[195]), .S(S[195]), .CO(C[196]) );
  FA_8810 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(B[196]), .CI(
        C[196]), .S(S[196]), .CO(C[197]) );
  FA_8809 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(B[197]), .CI(
        C[197]), .S(S[197]), .CO(C[198]) );
  FA_8808 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(B[198]), .CI(
        C[198]), .S(S[198]), .CO(C[199]) );
  FA_8807 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(B[199]), .CI(
        C[199]), .S(S[199]), .CO(C[200]) );
  FA_8806 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(B[200]), .CI(
        C[200]), .S(S[200]), .CO(C[201]) );
  FA_8805 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(B[201]), .CI(
        C[201]), .S(S[201]), .CO(C[202]) );
  FA_8804 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(B[202]), .CI(
        C[202]), .S(S[202]), .CO(C[203]) );
  FA_8803 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(B[203]), .CI(
        C[203]), .S(S[203]), .CO(C[204]) );
  FA_8802 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(B[204]), .CI(
        C[204]), .S(S[204]), .CO(C[205]) );
  FA_8801 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(B[205]), .CI(
        C[205]), .S(S[205]), .CO(C[206]) );
  FA_8800 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(B[206]), .CI(
        C[206]), .S(S[206]), .CO(C[207]) );
  FA_8799 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(B[207]), .CI(
        C[207]), .S(S[207]), .CO(C[208]) );
  FA_8798 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(B[208]), .CI(
        C[208]), .S(S[208]), .CO(C[209]) );
  FA_8797 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(B[209]), .CI(
        C[209]), .S(S[209]), .CO(C[210]) );
  FA_8796 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(B[210]), .CI(
        C[210]), .S(S[210]), .CO(C[211]) );
  FA_8795 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(B[211]), .CI(
        C[211]), .S(S[211]), .CO(C[212]) );
  FA_8794 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(B[212]), .CI(
        C[212]), .S(S[212]), .CO(C[213]) );
  FA_8793 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(B[213]), .CI(
        C[213]), .S(S[213]), .CO(C[214]) );
  FA_8792 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(B[214]), .CI(
        C[214]), .S(S[214]), .CO(C[215]) );
  FA_8791 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(B[215]), .CI(
        C[215]), .S(S[215]), .CO(C[216]) );
  FA_8790 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(B[216]), .CI(
        C[216]), .S(S[216]), .CO(C[217]) );
  FA_8789 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(B[217]), .CI(
        C[217]), .S(S[217]), .CO(C[218]) );
  FA_8788 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(B[218]), .CI(
        C[218]), .S(S[218]), .CO(C[219]) );
  FA_8787 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(B[219]), .CI(
        C[219]), .S(S[219]), .CO(C[220]) );
  FA_8786 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(B[220]), .CI(
        C[220]), .S(S[220]), .CO(C[221]) );
  FA_8785 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(B[221]), .CI(
        C[221]), .S(S[221]), .CO(C[222]) );
  FA_8784 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(B[222]), .CI(
        C[222]), .S(S[222]), .CO(C[223]) );
  FA_8783 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(B[223]), .CI(
        C[223]), .S(S[223]), .CO(C[224]) );
  FA_8782 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(B[224]), .CI(
        C[224]), .S(S[224]), .CO(C[225]) );
  FA_8781 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(B[225]), .CI(
        C[225]), .S(S[225]), .CO(C[226]) );
  FA_8780 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(B[226]), .CI(
        C[226]), .S(S[226]), .CO(C[227]) );
  FA_8779 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(B[227]), .CI(
        C[227]), .S(S[227]), .CO(C[228]) );
  FA_8778 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(B[228]), .CI(
        C[228]), .S(S[228]), .CO(C[229]) );
  FA_8777 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(B[229]), .CI(
        C[229]), .S(S[229]), .CO(C[230]) );
  FA_8776 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(B[230]), .CI(
        C[230]), .S(S[230]), .CO(C[231]) );
  FA_8775 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(B[231]), .CI(
        C[231]), .S(S[231]), .CO(C[232]) );
  FA_8774 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(B[232]), .CI(
        C[232]), .S(S[232]), .CO(C[233]) );
  FA_8773 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(B[233]), .CI(
        C[233]), .S(S[233]), .CO(C[234]) );
  FA_8772 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(B[234]), .CI(
        C[234]), .S(S[234]), .CO(C[235]) );
  FA_8771 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(B[235]), .CI(
        C[235]), .S(S[235]), .CO(C[236]) );
  FA_8770 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(B[236]), .CI(
        C[236]), .S(S[236]), .CO(C[237]) );
  FA_8769 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(B[237]), .CI(
        C[237]), .S(S[237]), .CO(C[238]) );
  FA_8768 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(B[238]), .CI(
        C[238]), .S(S[238]), .CO(C[239]) );
  FA_8767 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(B[239]), .CI(
        C[239]), .S(S[239]), .CO(C[240]) );
  FA_8766 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(B[240]), .CI(
        C[240]), .S(S[240]), .CO(C[241]) );
  FA_8765 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(B[241]), .CI(
        C[241]), .S(S[241]), .CO(C[242]) );
  FA_8764 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(B[242]), .CI(
        C[242]), .S(S[242]), .CO(C[243]) );
  FA_8763 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(B[243]), .CI(
        C[243]), .S(S[243]), .CO(C[244]) );
  FA_8762 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(B[244]), .CI(
        C[244]), .S(S[244]), .CO(C[245]) );
  FA_8761 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(B[245]), .CI(
        C[245]), .S(S[245]), .CO(C[246]) );
  FA_8760 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(B[246]), .CI(
        C[246]), .S(S[246]), .CO(C[247]) );
  FA_8759 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(B[247]), .CI(
        C[247]), .S(S[247]), .CO(C[248]) );
  FA_8758 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(B[248]), .CI(
        C[248]), .S(S[248]), .CO(C[249]) );
  FA_8757 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(B[249]), .CI(
        C[249]), .S(S[249]), .CO(C[250]) );
  FA_8756 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(B[250]), .CI(
        C[250]), .S(S[250]), .CO(C[251]) );
  FA_8755 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(B[251]), .CI(
        C[251]), .S(S[251]), .CO(C[252]) );
  FA_8754 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(B[252]), .CI(
        C[252]), .S(S[252]), .CO(C[253]) );
  FA_8753 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(B[253]), .CI(
        C[253]), .S(S[253]), .CO(C[254]) );
  FA_8752 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(B[254]), .CI(
        C[254]), .S(S[254]), .CO(C[255]) );
  FA_8751 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(B[255]), .CI(
        C[255]), .S(S[255]), .CO(C[256]) );
  FA_8750 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(B[256]), .CI(
        C[256]), .S(S[256]), .CO(C[257]) );
  FA_8749 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(B[257]), .CI(
        C[257]), .S(S[257]), .CO(C[258]) );
  FA_8748 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(B[258]), .CI(
        C[258]), .S(S[258]), .CO(C[259]) );
  FA_8747 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(B[259]), .CI(
        C[259]), .S(S[259]), .CO(C[260]) );
  FA_8746 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(B[260]), .CI(
        C[260]), .S(S[260]), .CO(C[261]) );
  FA_8745 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(B[261]), .CI(
        C[261]), .S(S[261]), .CO(C[262]) );
  FA_8744 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(B[262]), .CI(
        C[262]), .S(S[262]), .CO(C[263]) );
  FA_8743 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(B[263]), .CI(
        C[263]), .S(S[263]), .CO(C[264]) );
  FA_8742 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(B[264]), .CI(
        C[264]), .S(S[264]), .CO(C[265]) );
  FA_8741 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(B[265]), .CI(
        C[265]), .S(S[265]), .CO(C[266]) );
  FA_8740 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(B[266]), .CI(
        C[266]), .S(S[266]), .CO(C[267]) );
  FA_8739 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(B[267]), .CI(
        C[267]), .S(S[267]), .CO(C[268]) );
  FA_8738 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(B[268]), .CI(
        C[268]), .S(S[268]), .CO(C[269]) );
  FA_8737 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(B[269]), .CI(
        C[269]), .S(S[269]), .CO(C[270]) );
  FA_8736 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(B[270]), .CI(
        C[270]), .S(S[270]), .CO(C[271]) );
  FA_8735 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(B[271]), .CI(
        C[271]), .S(S[271]), .CO(C[272]) );
  FA_8734 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(B[272]), .CI(
        C[272]), .S(S[272]), .CO(C[273]) );
  FA_8733 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(B[273]), .CI(
        C[273]), .S(S[273]), .CO(C[274]) );
  FA_8732 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(B[274]), .CI(
        C[274]), .S(S[274]), .CO(C[275]) );
  FA_8731 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(B[275]), .CI(
        C[275]), .S(S[275]), .CO(C[276]) );
  FA_8730 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(B[276]), .CI(
        C[276]), .S(S[276]), .CO(C[277]) );
  FA_8729 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(B[277]), .CI(
        C[277]), .S(S[277]), .CO(C[278]) );
  FA_8728 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(B[278]), .CI(
        C[278]), .S(S[278]), .CO(C[279]) );
  FA_8727 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(B[279]), .CI(
        C[279]), .S(S[279]), .CO(C[280]) );
  FA_8726 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(B[280]), .CI(
        C[280]), .S(S[280]), .CO(C[281]) );
  FA_8725 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(B[281]), .CI(
        C[281]), .S(S[281]), .CO(C[282]) );
  FA_8724 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(B[282]), .CI(
        C[282]), .S(S[282]), .CO(C[283]) );
  FA_8723 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(B[283]), .CI(
        C[283]), .S(S[283]), .CO(C[284]) );
  FA_8722 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(B[284]), .CI(
        C[284]), .S(S[284]), .CO(C[285]) );
  FA_8721 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(B[285]), .CI(
        C[285]), .S(S[285]), .CO(C[286]) );
  FA_8720 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(B[286]), .CI(
        C[286]), .S(S[286]), .CO(C[287]) );
  FA_8719 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(B[287]), .CI(
        C[287]), .S(S[287]), .CO(C[288]) );
  FA_8718 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(B[288]), .CI(
        C[288]), .S(S[288]), .CO(C[289]) );
  FA_8717 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(B[289]), .CI(
        C[289]), .S(S[289]), .CO(C[290]) );
  FA_8716 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(B[290]), .CI(
        C[290]), .S(S[290]), .CO(C[291]) );
  FA_8715 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(B[291]), .CI(
        C[291]), .S(S[291]), .CO(C[292]) );
  FA_8714 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(B[292]), .CI(
        C[292]), .S(S[292]), .CO(C[293]) );
  FA_8713 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(B[293]), .CI(
        C[293]), .S(S[293]), .CO(C[294]) );
  FA_8712 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(B[294]), .CI(
        C[294]), .S(S[294]), .CO(C[295]) );
  FA_8711 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(B[295]), .CI(
        C[295]), .S(S[295]), .CO(C[296]) );
  FA_8710 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(B[296]), .CI(
        C[296]), .S(S[296]), .CO(C[297]) );
  FA_8709 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(B[297]), .CI(
        C[297]), .S(S[297]), .CO(C[298]) );
  FA_8708 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(B[298]), .CI(
        C[298]), .S(S[298]), .CO(C[299]) );
  FA_8707 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(B[299]), .CI(
        C[299]), .S(S[299]), .CO(C[300]) );
  FA_8706 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(B[300]), .CI(
        C[300]), .S(S[300]), .CO(C[301]) );
  FA_8705 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(B[301]), .CI(
        C[301]), .S(S[301]), .CO(C[302]) );
  FA_8704 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(B[302]), .CI(
        C[302]), .S(S[302]), .CO(C[303]) );
  FA_8703 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(B[303]), .CI(
        C[303]), .S(S[303]), .CO(C[304]) );
  FA_8702 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(B[304]), .CI(
        C[304]), .S(S[304]), .CO(C[305]) );
  FA_8701 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(B[305]), .CI(
        C[305]), .S(S[305]), .CO(C[306]) );
  FA_8700 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(B[306]), .CI(
        C[306]), .S(S[306]), .CO(C[307]) );
  FA_8699 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(B[307]), .CI(
        C[307]), .S(S[307]), .CO(C[308]) );
  FA_8698 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(B[308]), .CI(
        C[308]), .S(S[308]), .CO(C[309]) );
  FA_8697 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(B[309]), .CI(
        C[309]), .S(S[309]), .CO(C[310]) );
  FA_8696 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(B[310]), .CI(
        C[310]), .S(S[310]), .CO(C[311]) );
  FA_8695 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(B[311]), .CI(
        C[311]), .S(S[311]), .CO(C[312]) );
  FA_8694 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(B[312]), .CI(
        C[312]), .S(S[312]), .CO(C[313]) );
  FA_8693 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(B[313]), .CI(
        C[313]), .S(S[313]), .CO(C[314]) );
  FA_8692 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(B[314]), .CI(
        C[314]), .S(S[314]), .CO(C[315]) );
  FA_8691 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(B[315]), .CI(
        C[315]), .S(S[315]), .CO(C[316]) );
  FA_8690 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(B[316]), .CI(
        C[316]), .S(S[316]), .CO(C[317]) );
  FA_8689 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(B[317]), .CI(
        C[317]), .S(S[317]), .CO(C[318]) );
  FA_8688 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(B[318]), .CI(
        C[318]), .S(S[318]), .CO(C[319]) );
  FA_8687 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(B[319]), .CI(
        C[319]), .S(S[319]), .CO(C[320]) );
  FA_8686 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(B[320]), .CI(
        C[320]), .S(S[320]), .CO(C[321]) );
  FA_8685 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(B[321]), .CI(
        C[321]), .S(S[321]), .CO(C[322]) );
  FA_8684 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(B[322]), .CI(
        C[322]), .S(S[322]), .CO(C[323]) );
  FA_8683 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(B[323]), .CI(
        C[323]), .S(S[323]), .CO(C[324]) );
  FA_8682 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(B[324]), .CI(
        C[324]), .S(S[324]), .CO(C[325]) );
  FA_8681 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(B[325]), .CI(
        C[325]), .S(S[325]), .CO(C[326]) );
  FA_8680 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(B[326]), .CI(
        C[326]), .S(S[326]), .CO(C[327]) );
  FA_8679 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(B[327]), .CI(
        C[327]), .S(S[327]), .CO(C[328]) );
  FA_8678 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(B[328]), .CI(
        C[328]), .S(S[328]), .CO(C[329]) );
  FA_8677 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(B[329]), .CI(
        C[329]), .S(S[329]), .CO(C[330]) );
  FA_8676 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(B[330]), .CI(
        C[330]), .S(S[330]), .CO(C[331]) );
  FA_8675 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(B[331]), .CI(
        C[331]), .S(S[331]), .CO(C[332]) );
  FA_8674 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(B[332]), .CI(
        C[332]), .S(S[332]), .CO(C[333]) );
  FA_8673 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(B[333]), .CI(
        C[333]), .S(S[333]), .CO(C[334]) );
  FA_8672 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(B[334]), .CI(
        C[334]), .S(S[334]), .CO(C[335]) );
  FA_8671 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(B[335]), .CI(
        C[335]), .S(S[335]), .CO(C[336]) );
  FA_8670 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(B[336]), .CI(
        C[336]), .S(S[336]), .CO(C[337]) );
  FA_8669 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(B[337]), .CI(
        C[337]), .S(S[337]), .CO(C[338]) );
  FA_8668 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(B[338]), .CI(
        C[338]), .S(S[338]), .CO(C[339]) );
  FA_8667 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(B[339]), .CI(
        C[339]), .S(S[339]), .CO(C[340]) );
  FA_8666 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(B[340]), .CI(
        C[340]), .S(S[340]), .CO(C[341]) );
  FA_8665 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(B[341]), .CI(
        C[341]), .S(S[341]), .CO(C[342]) );
  FA_8664 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(B[342]), .CI(
        C[342]), .S(S[342]), .CO(C[343]) );
  FA_8663 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(B[343]), .CI(
        C[343]), .S(S[343]), .CO(C[344]) );
  FA_8662 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(B[344]), .CI(
        C[344]), .S(S[344]), .CO(C[345]) );
  FA_8661 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(B[345]), .CI(
        C[345]), .S(S[345]), .CO(C[346]) );
  FA_8660 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(B[346]), .CI(
        C[346]), .S(S[346]), .CO(C[347]) );
  FA_8659 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(B[347]), .CI(
        C[347]), .S(S[347]), .CO(C[348]) );
  FA_8658 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(B[348]), .CI(
        C[348]), .S(S[348]), .CO(C[349]) );
  FA_8657 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(B[349]), .CI(
        C[349]), .S(S[349]), .CO(C[350]) );
  FA_8656 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(B[350]), .CI(
        C[350]), .S(S[350]), .CO(C[351]) );
  FA_8655 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(B[351]), .CI(
        C[351]), .S(S[351]), .CO(C[352]) );
  FA_8654 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(B[352]), .CI(
        C[352]), .S(S[352]), .CO(C[353]) );
  FA_8653 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(B[353]), .CI(
        C[353]), .S(S[353]), .CO(C[354]) );
  FA_8652 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(B[354]), .CI(
        C[354]), .S(S[354]), .CO(C[355]) );
  FA_8651 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(B[355]), .CI(
        C[355]), .S(S[355]), .CO(C[356]) );
  FA_8650 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(B[356]), .CI(
        C[356]), .S(S[356]), .CO(C[357]) );
  FA_8649 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(B[357]), .CI(
        C[357]), .S(S[357]), .CO(C[358]) );
  FA_8648 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(B[358]), .CI(
        C[358]), .S(S[358]), .CO(C[359]) );
  FA_8647 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(B[359]), .CI(
        C[359]), .S(S[359]), .CO(C[360]) );
  FA_8646 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(B[360]), .CI(
        C[360]), .S(S[360]), .CO(C[361]) );
  FA_8645 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(B[361]), .CI(
        C[361]), .S(S[361]), .CO(C[362]) );
  FA_8644 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(B[362]), .CI(
        C[362]), .S(S[362]), .CO(C[363]) );
  FA_8643 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(B[363]), .CI(
        C[363]), .S(S[363]), .CO(C[364]) );
  FA_8642 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(B[364]), .CI(
        C[364]), .S(S[364]), .CO(C[365]) );
  FA_8641 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(B[365]), .CI(
        C[365]), .S(S[365]), .CO(C[366]) );
  FA_8640 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(B[366]), .CI(
        C[366]), .S(S[366]), .CO(C[367]) );
  FA_8639 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(B[367]), .CI(
        C[367]), .S(S[367]), .CO(C[368]) );
  FA_8638 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(B[368]), .CI(
        C[368]), .S(S[368]), .CO(C[369]) );
  FA_8637 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(B[369]), .CI(
        C[369]), .S(S[369]), .CO(C[370]) );
  FA_8636 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(B[370]), .CI(
        C[370]), .S(S[370]), .CO(C[371]) );
  FA_8635 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(B[371]), .CI(
        C[371]), .S(S[371]), .CO(C[372]) );
  FA_8634 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(B[372]), .CI(
        C[372]), .S(S[372]), .CO(C[373]) );
  FA_8633 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(B[373]), .CI(
        C[373]), .S(S[373]), .CO(C[374]) );
  FA_8632 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(B[374]), .CI(
        C[374]), .S(S[374]), .CO(C[375]) );
  FA_8631 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(B[375]), .CI(
        C[375]), .S(S[375]), .CO(C[376]) );
  FA_8630 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(B[376]), .CI(
        C[376]), .S(S[376]), .CO(C[377]) );
  FA_8629 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(B[377]), .CI(
        C[377]), .S(S[377]), .CO(C[378]) );
  FA_8628 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(B[378]), .CI(
        C[378]), .S(S[378]), .CO(C[379]) );
  FA_8627 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(B[379]), .CI(
        C[379]), .S(S[379]), .CO(C[380]) );
  FA_8626 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(B[380]), .CI(
        C[380]), .S(S[380]), .CO(C[381]) );
  FA_8625 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(B[381]), .CI(
        C[381]), .S(S[381]), .CO(C[382]) );
  FA_8624 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(B[382]), .CI(
        C[382]), .S(S[382]), .CO(C[383]) );
  FA_8623 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(B[383]), .CI(
        C[383]), .S(S[383]), .CO(C[384]) );
  FA_8622 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(B[384]), .CI(
        C[384]), .S(S[384]), .CO(C[385]) );
  FA_8621 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(B[385]), .CI(
        C[385]), .S(S[385]), .CO(C[386]) );
  FA_8620 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(B[386]), .CI(
        C[386]), .S(S[386]), .CO(C[387]) );
  FA_8619 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(B[387]), .CI(
        C[387]), .S(S[387]), .CO(C[388]) );
  FA_8618 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(B[388]), .CI(
        C[388]), .S(S[388]), .CO(C[389]) );
  FA_8617 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(B[389]), .CI(
        C[389]), .S(S[389]), .CO(C[390]) );
  FA_8616 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(B[390]), .CI(
        C[390]), .S(S[390]), .CO(C[391]) );
  FA_8615 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(B[391]), .CI(
        C[391]), .S(S[391]), .CO(C[392]) );
  FA_8614 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(B[392]), .CI(
        C[392]), .S(S[392]), .CO(C[393]) );
  FA_8613 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(B[393]), .CI(
        C[393]), .S(S[393]), .CO(C[394]) );
  FA_8612 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(B[394]), .CI(
        C[394]), .S(S[394]), .CO(C[395]) );
  FA_8611 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(B[395]), .CI(
        C[395]), .S(S[395]), .CO(C[396]) );
  FA_8610 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(B[396]), .CI(
        C[396]), .S(S[396]), .CO(C[397]) );
  FA_8609 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(B[397]), .CI(
        C[397]), .S(S[397]), .CO(C[398]) );
  FA_8608 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(B[398]), .CI(
        C[398]), .S(S[398]), .CO(C[399]) );
  FA_8607 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(B[399]), .CI(
        C[399]), .S(S[399]), .CO(C[400]) );
  FA_8606 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(B[400]), .CI(
        C[400]), .S(S[400]), .CO(C[401]) );
  FA_8605 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(B[401]), .CI(
        C[401]), .S(S[401]), .CO(C[402]) );
  FA_8604 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(B[402]), .CI(
        C[402]), .S(S[402]), .CO(C[403]) );
  FA_8603 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(B[403]), .CI(
        C[403]), .S(S[403]), .CO(C[404]) );
  FA_8602 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(B[404]), .CI(
        C[404]), .S(S[404]), .CO(C[405]) );
  FA_8601 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(B[405]), .CI(
        C[405]), .S(S[405]), .CO(C[406]) );
  FA_8600 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(B[406]), .CI(
        C[406]), .S(S[406]), .CO(C[407]) );
  FA_8599 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(B[407]), .CI(
        C[407]), .S(S[407]), .CO(C[408]) );
  FA_8598 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(B[408]), .CI(
        C[408]), .S(S[408]), .CO(C[409]) );
  FA_8597 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(B[409]), .CI(
        C[409]), .S(S[409]), .CO(C[410]) );
  FA_8596 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(B[410]), .CI(
        C[410]), .S(S[410]), .CO(C[411]) );
  FA_8595 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(B[411]), .CI(
        C[411]), .S(S[411]), .CO(C[412]) );
  FA_8594 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(B[412]), .CI(
        C[412]), .S(S[412]), .CO(C[413]) );
  FA_8593 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(B[413]), .CI(
        C[413]), .S(S[413]), .CO(C[414]) );
  FA_8592 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(B[414]), .CI(
        C[414]), .S(S[414]), .CO(C[415]) );
  FA_8591 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(B[415]), .CI(
        C[415]), .S(S[415]), .CO(C[416]) );
  FA_8590 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(B[416]), .CI(
        C[416]), .S(S[416]), .CO(C[417]) );
  FA_8589 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(B[417]), .CI(
        C[417]), .S(S[417]), .CO(C[418]) );
  FA_8588 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(B[418]), .CI(
        C[418]), .S(S[418]), .CO(C[419]) );
  FA_8587 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(B[419]), .CI(
        C[419]), .S(S[419]), .CO(C[420]) );
  FA_8586 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(B[420]), .CI(
        C[420]), .S(S[420]), .CO(C[421]) );
  FA_8585 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(B[421]), .CI(
        C[421]), .S(S[421]), .CO(C[422]) );
  FA_8584 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(B[422]), .CI(
        C[422]), .S(S[422]), .CO(C[423]) );
  FA_8583 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(B[423]), .CI(
        C[423]), .S(S[423]), .CO(C[424]) );
  FA_8582 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(B[424]), .CI(
        C[424]), .S(S[424]), .CO(C[425]) );
  FA_8581 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(B[425]), .CI(
        C[425]), .S(S[425]), .CO(C[426]) );
  FA_8580 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(B[426]), .CI(
        C[426]), .S(S[426]), .CO(C[427]) );
  FA_8579 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(B[427]), .CI(
        C[427]), .S(S[427]), .CO(C[428]) );
  FA_8578 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(B[428]), .CI(
        C[428]), .S(S[428]), .CO(C[429]) );
  FA_8577 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(B[429]), .CI(
        C[429]), .S(S[429]), .CO(C[430]) );
  FA_8576 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(B[430]), .CI(
        C[430]), .S(S[430]), .CO(C[431]) );
  FA_8575 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(B[431]), .CI(
        C[431]), .S(S[431]), .CO(C[432]) );
  FA_8574 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(B[432]), .CI(
        C[432]), .S(S[432]), .CO(C[433]) );
  FA_8573 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(B[433]), .CI(
        C[433]), .S(S[433]), .CO(C[434]) );
  FA_8572 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(B[434]), .CI(
        C[434]), .S(S[434]), .CO(C[435]) );
  FA_8571 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(B[435]), .CI(
        C[435]), .S(S[435]), .CO(C[436]) );
  FA_8570 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(B[436]), .CI(
        C[436]), .S(S[436]), .CO(C[437]) );
  FA_8569 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(B[437]), .CI(
        C[437]), .S(S[437]), .CO(C[438]) );
  FA_8568 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(B[438]), .CI(
        C[438]), .S(S[438]), .CO(C[439]) );
  FA_8567 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(B[439]), .CI(
        C[439]), .S(S[439]), .CO(C[440]) );
  FA_8566 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(B[440]), .CI(
        C[440]), .S(S[440]), .CO(C[441]) );
  FA_8565 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(B[441]), .CI(
        C[441]), .S(S[441]), .CO(C[442]) );
  FA_8564 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(B[442]), .CI(
        C[442]), .S(S[442]), .CO(C[443]) );
  FA_8563 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(B[443]), .CI(
        C[443]), .S(S[443]), .CO(C[444]) );
  FA_8562 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(B[444]), .CI(
        C[444]), .S(S[444]), .CO(C[445]) );
  FA_8561 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(B[445]), .CI(
        C[445]), .S(S[445]), .CO(C[446]) );
  FA_8560 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(B[446]), .CI(
        C[446]), .S(S[446]), .CO(C[447]) );
  FA_8559 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(B[447]), .CI(
        C[447]), .S(S[447]), .CO(C[448]) );
  FA_8558 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(B[448]), .CI(
        C[448]), .S(S[448]), .CO(C[449]) );
  FA_8557 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(B[449]), .CI(
        C[449]), .S(S[449]), .CO(C[450]) );
  FA_8556 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(B[450]), .CI(
        C[450]), .S(S[450]), .CO(C[451]) );
  FA_8555 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(B[451]), .CI(
        C[451]), .S(S[451]), .CO(C[452]) );
  FA_8554 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(B[452]), .CI(
        C[452]), .S(S[452]), .CO(C[453]) );
  FA_8553 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(B[453]), .CI(
        C[453]), .S(S[453]), .CO(C[454]) );
  FA_8552 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(B[454]), .CI(
        C[454]), .S(S[454]), .CO(C[455]) );
  FA_8551 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(B[455]), .CI(
        C[455]), .S(S[455]), .CO(C[456]) );
  FA_8550 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(B[456]), .CI(
        C[456]), .S(S[456]), .CO(C[457]) );
  FA_8549 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(B[457]), .CI(
        C[457]), .S(S[457]), .CO(C[458]) );
  FA_8548 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(B[458]), .CI(
        C[458]), .S(S[458]), .CO(C[459]) );
  FA_8547 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(B[459]), .CI(
        C[459]), .S(S[459]), .CO(C[460]) );
  FA_8546 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(B[460]), .CI(
        C[460]), .S(S[460]), .CO(C[461]) );
  FA_8545 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(B[461]), .CI(
        C[461]), .S(S[461]), .CO(C[462]) );
  FA_8544 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(B[462]), .CI(
        C[462]), .S(S[462]), .CO(C[463]) );
  FA_8543 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(B[463]), .CI(
        C[463]), .S(S[463]), .CO(C[464]) );
  FA_8542 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(B[464]), .CI(
        C[464]), .S(S[464]), .CO(C[465]) );
  FA_8541 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(B[465]), .CI(
        C[465]), .S(S[465]), .CO(C[466]) );
  FA_8540 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(B[466]), .CI(
        C[466]), .S(S[466]), .CO(C[467]) );
  FA_8539 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(B[467]), .CI(
        C[467]), .S(S[467]), .CO(C[468]) );
  FA_8538 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(B[468]), .CI(
        C[468]), .S(S[468]), .CO(C[469]) );
  FA_8537 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(B[469]), .CI(
        C[469]), .S(S[469]), .CO(C[470]) );
  FA_8536 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(B[470]), .CI(
        C[470]), .S(S[470]), .CO(C[471]) );
  FA_8535 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(B[471]), .CI(
        C[471]), .S(S[471]), .CO(C[472]) );
  FA_8534 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(B[472]), .CI(
        C[472]), .S(S[472]), .CO(C[473]) );
  FA_8533 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(B[473]), .CI(
        C[473]), .S(S[473]), .CO(C[474]) );
  FA_8532 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(B[474]), .CI(
        C[474]), .S(S[474]), .CO(C[475]) );
  FA_8531 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(B[475]), .CI(
        C[475]), .S(S[475]), .CO(C[476]) );
  FA_8530 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(B[476]), .CI(
        C[476]), .S(S[476]), .CO(C[477]) );
  FA_8529 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(B[477]), .CI(
        C[477]), .S(S[477]), .CO(C[478]) );
  FA_8528 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(B[478]), .CI(
        C[478]), .S(S[478]), .CO(C[479]) );
  FA_8527 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(B[479]), .CI(
        C[479]), .S(S[479]), .CO(C[480]) );
  FA_8526 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(B[480]), .CI(
        C[480]), .S(S[480]), .CO(C[481]) );
  FA_8525 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(B[481]), .CI(
        C[481]), .S(S[481]), .CO(C[482]) );
  FA_8524 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(B[482]), .CI(
        C[482]), .S(S[482]), .CO(C[483]) );
  FA_8523 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(B[483]), .CI(
        C[483]), .S(S[483]), .CO(C[484]) );
  FA_8522 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(B[484]), .CI(
        C[484]), .S(S[484]), .CO(C[485]) );
  FA_8521 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(B[485]), .CI(
        C[485]), .S(S[485]), .CO(C[486]) );
  FA_8520 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(B[486]), .CI(
        C[486]), .S(S[486]), .CO(C[487]) );
  FA_8519 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(B[487]), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_8518 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(B[488]), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_8517 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(B[489]), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_8516 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(B[490]), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_8515 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(B[491]), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_8514 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(B[492]), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_8513 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(B[493]), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_8512 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(B[494]), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_8511 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(B[495]), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_8510 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(B[496]), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_8509 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(B[497]), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_8508 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(B[498]), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_8507 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(B[499]), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_8506 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(B[500]), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_8505 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(B[501]), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_8504 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(B[502]), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_8503 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(B[503]), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_8502 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(B[504]), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_8501 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(B[505]), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_8500 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(B[506]), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_8499 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(B[507]), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_8498 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(B[508]), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_8497 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(B[509]), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_8496 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(B[510]), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_8495 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(B[511]), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_8494 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b0), .CI(C[512]), .S(S[512]), 
        .CO(C[513]) );
  FA_8493 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b0), .CI(C[513]), .S(S[513])
         );
endmodule


module FA_6951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_6952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(CI), .B(B), .Z(CO) );
endmodule


module FA_6953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_6999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N514_3 ( A, B, O );
  input [513:0] A;
  input [513:0] B;
  output O;
  wire   n516, n517, n518, n519, n520, n521, n522, n523, n524, n525, n526,
         n527, n528, n529, n530, n531, n532, n533, n534, n535, n536, n537,
         n538, n539, n540, n541, n542, n543, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
         n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570,
         n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, n581,
         n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592,
         n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
         n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614,
         n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
         n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636,
         n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647,
         n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
         n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669,
         n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
         n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
         n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702,
         n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713,
         n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
         n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735,
         n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
         n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
         n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768,
         n769, n770, n771, n772, n773, n774, n775, n776, n777, n778, n779,
         n780, n781, n782, n783, n784, n785, n786, n787, n788, n789, n790,
         n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
         n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812,
         n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, n823,
         n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834,
         n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845,
         n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
         n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867,
         n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
         n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889,
         n890, n891, n892, n893, n894, n895, n896, n897, n898, n899, n900,
         n901, n902, n903, n904, n905, n906, n907, n908, n909, n910, n911,
         n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
         n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n933,
         n934, n935, n936, n937, n938, n939, n940, n941, n942, n943, n944,
         n945, n946, n947, n948, n949, n950, n951, n952, n953, n954, n955,
         n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, n966,
         n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
         n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
         n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
         n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
         n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
         n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029;
  wire   [513:1] C;

  FA_7464 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n516), .CI(1'b1), 
        .CO(C[1]) );
  FA_7463 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n517), .CI(C[1]), 
        .CO(C[2]) );
  FA_7462 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n518), .CI(C[2]), 
        .CO(C[3]) );
  FA_7461 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n519), .CI(C[3]), 
        .CO(C[4]) );
  FA_7460 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n520), .CI(C[4]), 
        .CO(C[5]) );
  FA_7459 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n521), .CI(C[5]), 
        .CO(C[6]) );
  FA_7458 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n522), .CI(C[6]), 
        .CO(C[7]) );
  FA_7457 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n523), .CI(C[7]), 
        .CO(C[8]) );
  FA_7456 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n524), .CI(C[8]), 
        .CO(C[9]) );
  FA_7455 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n525), .CI(C[9]), 
        .CO(C[10]) );
  FA_7454 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n526), .CI(C[10]), 
        .CO(C[11]) );
  FA_7453 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n527), .CI(C[11]), 
        .CO(C[12]) );
  FA_7452 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n528), .CI(C[12]), 
        .CO(C[13]) );
  FA_7451 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n529), .CI(C[13]), 
        .CO(C[14]) );
  FA_7450 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n530), .CI(C[14]), 
        .CO(C[15]) );
  FA_7449 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n531), .CI(C[15]), 
        .CO(C[16]) );
  FA_7448 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n532), .CI(C[16]), 
        .CO(C[17]) );
  FA_7447 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n533), .CI(C[17]), 
        .CO(C[18]) );
  FA_7446 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n534), .CI(C[18]), 
        .CO(C[19]) );
  FA_7445 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n535), .CI(C[19]), 
        .CO(C[20]) );
  FA_7444 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n536), .CI(C[20]), 
        .CO(C[21]) );
  FA_7443 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n537), .CI(C[21]), 
        .CO(C[22]) );
  FA_7442 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n538), .CI(C[22]), 
        .CO(C[23]) );
  FA_7441 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n539), .CI(C[23]), 
        .CO(C[24]) );
  FA_7440 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n540), .CI(C[24]), 
        .CO(C[25]) );
  FA_7439 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n541), .CI(C[25]), 
        .CO(C[26]) );
  FA_7438 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n542), .CI(C[26]), 
        .CO(C[27]) );
  FA_7437 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n543), .CI(C[27]), 
        .CO(C[28]) );
  FA_7436 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n544), .CI(C[28]), 
        .CO(C[29]) );
  FA_7435 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n545), .CI(C[29]), 
        .CO(C[30]) );
  FA_7434 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n546), .CI(C[30]), 
        .CO(C[31]) );
  FA_7433 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n547), .CI(C[31]), 
        .CO(C[32]) );
  FA_7432 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n548), .CI(C[32]), 
        .CO(C[33]) );
  FA_7431 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n549), .CI(C[33]), 
        .CO(C[34]) );
  FA_7430 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n550), .CI(C[34]), 
        .CO(C[35]) );
  FA_7429 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n551), .CI(C[35]), 
        .CO(C[36]) );
  FA_7428 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n552), .CI(C[36]), 
        .CO(C[37]) );
  FA_7427 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n553), .CI(C[37]), 
        .CO(C[38]) );
  FA_7426 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n554), .CI(C[38]), 
        .CO(C[39]) );
  FA_7425 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n555), .CI(C[39]), 
        .CO(C[40]) );
  FA_7424 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n556), .CI(C[40]), 
        .CO(C[41]) );
  FA_7423 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n557), .CI(C[41]), 
        .CO(C[42]) );
  FA_7422 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n558), .CI(C[42]), 
        .CO(C[43]) );
  FA_7421 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n559), .CI(C[43]), 
        .CO(C[44]) );
  FA_7420 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n560), .CI(C[44]), 
        .CO(C[45]) );
  FA_7419 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n561), .CI(C[45]), 
        .CO(C[46]) );
  FA_7418 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n562), .CI(C[46]), 
        .CO(C[47]) );
  FA_7417 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n563), .CI(C[47]), 
        .CO(C[48]) );
  FA_7416 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n564), .CI(C[48]), 
        .CO(C[49]) );
  FA_7415 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n565), .CI(C[49]), 
        .CO(C[50]) );
  FA_7414 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n566), .CI(C[50]), 
        .CO(C[51]) );
  FA_7413 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n567), .CI(C[51]), 
        .CO(C[52]) );
  FA_7412 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n568), .CI(C[52]), 
        .CO(C[53]) );
  FA_7411 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n569), .CI(C[53]), 
        .CO(C[54]) );
  FA_7410 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n570), .CI(C[54]), 
        .CO(C[55]) );
  FA_7409 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n571), .CI(C[55]), 
        .CO(C[56]) );
  FA_7408 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n572), .CI(C[56]), 
        .CO(C[57]) );
  FA_7407 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n573), .CI(C[57]), 
        .CO(C[58]) );
  FA_7406 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n574), .CI(C[58]), 
        .CO(C[59]) );
  FA_7405 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n575), .CI(C[59]), 
        .CO(C[60]) );
  FA_7404 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n576), .CI(C[60]), 
        .CO(C[61]) );
  FA_7403 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n577), .CI(C[61]), 
        .CO(C[62]) );
  FA_7402 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n578), .CI(C[62]), 
        .CO(C[63]) );
  FA_7401 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n579), .CI(C[63]), 
        .CO(C[64]) );
  FA_7400 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n580), .CI(C[64]), 
        .CO(C[65]) );
  FA_7399 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n581), .CI(C[65]), 
        .CO(C[66]) );
  FA_7398 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n582), .CI(C[66]), 
        .CO(C[67]) );
  FA_7397 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n583), .CI(C[67]), 
        .CO(C[68]) );
  FA_7396 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n584), .CI(C[68]), 
        .CO(C[69]) );
  FA_7395 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n585), .CI(C[69]), 
        .CO(C[70]) );
  FA_7394 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n586), .CI(C[70]), 
        .CO(C[71]) );
  FA_7393 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n587), .CI(C[71]), 
        .CO(C[72]) );
  FA_7392 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n588), .CI(C[72]), 
        .CO(C[73]) );
  FA_7391 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n589), .CI(C[73]), 
        .CO(C[74]) );
  FA_7390 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n590), .CI(C[74]), 
        .CO(C[75]) );
  FA_7389 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n591), .CI(C[75]), 
        .CO(C[76]) );
  FA_7388 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n592), .CI(C[76]), 
        .CO(C[77]) );
  FA_7387 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n593), .CI(C[77]), 
        .CO(C[78]) );
  FA_7386 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n594), .CI(C[78]), 
        .CO(C[79]) );
  FA_7385 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n595), .CI(C[79]), 
        .CO(C[80]) );
  FA_7384 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n596), .CI(C[80]), 
        .CO(C[81]) );
  FA_7383 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n597), .CI(C[81]), 
        .CO(C[82]) );
  FA_7382 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n598), .CI(C[82]), 
        .CO(C[83]) );
  FA_7381 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n599), .CI(C[83]), 
        .CO(C[84]) );
  FA_7380 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n600), .CI(C[84]), 
        .CO(C[85]) );
  FA_7379 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n601), .CI(C[85]), 
        .CO(C[86]) );
  FA_7378 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n602), .CI(C[86]), 
        .CO(C[87]) );
  FA_7377 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n603), .CI(C[87]), 
        .CO(C[88]) );
  FA_7376 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n604), .CI(C[88]), 
        .CO(C[89]) );
  FA_7375 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n605), .CI(C[89]), 
        .CO(C[90]) );
  FA_7374 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n606), .CI(C[90]), 
        .CO(C[91]) );
  FA_7373 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n607), .CI(C[91]), 
        .CO(C[92]) );
  FA_7372 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n608), .CI(C[92]), 
        .CO(C[93]) );
  FA_7371 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n609), .CI(C[93]), 
        .CO(C[94]) );
  FA_7370 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n610), .CI(C[94]), 
        .CO(C[95]) );
  FA_7369 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n611), .CI(C[95]), 
        .CO(C[96]) );
  FA_7368 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n612), .CI(C[96]), 
        .CO(C[97]) );
  FA_7367 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n613), .CI(C[97]), 
        .CO(C[98]) );
  FA_7366 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n614), .CI(C[98]), 
        .CO(C[99]) );
  FA_7365 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n615), .CI(C[99]), 
        .CO(C[100]) );
  FA_7364 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n616), .CI(C[100]), .CO(C[101]) );
  FA_7363 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n617), .CI(C[101]), .CO(C[102]) );
  FA_7362 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n618), .CI(C[102]), .CO(C[103]) );
  FA_7361 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n619), .CI(C[103]), .CO(C[104]) );
  FA_7360 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n620), .CI(C[104]), .CO(C[105]) );
  FA_7359 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n621), .CI(C[105]), .CO(C[106]) );
  FA_7358 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n622), .CI(C[106]), .CO(C[107]) );
  FA_7357 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n623), .CI(C[107]), .CO(C[108]) );
  FA_7356 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n624), .CI(C[108]), .CO(C[109]) );
  FA_7355 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n625), .CI(C[109]), .CO(C[110]) );
  FA_7354 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n626), .CI(C[110]), .CO(C[111]) );
  FA_7353 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n627), .CI(C[111]), .CO(C[112]) );
  FA_7352 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n628), .CI(C[112]), .CO(C[113]) );
  FA_7351 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n629), .CI(C[113]), .CO(C[114]) );
  FA_7350 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n630), .CI(C[114]), .CO(C[115]) );
  FA_7349 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n631), .CI(C[115]), .CO(C[116]) );
  FA_7348 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n632), .CI(C[116]), .CO(C[117]) );
  FA_7347 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n633), .CI(C[117]), .CO(C[118]) );
  FA_7346 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n634), .CI(C[118]), .CO(C[119]) );
  FA_7345 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n635), .CI(C[119]), .CO(C[120]) );
  FA_7344 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n636), .CI(C[120]), .CO(C[121]) );
  FA_7343 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n637), .CI(C[121]), .CO(C[122]) );
  FA_7342 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n638), .CI(C[122]), .CO(C[123]) );
  FA_7341 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n639), .CI(C[123]), .CO(C[124]) );
  FA_7340 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n640), .CI(C[124]), .CO(C[125]) );
  FA_7339 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n641), .CI(C[125]), .CO(C[126]) );
  FA_7338 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n642), .CI(C[126]), .CO(C[127]) );
  FA_7337 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n643), .CI(C[127]), .CO(C[128]) );
  FA_7336 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n644), .CI(C[128]), .CO(C[129]) );
  FA_7335 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n645), .CI(C[129]), .CO(C[130]) );
  FA_7334 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n646), .CI(C[130]), .CO(C[131]) );
  FA_7333 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n647), .CI(C[131]), .CO(C[132]) );
  FA_7332 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n648), .CI(C[132]), .CO(C[133]) );
  FA_7331 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n649), .CI(C[133]), .CO(C[134]) );
  FA_7330 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n650), .CI(C[134]), .CO(C[135]) );
  FA_7329 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n651), .CI(C[135]), .CO(C[136]) );
  FA_7328 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n652), .CI(C[136]), .CO(C[137]) );
  FA_7327 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n653), .CI(C[137]), .CO(C[138]) );
  FA_7326 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n654), .CI(C[138]), .CO(C[139]) );
  FA_7325 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n655), .CI(C[139]), .CO(C[140]) );
  FA_7324 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n656), .CI(C[140]), .CO(C[141]) );
  FA_7323 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n657), .CI(C[141]), .CO(C[142]) );
  FA_7322 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n658), .CI(C[142]), .CO(C[143]) );
  FA_7321 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n659), .CI(C[143]), .CO(C[144]) );
  FA_7320 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n660), .CI(C[144]), .CO(C[145]) );
  FA_7319 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n661), .CI(C[145]), .CO(C[146]) );
  FA_7318 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n662), .CI(C[146]), .CO(C[147]) );
  FA_7317 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n663), .CI(C[147]), .CO(C[148]) );
  FA_7316 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n664), .CI(C[148]), .CO(C[149]) );
  FA_7315 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n665), .CI(C[149]), .CO(C[150]) );
  FA_7314 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n666), .CI(C[150]), .CO(C[151]) );
  FA_7313 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n667), .CI(C[151]), .CO(C[152]) );
  FA_7312 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n668), .CI(C[152]), .CO(C[153]) );
  FA_7311 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n669), .CI(C[153]), .CO(C[154]) );
  FA_7310 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n670), .CI(C[154]), .CO(C[155]) );
  FA_7309 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n671), .CI(C[155]), .CO(C[156]) );
  FA_7308 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n672), .CI(C[156]), .CO(C[157]) );
  FA_7307 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n673), .CI(C[157]), .CO(C[158]) );
  FA_7306 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n674), .CI(C[158]), .CO(C[159]) );
  FA_7305 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n675), .CI(C[159]), .CO(C[160]) );
  FA_7304 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n676), .CI(C[160]), .CO(C[161]) );
  FA_7303 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n677), .CI(C[161]), .CO(C[162]) );
  FA_7302 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n678), .CI(C[162]), .CO(C[163]) );
  FA_7301 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n679), .CI(C[163]), .CO(C[164]) );
  FA_7300 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n680), .CI(C[164]), .CO(C[165]) );
  FA_7299 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n681), .CI(C[165]), .CO(C[166]) );
  FA_7298 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n682), .CI(C[166]), .CO(C[167]) );
  FA_7297 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n683), .CI(C[167]), .CO(C[168]) );
  FA_7296 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n684), .CI(C[168]), .CO(C[169]) );
  FA_7295 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n685), .CI(C[169]), .CO(C[170]) );
  FA_7294 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n686), .CI(C[170]), .CO(C[171]) );
  FA_7293 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n687), .CI(C[171]), .CO(C[172]) );
  FA_7292 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n688), .CI(C[172]), .CO(C[173]) );
  FA_7291 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n689), .CI(C[173]), .CO(C[174]) );
  FA_7290 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n690), .CI(C[174]), .CO(C[175]) );
  FA_7289 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n691), .CI(C[175]), .CO(C[176]) );
  FA_7288 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n692), .CI(C[176]), .CO(C[177]) );
  FA_7287 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n693), .CI(C[177]), .CO(C[178]) );
  FA_7286 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n694), .CI(C[178]), .CO(C[179]) );
  FA_7285 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n695), .CI(C[179]), .CO(C[180]) );
  FA_7284 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n696), .CI(C[180]), .CO(C[181]) );
  FA_7283 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n697), .CI(C[181]), .CO(C[182]) );
  FA_7282 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n698), .CI(C[182]), .CO(C[183]) );
  FA_7281 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n699), .CI(C[183]), .CO(C[184]) );
  FA_7280 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n700), .CI(C[184]), .CO(C[185]) );
  FA_7279 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n701), .CI(C[185]), .CO(C[186]) );
  FA_7278 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n702), .CI(C[186]), .CO(C[187]) );
  FA_7277 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n703), .CI(C[187]), .CO(C[188]) );
  FA_7276 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n704), .CI(C[188]), .CO(C[189]) );
  FA_7275 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n705), .CI(C[189]), .CO(C[190]) );
  FA_7274 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n706), .CI(C[190]), .CO(C[191]) );
  FA_7273 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n707), .CI(C[191]), .CO(C[192]) );
  FA_7272 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n708), .CI(C[192]), .CO(C[193]) );
  FA_7271 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n709), .CI(C[193]), .CO(C[194]) );
  FA_7270 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n710), .CI(C[194]), .CO(C[195]) );
  FA_7269 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n711), .CI(C[195]), .CO(C[196]) );
  FA_7268 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n712), .CI(C[196]), .CO(C[197]) );
  FA_7267 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n713), .CI(C[197]), .CO(C[198]) );
  FA_7266 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n714), .CI(C[198]), .CO(C[199]) );
  FA_7265 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n715), .CI(C[199]), .CO(C[200]) );
  FA_7264 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n716), .CI(C[200]), .CO(C[201]) );
  FA_7263 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n717), .CI(C[201]), .CO(C[202]) );
  FA_7262 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n718), .CI(C[202]), .CO(C[203]) );
  FA_7261 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n719), .CI(C[203]), .CO(C[204]) );
  FA_7260 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n720), .CI(C[204]), .CO(C[205]) );
  FA_7259 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n721), .CI(C[205]), .CO(C[206]) );
  FA_7258 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n722), .CI(C[206]), .CO(C[207]) );
  FA_7257 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n723), .CI(C[207]), .CO(C[208]) );
  FA_7256 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n724), .CI(C[208]), .CO(C[209]) );
  FA_7255 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n725), .CI(C[209]), .CO(C[210]) );
  FA_7254 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n726), .CI(C[210]), .CO(C[211]) );
  FA_7253 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n727), .CI(C[211]), .CO(C[212]) );
  FA_7252 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n728), .CI(C[212]), .CO(C[213]) );
  FA_7251 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n729), .CI(C[213]), .CO(C[214]) );
  FA_7250 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n730), .CI(C[214]), .CO(C[215]) );
  FA_7249 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n731), .CI(C[215]), .CO(C[216]) );
  FA_7248 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n732), .CI(C[216]), .CO(C[217]) );
  FA_7247 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n733), .CI(C[217]), .CO(C[218]) );
  FA_7246 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n734), .CI(C[218]), .CO(C[219]) );
  FA_7245 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n735), .CI(C[219]), .CO(C[220]) );
  FA_7244 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n736), .CI(C[220]), .CO(C[221]) );
  FA_7243 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n737), .CI(C[221]), .CO(C[222]) );
  FA_7242 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n738), .CI(C[222]), .CO(C[223]) );
  FA_7241 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n739), .CI(C[223]), .CO(C[224]) );
  FA_7240 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n740), .CI(C[224]), .CO(C[225]) );
  FA_7239 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n741), .CI(C[225]), .CO(C[226]) );
  FA_7238 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n742), .CI(C[226]), .CO(C[227]) );
  FA_7237 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n743), .CI(C[227]), .CO(C[228]) );
  FA_7236 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n744), .CI(C[228]), .CO(C[229]) );
  FA_7235 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n745), .CI(C[229]), .CO(C[230]) );
  FA_7234 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n746), .CI(C[230]), .CO(C[231]) );
  FA_7233 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n747), .CI(C[231]), .CO(C[232]) );
  FA_7232 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n748), .CI(C[232]), .CO(C[233]) );
  FA_7231 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n749), .CI(C[233]), .CO(C[234]) );
  FA_7230 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n750), .CI(C[234]), .CO(C[235]) );
  FA_7229 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n751), .CI(C[235]), .CO(C[236]) );
  FA_7228 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n752), .CI(C[236]), .CO(C[237]) );
  FA_7227 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n753), .CI(C[237]), .CO(C[238]) );
  FA_7226 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n754), .CI(C[238]), .CO(C[239]) );
  FA_7225 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n755), .CI(C[239]), .CO(C[240]) );
  FA_7224 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n756), .CI(C[240]), .CO(C[241]) );
  FA_7223 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n757), .CI(C[241]), .CO(C[242]) );
  FA_7222 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n758), .CI(C[242]), .CO(C[243]) );
  FA_7221 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n759), .CI(C[243]), .CO(C[244]) );
  FA_7220 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n760), .CI(C[244]), .CO(C[245]) );
  FA_7219 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n761), .CI(C[245]), .CO(C[246]) );
  FA_7218 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n762), .CI(C[246]), .CO(C[247]) );
  FA_7217 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n763), .CI(C[247]), .CO(C[248]) );
  FA_7216 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n764), .CI(C[248]), .CO(C[249]) );
  FA_7215 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n765), .CI(C[249]), .CO(C[250]) );
  FA_7214 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n766), .CI(C[250]), .CO(C[251]) );
  FA_7213 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n767), .CI(C[251]), .CO(C[252]) );
  FA_7212 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n768), .CI(C[252]), .CO(C[253]) );
  FA_7211 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n769), .CI(C[253]), .CO(C[254]) );
  FA_7210 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n770), .CI(C[254]), .CO(C[255]) );
  FA_7209 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n771), .CI(C[255]), .CO(C[256]) );
  FA_7208 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n772), .CI(C[256]), .CO(C[257]) );
  FA_7207 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n773), .CI(C[257]), .CO(C[258]) );
  FA_7206 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n774), .CI(C[258]), .CO(C[259]) );
  FA_7205 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n775), .CI(C[259]), .CO(C[260]) );
  FA_7204 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n776), .CI(C[260]), .CO(C[261]) );
  FA_7203 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n777), .CI(C[261]), .CO(C[262]) );
  FA_7202 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n778), .CI(C[262]), .CO(C[263]) );
  FA_7201 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n779), .CI(C[263]), .CO(C[264]) );
  FA_7200 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n780), .CI(C[264]), .CO(C[265]) );
  FA_7199 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n781), .CI(C[265]), .CO(C[266]) );
  FA_7198 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n782), .CI(C[266]), .CO(C[267]) );
  FA_7197 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n783), .CI(C[267]), .CO(C[268]) );
  FA_7196 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n784), .CI(C[268]), .CO(C[269]) );
  FA_7195 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n785), .CI(C[269]), .CO(C[270]) );
  FA_7194 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n786), .CI(C[270]), .CO(C[271]) );
  FA_7193 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n787), .CI(C[271]), .CO(C[272]) );
  FA_7192 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n788), .CI(C[272]), .CO(C[273]) );
  FA_7191 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n789), .CI(C[273]), .CO(C[274]) );
  FA_7190 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n790), .CI(C[274]), .CO(C[275]) );
  FA_7189 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n791), .CI(C[275]), .CO(C[276]) );
  FA_7188 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n792), .CI(C[276]), .CO(C[277]) );
  FA_7187 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n793), .CI(C[277]), .CO(C[278]) );
  FA_7186 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n794), .CI(C[278]), .CO(C[279]) );
  FA_7185 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n795), .CI(C[279]), .CO(C[280]) );
  FA_7184 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n796), .CI(C[280]), .CO(C[281]) );
  FA_7183 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n797), .CI(C[281]), .CO(C[282]) );
  FA_7182 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n798), .CI(C[282]), .CO(C[283]) );
  FA_7181 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n799), .CI(C[283]), .CO(C[284]) );
  FA_7180 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n800), .CI(C[284]), .CO(C[285]) );
  FA_7179 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n801), .CI(C[285]), .CO(C[286]) );
  FA_7178 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n802), .CI(C[286]), .CO(C[287]) );
  FA_7177 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n803), .CI(C[287]), .CO(C[288]) );
  FA_7176 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n804), .CI(C[288]), .CO(C[289]) );
  FA_7175 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n805), .CI(C[289]), .CO(C[290]) );
  FA_7174 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n806), .CI(C[290]), .CO(C[291]) );
  FA_7173 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n807), .CI(C[291]), .CO(C[292]) );
  FA_7172 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n808), .CI(C[292]), .CO(C[293]) );
  FA_7171 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n809), .CI(C[293]), .CO(C[294]) );
  FA_7170 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n810), .CI(C[294]), .CO(C[295]) );
  FA_7169 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n811), .CI(C[295]), .CO(C[296]) );
  FA_7168 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n812), .CI(C[296]), .CO(C[297]) );
  FA_7167 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n813), .CI(C[297]), .CO(C[298]) );
  FA_7166 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n814), .CI(C[298]), .CO(C[299]) );
  FA_7165 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n815), .CI(C[299]), .CO(C[300]) );
  FA_7164 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n816), .CI(C[300]), .CO(C[301]) );
  FA_7163 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n817), .CI(C[301]), .CO(C[302]) );
  FA_7162 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n818), .CI(C[302]), .CO(C[303]) );
  FA_7161 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n819), .CI(C[303]), .CO(C[304]) );
  FA_7160 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n820), .CI(C[304]), .CO(C[305]) );
  FA_7159 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n821), .CI(C[305]), .CO(C[306]) );
  FA_7158 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n822), .CI(C[306]), .CO(C[307]) );
  FA_7157 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n823), .CI(C[307]), .CO(C[308]) );
  FA_7156 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n824), .CI(C[308]), .CO(C[309]) );
  FA_7155 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n825), .CI(C[309]), .CO(C[310]) );
  FA_7154 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n826), .CI(C[310]), .CO(C[311]) );
  FA_7153 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n827), .CI(C[311]), .CO(C[312]) );
  FA_7152 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n828), .CI(C[312]), .CO(C[313]) );
  FA_7151 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n829), .CI(C[313]), .CO(C[314]) );
  FA_7150 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n830), .CI(C[314]), .CO(C[315]) );
  FA_7149 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n831), .CI(C[315]), .CO(C[316]) );
  FA_7148 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n832), .CI(C[316]), .CO(C[317]) );
  FA_7147 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n833), .CI(C[317]), .CO(C[318]) );
  FA_7146 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n834), .CI(C[318]), .CO(C[319]) );
  FA_7145 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n835), .CI(C[319]), .CO(C[320]) );
  FA_7144 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n836), .CI(C[320]), .CO(C[321]) );
  FA_7143 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n837), .CI(C[321]), .CO(C[322]) );
  FA_7142 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n838), .CI(C[322]), .CO(C[323]) );
  FA_7141 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n839), .CI(C[323]), .CO(C[324]) );
  FA_7140 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n840), .CI(C[324]), .CO(C[325]) );
  FA_7139 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n841), .CI(C[325]), .CO(C[326]) );
  FA_7138 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n842), .CI(C[326]), .CO(C[327]) );
  FA_7137 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n843), .CI(C[327]), .CO(C[328]) );
  FA_7136 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n844), .CI(C[328]), .CO(C[329]) );
  FA_7135 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n845), .CI(C[329]), .CO(C[330]) );
  FA_7134 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n846), .CI(C[330]), .CO(C[331]) );
  FA_7133 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n847), .CI(C[331]), .CO(C[332]) );
  FA_7132 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n848), .CI(C[332]), .CO(C[333]) );
  FA_7131 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n849), .CI(C[333]), .CO(C[334]) );
  FA_7130 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n850), .CI(C[334]), .CO(C[335]) );
  FA_7129 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n851), .CI(C[335]), .CO(C[336]) );
  FA_7128 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n852), .CI(C[336]), .CO(C[337]) );
  FA_7127 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n853), .CI(C[337]), .CO(C[338]) );
  FA_7126 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n854), .CI(C[338]), .CO(C[339]) );
  FA_7125 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n855), .CI(C[339]), .CO(C[340]) );
  FA_7124 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n856), .CI(C[340]), .CO(C[341]) );
  FA_7123 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n857), .CI(C[341]), .CO(C[342]) );
  FA_7122 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n858), .CI(C[342]), .CO(C[343]) );
  FA_7121 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n859), .CI(C[343]), .CO(C[344]) );
  FA_7120 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n860), .CI(C[344]), .CO(C[345]) );
  FA_7119 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n861), .CI(C[345]), .CO(C[346]) );
  FA_7118 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n862), .CI(C[346]), .CO(C[347]) );
  FA_7117 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n863), .CI(C[347]), .CO(C[348]) );
  FA_7116 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n864), .CI(C[348]), .CO(C[349]) );
  FA_7115 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n865), .CI(C[349]), .CO(C[350]) );
  FA_7114 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n866), .CI(C[350]), .CO(C[351]) );
  FA_7113 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n867), .CI(C[351]), .CO(C[352]) );
  FA_7112 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n868), .CI(C[352]), .CO(C[353]) );
  FA_7111 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n869), .CI(C[353]), .CO(C[354]) );
  FA_7110 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n870), .CI(C[354]), .CO(C[355]) );
  FA_7109 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n871), .CI(C[355]), .CO(C[356]) );
  FA_7108 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n872), .CI(C[356]), .CO(C[357]) );
  FA_7107 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n873), .CI(C[357]), .CO(C[358]) );
  FA_7106 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n874), .CI(C[358]), .CO(C[359]) );
  FA_7105 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n875), .CI(C[359]), .CO(C[360]) );
  FA_7104 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n876), .CI(C[360]), .CO(C[361]) );
  FA_7103 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n877), .CI(C[361]), .CO(C[362]) );
  FA_7102 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n878), .CI(C[362]), .CO(C[363]) );
  FA_7101 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n879), .CI(C[363]), .CO(C[364]) );
  FA_7100 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n880), .CI(C[364]), .CO(C[365]) );
  FA_7099 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n881), .CI(C[365]), .CO(C[366]) );
  FA_7098 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n882), .CI(C[366]), .CO(C[367]) );
  FA_7097 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n883), .CI(C[367]), .CO(C[368]) );
  FA_7096 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n884), .CI(C[368]), .CO(C[369]) );
  FA_7095 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n885), .CI(C[369]), .CO(C[370]) );
  FA_7094 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n886), .CI(C[370]), .CO(C[371]) );
  FA_7093 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n887), .CI(C[371]), .CO(C[372]) );
  FA_7092 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n888), .CI(C[372]), .CO(C[373]) );
  FA_7091 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n889), .CI(C[373]), .CO(C[374]) );
  FA_7090 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n890), .CI(C[374]), .CO(C[375]) );
  FA_7089 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n891), .CI(C[375]), .CO(C[376]) );
  FA_7088 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n892), .CI(C[376]), .CO(C[377]) );
  FA_7087 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n893), .CI(C[377]), .CO(C[378]) );
  FA_7086 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n894), .CI(C[378]), .CO(C[379]) );
  FA_7085 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n895), .CI(C[379]), .CO(C[380]) );
  FA_7084 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n896), .CI(C[380]), .CO(C[381]) );
  FA_7083 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n897), .CI(C[381]), .CO(C[382]) );
  FA_7082 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n898), .CI(C[382]), .CO(C[383]) );
  FA_7081 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n899), .CI(C[383]), .CO(C[384]) );
  FA_7080 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n900), .CI(C[384]), .CO(C[385]) );
  FA_7079 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n901), .CI(C[385]), .CO(C[386]) );
  FA_7078 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n902), .CI(C[386]), .CO(C[387]) );
  FA_7077 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n903), .CI(C[387]), .CO(C[388]) );
  FA_7076 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n904), .CI(C[388]), .CO(C[389]) );
  FA_7075 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n905), .CI(C[389]), .CO(C[390]) );
  FA_7074 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n906), .CI(C[390]), .CO(C[391]) );
  FA_7073 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n907), .CI(C[391]), .CO(C[392]) );
  FA_7072 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n908), .CI(C[392]), .CO(C[393]) );
  FA_7071 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n909), .CI(C[393]), .CO(C[394]) );
  FA_7070 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n910), .CI(C[394]), .CO(C[395]) );
  FA_7069 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n911), .CI(C[395]), .CO(C[396]) );
  FA_7068 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n912), .CI(C[396]), .CO(C[397]) );
  FA_7067 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n913), .CI(C[397]), .CO(C[398]) );
  FA_7066 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n914), .CI(C[398]), .CO(C[399]) );
  FA_7065 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n915), .CI(C[399]), .CO(C[400]) );
  FA_7064 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n916), .CI(C[400]), .CO(C[401]) );
  FA_7063 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n917), .CI(C[401]), .CO(C[402]) );
  FA_7062 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n918), .CI(C[402]), .CO(C[403]) );
  FA_7061 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n919), .CI(C[403]), .CO(C[404]) );
  FA_7060 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n920), .CI(C[404]), .CO(C[405]) );
  FA_7059 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n921), .CI(C[405]), .CO(C[406]) );
  FA_7058 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n922), .CI(C[406]), .CO(C[407]) );
  FA_7057 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n923), .CI(C[407]), .CO(C[408]) );
  FA_7056 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n924), .CI(C[408]), .CO(C[409]) );
  FA_7055 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n925), .CI(C[409]), .CO(C[410]) );
  FA_7054 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n926), .CI(C[410]), .CO(C[411]) );
  FA_7053 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n927), .CI(C[411]), .CO(C[412]) );
  FA_7052 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n928), .CI(C[412]), .CO(C[413]) );
  FA_7051 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n929), .CI(C[413]), .CO(C[414]) );
  FA_7050 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n930), .CI(C[414]), .CO(C[415]) );
  FA_7049 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n931), .CI(C[415]), .CO(C[416]) );
  FA_7048 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n932), .CI(C[416]), .CO(C[417]) );
  FA_7047 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n933), .CI(C[417]), .CO(C[418]) );
  FA_7046 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n934), .CI(C[418]), .CO(C[419]) );
  FA_7045 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n935), .CI(C[419]), .CO(C[420]) );
  FA_7044 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n936), .CI(C[420]), .CO(C[421]) );
  FA_7043 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n937), .CI(C[421]), .CO(C[422]) );
  FA_7042 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n938), .CI(C[422]), .CO(C[423]) );
  FA_7041 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n939), .CI(C[423]), .CO(C[424]) );
  FA_7040 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n940), .CI(C[424]), .CO(C[425]) );
  FA_7039 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n941), .CI(C[425]), .CO(C[426]) );
  FA_7038 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n942), .CI(C[426]), .CO(C[427]) );
  FA_7037 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n943), .CI(C[427]), .CO(C[428]) );
  FA_7036 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n944), .CI(C[428]), .CO(C[429]) );
  FA_7035 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n945), .CI(C[429]), .CO(C[430]) );
  FA_7034 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n946), .CI(C[430]), .CO(C[431]) );
  FA_7033 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n947), .CI(C[431]), .CO(C[432]) );
  FA_7032 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n948), .CI(C[432]), .CO(C[433]) );
  FA_7031 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n949), .CI(C[433]), .CO(C[434]) );
  FA_7030 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n950), .CI(C[434]), .CO(C[435]) );
  FA_7029 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n951), .CI(C[435]), .CO(C[436]) );
  FA_7028 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n952), .CI(C[436]), .CO(C[437]) );
  FA_7027 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n953), .CI(C[437]), .CO(C[438]) );
  FA_7026 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n954), .CI(C[438]), .CO(C[439]) );
  FA_7025 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n955), .CI(C[439]), .CO(C[440]) );
  FA_7024 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n956), .CI(C[440]), .CO(C[441]) );
  FA_7023 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n957), .CI(C[441]), .CO(C[442]) );
  FA_7022 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n958), .CI(C[442]), .CO(C[443]) );
  FA_7021 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n959), .CI(C[443]), .CO(C[444]) );
  FA_7020 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n960), .CI(C[444]), .CO(C[445]) );
  FA_7019 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n961), .CI(C[445]), .CO(C[446]) );
  FA_7018 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n962), .CI(C[446]), .CO(C[447]) );
  FA_7017 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n963), .CI(C[447]), .CO(C[448]) );
  FA_7016 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n964), .CI(C[448]), .CO(C[449]) );
  FA_7015 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n965), .CI(C[449]), .CO(C[450]) );
  FA_7014 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n966), .CI(C[450]), .CO(C[451]) );
  FA_7013 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n967), .CI(C[451]), .CO(C[452]) );
  FA_7012 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n968), .CI(C[452]), .CO(C[453]) );
  FA_7011 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n969), .CI(C[453]), .CO(C[454]) );
  FA_7010 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n970), .CI(C[454]), .CO(C[455]) );
  FA_7009 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n971), .CI(C[455]), .CO(C[456]) );
  FA_7008 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n972), .CI(C[456]), .CO(C[457]) );
  FA_7007 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n973), .CI(C[457]), .CO(C[458]) );
  FA_7006 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n974), .CI(C[458]), .CO(C[459]) );
  FA_7005 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n975), .CI(C[459]), .CO(C[460]) );
  FA_7004 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n976), .CI(C[460]), .CO(C[461]) );
  FA_7003 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n977), .CI(C[461]), .CO(C[462]) );
  FA_7002 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n978), .CI(C[462]), .CO(C[463]) );
  FA_7001 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n979), .CI(C[463]), .CO(C[464]) );
  FA_7000 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n980), .CI(C[464]), .CO(C[465]) );
  FA_6999 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n981), .CI(C[465]), .CO(C[466]) );
  FA_6998 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n982), .CI(C[466]), .CO(C[467]) );
  FA_6997 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n983), .CI(C[467]), .CO(C[468]) );
  FA_6996 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n984), .CI(C[468]), .CO(C[469]) );
  FA_6995 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n985), .CI(C[469]), .CO(C[470]) );
  FA_6994 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n986), .CI(C[470]), .CO(C[471]) );
  FA_6993 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n987), .CI(C[471]), .CO(C[472]) );
  FA_6992 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n988), .CI(C[472]), .CO(C[473]) );
  FA_6991 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n989), .CI(C[473]), .CO(C[474]) );
  FA_6990 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n990), .CI(C[474]), .CO(C[475]) );
  FA_6989 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n991), .CI(C[475]), .CO(C[476]) );
  FA_6988 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n992), .CI(C[476]), .CO(C[477]) );
  FA_6987 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n993), .CI(C[477]), .CO(C[478]) );
  FA_6986 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n994), .CI(C[478]), .CO(C[479]) );
  FA_6985 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n995), .CI(C[479]), .CO(C[480]) );
  FA_6984 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n996), .CI(C[480]), .CO(C[481]) );
  FA_6983 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n997), .CI(C[481]), .CO(C[482]) );
  FA_6982 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n998), .CI(C[482]), .CO(C[483]) );
  FA_6981 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n999), .CI(C[483]), .CO(C[484]) );
  FA_6980 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n1000), .CI(
        C[484]), .CO(C[485]) );
  FA_6979 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n1001), .CI(
        C[485]), .CO(C[486]) );
  FA_6978 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n1002), .CI(
        C[486]), .CO(C[487]) );
  FA_6977 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1003), .CI(
        C[487]), .CO(C[488]) );
  FA_6976 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1004), .CI(
        C[488]), .CO(C[489]) );
  FA_6975 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1005), .CI(
        C[489]), .CO(C[490]) );
  FA_6974 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1006), .CI(
        C[490]), .CO(C[491]) );
  FA_6973 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1007), .CI(
        C[491]), .CO(C[492]) );
  FA_6972 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1008), .CI(
        C[492]), .CO(C[493]) );
  FA_6971 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1009), .CI(
        C[493]), .CO(C[494]) );
  FA_6970 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1010), .CI(
        C[494]), .CO(C[495]) );
  FA_6969 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1011), .CI(
        C[495]), .CO(C[496]) );
  FA_6968 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1012), .CI(
        C[496]), .CO(C[497]) );
  FA_6967 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1013), .CI(
        C[497]), .CO(C[498]) );
  FA_6966 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1014), .CI(
        C[498]), .CO(C[499]) );
  FA_6965 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1015), .CI(
        C[499]), .CO(C[500]) );
  FA_6964 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1016), .CI(
        C[500]), .CO(C[501]) );
  FA_6963 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1017), .CI(
        C[501]), .CO(C[502]) );
  FA_6962 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1018), .CI(
        C[502]), .CO(C[503]) );
  FA_6961 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1019), .CI(
        C[503]), .CO(C[504]) );
  FA_6960 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1020), .CI(
        C[504]), .CO(C[505]) );
  FA_6959 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1021), .CI(
        C[505]), .CO(C[506]) );
  FA_6958 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1022), .CI(
        C[506]), .CO(C[507]) );
  FA_6957 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1023), .CI(
        C[507]), .CO(C[508]) );
  FA_6956 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1024), .CI(
        C[508]), .CO(C[509]) );
  FA_6955 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1025), .CI(
        C[509]), .CO(C[510]) );
  FA_6954 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1026), .CI(
        C[510]), .CO(C[511]) );
  FA_6953 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1027), .CI(
        C[511]), .CO(C[512]) );
  FA_6952 \FA_INST_1[512].FA_  ( .A(1'b0), .B(n1028), .CI(C[512]), .CO(C[513])
         );
  FA_6951 \FA_INST_1[513].FA_  ( .A(1'b0), .B(n1029), .CI(C[513]), .CO(O) );
  IV U2 ( .A(B[415]), .Z(n931) );
  IV U3 ( .A(B[416]), .Z(n932) );
  IV U4 ( .A(B[417]), .Z(n933) );
  IV U5 ( .A(B[418]), .Z(n934) );
  IV U6 ( .A(B[419]), .Z(n935) );
  IV U7 ( .A(B[420]), .Z(n936) );
  IV U8 ( .A(B[421]), .Z(n937) );
  IV U9 ( .A(B[422]), .Z(n938) );
  IV U10 ( .A(B[423]), .Z(n939) );
  IV U11 ( .A(B[424]), .Z(n940) );
  IV U12 ( .A(B[505]), .Z(n1021) );
  IV U13 ( .A(B[425]), .Z(n941) );
  IV U14 ( .A(B[426]), .Z(n942) );
  IV U15 ( .A(B[427]), .Z(n943) );
  IV U16 ( .A(B[428]), .Z(n944) );
  IV U17 ( .A(B[429]), .Z(n945) );
  IV U18 ( .A(B[430]), .Z(n946) );
  IV U19 ( .A(B[431]), .Z(n947) );
  IV U20 ( .A(B[432]), .Z(n948) );
  IV U21 ( .A(B[433]), .Z(n949) );
  IV U22 ( .A(B[434]), .Z(n950) );
  IV U23 ( .A(B[506]), .Z(n1022) );
  IV U24 ( .A(B[435]), .Z(n951) );
  IV U25 ( .A(B[436]), .Z(n952) );
  IV U26 ( .A(B[437]), .Z(n953) );
  IV U27 ( .A(B[438]), .Z(n954) );
  IV U28 ( .A(B[439]), .Z(n955) );
  IV U29 ( .A(B[440]), .Z(n956) );
  IV U30 ( .A(B[441]), .Z(n957) );
  IV U31 ( .A(B[442]), .Z(n958) );
  IV U32 ( .A(B[443]), .Z(n959) );
  IV U33 ( .A(B[444]), .Z(n960) );
  IV U34 ( .A(B[507]), .Z(n1023) );
  IV U35 ( .A(B[445]), .Z(n961) );
  IV U36 ( .A(B[446]), .Z(n962) );
  IV U37 ( .A(B[447]), .Z(n963) );
  IV U38 ( .A(B[448]), .Z(n964) );
  IV U39 ( .A(B[449]), .Z(n965) );
  IV U40 ( .A(B[450]), .Z(n966) );
  IV U41 ( .A(B[451]), .Z(n967) );
  IV U42 ( .A(B[452]), .Z(n968) );
  IV U43 ( .A(B[453]), .Z(n969) );
  IV U44 ( .A(B[454]), .Z(n970) );
  IV U45 ( .A(B[508]), .Z(n1024) );
  IV U46 ( .A(B[455]), .Z(n971) );
  IV U47 ( .A(B[456]), .Z(n972) );
  IV U48 ( .A(B[457]), .Z(n973) );
  IV U49 ( .A(B[458]), .Z(n974) );
  IV U50 ( .A(B[459]), .Z(n975) );
  IV U51 ( .A(B[460]), .Z(n976) );
  IV U52 ( .A(B[461]), .Z(n977) );
  IV U53 ( .A(B[462]), .Z(n978) );
  IV U54 ( .A(B[0]), .Z(n516) );
  IV U55 ( .A(B[1]), .Z(n517) );
  IV U56 ( .A(B[2]), .Z(n518) );
  IV U57 ( .A(B[3]), .Z(n519) );
  IV U58 ( .A(B[4]), .Z(n520) );
  IV U59 ( .A(B[463]), .Z(n979) );
  IV U60 ( .A(B[5]), .Z(n521) );
  IV U61 ( .A(B[6]), .Z(n522) );
  IV U62 ( .A(B[7]), .Z(n523) );
  IV U63 ( .A(B[8]), .Z(n524) );
  IV U64 ( .A(B[9]), .Z(n525) );
  IV U65 ( .A(B[10]), .Z(n526) );
  IV U66 ( .A(B[11]), .Z(n527) );
  IV U67 ( .A(B[12]), .Z(n528) );
  IV U68 ( .A(B[13]), .Z(n529) );
  IV U69 ( .A(B[14]), .Z(n530) );
  IV U70 ( .A(B[464]), .Z(n980) );
  IV U71 ( .A(B[509]), .Z(n1025) );
  IV U72 ( .A(B[15]), .Z(n531) );
  IV U73 ( .A(B[16]), .Z(n532) );
  IV U74 ( .A(B[17]), .Z(n533) );
  IV U75 ( .A(B[18]), .Z(n534) );
  IV U76 ( .A(B[19]), .Z(n535) );
  IV U77 ( .A(B[20]), .Z(n536) );
  IV U78 ( .A(B[21]), .Z(n537) );
  IV U79 ( .A(B[22]), .Z(n538) );
  IV U80 ( .A(B[23]), .Z(n539) );
  IV U81 ( .A(B[24]), .Z(n540) );
  IV U82 ( .A(B[465]), .Z(n981) );
  IV U83 ( .A(B[25]), .Z(n541) );
  IV U84 ( .A(B[26]), .Z(n542) );
  IV U85 ( .A(B[27]), .Z(n543) );
  IV U86 ( .A(B[28]), .Z(n544) );
  IV U87 ( .A(B[29]), .Z(n545) );
  IV U88 ( .A(B[30]), .Z(n546) );
  IV U89 ( .A(B[31]), .Z(n547) );
  IV U90 ( .A(B[32]), .Z(n548) );
  IV U91 ( .A(B[33]), .Z(n549) );
  IV U92 ( .A(B[34]), .Z(n550) );
  IV U93 ( .A(B[466]), .Z(n982) );
  IV U94 ( .A(B[35]), .Z(n551) );
  IV U95 ( .A(B[36]), .Z(n552) );
  IV U96 ( .A(B[37]), .Z(n553) );
  IV U97 ( .A(B[38]), .Z(n554) );
  IV U98 ( .A(B[39]), .Z(n555) );
  IV U99 ( .A(B[40]), .Z(n556) );
  IV U100 ( .A(B[41]), .Z(n557) );
  IV U101 ( .A(B[42]), .Z(n558) );
  IV U102 ( .A(B[43]), .Z(n559) );
  IV U103 ( .A(B[44]), .Z(n560) );
  IV U104 ( .A(B[467]), .Z(n983) );
  IV U105 ( .A(B[45]), .Z(n561) );
  IV U106 ( .A(B[46]), .Z(n562) );
  IV U107 ( .A(B[47]), .Z(n563) );
  IV U108 ( .A(B[48]), .Z(n564) );
  IV U109 ( .A(B[49]), .Z(n565) );
  IV U110 ( .A(B[50]), .Z(n566) );
  IV U111 ( .A(B[51]), .Z(n567) );
  IV U112 ( .A(B[52]), .Z(n568) );
  IV U113 ( .A(B[53]), .Z(n569) );
  IV U114 ( .A(B[54]), .Z(n570) );
  IV U115 ( .A(B[468]), .Z(n984) );
  IV U116 ( .A(B[55]), .Z(n571) );
  IV U117 ( .A(B[56]), .Z(n572) );
  IV U118 ( .A(B[57]), .Z(n573) );
  IV U119 ( .A(B[58]), .Z(n574) );
  IV U120 ( .A(B[59]), .Z(n575) );
  IV U121 ( .A(B[60]), .Z(n576) );
  IV U122 ( .A(B[61]), .Z(n577) );
  IV U123 ( .A(B[62]), .Z(n578) );
  IV U124 ( .A(B[63]), .Z(n579) );
  IV U125 ( .A(B[64]), .Z(n580) );
  IV U126 ( .A(B[469]), .Z(n985) );
  IV U127 ( .A(B[65]), .Z(n581) );
  IV U128 ( .A(B[66]), .Z(n582) );
  IV U129 ( .A(B[67]), .Z(n583) );
  IV U130 ( .A(B[68]), .Z(n584) );
  IV U131 ( .A(B[69]), .Z(n585) );
  IV U132 ( .A(B[70]), .Z(n586) );
  IV U133 ( .A(B[71]), .Z(n587) );
  IV U134 ( .A(B[72]), .Z(n588) );
  IV U135 ( .A(B[73]), .Z(n589) );
  IV U136 ( .A(B[74]), .Z(n590) );
  IV U137 ( .A(B[470]), .Z(n986) );
  IV U138 ( .A(B[75]), .Z(n591) );
  IV U139 ( .A(B[76]), .Z(n592) );
  IV U140 ( .A(B[77]), .Z(n593) );
  IV U141 ( .A(B[78]), .Z(n594) );
  IV U142 ( .A(B[79]), .Z(n595) );
  IV U143 ( .A(B[80]), .Z(n596) );
  IV U144 ( .A(B[81]), .Z(n597) );
  IV U145 ( .A(B[82]), .Z(n598) );
  IV U146 ( .A(B[83]), .Z(n599) );
  IV U147 ( .A(B[84]), .Z(n600) );
  IV U148 ( .A(B[471]), .Z(n987) );
  IV U149 ( .A(B[85]), .Z(n601) );
  IV U150 ( .A(B[86]), .Z(n602) );
  IV U151 ( .A(B[87]), .Z(n603) );
  IV U152 ( .A(B[88]), .Z(n604) );
  IV U153 ( .A(B[89]), .Z(n605) );
  IV U154 ( .A(B[90]), .Z(n606) );
  IV U155 ( .A(B[91]), .Z(n607) );
  IV U156 ( .A(B[92]), .Z(n608) );
  IV U157 ( .A(B[93]), .Z(n609) );
  IV U158 ( .A(B[94]), .Z(n610) );
  IV U159 ( .A(B[472]), .Z(n988) );
  IV U160 ( .A(B[95]), .Z(n611) );
  IV U161 ( .A(B[96]), .Z(n612) );
  IV U162 ( .A(B[97]), .Z(n613) );
  IV U163 ( .A(B[98]), .Z(n614) );
  IV U164 ( .A(B[99]), .Z(n615) );
  IV U165 ( .A(B[100]), .Z(n616) );
  IV U166 ( .A(B[101]), .Z(n617) );
  IV U167 ( .A(B[102]), .Z(n618) );
  IV U168 ( .A(B[103]), .Z(n619) );
  IV U169 ( .A(B[104]), .Z(n620) );
  IV U170 ( .A(B[473]), .Z(n989) );
  IV U171 ( .A(B[105]), .Z(n621) );
  IV U172 ( .A(B[106]), .Z(n622) );
  IV U173 ( .A(B[107]), .Z(n623) );
  IV U174 ( .A(B[108]), .Z(n624) );
  IV U175 ( .A(B[109]), .Z(n625) );
  IV U176 ( .A(B[110]), .Z(n626) );
  IV U177 ( .A(B[111]), .Z(n627) );
  IV U178 ( .A(B[112]), .Z(n628) );
  IV U179 ( .A(B[113]), .Z(n629) );
  IV U180 ( .A(B[114]), .Z(n630) );
  IV U181 ( .A(B[474]), .Z(n990) );
  IV U182 ( .A(B[510]), .Z(n1026) );
  IV U183 ( .A(B[115]), .Z(n631) );
  IV U184 ( .A(B[116]), .Z(n632) );
  IV U185 ( .A(B[117]), .Z(n633) );
  IV U186 ( .A(B[118]), .Z(n634) );
  IV U187 ( .A(B[119]), .Z(n635) );
  IV U188 ( .A(B[120]), .Z(n636) );
  IV U189 ( .A(B[121]), .Z(n637) );
  IV U190 ( .A(B[122]), .Z(n638) );
  IV U191 ( .A(B[123]), .Z(n639) );
  IV U192 ( .A(B[124]), .Z(n640) );
  IV U193 ( .A(B[475]), .Z(n991) );
  IV U194 ( .A(B[125]), .Z(n641) );
  IV U195 ( .A(B[126]), .Z(n642) );
  IV U196 ( .A(B[127]), .Z(n643) );
  IV U197 ( .A(B[128]), .Z(n644) );
  IV U198 ( .A(B[129]), .Z(n645) );
  IV U199 ( .A(B[130]), .Z(n646) );
  IV U200 ( .A(B[131]), .Z(n647) );
  IV U201 ( .A(B[132]), .Z(n648) );
  IV U202 ( .A(B[133]), .Z(n649) );
  IV U203 ( .A(B[134]), .Z(n650) );
  IV U204 ( .A(B[476]), .Z(n992) );
  IV U205 ( .A(B[135]), .Z(n651) );
  IV U206 ( .A(B[136]), .Z(n652) );
  IV U207 ( .A(B[137]), .Z(n653) );
  IV U208 ( .A(B[138]), .Z(n654) );
  IV U209 ( .A(B[139]), .Z(n655) );
  IV U210 ( .A(B[140]), .Z(n656) );
  IV U211 ( .A(B[141]), .Z(n657) );
  IV U212 ( .A(B[142]), .Z(n658) );
  IV U213 ( .A(B[143]), .Z(n659) );
  IV U214 ( .A(B[144]), .Z(n660) );
  IV U215 ( .A(B[477]), .Z(n993) );
  IV U216 ( .A(B[145]), .Z(n661) );
  IV U217 ( .A(B[146]), .Z(n662) );
  IV U218 ( .A(B[147]), .Z(n663) );
  IV U219 ( .A(B[148]), .Z(n664) );
  IV U220 ( .A(B[149]), .Z(n665) );
  IV U221 ( .A(B[150]), .Z(n666) );
  IV U222 ( .A(B[151]), .Z(n667) );
  IV U223 ( .A(B[152]), .Z(n668) );
  IV U224 ( .A(B[153]), .Z(n669) );
  IV U225 ( .A(B[154]), .Z(n670) );
  IV U226 ( .A(B[478]), .Z(n994) );
  IV U227 ( .A(B[155]), .Z(n671) );
  IV U228 ( .A(B[156]), .Z(n672) );
  IV U229 ( .A(B[157]), .Z(n673) );
  IV U230 ( .A(B[158]), .Z(n674) );
  IV U231 ( .A(B[159]), .Z(n675) );
  IV U232 ( .A(B[160]), .Z(n676) );
  IV U233 ( .A(B[161]), .Z(n677) );
  IV U234 ( .A(B[162]), .Z(n678) );
  IV U235 ( .A(B[163]), .Z(n679) );
  IV U236 ( .A(B[164]), .Z(n680) );
  IV U237 ( .A(B[479]), .Z(n995) );
  IV U238 ( .A(B[165]), .Z(n681) );
  IV U239 ( .A(B[166]), .Z(n682) );
  IV U240 ( .A(B[167]), .Z(n683) );
  IV U241 ( .A(B[168]), .Z(n684) );
  IV U242 ( .A(B[169]), .Z(n685) );
  IV U243 ( .A(B[170]), .Z(n686) );
  IV U244 ( .A(B[171]), .Z(n687) );
  IV U245 ( .A(B[172]), .Z(n688) );
  IV U246 ( .A(B[173]), .Z(n689) );
  IV U247 ( .A(B[174]), .Z(n690) );
  IV U248 ( .A(B[480]), .Z(n996) );
  IV U249 ( .A(B[175]), .Z(n691) );
  IV U250 ( .A(B[176]), .Z(n692) );
  IV U251 ( .A(B[177]), .Z(n693) );
  IV U252 ( .A(B[178]), .Z(n694) );
  IV U253 ( .A(B[179]), .Z(n695) );
  IV U254 ( .A(B[180]), .Z(n696) );
  IV U255 ( .A(B[181]), .Z(n697) );
  IV U256 ( .A(B[182]), .Z(n698) );
  IV U257 ( .A(B[183]), .Z(n699) );
  IV U258 ( .A(B[184]), .Z(n700) );
  IV U259 ( .A(B[481]), .Z(n997) );
  IV U260 ( .A(B[185]), .Z(n701) );
  IV U261 ( .A(B[186]), .Z(n702) );
  IV U262 ( .A(B[187]), .Z(n703) );
  IV U263 ( .A(B[188]), .Z(n704) );
  IV U264 ( .A(B[189]), .Z(n705) );
  IV U265 ( .A(B[190]), .Z(n706) );
  IV U266 ( .A(B[191]), .Z(n707) );
  IV U267 ( .A(B[192]), .Z(n708) );
  IV U268 ( .A(B[193]), .Z(n709) );
  IV U269 ( .A(B[194]), .Z(n710) );
  IV U270 ( .A(B[482]), .Z(n998) );
  IV U271 ( .A(B[195]), .Z(n711) );
  IV U272 ( .A(B[196]), .Z(n712) );
  IV U273 ( .A(B[197]), .Z(n713) );
  IV U274 ( .A(B[198]), .Z(n714) );
  IV U275 ( .A(B[199]), .Z(n715) );
  IV U276 ( .A(B[200]), .Z(n716) );
  IV U277 ( .A(B[201]), .Z(n717) );
  IV U278 ( .A(B[202]), .Z(n718) );
  IV U279 ( .A(B[203]), .Z(n719) );
  IV U280 ( .A(B[204]), .Z(n720) );
  IV U281 ( .A(B[483]), .Z(n999) );
  IV U282 ( .A(B[205]), .Z(n721) );
  IV U283 ( .A(B[206]), .Z(n722) );
  IV U284 ( .A(B[207]), .Z(n723) );
  IV U285 ( .A(B[208]), .Z(n724) );
  IV U286 ( .A(B[209]), .Z(n725) );
  IV U287 ( .A(B[210]), .Z(n726) );
  IV U288 ( .A(B[211]), .Z(n727) );
  IV U289 ( .A(B[212]), .Z(n728) );
  IV U290 ( .A(B[213]), .Z(n729) );
  IV U291 ( .A(B[214]), .Z(n730) );
  IV U292 ( .A(B[484]), .Z(n1000) );
  IV U293 ( .A(B[511]), .Z(n1027) );
  IV U294 ( .A(B[215]), .Z(n731) );
  IV U295 ( .A(B[216]), .Z(n732) );
  IV U296 ( .A(B[217]), .Z(n733) );
  IV U297 ( .A(B[218]), .Z(n734) );
  IV U298 ( .A(B[219]), .Z(n735) );
  IV U299 ( .A(B[220]), .Z(n736) );
  IV U300 ( .A(B[221]), .Z(n737) );
  IV U301 ( .A(B[222]), .Z(n738) );
  IV U302 ( .A(B[223]), .Z(n739) );
  IV U303 ( .A(B[224]), .Z(n740) );
  IV U304 ( .A(B[485]), .Z(n1001) );
  IV U305 ( .A(B[225]), .Z(n741) );
  IV U306 ( .A(B[226]), .Z(n742) );
  IV U307 ( .A(B[227]), .Z(n743) );
  IV U308 ( .A(B[228]), .Z(n744) );
  IV U309 ( .A(B[229]), .Z(n745) );
  IV U310 ( .A(B[230]), .Z(n746) );
  IV U311 ( .A(B[231]), .Z(n747) );
  IV U312 ( .A(B[232]), .Z(n748) );
  IV U313 ( .A(B[233]), .Z(n749) );
  IV U314 ( .A(B[234]), .Z(n750) );
  IV U315 ( .A(B[486]), .Z(n1002) );
  IV U316 ( .A(B[235]), .Z(n751) );
  IV U317 ( .A(B[236]), .Z(n752) );
  IV U318 ( .A(B[237]), .Z(n753) );
  IV U319 ( .A(B[238]), .Z(n754) );
  IV U320 ( .A(B[239]), .Z(n755) );
  IV U321 ( .A(B[240]), .Z(n756) );
  IV U322 ( .A(B[241]), .Z(n757) );
  IV U323 ( .A(B[242]), .Z(n758) );
  IV U324 ( .A(B[243]), .Z(n759) );
  IV U325 ( .A(B[244]), .Z(n760) );
  IV U326 ( .A(B[487]), .Z(n1003) );
  IV U327 ( .A(B[245]), .Z(n761) );
  IV U328 ( .A(B[246]), .Z(n762) );
  IV U329 ( .A(B[247]), .Z(n763) );
  IV U330 ( .A(B[248]), .Z(n764) );
  IV U331 ( .A(B[249]), .Z(n765) );
  IV U332 ( .A(B[250]), .Z(n766) );
  IV U333 ( .A(B[251]), .Z(n767) );
  IV U334 ( .A(B[252]), .Z(n768) );
  IV U335 ( .A(B[253]), .Z(n769) );
  IV U336 ( .A(B[254]), .Z(n770) );
  IV U337 ( .A(B[488]), .Z(n1004) );
  IV U338 ( .A(B[255]), .Z(n771) );
  IV U339 ( .A(B[256]), .Z(n772) );
  IV U340 ( .A(B[257]), .Z(n773) );
  IV U341 ( .A(B[258]), .Z(n774) );
  IV U342 ( .A(B[259]), .Z(n775) );
  IV U343 ( .A(B[260]), .Z(n776) );
  IV U344 ( .A(B[261]), .Z(n777) );
  IV U345 ( .A(B[262]), .Z(n778) );
  IV U346 ( .A(B[263]), .Z(n779) );
  IV U347 ( .A(B[264]), .Z(n780) );
  IV U348 ( .A(B[489]), .Z(n1005) );
  IV U349 ( .A(B[265]), .Z(n781) );
  IV U350 ( .A(B[266]), .Z(n782) );
  IV U351 ( .A(B[267]), .Z(n783) );
  IV U352 ( .A(B[268]), .Z(n784) );
  IV U353 ( .A(B[269]), .Z(n785) );
  IV U354 ( .A(B[270]), .Z(n786) );
  IV U355 ( .A(B[271]), .Z(n787) );
  IV U356 ( .A(B[272]), .Z(n788) );
  IV U357 ( .A(B[273]), .Z(n789) );
  IV U358 ( .A(B[274]), .Z(n790) );
  IV U359 ( .A(B[490]), .Z(n1006) );
  IV U360 ( .A(B[275]), .Z(n791) );
  IV U361 ( .A(B[276]), .Z(n792) );
  IV U362 ( .A(B[277]), .Z(n793) );
  IV U363 ( .A(B[278]), .Z(n794) );
  IV U364 ( .A(B[279]), .Z(n795) );
  IV U365 ( .A(B[280]), .Z(n796) );
  IV U366 ( .A(B[281]), .Z(n797) );
  IV U367 ( .A(B[282]), .Z(n798) );
  IV U368 ( .A(B[283]), .Z(n799) );
  IV U369 ( .A(B[284]), .Z(n800) );
  IV U370 ( .A(B[491]), .Z(n1007) );
  IV U371 ( .A(B[285]), .Z(n801) );
  IV U372 ( .A(B[286]), .Z(n802) );
  IV U373 ( .A(B[287]), .Z(n803) );
  IV U374 ( .A(B[288]), .Z(n804) );
  IV U375 ( .A(B[289]), .Z(n805) );
  IV U376 ( .A(B[290]), .Z(n806) );
  IV U377 ( .A(B[291]), .Z(n807) );
  IV U378 ( .A(B[292]), .Z(n808) );
  IV U379 ( .A(B[293]), .Z(n809) );
  IV U380 ( .A(B[294]), .Z(n810) );
  IV U381 ( .A(B[492]), .Z(n1008) );
  IV U382 ( .A(B[295]), .Z(n811) );
  IV U383 ( .A(B[296]), .Z(n812) );
  IV U384 ( .A(B[297]), .Z(n813) );
  IV U385 ( .A(B[298]), .Z(n814) );
  IV U386 ( .A(B[299]), .Z(n815) );
  IV U387 ( .A(B[300]), .Z(n816) );
  IV U388 ( .A(B[301]), .Z(n817) );
  IV U389 ( .A(B[302]), .Z(n818) );
  IV U390 ( .A(B[303]), .Z(n819) );
  IV U391 ( .A(B[304]), .Z(n820) );
  IV U392 ( .A(B[493]), .Z(n1009) );
  IV U393 ( .A(B[305]), .Z(n821) );
  IV U394 ( .A(B[306]), .Z(n822) );
  IV U395 ( .A(B[307]), .Z(n823) );
  IV U396 ( .A(B[308]), .Z(n824) );
  IV U397 ( .A(B[309]), .Z(n825) );
  IV U398 ( .A(B[310]), .Z(n826) );
  IV U399 ( .A(B[311]), .Z(n827) );
  IV U400 ( .A(B[312]), .Z(n828) );
  IV U401 ( .A(B[313]), .Z(n829) );
  IV U402 ( .A(B[314]), .Z(n830) );
  IV U403 ( .A(B[494]), .Z(n1010) );
  IV U404 ( .A(B[512]), .Z(n1028) );
  IV U405 ( .A(B[315]), .Z(n831) );
  IV U406 ( .A(B[316]), .Z(n832) );
  IV U407 ( .A(B[317]), .Z(n833) );
  IV U408 ( .A(B[318]), .Z(n834) );
  IV U409 ( .A(B[319]), .Z(n835) );
  IV U410 ( .A(B[320]), .Z(n836) );
  IV U411 ( .A(B[321]), .Z(n837) );
  IV U412 ( .A(B[322]), .Z(n838) );
  IV U413 ( .A(B[323]), .Z(n839) );
  IV U414 ( .A(B[324]), .Z(n840) );
  IV U415 ( .A(B[495]), .Z(n1011) );
  IV U416 ( .A(B[325]), .Z(n841) );
  IV U417 ( .A(B[326]), .Z(n842) );
  IV U418 ( .A(B[327]), .Z(n843) );
  IV U419 ( .A(B[328]), .Z(n844) );
  IV U420 ( .A(B[329]), .Z(n845) );
  IV U421 ( .A(B[330]), .Z(n846) );
  IV U422 ( .A(B[331]), .Z(n847) );
  IV U423 ( .A(B[332]), .Z(n848) );
  IV U424 ( .A(B[333]), .Z(n849) );
  IV U425 ( .A(B[334]), .Z(n850) );
  IV U426 ( .A(B[496]), .Z(n1012) );
  IV U427 ( .A(B[335]), .Z(n851) );
  IV U428 ( .A(B[336]), .Z(n852) );
  IV U429 ( .A(B[337]), .Z(n853) );
  IV U430 ( .A(B[338]), .Z(n854) );
  IV U431 ( .A(B[339]), .Z(n855) );
  IV U432 ( .A(B[340]), .Z(n856) );
  IV U433 ( .A(B[341]), .Z(n857) );
  IV U434 ( .A(B[342]), .Z(n858) );
  IV U435 ( .A(B[343]), .Z(n859) );
  IV U436 ( .A(B[344]), .Z(n860) );
  IV U437 ( .A(B[497]), .Z(n1013) );
  IV U438 ( .A(B[345]), .Z(n861) );
  IV U439 ( .A(B[346]), .Z(n862) );
  IV U440 ( .A(B[347]), .Z(n863) );
  IV U441 ( .A(B[348]), .Z(n864) );
  IV U442 ( .A(B[349]), .Z(n865) );
  IV U443 ( .A(B[350]), .Z(n866) );
  IV U444 ( .A(B[351]), .Z(n867) );
  IV U445 ( .A(B[352]), .Z(n868) );
  IV U446 ( .A(B[353]), .Z(n869) );
  IV U447 ( .A(B[354]), .Z(n870) );
  IV U448 ( .A(B[498]), .Z(n1014) );
  IV U449 ( .A(B[355]), .Z(n871) );
  IV U450 ( .A(B[356]), .Z(n872) );
  IV U451 ( .A(B[357]), .Z(n873) );
  IV U452 ( .A(B[358]), .Z(n874) );
  IV U453 ( .A(B[359]), .Z(n875) );
  IV U454 ( .A(B[360]), .Z(n876) );
  IV U455 ( .A(B[361]), .Z(n877) );
  IV U456 ( .A(B[362]), .Z(n878) );
  IV U457 ( .A(B[363]), .Z(n879) );
  IV U458 ( .A(B[364]), .Z(n880) );
  IV U459 ( .A(B[499]), .Z(n1015) );
  IV U460 ( .A(B[365]), .Z(n881) );
  IV U461 ( .A(B[366]), .Z(n882) );
  IV U462 ( .A(B[367]), .Z(n883) );
  IV U463 ( .A(B[368]), .Z(n884) );
  IV U464 ( .A(B[369]), .Z(n885) );
  IV U465 ( .A(B[370]), .Z(n886) );
  IV U466 ( .A(B[371]), .Z(n887) );
  IV U467 ( .A(B[372]), .Z(n888) );
  IV U468 ( .A(B[373]), .Z(n889) );
  IV U469 ( .A(B[374]), .Z(n890) );
  IV U470 ( .A(B[500]), .Z(n1016) );
  IV U471 ( .A(B[375]), .Z(n891) );
  IV U472 ( .A(B[376]), .Z(n892) );
  IV U473 ( .A(B[377]), .Z(n893) );
  IV U474 ( .A(B[378]), .Z(n894) );
  IV U475 ( .A(B[379]), .Z(n895) );
  IV U476 ( .A(B[380]), .Z(n896) );
  IV U477 ( .A(B[381]), .Z(n897) );
  IV U478 ( .A(B[382]), .Z(n898) );
  IV U479 ( .A(B[383]), .Z(n899) );
  IV U480 ( .A(B[384]), .Z(n900) );
  IV U481 ( .A(B[501]), .Z(n1017) );
  IV U482 ( .A(B[385]), .Z(n901) );
  IV U483 ( .A(B[386]), .Z(n902) );
  IV U484 ( .A(B[387]), .Z(n903) );
  IV U485 ( .A(B[388]), .Z(n904) );
  IV U486 ( .A(B[389]), .Z(n905) );
  IV U487 ( .A(B[390]), .Z(n906) );
  IV U488 ( .A(B[391]), .Z(n907) );
  IV U489 ( .A(B[392]), .Z(n908) );
  IV U490 ( .A(B[393]), .Z(n909) );
  IV U491 ( .A(B[394]), .Z(n910) );
  IV U492 ( .A(B[502]), .Z(n1018) );
  IV U493 ( .A(B[395]), .Z(n911) );
  IV U494 ( .A(B[396]), .Z(n912) );
  IV U495 ( .A(B[397]), .Z(n913) );
  IV U496 ( .A(B[398]), .Z(n914) );
  IV U497 ( .A(B[399]), .Z(n915) );
  IV U498 ( .A(B[400]), .Z(n916) );
  IV U499 ( .A(B[401]), .Z(n917) );
  IV U500 ( .A(B[402]), .Z(n918) );
  IV U501 ( .A(B[403]), .Z(n919) );
  IV U502 ( .A(B[404]), .Z(n920) );
  IV U503 ( .A(B[503]), .Z(n1019) );
  IV U504 ( .A(B[405]), .Z(n921) );
  IV U505 ( .A(B[406]), .Z(n922) );
  IV U506 ( .A(B[407]), .Z(n923) );
  IV U507 ( .A(B[408]), .Z(n924) );
  IV U508 ( .A(B[409]), .Z(n925) );
  IV U509 ( .A(B[410]), .Z(n926) );
  IV U510 ( .A(B[411]), .Z(n927) );
  IV U511 ( .A(B[412]), .Z(n928) );
  IV U512 ( .A(B[413]), .Z(n929) );
  IV U513 ( .A(B[414]), .Z(n930) );
  IV U514 ( .A(B[504]), .Z(n1020) );
  IV U515 ( .A(B[513]), .Z(n1029) );
endmodule


module FA_7979 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_7980 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(CI), .B(A), .Z(CO) );
endmodule


module FA_7981 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7982 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7983 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7984 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7985 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7986 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7987 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7988 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7989 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7990 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7991 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7992 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7993 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7994 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7995 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7996 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7997 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7998 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_7999 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8000 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8001 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8002 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8003 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8004 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8005 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8006 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8007 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8008 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8009 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8010 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8011 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8012 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8013 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8014 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8015 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8016 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8017 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8018 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8019 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8020 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8021 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8022 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8023 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8024 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8025 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8026 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8027 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8028 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8029 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8030 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8031 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8032 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8033 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8034 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8035 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8036 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8037 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8038 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8039 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8040 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8041 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8042 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8043 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8044 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8045 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8046 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8047 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8048 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8049 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8050 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8051 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8052 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8053 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8054 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8055 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8056 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8057 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8058 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8059 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8060 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8061 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8062 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8063 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8064 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8065 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8066 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8067 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8068 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8069 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8070 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8071 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8072 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8073 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8074 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8075 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8076 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8077 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8078 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8079 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8080 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8081 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8082 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8083 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8084 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8085 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8086 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8087 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8088 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8089 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8090 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8091 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8092 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8093 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8094 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8095 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8096 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8097 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8098 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8099 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8100 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8101 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8102 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8103 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8104 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8105 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8106 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8107 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8108 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8109 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8110 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8111 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8112 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8113 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8114 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8115 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8116 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8117 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8118 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8119 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8120 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8121 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8122 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8123 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8124 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8125 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8126 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8127 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8128 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8129 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8130 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8131 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8132 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8133 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8134 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8135 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8136 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8137 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8138 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8139 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8140 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8141 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8142 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8143 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8144 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8145 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8146 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8147 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8148 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8149 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8150 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8151 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8152 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8153 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8154 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8155 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8156 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8157 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8158 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8159 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8160 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8161 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8162 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8163 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8164 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8165 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8166 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8167 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8168 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8169 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8170 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8171 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8172 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8173 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8174 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8175 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8176 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8177 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8178 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8179 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8180 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8181 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8182 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8183 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8184 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8185 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8186 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8187 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8188 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8189 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8190 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8191 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8192 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8193 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8194 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8195 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8196 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8197 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8198 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8199 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8200 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8201 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8202 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8203 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8204 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8205 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8206 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8207 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8208 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8209 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8210 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8211 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8212 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8213 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8214 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8215 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8216 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8217 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8218 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8219 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8220 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8221 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8222 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8223 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8224 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8225 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8226 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8227 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8228 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8229 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8230 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8231 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8232 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8233 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8234 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8235 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8236 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8237 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8238 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8239 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8240 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8241 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8242 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8243 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8244 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8245 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8246 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8247 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8248 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8249 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8250 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8251 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8252 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8253 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8254 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8255 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XOR U1 ( .A(CI), .B(n1), .Z(CO) );
  AND U2 ( .A(n2), .B(n3), .Z(n1) );
  XOR U3 ( .A(CI), .B(A), .Z(n3) );
  XOR U4 ( .A(CI), .B(B), .Z(n2) );
endmodule


module FA_8492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  OR U1 ( .A(B), .B(A), .Z(CO) );
endmodule


module COMP_N514_4 ( A, B, O );
  input [513:0] A;
  input [513:0] B;
  output O;
  wire   n2, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  wire   [513:1] C;

  FA_8492 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .CO(
        C[1]) );
  FA_8491 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n514), .CI(C[1]), 
        .CO(C[2]) );
  FA_8490 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n515), .CI(C[2]), 
        .CO(C[3]) );
  FA_8489 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n516), .CI(C[3]), 
        .CO(C[4]) );
  FA_8488 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n517), .CI(C[4]), 
        .CO(C[5]) );
  FA_8487 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n518), .CI(C[5]), 
        .CO(C[6]) );
  FA_8486 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n519), .CI(C[6]), 
        .CO(C[7]) );
  FA_8485 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n520), .CI(C[7]), 
        .CO(C[8]) );
  FA_8484 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n521), .CI(C[8]), 
        .CO(C[9]) );
  FA_8483 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n522), .CI(C[9]), 
        .CO(C[10]) );
  FA_8482 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n523), .CI(C[10]), 
        .CO(C[11]) );
  FA_8481 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n524), .CI(C[11]), 
        .CO(C[12]) );
  FA_8480 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n525), .CI(C[12]), 
        .CO(C[13]) );
  FA_8479 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n526), .CI(C[13]), 
        .CO(C[14]) );
  FA_8478 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n527), .CI(C[14]), 
        .CO(C[15]) );
  FA_8477 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n528), .CI(C[15]), 
        .CO(C[16]) );
  FA_8476 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n529), .CI(C[16]), 
        .CO(C[17]) );
  FA_8475 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n530), .CI(C[17]), 
        .CO(C[18]) );
  FA_8474 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n531), .CI(C[18]), 
        .CO(C[19]) );
  FA_8473 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n532), .CI(C[19]), 
        .CO(C[20]) );
  FA_8472 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n533), .CI(C[20]), 
        .CO(C[21]) );
  FA_8471 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n534), .CI(C[21]), 
        .CO(C[22]) );
  FA_8470 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n535), .CI(C[22]), 
        .CO(C[23]) );
  FA_8469 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n536), .CI(C[23]), 
        .CO(C[24]) );
  FA_8468 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n537), .CI(C[24]), 
        .CO(C[25]) );
  FA_8467 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n538), .CI(C[25]), 
        .CO(C[26]) );
  FA_8466 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n539), .CI(C[26]), 
        .CO(C[27]) );
  FA_8465 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n540), .CI(C[27]), 
        .CO(C[28]) );
  FA_8464 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n541), .CI(C[28]), 
        .CO(C[29]) );
  FA_8463 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n542), .CI(C[29]), 
        .CO(C[30]) );
  FA_8462 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n543), .CI(C[30]), 
        .CO(C[31]) );
  FA_8461 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n544), .CI(C[31]), 
        .CO(C[32]) );
  FA_8460 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n545), .CI(C[32]), 
        .CO(C[33]) );
  FA_8459 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n546), .CI(C[33]), 
        .CO(C[34]) );
  FA_8458 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n547), .CI(C[34]), 
        .CO(C[35]) );
  FA_8457 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n548), .CI(C[35]), 
        .CO(C[36]) );
  FA_8456 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n549), .CI(C[36]), 
        .CO(C[37]) );
  FA_8455 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n550), .CI(C[37]), 
        .CO(C[38]) );
  FA_8454 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n551), .CI(C[38]), 
        .CO(C[39]) );
  FA_8453 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n552), .CI(C[39]), 
        .CO(C[40]) );
  FA_8452 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n553), .CI(C[40]), 
        .CO(C[41]) );
  FA_8451 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n554), .CI(C[41]), 
        .CO(C[42]) );
  FA_8450 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n555), .CI(C[42]), 
        .CO(C[43]) );
  FA_8449 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n556), .CI(C[43]), 
        .CO(C[44]) );
  FA_8448 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n557), .CI(C[44]), 
        .CO(C[45]) );
  FA_8447 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n558), .CI(C[45]), 
        .CO(C[46]) );
  FA_8446 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n559), .CI(C[46]), 
        .CO(C[47]) );
  FA_8445 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n560), .CI(C[47]), 
        .CO(C[48]) );
  FA_8444 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n561), .CI(C[48]), 
        .CO(C[49]) );
  FA_8443 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n562), .CI(C[49]), 
        .CO(C[50]) );
  FA_8442 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n563), .CI(C[50]), 
        .CO(C[51]) );
  FA_8441 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n564), .CI(C[51]), 
        .CO(C[52]) );
  FA_8440 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n565), .CI(C[52]), 
        .CO(C[53]) );
  FA_8439 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n566), .CI(C[53]), 
        .CO(C[54]) );
  FA_8438 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n567), .CI(C[54]), 
        .CO(C[55]) );
  FA_8437 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n568), .CI(C[55]), 
        .CO(C[56]) );
  FA_8436 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n569), .CI(C[56]), 
        .CO(C[57]) );
  FA_8435 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n570), .CI(C[57]), 
        .CO(C[58]) );
  FA_8434 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n571), .CI(C[58]), 
        .CO(C[59]) );
  FA_8433 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n572), .CI(C[59]), 
        .CO(C[60]) );
  FA_8432 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n573), .CI(C[60]), 
        .CO(C[61]) );
  FA_8431 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n574), .CI(C[61]), 
        .CO(C[62]) );
  FA_8430 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n575), .CI(C[62]), 
        .CO(C[63]) );
  FA_8429 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n576), .CI(C[63]), 
        .CO(C[64]) );
  FA_8428 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n577), .CI(C[64]), 
        .CO(C[65]) );
  FA_8427 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n578), .CI(C[65]), 
        .CO(C[66]) );
  FA_8426 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n579), .CI(C[66]), 
        .CO(C[67]) );
  FA_8425 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n580), .CI(C[67]), 
        .CO(C[68]) );
  FA_8424 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n581), .CI(C[68]), 
        .CO(C[69]) );
  FA_8423 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n582), .CI(C[69]), 
        .CO(C[70]) );
  FA_8422 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n583), .CI(C[70]), 
        .CO(C[71]) );
  FA_8421 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n584), .CI(C[71]), 
        .CO(C[72]) );
  FA_8420 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n585), .CI(C[72]), 
        .CO(C[73]) );
  FA_8419 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n586), .CI(C[73]), 
        .CO(C[74]) );
  FA_8418 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n587), .CI(C[74]), 
        .CO(C[75]) );
  FA_8417 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n588), .CI(C[75]), 
        .CO(C[76]) );
  FA_8416 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n589), .CI(C[76]), 
        .CO(C[77]) );
  FA_8415 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n590), .CI(C[77]), 
        .CO(C[78]) );
  FA_8414 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n591), .CI(C[78]), 
        .CO(C[79]) );
  FA_8413 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n592), .CI(C[79]), 
        .CO(C[80]) );
  FA_8412 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n593), .CI(C[80]), 
        .CO(C[81]) );
  FA_8411 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n594), .CI(C[81]), 
        .CO(C[82]) );
  FA_8410 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n595), .CI(C[82]), 
        .CO(C[83]) );
  FA_8409 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n596), .CI(C[83]), 
        .CO(C[84]) );
  FA_8408 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n597), .CI(C[84]), 
        .CO(C[85]) );
  FA_8407 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n598), .CI(C[85]), 
        .CO(C[86]) );
  FA_8406 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n599), .CI(C[86]), 
        .CO(C[87]) );
  FA_8405 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n600), .CI(C[87]), 
        .CO(C[88]) );
  FA_8404 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n601), .CI(C[88]), 
        .CO(C[89]) );
  FA_8403 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n602), .CI(C[89]), 
        .CO(C[90]) );
  FA_8402 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n603), .CI(C[90]), 
        .CO(C[91]) );
  FA_8401 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n604), .CI(C[91]), 
        .CO(C[92]) );
  FA_8400 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n605), .CI(C[92]), 
        .CO(C[93]) );
  FA_8399 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n606), .CI(C[93]), 
        .CO(C[94]) );
  FA_8398 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n607), .CI(C[94]), 
        .CO(C[95]) );
  FA_8397 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n608), .CI(C[95]), 
        .CO(C[96]) );
  FA_8396 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n609), .CI(C[96]), 
        .CO(C[97]) );
  FA_8395 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n610), .CI(C[97]), 
        .CO(C[98]) );
  FA_8394 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n611), .CI(C[98]), 
        .CO(C[99]) );
  FA_8393 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n612), .CI(C[99]), 
        .CO(C[100]) );
  FA_8392 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n613), .CI(C[100]), .CO(C[101]) );
  FA_8391 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n614), .CI(C[101]), .CO(C[102]) );
  FA_8390 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n615), .CI(C[102]), .CO(C[103]) );
  FA_8389 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n616), .CI(C[103]), .CO(C[104]) );
  FA_8388 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n617), .CI(C[104]), .CO(C[105]) );
  FA_8387 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n618), .CI(C[105]), .CO(C[106]) );
  FA_8386 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n619), .CI(C[106]), .CO(C[107]) );
  FA_8385 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n620), .CI(C[107]), .CO(C[108]) );
  FA_8384 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n621), .CI(C[108]), .CO(C[109]) );
  FA_8383 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n622), .CI(C[109]), .CO(C[110]) );
  FA_8382 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n623), .CI(C[110]), .CO(C[111]) );
  FA_8381 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n624), .CI(C[111]), .CO(C[112]) );
  FA_8380 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n625), .CI(C[112]), .CO(C[113]) );
  FA_8379 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n626), .CI(C[113]), .CO(C[114]) );
  FA_8378 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n627), .CI(C[114]), .CO(C[115]) );
  FA_8377 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n628), .CI(C[115]), .CO(C[116]) );
  FA_8376 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n629), .CI(C[116]), .CO(C[117]) );
  FA_8375 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n630), .CI(C[117]), .CO(C[118]) );
  FA_8374 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n631), .CI(C[118]), .CO(C[119]) );
  FA_8373 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n632), .CI(C[119]), .CO(C[120]) );
  FA_8372 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n633), .CI(C[120]), .CO(C[121]) );
  FA_8371 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n634), .CI(C[121]), .CO(C[122]) );
  FA_8370 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n635), .CI(C[122]), .CO(C[123]) );
  FA_8369 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n636), .CI(C[123]), .CO(C[124]) );
  FA_8368 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n637), .CI(C[124]), .CO(C[125]) );
  FA_8367 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n638), .CI(C[125]), .CO(C[126]) );
  FA_8366 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n639), .CI(C[126]), .CO(C[127]) );
  FA_8365 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n640), .CI(C[127]), .CO(C[128]) );
  FA_8364 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n641), .CI(C[128]), .CO(C[129]) );
  FA_8363 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n642), .CI(C[129]), .CO(C[130]) );
  FA_8362 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n643), .CI(C[130]), .CO(C[131]) );
  FA_8361 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n644), .CI(C[131]), .CO(C[132]) );
  FA_8360 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n645), .CI(C[132]), .CO(C[133]) );
  FA_8359 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n646), .CI(C[133]), .CO(C[134]) );
  FA_8358 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n647), .CI(C[134]), .CO(C[135]) );
  FA_8357 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n648), .CI(C[135]), .CO(C[136]) );
  FA_8356 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n649), .CI(C[136]), .CO(C[137]) );
  FA_8355 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n650), .CI(C[137]), .CO(C[138]) );
  FA_8354 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n651), .CI(C[138]), .CO(C[139]) );
  FA_8353 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n652), .CI(C[139]), .CO(C[140]) );
  FA_8352 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n653), .CI(C[140]), .CO(C[141]) );
  FA_8351 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n654), .CI(C[141]), .CO(C[142]) );
  FA_8350 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n655), .CI(C[142]), .CO(C[143]) );
  FA_8349 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n656), .CI(C[143]), .CO(C[144]) );
  FA_8348 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n657), .CI(C[144]), .CO(C[145]) );
  FA_8347 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n658), .CI(C[145]), .CO(C[146]) );
  FA_8346 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n659), .CI(C[146]), .CO(C[147]) );
  FA_8345 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n660), .CI(C[147]), .CO(C[148]) );
  FA_8344 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n661), .CI(C[148]), .CO(C[149]) );
  FA_8343 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n662), .CI(C[149]), .CO(C[150]) );
  FA_8342 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n663), .CI(C[150]), .CO(C[151]) );
  FA_8341 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n664), .CI(C[151]), .CO(C[152]) );
  FA_8340 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n665), .CI(C[152]), .CO(C[153]) );
  FA_8339 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n666), .CI(C[153]), .CO(C[154]) );
  FA_8338 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n667), .CI(C[154]), .CO(C[155]) );
  FA_8337 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n668), .CI(C[155]), .CO(C[156]) );
  FA_8336 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n669), .CI(C[156]), .CO(C[157]) );
  FA_8335 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n670), .CI(C[157]), .CO(C[158]) );
  FA_8334 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n671), .CI(C[158]), .CO(C[159]) );
  FA_8333 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n672), .CI(C[159]), .CO(C[160]) );
  FA_8332 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n673), .CI(C[160]), .CO(C[161]) );
  FA_8331 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n674), .CI(C[161]), .CO(C[162]) );
  FA_8330 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n675), .CI(C[162]), .CO(C[163]) );
  FA_8329 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n676), .CI(C[163]), .CO(C[164]) );
  FA_8328 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n677), .CI(C[164]), .CO(C[165]) );
  FA_8327 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n678), .CI(C[165]), .CO(C[166]) );
  FA_8326 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n679), .CI(C[166]), .CO(C[167]) );
  FA_8325 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n680), .CI(C[167]), .CO(C[168]) );
  FA_8324 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n681), .CI(C[168]), .CO(C[169]) );
  FA_8323 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n682), .CI(C[169]), .CO(C[170]) );
  FA_8322 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n683), .CI(C[170]), .CO(C[171]) );
  FA_8321 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n684), .CI(C[171]), .CO(C[172]) );
  FA_8320 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n685), .CI(C[172]), .CO(C[173]) );
  FA_8319 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n686), .CI(C[173]), .CO(C[174]) );
  FA_8318 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n687), .CI(C[174]), .CO(C[175]) );
  FA_8317 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n688), .CI(C[175]), .CO(C[176]) );
  FA_8316 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n689), .CI(C[176]), .CO(C[177]) );
  FA_8315 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n690), .CI(C[177]), .CO(C[178]) );
  FA_8314 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n691), .CI(C[178]), .CO(C[179]) );
  FA_8313 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n692), .CI(C[179]), .CO(C[180]) );
  FA_8312 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n693), .CI(C[180]), .CO(C[181]) );
  FA_8311 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n694), .CI(C[181]), .CO(C[182]) );
  FA_8310 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n695), .CI(C[182]), .CO(C[183]) );
  FA_8309 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n696), .CI(C[183]), .CO(C[184]) );
  FA_8308 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n697), .CI(C[184]), .CO(C[185]) );
  FA_8307 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n698), .CI(C[185]), .CO(C[186]) );
  FA_8306 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n699), .CI(C[186]), .CO(C[187]) );
  FA_8305 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n700), .CI(C[187]), .CO(C[188]) );
  FA_8304 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n701), .CI(C[188]), .CO(C[189]) );
  FA_8303 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n702), .CI(C[189]), .CO(C[190]) );
  FA_8302 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n703), .CI(C[190]), .CO(C[191]) );
  FA_8301 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n704), .CI(C[191]), .CO(C[192]) );
  FA_8300 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n705), .CI(C[192]), .CO(C[193]) );
  FA_8299 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n706), .CI(C[193]), .CO(C[194]) );
  FA_8298 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n707), .CI(C[194]), .CO(C[195]) );
  FA_8297 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n708), .CI(C[195]), .CO(C[196]) );
  FA_8296 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n709), .CI(C[196]), .CO(C[197]) );
  FA_8295 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n710), .CI(C[197]), .CO(C[198]) );
  FA_8294 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n711), .CI(C[198]), .CO(C[199]) );
  FA_8293 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n712), .CI(C[199]), .CO(C[200]) );
  FA_8292 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n713), .CI(C[200]), .CO(C[201]) );
  FA_8291 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n714), .CI(C[201]), .CO(C[202]) );
  FA_8290 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n715), .CI(C[202]), .CO(C[203]) );
  FA_8289 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n716), .CI(C[203]), .CO(C[204]) );
  FA_8288 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n717), .CI(C[204]), .CO(C[205]) );
  FA_8287 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n718), .CI(C[205]), .CO(C[206]) );
  FA_8286 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n719), .CI(C[206]), .CO(C[207]) );
  FA_8285 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n720), .CI(C[207]), .CO(C[208]) );
  FA_8284 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n721), .CI(C[208]), .CO(C[209]) );
  FA_8283 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n722), .CI(C[209]), .CO(C[210]) );
  FA_8282 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n723), .CI(C[210]), .CO(C[211]) );
  FA_8281 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n724), .CI(C[211]), .CO(C[212]) );
  FA_8280 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n725), .CI(C[212]), .CO(C[213]) );
  FA_8279 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n726), .CI(C[213]), .CO(C[214]) );
  FA_8278 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n727), .CI(C[214]), .CO(C[215]) );
  FA_8277 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n728), .CI(C[215]), .CO(C[216]) );
  FA_8276 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n729), .CI(C[216]), .CO(C[217]) );
  FA_8275 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n730), .CI(C[217]), .CO(C[218]) );
  FA_8274 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n731), .CI(C[218]), .CO(C[219]) );
  FA_8273 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n732), .CI(C[219]), .CO(C[220]) );
  FA_8272 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n733), .CI(C[220]), .CO(C[221]) );
  FA_8271 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n734), .CI(C[221]), .CO(C[222]) );
  FA_8270 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n735), .CI(C[222]), .CO(C[223]) );
  FA_8269 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n736), .CI(C[223]), .CO(C[224]) );
  FA_8268 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n737), .CI(C[224]), .CO(C[225]) );
  FA_8267 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n738), .CI(C[225]), .CO(C[226]) );
  FA_8266 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n739), .CI(C[226]), .CO(C[227]) );
  FA_8265 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n740), .CI(C[227]), .CO(C[228]) );
  FA_8264 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n741), .CI(C[228]), .CO(C[229]) );
  FA_8263 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n742), .CI(C[229]), .CO(C[230]) );
  FA_8262 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n743), .CI(C[230]), .CO(C[231]) );
  FA_8261 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n744), .CI(C[231]), .CO(C[232]) );
  FA_8260 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n745), .CI(C[232]), .CO(C[233]) );
  FA_8259 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n746), .CI(C[233]), .CO(C[234]) );
  FA_8258 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n747), .CI(C[234]), .CO(C[235]) );
  FA_8257 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n748), .CI(C[235]), .CO(C[236]) );
  FA_8256 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n749), .CI(C[236]), .CO(C[237]) );
  FA_8255 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n750), .CI(C[237]), .CO(C[238]) );
  FA_8254 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n751), .CI(C[238]), .CO(C[239]) );
  FA_8253 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n752), .CI(C[239]), .CO(C[240]) );
  FA_8252 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n753), .CI(C[240]), .CO(C[241]) );
  FA_8251 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n754), .CI(C[241]), .CO(C[242]) );
  FA_8250 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n755), .CI(C[242]), .CO(C[243]) );
  FA_8249 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n756), .CI(C[243]), .CO(C[244]) );
  FA_8248 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n757), .CI(C[244]), .CO(C[245]) );
  FA_8247 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n758), .CI(C[245]), .CO(C[246]) );
  FA_8246 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n759), .CI(C[246]), .CO(C[247]) );
  FA_8245 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n760), .CI(C[247]), .CO(C[248]) );
  FA_8244 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n761), .CI(C[248]), .CO(C[249]) );
  FA_8243 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n762), .CI(C[249]), .CO(C[250]) );
  FA_8242 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n763), .CI(C[250]), .CO(C[251]) );
  FA_8241 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n764), .CI(C[251]), .CO(C[252]) );
  FA_8240 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n765), .CI(C[252]), .CO(C[253]) );
  FA_8239 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n766), .CI(C[253]), .CO(C[254]) );
  FA_8238 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n767), .CI(C[254]), .CO(C[255]) );
  FA_8237 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n768), .CI(C[255]), .CO(C[256]) );
  FA_8236 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n769), .CI(C[256]), .CO(C[257]) );
  FA_8235 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n770), .CI(C[257]), .CO(C[258]) );
  FA_8234 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n771), .CI(C[258]), .CO(C[259]) );
  FA_8233 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n772), .CI(C[259]), .CO(C[260]) );
  FA_8232 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n773), .CI(C[260]), .CO(C[261]) );
  FA_8231 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n774), .CI(C[261]), .CO(C[262]) );
  FA_8230 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n775), .CI(C[262]), .CO(C[263]) );
  FA_8229 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n776), .CI(C[263]), .CO(C[264]) );
  FA_8228 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n777), .CI(C[264]), .CO(C[265]) );
  FA_8227 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n778), .CI(C[265]), .CO(C[266]) );
  FA_8226 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n779), .CI(C[266]), .CO(C[267]) );
  FA_8225 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n780), .CI(C[267]), .CO(C[268]) );
  FA_8224 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n781), .CI(C[268]), .CO(C[269]) );
  FA_8223 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n782), .CI(C[269]), .CO(C[270]) );
  FA_8222 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n783), .CI(C[270]), .CO(C[271]) );
  FA_8221 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n784), .CI(C[271]), .CO(C[272]) );
  FA_8220 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n785), .CI(C[272]), .CO(C[273]) );
  FA_8219 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n786), .CI(C[273]), .CO(C[274]) );
  FA_8218 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n787), .CI(C[274]), .CO(C[275]) );
  FA_8217 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n788), .CI(C[275]), .CO(C[276]) );
  FA_8216 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n789), .CI(C[276]), .CO(C[277]) );
  FA_8215 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n790), .CI(C[277]), .CO(C[278]) );
  FA_8214 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n791), .CI(C[278]), .CO(C[279]) );
  FA_8213 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n792), .CI(C[279]), .CO(C[280]) );
  FA_8212 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n793), .CI(C[280]), .CO(C[281]) );
  FA_8211 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n794), .CI(C[281]), .CO(C[282]) );
  FA_8210 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n795), .CI(C[282]), .CO(C[283]) );
  FA_8209 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n796), .CI(C[283]), .CO(C[284]) );
  FA_8208 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n797), .CI(C[284]), .CO(C[285]) );
  FA_8207 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n798), .CI(C[285]), .CO(C[286]) );
  FA_8206 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n799), .CI(C[286]), .CO(C[287]) );
  FA_8205 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n800), .CI(C[287]), .CO(C[288]) );
  FA_8204 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n801), .CI(C[288]), .CO(C[289]) );
  FA_8203 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n802), .CI(C[289]), .CO(C[290]) );
  FA_8202 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n803), .CI(C[290]), .CO(C[291]) );
  FA_8201 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n804), .CI(C[291]), .CO(C[292]) );
  FA_8200 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n805), .CI(C[292]), .CO(C[293]) );
  FA_8199 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n806), .CI(C[293]), .CO(C[294]) );
  FA_8198 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n807), .CI(C[294]), .CO(C[295]) );
  FA_8197 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n808), .CI(C[295]), .CO(C[296]) );
  FA_8196 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n809), .CI(C[296]), .CO(C[297]) );
  FA_8195 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n810), .CI(C[297]), .CO(C[298]) );
  FA_8194 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n811), .CI(C[298]), .CO(C[299]) );
  FA_8193 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n812), .CI(C[299]), .CO(C[300]) );
  FA_8192 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n813), .CI(C[300]), .CO(C[301]) );
  FA_8191 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n814), .CI(C[301]), .CO(C[302]) );
  FA_8190 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n815), .CI(C[302]), .CO(C[303]) );
  FA_8189 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n816), .CI(C[303]), .CO(C[304]) );
  FA_8188 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n817), .CI(C[304]), .CO(C[305]) );
  FA_8187 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n818), .CI(C[305]), .CO(C[306]) );
  FA_8186 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n819), .CI(C[306]), .CO(C[307]) );
  FA_8185 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n820), .CI(C[307]), .CO(C[308]) );
  FA_8184 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n821), .CI(C[308]), .CO(C[309]) );
  FA_8183 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n822), .CI(C[309]), .CO(C[310]) );
  FA_8182 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n823), .CI(C[310]), .CO(C[311]) );
  FA_8181 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n824), .CI(C[311]), .CO(C[312]) );
  FA_8180 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n825), .CI(C[312]), .CO(C[313]) );
  FA_8179 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n826), .CI(C[313]), .CO(C[314]) );
  FA_8178 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n827), .CI(C[314]), .CO(C[315]) );
  FA_8177 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n828), .CI(C[315]), .CO(C[316]) );
  FA_8176 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n829), .CI(C[316]), .CO(C[317]) );
  FA_8175 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n830), .CI(C[317]), .CO(C[318]) );
  FA_8174 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n831), .CI(C[318]), .CO(C[319]) );
  FA_8173 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n832), .CI(C[319]), .CO(C[320]) );
  FA_8172 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n833), .CI(C[320]), .CO(C[321]) );
  FA_8171 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n834), .CI(C[321]), .CO(C[322]) );
  FA_8170 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n835), .CI(C[322]), .CO(C[323]) );
  FA_8169 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n836), .CI(C[323]), .CO(C[324]) );
  FA_8168 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n837), .CI(C[324]), .CO(C[325]) );
  FA_8167 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n838), .CI(C[325]), .CO(C[326]) );
  FA_8166 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n839), .CI(C[326]), .CO(C[327]) );
  FA_8165 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n840), .CI(C[327]), .CO(C[328]) );
  FA_8164 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n841), .CI(C[328]), .CO(C[329]) );
  FA_8163 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n842), .CI(C[329]), .CO(C[330]) );
  FA_8162 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n843), .CI(C[330]), .CO(C[331]) );
  FA_8161 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n844), .CI(C[331]), .CO(C[332]) );
  FA_8160 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n845), .CI(C[332]), .CO(C[333]) );
  FA_8159 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n846), .CI(C[333]), .CO(C[334]) );
  FA_8158 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n847), .CI(C[334]), .CO(C[335]) );
  FA_8157 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n848), .CI(C[335]), .CO(C[336]) );
  FA_8156 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n849), .CI(C[336]), .CO(C[337]) );
  FA_8155 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n850), .CI(C[337]), .CO(C[338]) );
  FA_8154 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n851), .CI(C[338]), .CO(C[339]) );
  FA_8153 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n852), .CI(C[339]), .CO(C[340]) );
  FA_8152 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n853), .CI(C[340]), .CO(C[341]) );
  FA_8151 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n854), .CI(C[341]), .CO(C[342]) );
  FA_8150 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n855), .CI(C[342]), .CO(C[343]) );
  FA_8149 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n856), .CI(C[343]), .CO(C[344]) );
  FA_8148 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n857), .CI(C[344]), .CO(C[345]) );
  FA_8147 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n858), .CI(C[345]), .CO(C[346]) );
  FA_8146 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n859), .CI(C[346]), .CO(C[347]) );
  FA_8145 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n860), .CI(C[347]), .CO(C[348]) );
  FA_8144 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n861), .CI(C[348]), .CO(C[349]) );
  FA_8143 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n862), .CI(C[349]), .CO(C[350]) );
  FA_8142 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n863), .CI(C[350]), .CO(C[351]) );
  FA_8141 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n864), .CI(C[351]), .CO(C[352]) );
  FA_8140 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n865), .CI(C[352]), .CO(C[353]) );
  FA_8139 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n866), .CI(C[353]), .CO(C[354]) );
  FA_8138 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n867), .CI(C[354]), .CO(C[355]) );
  FA_8137 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n868), .CI(C[355]), .CO(C[356]) );
  FA_8136 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n869), .CI(C[356]), .CO(C[357]) );
  FA_8135 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n870), .CI(C[357]), .CO(C[358]) );
  FA_8134 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n871), .CI(C[358]), .CO(C[359]) );
  FA_8133 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n872), .CI(C[359]), .CO(C[360]) );
  FA_8132 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n873), .CI(C[360]), .CO(C[361]) );
  FA_8131 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n874), .CI(C[361]), .CO(C[362]) );
  FA_8130 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n875), .CI(C[362]), .CO(C[363]) );
  FA_8129 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n876), .CI(C[363]), .CO(C[364]) );
  FA_8128 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n877), .CI(C[364]), .CO(C[365]) );
  FA_8127 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n878), .CI(C[365]), .CO(C[366]) );
  FA_8126 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n879), .CI(C[366]), .CO(C[367]) );
  FA_8125 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n880), .CI(C[367]), .CO(C[368]) );
  FA_8124 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n881), .CI(C[368]), .CO(C[369]) );
  FA_8123 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n882), .CI(C[369]), .CO(C[370]) );
  FA_8122 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n883), .CI(C[370]), .CO(C[371]) );
  FA_8121 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n884), .CI(C[371]), .CO(C[372]) );
  FA_8120 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n885), .CI(C[372]), .CO(C[373]) );
  FA_8119 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n886), .CI(C[373]), .CO(C[374]) );
  FA_8118 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n887), .CI(C[374]), .CO(C[375]) );
  FA_8117 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n888), .CI(C[375]), .CO(C[376]) );
  FA_8116 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n889), .CI(C[376]), .CO(C[377]) );
  FA_8115 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n890), .CI(C[377]), .CO(C[378]) );
  FA_8114 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n891), .CI(C[378]), .CO(C[379]) );
  FA_8113 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n892), .CI(C[379]), .CO(C[380]) );
  FA_8112 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n893), .CI(C[380]), .CO(C[381]) );
  FA_8111 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n894), .CI(C[381]), .CO(C[382]) );
  FA_8110 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n895), .CI(C[382]), .CO(C[383]) );
  FA_8109 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n896), .CI(C[383]), .CO(C[384]) );
  FA_8108 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n897), .CI(C[384]), .CO(C[385]) );
  FA_8107 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n898), .CI(C[385]), .CO(C[386]) );
  FA_8106 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n899), .CI(C[386]), .CO(C[387]) );
  FA_8105 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n900), .CI(C[387]), .CO(C[388]) );
  FA_8104 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n901), .CI(C[388]), .CO(C[389]) );
  FA_8103 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n902), .CI(C[389]), .CO(C[390]) );
  FA_8102 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n903), .CI(C[390]), .CO(C[391]) );
  FA_8101 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n904), .CI(C[391]), .CO(C[392]) );
  FA_8100 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n905), .CI(C[392]), .CO(C[393]) );
  FA_8099 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n906), .CI(C[393]), .CO(C[394]) );
  FA_8098 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n907), .CI(C[394]), .CO(C[395]) );
  FA_8097 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n908), .CI(C[395]), .CO(C[396]) );
  FA_8096 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n909), .CI(C[396]), .CO(C[397]) );
  FA_8095 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n910), .CI(C[397]), .CO(C[398]) );
  FA_8094 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n911), .CI(C[398]), .CO(C[399]) );
  FA_8093 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n912), .CI(C[399]), .CO(C[400]) );
  FA_8092 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n913), .CI(C[400]), .CO(C[401]) );
  FA_8091 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n914), .CI(C[401]), .CO(C[402]) );
  FA_8090 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n915), .CI(C[402]), .CO(C[403]) );
  FA_8089 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n916), .CI(C[403]), .CO(C[404]) );
  FA_8088 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n917), .CI(C[404]), .CO(C[405]) );
  FA_8087 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n918), .CI(C[405]), .CO(C[406]) );
  FA_8086 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n919), .CI(C[406]), .CO(C[407]) );
  FA_8085 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n920), .CI(C[407]), .CO(C[408]) );
  FA_8084 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n921), .CI(C[408]), .CO(C[409]) );
  FA_8083 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n922), .CI(C[409]), .CO(C[410]) );
  FA_8082 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n923), .CI(C[410]), .CO(C[411]) );
  FA_8081 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n924), .CI(C[411]), .CO(C[412]) );
  FA_8080 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n925), .CI(C[412]), .CO(C[413]) );
  FA_8079 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n926), .CI(C[413]), .CO(C[414]) );
  FA_8078 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n927), .CI(C[414]), .CO(C[415]) );
  FA_8077 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n928), .CI(C[415]), .CO(C[416]) );
  FA_8076 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n929), .CI(C[416]), .CO(C[417]) );
  FA_8075 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n930), .CI(C[417]), .CO(C[418]) );
  FA_8074 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n931), .CI(C[418]), .CO(C[419]) );
  FA_8073 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n932), .CI(C[419]), .CO(C[420]) );
  FA_8072 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n933), .CI(C[420]), .CO(C[421]) );
  FA_8071 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n934), .CI(C[421]), .CO(C[422]) );
  FA_8070 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n935), .CI(C[422]), .CO(C[423]) );
  FA_8069 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n936), .CI(C[423]), .CO(C[424]) );
  FA_8068 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n937), .CI(C[424]), .CO(C[425]) );
  FA_8067 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n938), .CI(C[425]), .CO(C[426]) );
  FA_8066 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n939), .CI(C[426]), .CO(C[427]) );
  FA_8065 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n940), .CI(C[427]), .CO(C[428]) );
  FA_8064 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n941), .CI(C[428]), .CO(C[429]) );
  FA_8063 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n942), .CI(C[429]), .CO(C[430]) );
  FA_8062 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n943), .CI(C[430]), .CO(C[431]) );
  FA_8061 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n944), .CI(C[431]), .CO(C[432]) );
  FA_8060 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n945), .CI(C[432]), .CO(C[433]) );
  FA_8059 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n946), .CI(C[433]), .CO(C[434]) );
  FA_8058 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n947), .CI(C[434]), .CO(C[435]) );
  FA_8057 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n948), .CI(C[435]), .CO(C[436]) );
  FA_8056 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n949), .CI(C[436]), .CO(C[437]) );
  FA_8055 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n950), .CI(C[437]), .CO(C[438]) );
  FA_8054 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n951), .CI(C[438]), .CO(C[439]) );
  FA_8053 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n952), .CI(C[439]), .CO(C[440]) );
  FA_8052 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n953), .CI(C[440]), .CO(C[441]) );
  FA_8051 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n954), .CI(C[441]), .CO(C[442]) );
  FA_8050 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n955), .CI(C[442]), .CO(C[443]) );
  FA_8049 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n956), .CI(C[443]), .CO(C[444]) );
  FA_8048 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n957), .CI(C[444]), .CO(C[445]) );
  FA_8047 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n958), .CI(C[445]), .CO(C[446]) );
  FA_8046 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n959), .CI(C[446]), .CO(C[447]) );
  FA_8045 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n960), .CI(C[447]), .CO(C[448]) );
  FA_8044 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n961), .CI(C[448]), .CO(C[449]) );
  FA_8043 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n962), .CI(C[449]), .CO(C[450]) );
  FA_8042 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n963), .CI(C[450]), .CO(C[451]) );
  FA_8041 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n964), .CI(C[451]), .CO(C[452]) );
  FA_8040 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n965), .CI(C[452]), .CO(C[453]) );
  FA_8039 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n966), .CI(C[453]), .CO(C[454]) );
  FA_8038 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n967), .CI(C[454]), .CO(C[455]) );
  FA_8037 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n968), .CI(C[455]), .CO(C[456]) );
  FA_8036 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n969), .CI(C[456]), .CO(C[457]) );
  FA_8035 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n970), .CI(C[457]), .CO(C[458]) );
  FA_8034 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n971), .CI(C[458]), .CO(C[459]) );
  FA_8033 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n972), .CI(C[459]), .CO(C[460]) );
  FA_8032 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n973), .CI(C[460]), .CO(C[461]) );
  FA_8031 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n974), .CI(C[461]), .CO(C[462]) );
  FA_8030 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n975), .CI(C[462]), .CO(C[463]) );
  FA_8029 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n976), .CI(C[463]), .CO(C[464]) );
  FA_8028 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n977), .CI(C[464]), .CO(C[465]) );
  FA_8027 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n978), .CI(C[465]), .CO(C[466]) );
  FA_8026 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n979), .CI(C[466]), .CO(C[467]) );
  FA_8025 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n980), .CI(C[467]), .CO(C[468]) );
  FA_8024 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n981), .CI(C[468]), .CO(C[469]) );
  FA_8023 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n982), .CI(C[469]), .CO(C[470]) );
  FA_8022 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n983), .CI(C[470]), .CO(C[471]) );
  FA_8021 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n984), .CI(C[471]), .CO(C[472]) );
  FA_8020 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n985), .CI(C[472]), .CO(C[473]) );
  FA_8019 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n986), .CI(C[473]), .CO(C[474]) );
  FA_8018 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n987), .CI(C[474]), .CO(C[475]) );
  FA_8017 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n988), .CI(C[475]), .CO(C[476]) );
  FA_8016 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n989), .CI(C[476]), .CO(C[477]) );
  FA_8015 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n990), .CI(C[477]), .CO(C[478]) );
  FA_8014 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n991), .CI(C[478]), .CO(C[479]) );
  FA_8013 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n992), .CI(C[479]), .CO(C[480]) );
  FA_8012 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n993), .CI(C[480]), .CO(C[481]) );
  FA_8011 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n994), .CI(C[481]), .CO(C[482]) );
  FA_8010 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n995), .CI(C[482]), .CO(C[483]) );
  FA_8009 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n996), .CI(C[483]), .CO(C[484]) );
  FA_8008 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n997), .CI(C[484]), .CO(C[485]) );
  FA_8007 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n998), .CI(C[485]), .CO(C[486]) );
  FA_8006 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n999), .CI(C[486]), .CO(C[487]) );
  FA_8005 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1000), .CI(
        C[487]), .CO(C[488]) );
  FA_8004 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1001), .CI(
        C[488]), .CO(C[489]) );
  FA_8003 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1002), .CI(
        C[489]), .CO(C[490]) );
  FA_8002 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1003), .CI(
        C[490]), .CO(C[491]) );
  FA_8001 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1004), .CI(
        C[491]), .CO(C[492]) );
  FA_8000 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1005), .CI(
        C[492]), .CO(C[493]) );
  FA_7999 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1006), .CI(
        C[493]), .CO(C[494]) );
  FA_7998 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1007), .CI(
        C[494]), .CO(C[495]) );
  FA_7997 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1008), .CI(
        C[495]), .CO(C[496]) );
  FA_7996 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1009), .CI(
        C[496]), .CO(C[497]) );
  FA_7995 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1010), .CI(
        C[497]), .CO(C[498]) );
  FA_7994 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1011), .CI(
        C[498]), .CO(C[499]) );
  FA_7993 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1012), .CI(
        C[499]), .CO(C[500]) );
  FA_7992 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1013), .CI(
        C[500]), .CO(C[501]) );
  FA_7991 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1014), .CI(
        C[501]), .CO(C[502]) );
  FA_7990 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1015), .CI(
        C[502]), .CO(C[503]) );
  FA_7989 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1016), .CI(
        C[503]), .CO(C[504]) );
  FA_7988 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1017), .CI(
        C[504]), .CO(C[505]) );
  FA_7987 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1018), .CI(
        C[505]), .CO(C[506]) );
  FA_7986 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1019), .CI(
        C[506]), .CO(C[507]) );
  FA_7985 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1020), .CI(
        C[507]), .CO(C[508]) );
  FA_7984 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1021), .CI(
        C[508]), .CO(C[509]) );
  FA_7983 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1022), .CI(
        C[509]), .CO(C[510]) );
  FA_7982 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1023), .CI(
        C[510]), .CO(C[511]) );
  FA_7981 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1024), .CI(
        C[511]), .CO(C[512]) );
  FA_7980 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .CO(C[513]) );
  FA_7979 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b1), .CI(C[513]), .CO(O) );
  IV U2 ( .A(B[415]), .Z(n928) );
  IV U3 ( .A(B[416]), .Z(n929) );
  IV U4 ( .A(B[417]), .Z(n930) );
  IV U5 ( .A(B[418]), .Z(n931) );
  IV U6 ( .A(B[419]), .Z(n932) );
  IV U7 ( .A(B[420]), .Z(n933) );
  IV U8 ( .A(B[421]), .Z(n934) );
  IV U9 ( .A(B[422]), .Z(n935) );
  IV U10 ( .A(B[423]), .Z(n936) );
  IV U11 ( .A(B[424]), .Z(n937) );
  IV U12 ( .A(B[505]), .Z(n1018) );
  IV U13 ( .A(B[425]), .Z(n938) );
  IV U14 ( .A(B[426]), .Z(n939) );
  IV U15 ( .A(B[427]), .Z(n940) );
  IV U16 ( .A(B[428]), .Z(n941) );
  IV U17 ( .A(B[429]), .Z(n942) );
  IV U18 ( .A(B[430]), .Z(n943) );
  IV U19 ( .A(B[431]), .Z(n944) );
  IV U20 ( .A(B[432]), .Z(n945) );
  IV U21 ( .A(B[433]), .Z(n946) );
  IV U22 ( .A(B[434]), .Z(n947) );
  IV U23 ( .A(B[506]), .Z(n1019) );
  IV U24 ( .A(B[435]), .Z(n948) );
  IV U25 ( .A(B[436]), .Z(n949) );
  IV U26 ( .A(B[437]), .Z(n950) );
  IV U27 ( .A(B[438]), .Z(n951) );
  IV U28 ( .A(B[439]), .Z(n952) );
  IV U29 ( .A(B[440]), .Z(n953) );
  IV U30 ( .A(B[441]), .Z(n954) );
  IV U31 ( .A(B[442]), .Z(n955) );
  IV U32 ( .A(B[443]), .Z(n956) );
  IV U33 ( .A(B[444]), .Z(n957) );
  IV U34 ( .A(B[507]), .Z(n1020) );
  IV U35 ( .A(B[445]), .Z(n958) );
  IV U36 ( .A(B[446]), .Z(n959) );
  IV U37 ( .A(B[447]), .Z(n960) );
  IV U38 ( .A(B[448]), .Z(n961) );
  IV U39 ( .A(B[449]), .Z(n962) );
  IV U40 ( .A(B[450]), .Z(n963) );
  IV U41 ( .A(B[451]), .Z(n964) );
  IV U42 ( .A(B[452]), .Z(n965) );
  IV U43 ( .A(B[453]), .Z(n966) );
  IV U44 ( .A(B[454]), .Z(n967) );
  IV U45 ( .A(B[508]), .Z(n1021) );
  IV U46 ( .A(B[455]), .Z(n968) );
  IV U47 ( .A(B[456]), .Z(n969) );
  IV U48 ( .A(B[457]), .Z(n970) );
  IV U49 ( .A(B[458]), .Z(n971) );
  IV U50 ( .A(B[459]), .Z(n972) );
  IV U51 ( .A(B[460]), .Z(n973) );
  IV U52 ( .A(B[461]), .Z(n974) );
  IV U53 ( .A(B[462]), .Z(n975) );
  IV U54 ( .A(B[0]), .Z(n2) );
  IV U55 ( .A(B[1]), .Z(n514) );
  IV U56 ( .A(B[2]), .Z(n515) );
  IV U57 ( .A(B[3]), .Z(n516) );
  IV U58 ( .A(B[4]), .Z(n517) );
  IV U59 ( .A(B[463]), .Z(n976) );
  IV U60 ( .A(B[5]), .Z(n518) );
  IV U61 ( .A(B[6]), .Z(n519) );
  IV U62 ( .A(B[7]), .Z(n520) );
  IV U63 ( .A(B[8]), .Z(n521) );
  IV U64 ( .A(B[9]), .Z(n522) );
  IV U65 ( .A(B[10]), .Z(n523) );
  IV U66 ( .A(B[11]), .Z(n524) );
  IV U67 ( .A(B[12]), .Z(n525) );
  IV U68 ( .A(B[13]), .Z(n526) );
  IV U69 ( .A(B[14]), .Z(n527) );
  IV U70 ( .A(B[464]), .Z(n977) );
  IV U71 ( .A(B[509]), .Z(n1022) );
  IV U72 ( .A(B[15]), .Z(n528) );
  IV U73 ( .A(B[16]), .Z(n529) );
  IV U74 ( .A(B[17]), .Z(n530) );
  IV U75 ( .A(B[18]), .Z(n531) );
  IV U76 ( .A(B[19]), .Z(n532) );
  IV U77 ( .A(B[20]), .Z(n533) );
  IV U78 ( .A(B[21]), .Z(n534) );
  IV U79 ( .A(B[22]), .Z(n535) );
  IV U80 ( .A(B[23]), .Z(n536) );
  IV U81 ( .A(B[24]), .Z(n537) );
  IV U82 ( .A(B[465]), .Z(n978) );
  IV U83 ( .A(B[25]), .Z(n538) );
  IV U84 ( .A(B[26]), .Z(n539) );
  IV U85 ( .A(B[27]), .Z(n540) );
  IV U86 ( .A(B[28]), .Z(n541) );
  IV U87 ( .A(B[29]), .Z(n542) );
  IV U88 ( .A(B[30]), .Z(n543) );
  IV U89 ( .A(B[31]), .Z(n544) );
  IV U90 ( .A(B[32]), .Z(n545) );
  IV U91 ( .A(B[33]), .Z(n546) );
  IV U92 ( .A(B[34]), .Z(n547) );
  IV U93 ( .A(B[466]), .Z(n979) );
  IV U94 ( .A(B[35]), .Z(n548) );
  IV U95 ( .A(B[36]), .Z(n549) );
  IV U96 ( .A(B[37]), .Z(n550) );
  IV U97 ( .A(B[38]), .Z(n551) );
  IV U98 ( .A(B[39]), .Z(n552) );
  IV U99 ( .A(B[40]), .Z(n553) );
  IV U100 ( .A(B[41]), .Z(n554) );
  IV U101 ( .A(B[42]), .Z(n555) );
  IV U102 ( .A(B[43]), .Z(n556) );
  IV U103 ( .A(B[44]), .Z(n557) );
  IV U104 ( .A(B[467]), .Z(n980) );
  IV U105 ( .A(B[45]), .Z(n558) );
  IV U106 ( .A(B[46]), .Z(n559) );
  IV U107 ( .A(B[47]), .Z(n560) );
  IV U108 ( .A(B[48]), .Z(n561) );
  IV U109 ( .A(B[49]), .Z(n562) );
  IV U110 ( .A(B[50]), .Z(n563) );
  IV U111 ( .A(B[51]), .Z(n564) );
  IV U112 ( .A(B[52]), .Z(n565) );
  IV U113 ( .A(B[53]), .Z(n566) );
  IV U114 ( .A(B[54]), .Z(n567) );
  IV U115 ( .A(B[468]), .Z(n981) );
  IV U116 ( .A(B[55]), .Z(n568) );
  IV U117 ( .A(B[56]), .Z(n569) );
  IV U118 ( .A(B[57]), .Z(n570) );
  IV U119 ( .A(B[58]), .Z(n571) );
  IV U120 ( .A(B[59]), .Z(n572) );
  IV U121 ( .A(B[60]), .Z(n573) );
  IV U122 ( .A(B[61]), .Z(n574) );
  IV U123 ( .A(B[62]), .Z(n575) );
  IV U124 ( .A(B[63]), .Z(n576) );
  IV U125 ( .A(B[64]), .Z(n577) );
  IV U126 ( .A(B[469]), .Z(n982) );
  IV U127 ( .A(B[65]), .Z(n578) );
  IV U128 ( .A(B[66]), .Z(n579) );
  IV U129 ( .A(B[67]), .Z(n580) );
  IV U130 ( .A(B[68]), .Z(n581) );
  IV U131 ( .A(B[69]), .Z(n582) );
  IV U132 ( .A(B[70]), .Z(n583) );
  IV U133 ( .A(B[71]), .Z(n584) );
  IV U134 ( .A(B[72]), .Z(n585) );
  IV U135 ( .A(B[73]), .Z(n586) );
  IV U136 ( .A(B[74]), .Z(n587) );
  IV U137 ( .A(B[470]), .Z(n983) );
  IV U138 ( .A(B[75]), .Z(n588) );
  IV U139 ( .A(B[76]), .Z(n589) );
  IV U140 ( .A(B[77]), .Z(n590) );
  IV U141 ( .A(B[78]), .Z(n591) );
  IV U142 ( .A(B[79]), .Z(n592) );
  IV U143 ( .A(B[80]), .Z(n593) );
  IV U144 ( .A(B[81]), .Z(n594) );
  IV U145 ( .A(B[82]), .Z(n595) );
  IV U146 ( .A(B[83]), .Z(n596) );
  IV U147 ( .A(B[84]), .Z(n597) );
  IV U148 ( .A(B[471]), .Z(n984) );
  IV U149 ( .A(B[85]), .Z(n598) );
  IV U150 ( .A(B[86]), .Z(n599) );
  IV U151 ( .A(B[87]), .Z(n600) );
  IV U152 ( .A(B[88]), .Z(n601) );
  IV U153 ( .A(B[89]), .Z(n602) );
  IV U154 ( .A(B[90]), .Z(n603) );
  IV U155 ( .A(B[91]), .Z(n604) );
  IV U156 ( .A(B[92]), .Z(n605) );
  IV U157 ( .A(B[93]), .Z(n606) );
  IV U158 ( .A(B[94]), .Z(n607) );
  IV U159 ( .A(B[472]), .Z(n985) );
  IV U160 ( .A(B[95]), .Z(n608) );
  IV U161 ( .A(B[96]), .Z(n609) );
  IV U162 ( .A(B[97]), .Z(n610) );
  IV U163 ( .A(B[98]), .Z(n611) );
  IV U164 ( .A(B[99]), .Z(n612) );
  IV U165 ( .A(B[100]), .Z(n613) );
  IV U166 ( .A(B[101]), .Z(n614) );
  IV U167 ( .A(B[102]), .Z(n615) );
  IV U168 ( .A(B[103]), .Z(n616) );
  IV U169 ( .A(B[104]), .Z(n617) );
  IV U170 ( .A(B[473]), .Z(n986) );
  IV U171 ( .A(B[105]), .Z(n618) );
  IV U172 ( .A(B[106]), .Z(n619) );
  IV U173 ( .A(B[107]), .Z(n620) );
  IV U174 ( .A(B[108]), .Z(n621) );
  IV U175 ( .A(B[109]), .Z(n622) );
  IV U176 ( .A(B[110]), .Z(n623) );
  IV U177 ( .A(B[111]), .Z(n624) );
  IV U178 ( .A(B[112]), .Z(n625) );
  IV U179 ( .A(B[113]), .Z(n626) );
  IV U180 ( .A(B[114]), .Z(n627) );
  IV U181 ( .A(B[474]), .Z(n987) );
  IV U182 ( .A(B[510]), .Z(n1023) );
  IV U183 ( .A(B[115]), .Z(n628) );
  IV U184 ( .A(B[116]), .Z(n629) );
  IV U185 ( .A(B[117]), .Z(n630) );
  IV U186 ( .A(B[118]), .Z(n631) );
  IV U187 ( .A(B[119]), .Z(n632) );
  IV U188 ( .A(B[120]), .Z(n633) );
  IV U189 ( .A(B[121]), .Z(n634) );
  IV U190 ( .A(B[122]), .Z(n635) );
  IV U191 ( .A(B[123]), .Z(n636) );
  IV U192 ( .A(B[124]), .Z(n637) );
  IV U193 ( .A(B[475]), .Z(n988) );
  IV U194 ( .A(B[125]), .Z(n638) );
  IV U195 ( .A(B[126]), .Z(n639) );
  IV U196 ( .A(B[127]), .Z(n640) );
  IV U197 ( .A(B[128]), .Z(n641) );
  IV U198 ( .A(B[129]), .Z(n642) );
  IV U199 ( .A(B[130]), .Z(n643) );
  IV U200 ( .A(B[131]), .Z(n644) );
  IV U201 ( .A(B[132]), .Z(n645) );
  IV U202 ( .A(B[133]), .Z(n646) );
  IV U203 ( .A(B[134]), .Z(n647) );
  IV U204 ( .A(B[476]), .Z(n989) );
  IV U205 ( .A(B[135]), .Z(n648) );
  IV U206 ( .A(B[136]), .Z(n649) );
  IV U207 ( .A(B[137]), .Z(n650) );
  IV U208 ( .A(B[138]), .Z(n651) );
  IV U209 ( .A(B[139]), .Z(n652) );
  IV U210 ( .A(B[140]), .Z(n653) );
  IV U211 ( .A(B[141]), .Z(n654) );
  IV U212 ( .A(B[142]), .Z(n655) );
  IV U213 ( .A(B[143]), .Z(n656) );
  IV U214 ( .A(B[144]), .Z(n657) );
  IV U215 ( .A(B[477]), .Z(n990) );
  IV U216 ( .A(B[145]), .Z(n658) );
  IV U217 ( .A(B[146]), .Z(n659) );
  IV U218 ( .A(B[147]), .Z(n660) );
  IV U219 ( .A(B[148]), .Z(n661) );
  IV U220 ( .A(B[149]), .Z(n662) );
  IV U221 ( .A(B[150]), .Z(n663) );
  IV U222 ( .A(B[151]), .Z(n664) );
  IV U223 ( .A(B[152]), .Z(n665) );
  IV U224 ( .A(B[153]), .Z(n666) );
  IV U225 ( .A(B[154]), .Z(n667) );
  IV U226 ( .A(B[478]), .Z(n991) );
  IV U227 ( .A(B[155]), .Z(n668) );
  IV U228 ( .A(B[156]), .Z(n669) );
  IV U229 ( .A(B[157]), .Z(n670) );
  IV U230 ( .A(B[158]), .Z(n671) );
  IV U231 ( .A(B[159]), .Z(n672) );
  IV U232 ( .A(B[160]), .Z(n673) );
  IV U233 ( .A(B[161]), .Z(n674) );
  IV U234 ( .A(B[162]), .Z(n675) );
  IV U235 ( .A(B[163]), .Z(n676) );
  IV U236 ( .A(B[164]), .Z(n677) );
  IV U237 ( .A(B[479]), .Z(n992) );
  IV U238 ( .A(B[165]), .Z(n678) );
  IV U239 ( .A(B[166]), .Z(n679) );
  IV U240 ( .A(B[167]), .Z(n680) );
  IV U241 ( .A(B[168]), .Z(n681) );
  IV U242 ( .A(B[169]), .Z(n682) );
  IV U243 ( .A(B[170]), .Z(n683) );
  IV U244 ( .A(B[171]), .Z(n684) );
  IV U245 ( .A(B[172]), .Z(n685) );
  IV U246 ( .A(B[173]), .Z(n686) );
  IV U247 ( .A(B[174]), .Z(n687) );
  IV U248 ( .A(B[480]), .Z(n993) );
  IV U249 ( .A(B[175]), .Z(n688) );
  IV U250 ( .A(B[176]), .Z(n689) );
  IV U251 ( .A(B[177]), .Z(n690) );
  IV U252 ( .A(B[178]), .Z(n691) );
  IV U253 ( .A(B[179]), .Z(n692) );
  IV U254 ( .A(B[180]), .Z(n693) );
  IV U255 ( .A(B[181]), .Z(n694) );
  IV U256 ( .A(B[182]), .Z(n695) );
  IV U257 ( .A(B[183]), .Z(n696) );
  IV U258 ( .A(B[184]), .Z(n697) );
  IV U259 ( .A(B[481]), .Z(n994) );
  IV U260 ( .A(B[185]), .Z(n698) );
  IV U261 ( .A(B[186]), .Z(n699) );
  IV U262 ( .A(B[187]), .Z(n700) );
  IV U263 ( .A(B[188]), .Z(n701) );
  IV U264 ( .A(B[189]), .Z(n702) );
  IV U265 ( .A(B[190]), .Z(n703) );
  IV U266 ( .A(B[191]), .Z(n704) );
  IV U267 ( .A(B[192]), .Z(n705) );
  IV U268 ( .A(B[193]), .Z(n706) );
  IV U269 ( .A(B[194]), .Z(n707) );
  IV U270 ( .A(B[482]), .Z(n995) );
  IV U271 ( .A(B[195]), .Z(n708) );
  IV U272 ( .A(B[196]), .Z(n709) );
  IV U273 ( .A(B[197]), .Z(n710) );
  IV U274 ( .A(B[198]), .Z(n711) );
  IV U275 ( .A(B[199]), .Z(n712) );
  IV U276 ( .A(B[200]), .Z(n713) );
  IV U277 ( .A(B[201]), .Z(n714) );
  IV U278 ( .A(B[202]), .Z(n715) );
  IV U279 ( .A(B[203]), .Z(n716) );
  IV U280 ( .A(B[204]), .Z(n717) );
  IV U281 ( .A(B[483]), .Z(n996) );
  IV U282 ( .A(B[205]), .Z(n718) );
  IV U283 ( .A(B[206]), .Z(n719) );
  IV U284 ( .A(B[207]), .Z(n720) );
  IV U285 ( .A(B[208]), .Z(n721) );
  IV U286 ( .A(B[209]), .Z(n722) );
  IV U287 ( .A(B[210]), .Z(n723) );
  IV U288 ( .A(B[211]), .Z(n724) );
  IV U289 ( .A(B[212]), .Z(n725) );
  IV U290 ( .A(B[213]), .Z(n726) );
  IV U291 ( .A(B[214]), .Z(n727) );
  IV U292 ( .A(B[484]), .Z(n997) );
  IV U293 ( .A(B[511]), .Z(n1024) );
  IV U294 ( .A(B[215]), .Z(n728) );
  IV U295 ( .A(B[216]), .Z(n729) );
  IV U296 ( .A(B[217]), .Z(n730) );
  IV U297 ( .A(B[218]), .Z(n731) );
  IV U298 ( .A(B[219]), .Z(n732) );
  IV U299 ( .A(B[220]), .Z(n733) );
  IV U300 ( .A(B[221]), .Z(n734) );
  IV U301 ( .A(B[222]), .Z(n735) );
  IV U302 ( .A(B[223]), .Z(n736) );
  IV U303 ( .A(B[224]), .Z(n737) );
  IV U304 ( .A(B[485]), .Z(n998) );
  IV U305 ( .A(B[225]), .Z(n738) );
  IV U306 ( .A(B[226]), .Z(n739) );
  IV U307 ( .A(B[227]), .Z(n740) );
  IV U308 ( .A(B[228]), .Z(n741) );
  IV U309 ( .A(B[229]), .Z(n742) );
  IV U310 ( .A(B[230]), .Z(n743) );
  IV U311 ( .A(B[231]), .Z(n744) );
  IV U312 ( .A(B[232]), .Z(n745) );
  IV U313 ( .A(B[233]), .Z(n746) );
  IV U314 ( .A(B[234]), .Z(n747) );
  IV U315 ( .A(B[486]), .Z(n999) );
  IV U316 ( .A(B[235]), .Z(n748) );
  IV U317 ( .A(B[236]), .Z(n749) );
  IV U318 ( .A(B[237]), .Z(n750) );
  IV U319 ( .A(B[238]), .Z(n751) );
  IV U320 ( .A(B[239]), .Z(n752) );
  IV U321 ( .A(B[240]), .Z(n753) );
  IV U322 ( .A(B[241]), .Z(n754) );
  IV U323 ( .A(B[242]), .Z(n755) );
  IV U324 ( .A(B[243]), .Z(n756) );
  IV U325 ( .A(B[244]), .Z(n757) );
  IV U326 ( .A(B[487]), .Z(n1000) );
  IV U327 ( .A(B[245]), .Z(n758) );
  IV U328 ( .A(B[246]), .Z(n759) );
  IV U329 ( .A(B[247]), .Z(n760) );
  IV U330 ( .A(B[248]), .Z(n761) );
  IV U331 ( .A(B[249]), .Z(n762) );
  IV U332 ( .A(B[250]), .Z(n763) );
  IV U333 ( .A(B[251]), .Z(n764) );
  IV U334 ( .A(B[252]), .Z(n765) );
  IV U335 ( .A(B[253]), .Z(n766) );
  IV U336 ( .A(B[254]), .Z(n767) );
  IV U337 ( .A(B[488]), .Z(n1001) );
  IV U338 ( .A(B[255]), .Z(n768) );
  IV U339 ( .A(B[256]), .Z(n769) );
  IV U340 ( .A(B[257]), .Z(n770) );
  IV U341 ( .A(B[258]), .Z(n771) );
  IV U342 ( .A(B[259]), .Z(n772) );
  IV U343 ( .A(B[260]), .Z(n773) );
  IV U344 ( .A(B[261]), .Z(n774) );
  IV U345 ( .A(B[262]), .Z(n775) );
  IV U346 ( .A(B[263]), .Z(n776) );
  IV U347 ( .A(B[264]), .Z(n777) );
  IV U348 ( .A(B[489]), .Z(n1002) );
  IV U349 ( .A(B[265]), .Z(n778) );
  IV U350 ( .A(B[266]), .Z(n779) );
  IV U351 ( .A(B[267]), .Z(n780) );
  IV U352 ( .A(B[268]), .Z(n781) );
  IV U353 ( .A(B[269]), .Z(n782) );
  IV U354 ( .A(B[270]), .Z(n783) );
  IV U355 ( .A(B[271]), .Z(n784) );
  IV U356 ( .A(B[272]), .Z(n785) );
  IV U357 ( .A(B[273]), .Z(n786) );
  IV U358 ( .A(B[274]), .Z(n787) );
  IV U359 ( .A(B[490]), .Z(n1003) );
  IV U360 ( .A(B[275]), .Z(n788) );
  IV U361 ( .A(B[276]), .Z(n789) );
  IV U362 ( .A(B[277]), .Z(n790) );
  IV U363 ( .A(B[278]), .Z(n791) );
  IV U364 ( .A(B[279]), .Z(n792) );
  IV U365 ( .A(B[280]), .Z(n793) );
  IV U366 ( .A(B[281]), .Z(n794) );
  IV U367 ( .A(B[282]), .Z(n795) );
  IV U368 ( .A(B[283]), .Z(n796) );
  IV U369 ( .A(B[284]), .Z(n797) );
  IV U370 ( .A(B[491]), .Z(n1004) );
  IV U371 ( .A(B[285]), .Z(n798) );
  IV U372 ( .A(B[286]), .Z(n799) );
  IV U373 ( .A(B[287]), .Z(n800) );
  IV U374 ( .A(B[288]), .Z(n801) );
  IV U375 ( .A(B[289]), .Z(n802) );
  IV U376 ( .A(B[290]), .Z(n803) );
  IV U377 ( .A(B[291]), .Z(n804) );
  IV U378 ( .A(B[292]), .Z(n805) );
  IV U379 ( .A(B[293]), .Z(n806) );
  IV U380 ( .A(B[294]), .Z(n807) );
  IV U381 ( .A(B[492]), .Z(n1005) );
  IV U382 ( .A(B[295]), .Z(n808) );
  IV U383 ( .A(B[296]), .Z(n809) );
  IV U384 ( .A(B[297]), .Z(n810) );
  IV U385 ( .A(B[298]), .Z(n811) );
  IV U386 ( .A(B[299]), .Z(n812) );
  IV U387 ( .A(B[300]), .Z(n813) );
  IV U388 ( .A(B[301]), .Z(n814) );
  IV U389 ( .A(B[302]), .Z(n815) );
  IV U390 ( .A(B[303]), .Z(n816) );
  IV U391 ( .A(B[304]), .Z(n817) );
  IV U392 ( .A(B[493]), .Z(n1006) );
  IV U393 ( .A(B[305]), .Z(n818) );
  IV U394 ( .A(B[306]), .Z(n819) );
  IV U395 ( .A(B[307]), .Z(n820) );
  IV U396 ( .A(B[308]), .Z(n821) );
  IV U397 ( .A(B[309]), .Z(n822) );
  IV U398 ( .A(B[310]), .Z(n823) );
  IV U399 ( .A(B[311]), .Z(n824) );
  IV U400 ( .A(B[312]), .Z(n825) );
  IV U401 ( .A(B[313]), .Z(n826) );
  IV U402 ( .A(B[314]), .Z(n827) );
  IV U403 ( .A(B[494]), .Z(n1007) );
  IV U404 ( .A(B[315]), .Z(n828) );
  IV U405 ( .A(B[316]), .Z(n829) );
  IV U406 ( .A(B[317]), .Z(n830) );
  IV U407 ( .A(B[318]), .Z(n831) );
  IV U408 ( .A(B[319]), .Z(n832) );
  IV U409 ( .A(B[320]), .Z(n833) );
  IV U410 ( .A(B[321]), .Z(n834) );
  IV U411 ( .A(B[322]), .Z(n835) );
  IV U412 ( .A(B[323]), .Z(n836) );
  IV U413 ( .A(B[324]), .Z(n837) );
  IV U414 ( .A(B[495]), .Z(n1008) );
  IV U415 ( .A(B[325]), .Z(n838) );
  IV U416 ( .A(B[326]), .Z(n839) );
  IV U417 ( .A(B[327]), .Z(n840) );
  IV U418 ( .A(B[328]), .Z(n841) );
  IV U419 ( .A(B[329]), .Z(n842) );
  IV U420 ( .A(B[330]), .Z(n843) );
  IV U421 ( .A(B[331]), .Z(n844) );
  IV U422 ( .A(B[332]), .Z(n845) );
  IV U423 ( .A(B[333]), .Z(n846) );
  IV U424 ( .A(B[334]), .Z(n847) );
  IV U425 ( .A(B[496]), .Z(n1009) );
  IV U426 ( .A(B[335]), .Z(n848) );
  IV U427 ( .A(B[336]), .Z(n849) );
  IV U428 ( .A(B[337]), .Z(n850) );
  IV U429 ( .A(B[338]), .Z(n851) );
  IV U430 ( .A(B[339]), .Z(n852) );
  IV U431 ( .A(B[340]), .Z(n853) );
  IV U432 ( .A(B[341]), .Z(n854) );
  IV U433 ( .A(B[342]), .Z(n855) );
  IV U434 ( .A(B[343]), .Z(n856) );
  IV U435 ( .A(B[344]), .Z(n857) );
  IV U436 ( .A(B[497]), .Z(n1010) );
  IV U437 ( .A(B[345]), .Z(n858) );
  IV U438 ( .A(B[346]), .Z(n859) );
  IV U439 ( .A(B[347]), .Z(n860) );
  IV U440 ( .A(B[348]), .Z(n861) );
  IV U441 ( .A(B[349]), .Z(n862) );
  IV U442 ( .A(B[350]), .Z(n863) );
  IV U443 ( .A(B[351]), .Z(n864) );
  IV U444 ( .A(B[352]), .Z(n865) );
  IV U445 ( .A(B[353]), .Z(n866) );
  IV U446 ( .A(B[354]), .Z(n867) );
  IV U447 ( .A(B[498]), .Z(n1011) );
  IV U448 ( .A(B[355]), .Z(n868) );
  IV U449 ( .A(B[356]), .Z(n869) );
  IV U450 ( .A(B[357]), .Z(n870) );
  IV U451 ( .A(B[358]), .Z(n871) );
  IV U452 ( .A(B[359]), .Z(n872) );
  IV U453 ( .A(B[360]), .Z(n873) );
  IV U454 ( .A(B[361]), .Z(n874) );
  IV U455 ( .A(B[362]), .Z(n875) );
  IV U456 ( .A(B[363]), .Z(n876) );
  IV U457 ( .A(B[364]), .Z(n877) );
  IV U458 ( .A(B[499]), .Z(n1012) );
  IV U459 ( .A(B[365]), .Z(n878) );
  IV U460 ( .A(B[366]), .Z(n879) );
  IV U461 ( .A(B[367]), .Z(n880) );
  IV U462 ( .A(B[368]), .Z(n881) );
  IV U463 ( .A(B[369]), .Z(n882) );
  IV U464 ( .A(B[370]), .Z(n883) );
  IV U465 ( .A(B[371]), .Z(n884) );
  IV U466 ( .A(B[372]), .Z(n885) );
  IV U467 ( .A(B[373]), .Z(n886) );
  IV U468 ( .A(B[374]), .Z(n887) );
  IV U469 ( .A(B[500]), .Z(n1013) );
  IV U470 ( .A(B[375]), .Z(n888) );
  IV U471 ( .A(B[376]), .Z(n889) );
  IV U472 ( .A(B[377]), .Z(n890) );
  IV U473 ( .A(B[378]), .Z(n891) );
  IV U474 ( .A(B[379]), .Z(n892) );
  IV U475 ( .A(B[380]), .Z(n893) );
  IV U476 ( .A(B[381]), .Z(n894) );
  IV U477 ( .A(B[382]), .Z(n895) );
  IV U478 ( .A(B[383]), .Z(n896) );
  IV U479 ( .A(B[384]), .Z(n897) );
  IV U480 ( .A(B[501]), .Z(n1014) );
  IV U481 ( .A(B[385]), .Z(n898) );
  IV U482 ( .A(B[386]), .Z(n899) );
  IV U483 ( .A(B[387]), .Z(n900) );
  IV U484 ( .A(B[388]), .Z(n901) );
  IV U485 ( .A(B[389]), .Z(n902) );
  IV U486 ( .A(B[390]), .Z(n903) );
  IV U487 ( .A(B[391]), .Z(n904) );
  IV U488 ( .A(B[392]), .Z(n905) );
  IV U489 ( .A(B[393]), .Z(n906) );
  IV U490 ( .A(B[394]), .Z(n907) );
  IV U491 ( .A(B[502]), .Z(n1015) );
  IV U492 ( .A(B[395]), .Z(n908) );
  IV U493 ( .A(B[396]), .Z(n909) );
  IV U494 ( .A(B[397]), .Z(n910) );
  IV U495 ( .A(B[398]), .Z(n911) );
  IV U496 ( .A(B[399]), .Z(n912) );
  IV U497 ( .A(B[400]), .Z(n913) );
  IV U498 ( .A(B[401]), .Z(n914) );
  IV U499 ( .A(B[402]), .Z(n915) );
  IV U500 ( .A(B[403]), .Z(n916) );
  IV U501 ( .A(B[404]), .Z(n917) );
  IV U502 ( .A(B[503]), .Z(n1016) );
  IV U503 ( .A(B[405]), .Z(n918) );
  IV U504 ( .A(B[406]), .Z(n919) );
  IV U505 ( .A(B[407]), .Z(n920) );
  IV U506 ( .A(B[408]), .Z(n921) );
  IV U507 ( .A(B[409]), .Z(n922) );
  IV U508 ( .A(B[410]), .Z(n923) );
  IV U509 ( .A(B[411]), .Z(n924) );
  IV U510 ( .A(B[412]), .Z(n925) );
  IV U511 ( .A(B[413]), .Z(n926) );
  IV U512 ( .A(B[414]), .Z(n927) );
  IV U513 ( .A(B[504]), .Z(n1017) );
endmodule


module FA_6438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_6439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_6950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N514_3 ( A, B, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  output CO;
  wire   n2, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  wire   [513:1] C;

  FA_6950 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(
        S[0]), .CO(C[1]) );
  FA_6949 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n514), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_6948 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n515), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_6947 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n516), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_6946 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n517), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_6945 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n518), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_6944 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n519), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_6943 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n520), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_6942 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n521), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_6941 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n522), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_6940 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n523), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_6939 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n524), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_6938 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n525), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_6937 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n526), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_6936 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n527), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_6935 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n528), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_6934 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n529), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_6933 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n530), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_6932 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n531), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_6931 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n532), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_6930 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n533), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_6929 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n534), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_6928 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n535), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_6927 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n536), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_6926 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n537), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_6925 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n538), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_6924 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n539), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_6923 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n540), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_6922 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n541), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_6921 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n542), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_6920 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n543), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_6919 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n544), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_6918 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n545), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_6917 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n546), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_6916 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n547), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_6915 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n548), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_6914 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n549), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_6913 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n550), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_6912 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n551), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_6911 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n552), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_6910 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n553), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_6909 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n554), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_6908 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n555), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_6907 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n556), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_6906 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n557), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_6905 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n558), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_6904 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n559), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_6903 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n560), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_6902 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n561), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_6901 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n562), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_6900 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n563), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_6899 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n564), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_6898 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n565), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_6897 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n566), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_6896 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n567), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_6895 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n568), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_6894 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n569), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_6893 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n570), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_6892 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n571), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_6891 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n572), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_6890 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n573), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_6889 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n574), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_6888 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n575), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_6887 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n576), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_6886 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n577), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_6885 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n578), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_6884 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n579), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_6883 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n580), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_6882 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n581), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_6881 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n582), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_6880 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n583), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_6879 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n584), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_6878 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n585), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_6877 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n586), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_6876 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n587), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_6875 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n588), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_6874 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n589), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_6873 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n590), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_6872 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n591), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_6871 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n592), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_6870 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n593), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_6869 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n594), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_6868 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n595), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_6867 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n596), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_6866 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n597), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_6865 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n598), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_6864 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n599), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_6863 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n600), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_6862 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n601), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_6861 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n602), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_6860 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n603), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_6859 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n604), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_6858 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n605), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_6857 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n606), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_6856 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n607), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_6855 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n608), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_6854 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n609), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_6853 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n610), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_6852 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n611), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_6851 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n612), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_6850 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n613), .CI(C[100]), .S(S[100]), .CO(C[101]) );
  FA_6849 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n614), .CI(C[101]), .S(S[101]), .CO(C[102]) );
  FA_6848 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n615), .CI(C[102]), .S(S[102]), .CO(C[103]) );
  FA_6847 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n616), .CI(C[103]), .S(S[103]), .CO(C[104]) );
  FA_6846 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n617), .CI(C[104]), .S(S[104]), .CO(C[105]) );
  FA_6845 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n618), .CI(C[105]), .S(S[105]), .CO(C[106]) );
  FA_6844 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n619), .CI(C[106]), .S(S[106]), .CO(C[107]) );
  FA_6843 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n620), .CI(C[107]), .S(S[107]), .CO(C[108]) );
  FA_6842 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n621), .CI(C[108]), .S(S[108]), .CO(C[109]) );
  FA_6841 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n622), .CI(C[109]), .S(S[109]), .CO(C[110]) );
  FA_6840 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n623), .CI(C[110]), .S(S[110]), .CO(C[111]) );
  FA_6839 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n624), .CI(C[111]), .S(S[111]), .CO(C[112]) );
  FA_6838 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n625), .CI(C[112]), .S(S[112]), .CO(C[113]) );
  FA_6837 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n626), .CI(C[113]), .S(S[113]), .CO(C[114]) );
  FA_6836 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n627), .CI(C[114]), .S(S[114]), .CO(C[115]) );
  FA_6835 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n628), .CI(C[115]), .S(S[115]), .CO(C[116]) );
  FA_6834 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n629), .CI(C[116]), .S(S[116]), .CO(C[117]) );
  FA_6833 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n630), .CI(C[117]), .S(S[117]), .CO(C[118]) );
  FA_6832 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n631), .CI(C[118]), .S(S[118]), .CO(C[119]) );
  FA_6831 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n632), .CI(C[119]), .S(S[119]), .CO(C[120]) );
  FA_6830 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n633), .CI(C[120]), .S(S[120]), .CO(C[121]) );
  FA_6829 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n634), .CI(C[121]), .S(S[121]), .CO(C[122]) );
  FA_6828 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n635), .CI(C[122]), .S(S[122]), .CO(C[123]) );
  FA_6827 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n636), .CI(C[123]), .S(S[123]), .CO(C[124]) );
  FA_6826 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n637), .CI(C[124]), .S(S[124]), .CO(C[125]) );
  FA_6825 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n638), .CI(C[125]), .S(S[125]), .CO(C[126]) );
  FA_6824 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n639), .CI(C[126]), .S(S[126]), .CO(C[127]) );
  FA_6823 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n640), .CI(C[127]), .S(S[127]), .CO(C[128]) );
  FA_6822 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n641), .CI(C[128]), .S(S[128]), .CO(C[129]) );
  FA_6821 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n642), .CI(C[129]), .S(S[129]), .CO(C[130]) );
  FA_6820 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n643), .CI(C[130]), .S(S[130]), .CO(C[131]) );
  FA_6819 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n644), .CI(C[131]), .S(S[131]), .CO(C[132]) );
  FA_6818 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n645), .CI(C[132]), .S(S[132]), .CO(C[133]) );
  FA_6817 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n646), .CI(C[133]), .S(S[133]), .CO(C[134]) );
  FA_6816 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n647), .CI(C[134]), .S(S[134]), .CO(C[135]) );
  FA_6815 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n648), .CI(C[135]), .S(S[135]), .CO(C[136]) );
  FA_6814 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n649), .CI(C[136]), .S(S[136]), .CO(C[137]) );
  FA_6813 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n650), .CI(C[137]), .S(S[137]), .CO(C[138]) );
  FA_6812 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n651), .CI(C[138]), .S(S[138]), .CO(C[139]) );
  FA_6811 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n652), .CI(C[139]), .S(S[139]), .CO(C[140]) );
  FA_6810 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n653), .CI(C[140]), .S(S[140]), .CO(C[141]) );
  FA_6809 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n654), .CI(C[141]), .S(S[141]), .CO(C[142]) );
  FA_6808 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n655), .CI(C[142]), .S(S[142]), .CO(C[143]) );
  FA_6807 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n656), .CI(C[143]), .S(S[143]), .CO(C[144]) );
  FA_6806 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n657), .CI(C[144]), .S(S[144]), .CO(C[145]) );
  FA_6805 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n658), .CI(C[145]), .S(S[145]), .CO(C[146]) );
  FA_6804 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n659), .CI(C[146]), .S(S[146]), .CO(C[147]) );
  FA_6803 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n660), .CI(C[147]), .S(S[147]), .CO(C[148]) );
  FA_6802 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n661), .CI(C[148]), .S(S[148]), .CO(C[149]) );
  FA_6801 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n662), .CI(C[149]), .S(S[149]), .CO(C[150]) );
  FA_6800 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n663), .CI(C[150]), .S(S[150]), .CO(C[151]) );
  FA_6799 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n664), .CI(C[151]), .S(S[151]), .CO(C[152]) );
  FA_6798 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n665), .CI(C[152]), .S(S[152]), .CO(C[153]) );
  FA_6797 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n666), .CI(C[153]), .S(S[153]), .CO(C[154]) );
  FA_6796 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n667), .CI(C[154]), .S(S[154]), .CO(C[155]) );
  FA_6795 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n668), .CI(C[155]), .S(S[155]), .CO(C[156]) );
  FA_6794 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n669), .CI(C[156]), .S(S[156]), .CO(C[157]) );
  FA_6793 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n670), .CI(C[157]), .S(S[157]), .CO(C[158]) );
  FA_6792 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n671), .CI(C[158]), .S(S[158]), .CO(C[159]) );
  FA_6791 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n672), .CI(C[159]), .S(S[159]), .CO(C[160]) );
  FA_6790 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n673), .CI(C[160]), .S(S[160]), .CO(C[161]) );
  FA_6789 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n674), .CI(C[161]), .S(S[161]), .CO(C[162]) );
  FA_6788 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n675), .CI(C[162]), .S(S[162]), .CO(C[163]) );
  FA_6787 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n676), .CI(C[163]), .S(S[163]), .CO(C[164]) );
  FA_6786 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n677), .CI(C[164]), .S(S[164]), .CO(C[165]) );
  FA_6785 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n678), .CI(C[165]), .S(S[165]), .CO(C[166]) );
  FA_6784 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n679), .CI(C[166]), .S(S[166]), .CO(C[167]) );
  FA_6783 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n680), .CI(C[167]), .S(S[167]), .CO(C[168]) );
  FA_6782 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n681), .CI(C[168]), .S(S[168]), .CO(C[169]) );
  FA_6781 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n682), .CI(C[169]), .S(S[169]), .CO(C[170]) );
  FA_6780 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n683), .CI(C[170]), .S(S[170]), .CO(C[171]) );
  FA_6779 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n684), .CI(C[171]), .S(S[171]), .CO(C[172]) );
  FA_6778 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n685), .CI(C[172]), .S(S[172]), .CO(C[173]) );
  FA_6777 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n686), .CI(C[173]), .S(S[173]), .CO(C[174]) );
  FA_6776 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n687), .CI(C[174]), .S(S[174]), .CO(C[175]) );
  FA_6775 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n688), .CI(C[175]), .S(S[175]), .CO(C[176]) );
  FA_6774 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n689), .CI(C[176]), .S(S[176]), .CO(C[177]) );
  FA_6773 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n690), .CI(C[177]), .S(S[177]), .CO(C[178]) );
  FA_6772 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n691), .CI(C[178]), .S(S[178]), .CO(C[179]) );
  FA_6771 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n692), .CI(C[179]), .S(S[179]), .CO(C[180]) );
  FA_6770 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n693), .CI(C[180]), .S(S[180]), .CO(C[181]) );
  FA_6769 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n694), .CI(C[181]), .S(S[181]), .CO(C[182]) );
  FA_6768 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n695), .CI(C[182]), .S(S[182]), .CO(C[183]) );
  FA_6767 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n696), .CI(C[183]), .S(S[183]), .CO(C[184]) );
  FA_6766 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n697), .CI(C[184]), .S(S[184]), .CO(C[185]) );
  FA_6765 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n698), .CI(C[185]), .S(S[185]), .CO(C[186]) );
  FA_6764 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n699), .CI(C[186]), .S(S[186]), .CO(C[187]) );
  FA_6763 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n700), .CI(C[187]), .S(S[187]), .CO(C[188]) );
  FA_6762 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n701), .CI(C[188]), .S(S[188]), .CO(C[189]) );
  FA_6761 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n702), .CI(C[189]), .S(S[189]), .CO(C[190]) );
  FA_6760 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n703), .CI(C[190]), .S(S[190]), .CO(C[191]) );
  FA_6759 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n704), .CI(C[191]), .S(S[191]), .CO(C[192]) );
  FA_6758 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n705), .CI(C[192]), .S(S[192]), .CO(C[193]) );
  FA_6757 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n706), .CI(C[193]), .S(S[193]), .CO(C[194]) );
  FA_6756 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n707), .CI(C[194]), .S(S[194]), .CO(C[195]) );
  FA_6755 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n708), .CI(C[195]), .S(S[195]), .CO(C[196]) );
  FA_6754 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n709), .CI(C[196]), .S(S[196]), .CO(C[197]) );
  FA_6753 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n710), .CI(C[197]), .S(S[197]), .CO(C[198]) );
  FA_6752 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n711), .CI(C[198]), .S(S[198]), .CO(C[199]) );
  FA_6751 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n712), .CI(C[199]), .S(S[199]), .CO(C[200]) );
  FA_6750 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n713), .CI(C[200]), .S(S[200]), .CO(C[201]) );
  FA_6749 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n714), .CI(C[201]), .S(S[201]), .CO(C[202]) );
  FA_6748 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n715), .CI(C[202]), .S(S[202]), .CO(C[203]) );
  FA_6747 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n716), .CI(C[203]), .S(S[203]), .CO(C[204]) );
  FA_6746 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n717), .CI(C[204]), .S(S[204]), .CO(C[205]) );
  FA_6745 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n718), .CI(C[205]), .S(S[205]), .CO(C[206]) );
  FA_6744 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n719), .CI(C[206]), .S(S[206]), .CO(C[207]) );
  FA_6743 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n720), .CI(C[207]), .S(S[207]), .CO(C[208]) );
  FA_6742 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n721), .CI(C[208]), .S(S[208]), .CO(C[209]) );
  FA_6741 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n722), .CI(C[209]), .S(S[209]), .CO(C[210]) );
  FA_6740 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n723), .CI(C[210]), .S(S[210]), .CO(C[211]) );
  FA_6739 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n724), .CI(C[211]), .S(S[211]), .CO(C[212]) );
  FA_6738 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n725), .CI(C[212]), .S(S[212]), .CO(C[213]) );
  FA_6737 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n726), .CI(C[213]), .S(S[213]), .CO(C[214]) );
  FA_6736 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n727), .CI(C[214]), .S(S[214]), .CO(C[215]) );
  FA_6735 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n728), .CI(C[215]), .S(S[215]), .CO(C[216]) );
  FA_6734 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n729), .CI(C[216]), .S(S[216]), .CO(C[217]) );
  FA_6733 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n730), .CI(C[217]), .S(S[217]), .CO(C[218]) );
  FA_6732 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n731), .CI(C[218]), .S(S[218]), .CO(C[219]) );
  FA_6731 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n732), .CI(C[219]), .S(S[219]), .CO(C[220]) );
  FA_6730 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n733), .CI(C[220]), .S(S[220]), .CO(C[221]) );
  FA_6729 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n734), .CI(C[221]), .S(S[221]), .CO(C[222]) );
  FA_6728 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n735), .CI(C[222]), .S(S[222]), .CO(C[223]) );
  FA_6727 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n736), .CI(C[223]), .S(S[223]), .CO(C[224]) );
  FA_6726 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n737), .CI(C[224]), .S(S[224]), .CO(C[225]) );
  FA_6725 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n738), .CI(C[225]), .S(S[225]), .CO(C[226]) );
  FA_6724 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n739), .CI(C[226]), .S(S[226]), .CO(C[227]) );
  FA_6723 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n740), .CI(C[227]), .S(S[227]), .CO(C[228]) );
  FA_6722 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n741), .CI(C[228]), .S(S[228]), .CO(C[229]) );
  FA_6721 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n742), .CI(C[229]), .S(S[229]), .CO(C[230]) );
  FA_6720 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n743), .CI(C[230]), .S(S[230]), .CO(C[231]) );
  FA_6719 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n744), .CI(C[231]), .S(S[231]), .CO(C[232]) );
  FA_6718 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n745), .CI(C[232]), .S(S[232]), .CO(C[233]) );
  FA_6717 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n746), .CI(C[233]), .S(S[233]), .CO(C[234]) );
  FA_6716 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n747), .CI(C[234]), .S(S[234]), .CO(C[235]) );
  FA_6715 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n748), .CI(C[235]), .S(S[235]), .CO(C[236]) );
  FA_6714 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n749), .CI(C[236]), .S(S[236]), .CO(C[237]) );
  FA_6713 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n750), .CI(C[237]), .S(S[237]), .CO(C[238]) );
  FA_6712 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n751), .CI(C[238]), .S(S[238]), .CO(C[239]) );
  FA_6711 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n752), .CI(C[239]), .S(S[239]), .CO(C[240]) );
  FA_6710 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n753), .CI(C[240]), .S(S[240]), .CO(C[241]) );
  FA_6709 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n754), .CI(C[241]), .S(S[241]), .CO(C[242]) );
  FA_6708 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n755), .CI(C[242]), .S(S[242]), .CO(C[243]) );
  FA_6707 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n756), .CI(C[243]), .S(S[243]), .CO(C[244]) );
  FA_6706 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n757), .CI(C[244]), .S(S[244]), .CO(C[245]) );
  FA_6705 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n758), .CI(C[245]), .S(S[245]), .CO(C[246]) );
  FA_6704 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n759), .CI(C[246]), .S(S[246]), .CO(C[247]) );
  FA_6703 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n760), .CI(C[247]), .S(S[247]), .CO(C[248]) );
  FA_6702 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n761), .CI(C[248]), .S(S[248]), .CO(C[249]) );
  FA_6701 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n762), .CI(C[249]), .S(S[249]), .CO(C[250]) );
  FA_6700 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n763), .CI(C[250]), .S(S[250]), .CO(C[251]) );
  FA_6699 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n764), .CI(C[251]), .S(S[251]), .CO(C[252]) );
  FA_6698 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n765), .CI(C[252]), .S(S[252]), .CO(C[253]) );
  FA_6697 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n766), .CI(C[253]), .S(S[253]), .CO(C[254]) );
  FA_6696 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n767), .CI(C[254]), .S(S[254]), .CO(C[255]) );
  FA_6695 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n768), .CI(C[255]), .S(S[255]), .CO(C[256]) );
  FA_6694 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n769), .CI(C[256]), .S(S[256]), .CO(C[257]) );
  FA_6693 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n770), .CI(C[257]), .S(S[257]), .CO(C[258]) );
  FA_6692 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n771), .CI(C[258]), .S(S[258]), .CO(C[259]) );
  FA_6691 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n772), .CI(C[259]), .S(S[259]), .CO(C[260]) );
  FA_6690 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n773), .CI(C[260]), .S(S[260]), .CO(C[261]) );
  FA_6689 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n774), .CI(C[261]), .S(S[261]), .CO(C[262]) );
  FA_6688 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n775), .CI(C[262]), .S(S[262]), .CO(C[263]) );
  FA_6687 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n776), .CI(C[263]), .S(S[263]), .CO(C[264]) );
  FA_6686 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n777), .CI(C[264]), .S(S[264]), .CO(C[265]) );
  FA_6685 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n778), .CI(C[265]), .S(S[265]), .CO(C[266]) );
  FA_6684 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n779), .CI(C[266]), .S(S[266]), .CO(C[267]) );
  FA_6683 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n780), .CI(C[267]), .S(S[267]), .CO(C[268]) );
  FA_6682 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n781), .CI(C[268]), .S(S[268]), .CO(C[269]) );
  FA_6681 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n782), .CI(C[269]), .S(S[269]), .CO(C[270]) );
  FA_6680 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n783), .CI(C[270]), .S(S[270]), .CO(C[271]) );
  FA_6679 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n784), .CI(C[271]), .S(S[271]), .CO(C[272]) );
  FA_6678 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n785), .CI(C[272]), .S(S[272]), .CO(C[273]) );
  FA_6677 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n786), .CI(C[273]), .S(S[273]), .CO(C[274]) );
  FA_6676 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n787), .CI(C[274]), .S(S[274]), .CO(C[275]) );
  FA_6675 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n788), .CI(C[275]), .S(S[275]), .CO(C[276]) );
  FA_6674 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n789), .CI(C[276]), .S(S[276]), .CO(C[277]) );
  FA_6673 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n790), .CI(C[277]), .S(S[277]), .CO(C[278]) );
  FA_6672 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n791), .CI(C[278]), .S(S[278]), .CO(C[279]) );
  FA_6671 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n792), .CI(C[279]), .S(S[279]), .CO(C[280]) );
  FA_6670 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n793), .CI(C[280]), .S(S[280]), .CO(C[281]) );
  FA_6669 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n794), .CI(C[281]), .S(S[281]), .CO(C[282]) );
  FA_6668 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n795), .CI(C[282]), .S(S[282]), .CO(C[283]) );
  FA_6667 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n796), .CI(C[283]), .S(S[283]), .CO(C[284]) );
  FA_6666 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n797), .CI(C[284]), .S(S[284]), .CO(C[285]) );
  FA_6665 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n798), .CI(C[285]), .S(S[285]), .CO(C[286]) );
  FA_6664 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n799), .CI(C[286]), .S(S[286]), .CO(C[287]) );
  FA_6663 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n800), .CI(C[287]), .S(S[287]), .CO(C[288]) );
  FA_6662 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n801), .CI(C[288]), .S(S[288]), .CO(C[289]) );
  FA_6661 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n802), .CI(C[289]), .S(S[289]), .CO(C[290]) );
  FA_6660 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n803), .CI(C[290]), .S(S[290]), .CO(C[291]) );
  FA_6659 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n804), .CI(C[291]), .S(S[291]), .CO(C[292]) );
  FA_6658 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n805), .CI(C[292]), .S(S[292]), .CO(C[293]) );
  FA_6657 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n806), .CI(C[293]), .S(S[293]), .CO(C[294]) );
  FA_6656 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n807), .CI(C[294]), .S(S[294]), .CO(C[295]) );
  FA_6655 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n808), .CI(C[295]), .S(S[295]), .CO(C[296]) );
  FA_6654 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n809), .CI(C[296]), .S(S[296]), .CO(C[297]) );
  FA_6653 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n810), .CI(C[297]), .S(S[297]), .CO(C[298]) );
  FA_6652 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n811), .CI(C[298]), .S(S[298]), .CO(C[299]) );
  FA_6651 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n812), .CI(C[299]), .S(S[299]), .CO(C[300]) );
  FA_6650 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n813), .CI(C[300]), .S(S[300]), .CO(C[301]) );
  FA_6649 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n814), .CI(C[301]), .S(S[301]), .CO(C[302]) );
  FA_6648 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n815), .CI(C[302]), .S(S[302]), .CO(C[303]) );
  FA_6647 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n816), .CI(C[303]), .S(S[303]), .CO(C[304]) );
  FA_6646 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n817), .CI(C[304]), .S(S[304]), .CO(C[305]) );
  FA_6645 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n818), .CI(C[305]), .S(S[305]), .CO(C[306]) );
  FA_6644 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n819), .CI(C[306]), .S(S[306]), .CO(C[307]) );
  FA_6643 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n820), .CI(C[307]), .S(S[307]), .CO(C[308]) );
  FA_6642 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n821), .CI(C[308]), .S(S[308]), .CO(C[309]) );
  FA_6641 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n822), .CI(C[309]), .S(S[309]), .CO(C[310]) );
  FA_6640 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n823), .CI(C[310]), .S(S[310]), .CO(C[311]) );
  FA_6639 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n824), .CI(C[311]), .S(S[311]), .CO(C[312]) );
  FA_6638 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n825), .CI(C[312]), .S(S[312]), .CO(C[313]) );
  FA_6637 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n826), .CI(C[313]), .S(S[313]), .CO(C[314]) );
  FA_6636 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n827), .CI(C[314]), .S(S[314]), .CO(C[315]) );
  FA_6635 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n828), .CI(C[315]), .S(S[315]), .CO(C[316]) );
  FA_6634 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n829), .CI(C[316]), .S(S[316]), .CO(C[317]) );
  FA_6633 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n830), .CI(C[317]), .S(S[317]), .CO(C[318]) );
  FA_6632 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n831), .CI(C[318]), .S(S[318]), .CO(C[319]) );
  FA_6631 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n832), .CI(C[319]), .S(S[319]), .CO(C[320]) );
  FA_6630 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n833), .CI(C[320]), .S(S[320]), .CO(C[321]) );
  FA_6629 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n834), .CI(C[321]), .S(S[321]), .CO(C[322]) );
  FA_6628 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n835), .CI(C[322]), .S(S[322]), .CO(C[323]) );
  FA_6627 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n836), .CI(C[323]), .S(S[323]), .CO(C[324]) );
  FA_6626 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n837), .CI(C[324]), .S(S[324]), .CO(C[325]) );
  FA_6625 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n838), .CI(C[325]), .S(S[325]), .CO(C[326]) );
  FA_6624 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n839), .CI(C[326]), .S(S[326]), .CO(C[327]) );
  FA_6623 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n840), .CI(C[327]), .S(S[327]), .CO(C[328]) );
  FA_6622 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n841), .CI(C[328]), .S(S[328]), .CO(C[329]) );
  FA_6621 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n842), .CI(C[329]), .S(S[329]), .CO(C[330]) );
  FA_6620 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n843), .CI(C[330]), .S(S[330]), .CO(C[331]) );
  FA_6619 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n844), .CI(C[331]), .S(S[331]), .CO(C[332]) );
  FA_6618 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n845), .CI(C[332]), .S(S[332]), .CO(C[333]) );
  FA_6617 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n846), .CI(C[333]), .S(S[333]), .CO(C[334]) );
  FA_6616 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n847), .CI(C[334]), .S(S[334]), .CO(C[335]) );
  FA_6615 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n848), .CI(C[335]), .S(S[335]), .CO(C[336]) );
  FA_6614 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n849), .CI(C[336]), .S(S[336]), .CO(C[337]) );
  FA_6613 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n850), .CI(C[337]), .S(S[337]), .CO(C[338]) );
  FA_6612 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n851), .CI(C[338]), .S(S[338]), .CO(C[339]) );
  FA_6611 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n852), .CI(C[339]), .S(S[339]), .CO(C[340]) );
  FA_6610 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n853), .CI(C[340]), .S(S[340]), .CO(C[341]) );
  FA_6609 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n854), .CI(C[341]), .S(S[341]), .CO(C[342]) );
  FA_6608 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n855), .CI(C[342]), .S(S[342]), .CO(C[343]) );
  FA_6607 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n856), .CI(C[343]), .S(S[343]), .CO(C[344]) );
  FA_6606 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n857), .CI(C[344]), .S(S[344]), .CO(C[345]) );
  FA_6605 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n858), .CI(C[345]), .S(S[345]), .CO(C[346]) );
  FA_6604 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n859), .CI(C[346]), .S(S[346]), .CO(C[347]) );
  FA_6603 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n860), .CI(C[347]), .S(S[347]), .CO(C[348]) );
  FA_6602 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n861), .CI(C[348]), .S(S[348]), .CO(C[349]) );
  FA_6601 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n862), .CI(C[349]), .S(S[349]), .CO(C[350]) );
  FA_6600 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n863), .CI(C[350]), .S(S[350]), .CO(C[351]) );
  FA_6599 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n864), .CI(C[351]), .S(S[351]), .CO(C[352]) );
  FA_6598 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n865), .CI(C[352]), .S(S[352]), .CO(C[353]) );
  FA_6597 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n866), .CI(C[353]), .S(S[353]), .CO(C[354]) );
  FA_6596 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n867), .CI(C[354]), .S(S[354]), .CO(C[355]) );
  FA_6595 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n868), .CI(C[355]), .S(S[355]), .CO(C[356]) );
  FA_6594 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n869), .CI(C[356]), .S(S[356]), .CO(C[357]) );
  FA_6593 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n870), .CI(C[357]), .S(S[357]), .CO(C[358]) );
  FA_6592 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n871), .CI(C[358]), .S(S[358]), .CO(C[359]) );
  FA_6591 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n872), .CI(C[359]), .S(S[359]), .CO(C[360]) );
  FA_6590 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n873), .CI(C[360]), .S(S[360]), .CO(C[361]) );
  FA_6589 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n874), .CI(C[361]), .S(S[361]), .CO(C[362]) );
  FA_6588 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n875), .CI(C[362]), .S(S[362]), .CO(C[363]) );
  FA_6587 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n876), .CI(C[363]), .S(S[363]), .CO(C[364]) );
  FA_6586 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n877), .CI(C[364]), .S(S[364]), .CO(C[365]) );
  FA_6585 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n878), .CI(C[365]), .S(S[365]), .CO(C[366]) );
  FA_6584 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n879), .CI(C[366]), .S(S[366]), .CO(C[367]) );
  FA_6583 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n880), .CI(C[367]), .S(S[367]), .CO(C[368]) );
  FA_6582 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n881), .CI(C[368]), .S(S[368]), .CO(C[369]) );
  FA_6581 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n882), .CI(C[369]), .S(S[369]), .CO(C[370]) );
  FA_6580 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n883), .CI(C[370]), .S(S[370]), .CO(C[371]) );
  FA_6579 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n884), .CI(C[371]), .S(S[371]), .CO(C[372]) );
  FA_6578 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n885), .CI(C[372]), .S(S[372]), .CO(C[373]) );
  FA_6577 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n886), .CI(C[373]), .S(S[373]), .CO(C[374]) );
  FA_6576 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n887), .CI(C[374]), .S(S[374]), .CO(C[375]) );
  FA_6575 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n888), .CI(C[375]), .S(S[375]), .CO(C[376]) );
  FA_6574 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n889), .CI(C[376]), .S(S[376]), .CO(C[377]) );
  FA_6573 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n890), .CI(C[377]), .S(S[377]), .CO(C[378]) );
  FA_6572 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n891), .CI(C[378]), .S(S[378]), .CO(C[379]) );
  FA_6571 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n892), .CI(C[379]), .S(S[379]), .CO(C[380]) );
  FA_6570 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n893), .CI(C[380]), .S(S[380]), .CO(C[381]) );
  FA_6569 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n894), .CI(C[381]), .S(S[381]), .CO(C[382]) );
  FA_6568 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n895), .CI(C[382]), .S(S[382]), .CO(C[383]) );
  FA_6567 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n896), .CI(C[383]), .S(S[383]), .CO(C[384]) );
  FA_6566 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n897), .CI(C[384]), .S(S[384]), .CO(C[385]) );
  FA_6565 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n898), .CI(C[385]), .S(S[385]), .CO(C[386]) );
  FA_6564 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n899), .CI(C[386]), .S(S[386]), .CO(C[387]) );
  FA_6563 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n900), .CI(C[387]), .S(S[387]), .CO(C[388]) );
  FA_6562 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n901), .CI(C[388]), .S(S[388]), .CO(C[389]) );
  FA_6561 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n902), .CI(C[389]), .S(S[389]), .CO(C[390]) );
  FA_6560 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n903), .CI(C[390]), .S(S[390]), .CO(C[391]) );
  FA_6559 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n904), .CI(C[391]), .S(S[391]), .CO(C[392]) );
  FA_6558 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n905), .CI(C[392]), .S(S[392]), .CO(C[393]) );
  FA_6557 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n906), .CI(C[393]), .S(S[393]), .CO(C[394]) );
  FA_6556 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n907), .CI(C[394]), .S(S[394]), .CO(C[395]) );
  FA_6555 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n908), .CI(C[395]), .S(S[395]), .CO(C[396]) );
  FA_6554 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n909), .CI(C[396]), .S(S[396]), .CO(C[397]) );
  FA_6553 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n910), .CI(C[397]), .S(S[397]), .CO(C[398]) );
  FA_6552 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n911), .CI(C[398]), .S(S[398]), .CO(C[399]) );
  FA_6551 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n912), .CI(C[399]), .S(S[399]), .CO(C[400]) );
  FA_6550 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n913), .CI(C[400]), .S(S[400]), .CO(C[401]) );
  FA_6549 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n914), .CI(C[401]), .S(S[401]), .CO(C[402]) );
  FA_6548 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n915), .CI(C[402]), .S(S[402]), .CO(C[403]) );
  FA_6547 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n916), .CI(C[403]), .S(S[403]), .CO(C[404]) );
  FA_6546 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n917), .CI(C[404]), .S(S[404]), .CO(C[405]) );
  FA_6545 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n918), .CI(C[405]), .S(S[405]), .CO(C[406]) );
  FA_6544 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n919), .CI(C[406]), .S(S[406]), .CO(C[407]) );
  FA_6543 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n920), .CI(C[407]), .S(S[407]), .CO(C[408]) );
  FA_6542 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n921), .CI(C[408]), .S(S[408]), .CO(C[409]) );
  FA_6541 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n922), .CI(C[409]), .S(S[409]), .CO(C[410]) );
  FA_6540 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n923), .CI(C[410]), .S(S[410]), .CO(C[411]) );
  FA_6539 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n924), .CI(C[411]), .S(S[411]), .CO(C[412]) );
  FA_6538 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n925), .CI(C[412]), .S(S[412]), .CO(C[413]) );
  FA_6537 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n926), .CI(C[413]), .S(S[413]), .CO(C[414]) );
  FA_6536 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n927), .CI(C[414]), .S(S[414]), .CO(C[415]) );
  FA_6535 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n928), .CI(C[415]), .S(S[415]), .CO(C[416]) );
  FA_6534 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n929), .CI(C[416]), .S(S[416]), .CO(C[417]) );
  FA_6533 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n930), .CI(C[417]), .S(S[417]), .CO(C[418]) );
  FA_6532 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n931), .CI(C[418]), .S(S[418]), .CO(C[419]) );
  FA_6531 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n932), .CI(C[419]), .S(S[419]), .CO(C[420]) );
  FA_6530 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n933), .CI(C[420]), .S(S[420]), .CO(C[421]) );
  FA_6529 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n934), .CI(C[421]), .S(S[421]), .CO(C[422]) );
  FA_6528 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n935), .CI(C[422]), .S(S[422]), .CO(C[423]) );
  FA_6527 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n936), .CI(C[423]), .S(S[423]), .CO(C[424]) );
  FA_6526 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n937), .CI(C[424]), .S(S[424]), .CO(C[425]) );
  FA_6525 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n938), .CI(C[425]), .S(S[425]), .CO(C[426]) );
  FA_6524 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n939), .CI(C[426]), .S(S[426]), .CO(C[427]) );
  FA_6523 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n940), .CI(C[427]), .S(S[427]), .CO(C[428]) );
  FA_6522 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n941), .CI(C[428]), .S(S[428]), .CO(C[429]) );
  FA_6521 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n942), .CI(C[429]), .S(S[429]), .CO(C[430]) );
  FA_6520 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n943), .CI(C[430]), .S(S[430]), .CO(C[431]) );
  FA_6519 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n944), .CI(C[431]), .S(S[431]), .CO(C[432]) );
  FA_6518 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n945), .CI(C[432]), .S(S[432]), .CO(C[433]) );
  FA_6517 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n946), .CI(C[433]), .S(S[433]), .CO(C[434]) );
  FA_6516 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n947), .CI(C[434]), .S(S[434]), .CO(C[435]) );
  FA_6515 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n948), .CI(C[435]), .S(S[435]), .CO(C[436]) );
  FA_6514 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n949), .CI(C[436]), .S(S[436]), .CO(C[437]) );
  FA_6513 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n950), .CI(C[437]), .S(S[437]), .CO(C[438]) );
  FA_6512 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n951), .CI(C[438]), .S(S[438]), .CO(C[439]) );
  FA_6511 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n952), .CI(C[439]), .S(S[439]), .CO(C[440]) );
  FA_6510 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n953), .CI(C[440]), .S(S[440]), .CO(C[441]) );
  FA_6509 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n954), .CI(C[441]), .S(S[441]), .CO(C[442]) );
  FA_6508 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n955), .CI(C[442]), .S(S[442]), .CO(C[443]) );
  FA_6507 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n956), .CI(C[443]), .S(S[443]), .CO(C[444]) );
  FA_6506 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n957), .CI(C[444]), .S(S[444]), .CO(C[445]) );
  FA_6505 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n958), .CI(C[445]), .S(S[445]), .CO(C[446]) );
  FA_6504 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n959), .CI(C[446]), .S(S[446]), .CO(C[447]) );
  FA_6503 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n960), .CI(C[447]), .S(S[447]), .CO(C[448]) );
  FA_6502 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n961), .CI(C[448]), .S(S[448]), .CO(C[449]) );
  FA_6501 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n962), .CI(C[449]), .S(S[449]), .CO(C[450]) );
  FA_6500 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n963), .CI(C[450]), .S(S[450]), .CO(C[451]) );
  FA_6499 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n964), .CI(C[451]), .S(S[451]), .CO(C[452]) );
  FA_6498 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n965), .CI(C[452]), .S(S[452]), .CO(C[453]) );
  FA_6497 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n966), .CI(C[453]), .S(S[453]), .CO(C[454]) );
  FA_6496 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n967), .CI(C[454]), .S(S[454]), .CO(C[455]) );
  FA_6495 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n968), .CI(C[455]), .S(S[455]), .CO(C[456]) );
  FA_6494 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n969), .CI(C[456]), .S(S[456]), .CO(C[457]) );
  FA_6493 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n970), .CI(C[457]), .S(S[457]), .CO(C[458]) );
  FA_6492 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n971), .CI(C[458]), .S(S[458]), .CO(C[459]) );
  FA_6491 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n972), .CI(C[459]), .S(S[459]), .CO(C[460]) );
  FA_6490 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n973), .CI(C[460]), .S(S[460]), .CO(C[461]) );
  FA_6489 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n974), .CI(C[461]), .S(S[461]), .CO(C[462]) );
  FA_6488 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n975), .CI(C[462]), .S(S[462]), .CO(C[463]) );
  FA_6487 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n976), .CI(C[463]), .S(S[463]), .CO(C[464]) );
  FA_6486 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n977), .CI(C[464]), .S(S[464]), .CO(C[465]) );
  FA_6485 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n978), .CI(C[465]), .S(S[465]), .CO(C[466]) );
  FA_6484 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n979), .CI(C[466]), .S(S[466]), .CO(C[467]) );
  FA_6483 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n980), .CI(C[467]), .S(S[467]), .CO(C[468]) );
  FA_6482 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n981), .CI(C[468]), .S(S[468]), .CO(C[469]) );
  FA_6481 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n982), .CI(C[469]), .S(S[469]), .CO(C[470]) );
  FA_6480 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n983), .CI(C[470]), .S(S[470]), .CO(C[471]) );
  FA_6479 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n984), .CI(C[471]), .S(S[471]), .CO(C[472]) );
  FA_6478 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n985), .CI(C[472]), .S(S[472]), .CO(C[473]) );
  FA_6477 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n986), .CI(C[473]), .S(S[473]), .CO(C[474]) );
  FA_6476 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n987), .CI(C[474]), .S(S[474]), .CO(C[475]) );
  FA_6475 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n988), .CI(C[475]), .S(S[475]), .CO(C[476]) );
  FA_6474 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n989), .CI(C[476]), .S(S[476]), .CO(C[477]) );
  FA_6473 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n990), .CI(C[477]), .S(S[477]), .CO(C[478]) );
  FA_6472 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n991), .CI(C[478]), .S(S[478]), .CO(C[479]) );
  FA_6471 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n992), .CI(C[479]), .S(S[479]), .CO(C[480]) );
  FA_6470 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n993), .CI(C[480]), .S(S[480]), .CO(C[481]) );
  FA_6469 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n994), .CI(C[481]), .S(S[481]), .CO(C[482]) );
  FA_6468 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n995), .CI(C[482]), .S(S[482]), .CO(C[483]) );
  FA_6467 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n996), .CI(C[483]), .S(S[483]), .CO(C[484]) );
  FA_6466 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n997), .CI(C[484]), .S(S[484]), .CO(C[485]) );
  FA_6465 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n998), .CI(C[485]), .S(S[485]), .CO(C[486]) );
  FA_6464 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n999), .CI(C[486]), .S(S[486]), .CO(C[487]) );
  FA_6463 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1000), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_6462 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1001), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_6461 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1002), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_6460 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1003), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_6459 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1004), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_6458 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1005), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_6457 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1006), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_6456 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1007), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_6455 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1008), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_6454 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1009), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_6453 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1010), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_6452 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1011), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_6451 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1012), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_6450 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1013), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_6449 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1014), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_6448 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1015), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_6447 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1016), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_6446 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1017), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_6445 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1018), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_6444 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1019), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_6443 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1020), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_6442 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1021), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_6441 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1022), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_6440 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1023), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_6439 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1024), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_6438 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .S(S[512])
         );
  IV U2 ( .A(B[415]), .Z(n928) );
  IV U3 ( .A(B[416]), .Z(n929) );
  IV U4 ( .A(B[417]), .Z(n930) );
  IV U5 ( .A(B[418]), .Z(n931) );
  IV U6 ( .A(B[419]), .Z(n932) );
  IV U7 ( .A(B[420]), .Z(n933) );
  IV U8 ( .A(B[421]), .Z(n934) );
  IV U9 ( .A(B[422]), .Z(n935) );
  IV U10 ( .A(B[423]), .Z(n936) );
  IV U11 ( .A(B[424]), .Z(n937) );
  IV U12 ( .A(B[505]), .Z(n1018) );
  IV U13 ( .A(B[425]), .Z(n938) );
  IV U14 ( .A(B[426]), .Z(n939) );
  IV U15 ( .A(B[427]), .Z(n940) );
  IV U16 ( .A(B[428]), .Z(n941) );
  IV U17 ( .A(B[429]), .Z(n942) );
  IV U18 ( .A(B[430]), .Z(n943) );
  IV U19 ( .A(B[431]), .Z(n944) );
  IV U20 ( .A(B[432]), .Z(n945) );
  IV U21 ( .A(B[433]), .Z(n946) );
  IV U22 ( .A(B[434]), .Z(n947) );
  IV U23 ( .A(B[506]), .Z(n1019) );
  IV U24 ( .A(B[435]), .Z(n948) );
  IV U25 ( .A(B[436]), .Z(n949) );
  IV U26 ( .A(B[437]), .Z(n950) );
  IV U27 ( .A(B[438]), .Z(n951) );
  IV U28 ( .A(B[439]), .Z(n952) );
  IV U29 ( .A(B[440]), .Z(n953) );
  IV U30 ( .A(B[441]), .Z(n954) );
  IV U31 ( .A(B[442]), .Z(n955) );
  IV U32 ( .A(B[443]), .Z(n956) );
  IV U33 ( .A(B[444]), .Z(n957) );
  IV U34 ( .A(B[507]), .Z(n1020) );
  IV U35 ( .A(B[445]), .Z(n958) );
  IV U36 ( .A(B[446]), .Z(n959) );
  IV U37 ( .A(B[447]), .Z(n960) );
  IV U38 ( .A(B[448]), .Z(n961) );
  IV U39 ( .A(B[449]), .Z(n962) );
  IV U40 ( .A(B[450]), .Z(n963) );
  IV U41 ( .A(B[451]), .Z(n964) );
  IV U42 ( .A(B[452]), .Z(n965) );
  IV U43 ( .A(B[453]), .Z(n966) );
  IV U44 ( .A(B[454]), .Z(n967) );
  IV U45 ( .A(B[508]), .Z(n1021) );
  IV U46 ( .A(B[455]), .Z(n968) );
  IV U47 ( .A(B[456]), .Z(n969) );
  IV U48 ( .A(B[457]), .Z(n970) );
  IV U49 ( .A(B[458]), .Z(n971) );
  IV U50 ( .A(B[459]), .Z(n972) );
  IV U51 ( .A(B[460]), .Z(n973) );
  IV U52 ( .A(B[461]), .Z(n974) );
  IV U53 ( .A(B[462]), .Z(n975) );
  IV U54 ( .A(B[0]), .Z(n2) );
  IV U55 ( .A(B[1]), .Z(n514) );
  IV U56 ( .A(B[2]), .Z(n515) );
  IV U57 ( .A(B[3]), .Z(n516) );
  IV U58 ( .A(B[4]), .Z(n517) );
  IV U59 ( .A(B[463]), .Z(n976) );
  IV U60 ( .A(B[5]), .Z(n518) );
  IV U61 ( .A(B[6]), .Z(n519) );
  IV U62 ( .A(B[7]), .Z(n520) );
  IV U63 ( .A(B[8]), .Z(n521) );
  IV U64 ( .A(B[9]), .Z(n522) );
  IV U65 ( .A(B[10]), .Z(n523) );
  IV U66 ( .A(B[11]), .Z(n524) );
  IV U67 ( .A(B[12]), .Z(n525) );
  IV U68 ( .A(B[13]), .Z(n526) );
  IV U69 ( .A(B[14]), .Z(n527) );
  IV U70 ( .A(B[464]), .Z(n977) );
  IV U71 ( .A(B[509]), .Z(n1022) );
  IV U72 ( .A(B[15]), .Z(n528) );
  IV U73 ( .A(B[16]), .Z(n529) );
  IV U74 ( .A(B[17]), .Z(n530) );
  IV U75 ( .A(B[18]), .Z(n531) );
  IV U76 ( .A(B[19]), .Z(n532) );
  IV U77 ( .A(B[20]), .Z(n533) );
  IV U78 ( .A(B[21]), .Z(n534) );
  IV U79 ( .A(B[22]), .Z(n535) );
  IV U80 ( .A(B[23]), .Z(n536) );
  IV U81 ( .A(B[24]), .Z(n537) );
  IV U82 ( .A(B[465]), .Z(n978) );
  IV U83 ( .A(B[25]), .Z(n538) );
  IV U84 ( .A(B[26]), .Z(n539) );
  IV U85 ( .A(B[27]), .Z(n540) );
  IV U86 ( .A(B[28]), .Z(n541) );
  IV U87 ( .A(B[29]), .Z(n542) );
  IV U88 ( .A(B[30]), .Z(n543) );
  IV U89 ( .A(B[31]), .Z(n544) );
  IV U90 ( .A(B[32]), .Z(n545) );
  IV U91 ( .A(B[33]), .Z(n546) );
  IV U92 ( .A(B[34]), .Z(n547) );
  IV U93 ( .A(B[466]), .Z(n979) );
  IV U94 ( .A(B[35]), .Z(n548) );
  IV U95 ( .A(B[36]), .Z(n549) );
  IV U96 ( .A(B[37]), .Z(n550) );
  IV U97 ( .A(B[38]), .Z(n551) );
  IV U98 ( .A(B[39]), .Z(n552) );
  IV U99 ( .A(B[40]), .Z(n553) );
  IV U100 ( .A(B[41]), .Z(n554) );
  IV U101 ( .A(B[42]), .Z(n555) );
  IV U102 ( .A(B[43]), .Z(n556) );
  IV U103 ( .A(B[44]), .Z(n557) );
  IV U104 ( .A(B[467]), .Z(n980) );
  IV U105 ( .A(B[45]), .Z(n558) );
  IV U106 ( .A(B[46]), .Z(n559) );
  IV U107 ( .A(B[47]), .Z(n560) );
  IV U108 ( .A(B[48]), .Z(n561) );
  IV U109 ( .A(B[49]), .Z(n562) );
  IV U110 ( .A(B[50]), .Z(n563) );
  IV U111 ( .A(B[51]), .Z(n564) );
  IV U112 ( .A(B[52]), .Z(n565) );
  IV U113 ( .A(B[53]), .Z(n566) );
  IV U114 ( .A(B[54]), .Z(n567) );
  IV U115 ( .A(B[468]), .Z(n981) );
  IV U116 ( .A(B[55]), .Z(n568) );
  IV U117 ( .A(B[56]), .Z(n569) );
  IV U118 ( .A(B[57]), .Z(n570) );
  IV U119 ( .A(B[58]), .Z(n571) );
  IV U120 ( .A(B[59]), .Z(n572) );
  IV U121 ( .A(B[60]), .Z(n573) );
  IV U122 ( .A(B[61]), .Z(n574) );
  IV U123 ( .A(B[62]), .Z(n575) );
  IV U124 ( .A(B[63]), .Z(n576) );
  IV U125 ( .A(B[64]), .Z(n577) );
  IV U126 ( .A(B[469]), .Z(n982) );
  IV U127 ( .A(B[65]), .Z(n578) );
  IV U128 ( .A(B[66]), .Z(n579) );
  IV U129 ( .A(B[67]), .Z(n580) );
  IV U130 ( .A(B[68]), .Z(n581) );
  IV U131 ( .A(B[69]), .Z(n582) );
  IV U132 ( .A(B[70]), .Z(n583) );
  IV U133 ( .A(B[71]), .Z(n584) );
  IV U134 ( .A(B[72]), .Z(n585) );
  IV U135 ( .A(B[73]), .Z(n586) );
  IV U136 ( .A(B[74]), .Z(n587) );
  IV U137 ( .A(B[470]), .Z(n983) );
  IV U138 ( .A(B[75]), .Z(n588) );
  IV U139 ( .A(B[76]), .Z(n589) );
  IV U140 ( .A(B[77]), .Z(n590) );
  IV U141 ( .A(B[78]), .Z(n591) );
  IV U142 ( .A(B[79]), .Z(n592) );
  IV U143 ( .A(B[80]), .Z(n593) );
  IV U144 ( .A(B[81]), .Z(n594) );
  IV U145 ( .A(B[82]), .Z(n595) );
  IV U146 ( .A(B[83]), .Z(n596) );
  IV U147 ( .A(B[84]), .Z(n597) );
  IV U148 ( .A(B[471]), .Z(n984) );
  IV U149 ( .A(B[85]), .Z(n598) );
  IV U150 ( .A(B[86]), .Z(n599) );
  IV U151 ( .A(B[87]), .Z(n600) );
  IV U152 ( .A(B[88]), .Z(n601) );
  IV U153 ( .A(B[89]), .Z(n602) );
  IV U154 ( .A(B[90]), .Z(n603) );
  IV U155 ( .A(B[91]), .Z(n604) );
  IV U156 ( .A(B[92]), .Z(n605) );
  IV U157 ( .A(B[93]), .Z(n606) );
  IV U158 ( .A(B[94]), .Z(n607) );
  IV U159 ( .A(B[472]), .Z(n985) );
  IV U160 ( .A(B[95]), .Z(n608) );
  IV U161 ( .A(B[96]), .Z(n609) );
  IV U162 ( .A(B[97]), .Z(n610) );
  IV U163 ( .A(B[98]), .Z(n611) );
  IV U164 ( .A(B[99]), .Z(n612) );
  IV U165 ( .A(B[100]), .Z(n613) );
  IV U166 ( .A(B[101]), .Z(n614) );
  IV U167 ( .A(B[102]), .Z(n615) );
  IV U168 ( .A(B[103]), .Z(n616) );
  IV U169 ( .A(B[104]), .Z(n617) );
  IV U170 ( .A(B[473]), .Z(n986) );
  IV U171 ( .A(B[105]), .Z(n618) );
  IV U172 ( .A(B[106]), .Z(n619) );
  IV U173 ( .A(B[107]), .Z(n620) );
  IV U174 ( .A(B[108]), .Z(n621) );
  IV U175 ( .A(B[109]), .Z(n622) );
  IV U176 ( .A(B[110]), .Z(n623) );
  IV U177 ( .A(B[111]), .Z(n624) );
  IV U178 ( .A(B[112]), .Z(n625) );
  IV U179 ( .A(B[113]), .Z(n626) );
  IV U180 ( .A(B[114]), .Z(n627) );
  IV U181 ( .A(B[474]), .Z(n987) );
  IV U182 ( .A(B[510]), .Z(n1023) );
  IV U183 ( .A(B[115]), .Z(n628) );
  IV U184 ( .A(B[116]), .Z(n629) );
  IV U185 ( .A(B[117]), .Z(n630) );
  IV U186 ( .A(B[118]), .Z(n631) );
  IV U187 ( .A(B[119]), .Z(n632) );
  IV U188 ( .A(B[120]), .Z(n633) );
  IV U189 ( .A(B[121]), .Z(n634) );
  IV U190 ( .A(B[122]), .Z(n635) );
  IV U191 ( .A(B[123]), .Z(n636) );
  IV U192 ( .A(B[124]), .Z(n637) );
  IV U193 ( .A(B[475]), .Z(n988) );
  IV U194 ( .A(B[125]), .Z(n638) );
  IV U195 ( .A(B[126]), .Z(n639) );
  IV U196 ( .A(B[127]), .Z(n640) );
  IV U197 ( .A(B[128]), .Z(n641) );
  IV U198 ( .A(B[129]), .Z(n642) );
  IV U199 ( .A(B[130]), .Z(n643) );
  IV U200 ( .A(B[131]), .Z(n644) );
  IV U201 ( .A(B[132]), .Z(n645) );
  IV U202 ( .A(B[133]), .Z(n646) );
  IV U203 ( .A(B[134]), .Z(n647) );
  IV U204 ( .A(B[476]), .Z(n989) );
  IV U205 ( .A(B[135]), .Z(n648) );
  IV U206 ( .A(B[136]), .Z(n649) );
  IV U207 ( .A(B[137]), .Z(n650) );
  IV U208 ( .A(B[138]), .Z(n651) );
  IV U209 ( .A(B[139]), .Z(n652) );
  IV U210 ( .A(B[140]), .Z(n653) );
  IV U211 ( .A(B[141]), .Z(n654) );
  IV U212 ( .A(B[142]), .Z(n655) );
  IV U213 ( .A(B[143]), .Z(n656) );
  IV U214 ( .A(B[144]), .Z(n657) );
  IV U215 ( .A(B[477]), .Z(n990) );
  IV U216 ( .A(B[145]), .Z(n658) );
  IV U217 ( .A(B[146]), .Z(n659) );
  IV U218 ( .A(B[147]), .Z(n660) );
  IV U219 ( .A(B[148]), .Z(n661) );
  IV U220 ( .A(B[149]), .Z(n662) );
  IV U221 ( .A(B[150]), .Z(n663) );
  IV U222 ( .A(B[151]), .Z(n664) );
  IV U223 ( .A(B[152]), .Z(n665) );
  IV U224 ( .A(B[153]), .Z(n666) );
  IV U225 ( .A(B[154]), .Z(n667) );
  IV U226 ( .A(B[478]), .Z(n991) );
  IV U227 ( .A(B[155]), .Z(n668) );
  IV U228 ( .A(B[156]), .Z(n669) );
  IV U229 ( .A(B[157]), .Z(n670) );
  IV U230 ( .A(B[158]), .Z(n671) );
  IV U231 ( .A(B[159]), .Z(n672) );
  IV U232 ( .A(B[160]), .Z(n673) );
  IV U233 ( .A(B[161]), .Z(n674) );
  IV U234 ( .A(B[162]), .Z(n675) );
  IV U235 ( .A(B[163]), .Z(n676) );
  IV U236 ( .A(B[164]), .Z(n677) );
  IV U237 ( .A(B[479]), .Z(n992) );
  IV U238 ( .A(B[165]), .Z(n678) );
  IV U239 ( .A(B[166]), .Z(n679) );
  IV U240 ( .A(B[167]), .Z(n680) );
  IV U241 ( .A(B[168]), .Z(n681) );
  IV U242 ( .A(B[169]), .Z(n682) );
  IV U243 ( .A(B[170]), .Z(n683) );
  IV U244 ( .A(B[171]), .Z(n684) );
  IV U245 ( .A(B[172]), .Z(n685) );
  IV U246 ( .A(B[173]), .Z(n686) );
  IV U247 ( .A(B[174]), .Z(n687) );
  IV U248 ( .A(B[480]), .Z(n993) );
  IV U249 ( .A(B[175]), .Z(n688) );
  IV U250 ( .A(B[176]), .Z(n689) );
  IV U251 ( .A(B[177]), .Z(n690) );
  IV U252 ( .A(B[178]), .Z(n691) );
  IV U253 ( .A(B[179]), .Z(n692) );
  IV U254 ( .A(B[180]), .Z(n693) );
  IV U255 ( .A(B[181]), .Z(n694) );
  IV U256 ( .A(B[182]), .Z(n695) );
  IV U257 ( .A(B[183]), .Z(n696) );
  IV U258 ( .A(B[184]), .Z(n697) );
  IV U259 ( .A(B[481]), .Z(n994) );
  IV U260 ( .A(B[185]), .Z(n698) );
  IV U261 ( .A(B[186]), .Z(n699) );
  IV U262 ( .A(B[187]), .Z(n700) );
  IV U263 ( .A(B[188]), .Z(n701) );
  IV U264 ( .A(B[189]), .Z(n702) );
  IV U265 ( .A(B[190]), .Z(n703) );
  IV U266 ( .A(B[191]), .Z(n704) );
  IV U267 ( .A(B[192]), .Z(n705) );
  IV U268 ( .A(B[193]), .Z(n706) );
  IV U269 ( .A(B[194]), .Z(n707) );
  IV U270 ( .A(B[482]), .Z(n995) );
  IV U271 ( .A(B[195]), .Z(n708) );
  IV U272 ( .A(B[196]), .Z(n709) );
  IV U273 ( .A(B[197]), .Z(n710) );
  IV U274 ( .A(B[198]), .Z(n711) );
  IV U275 ( .A(B[199]), .Z(n712) );
  IV U276 ( .A(B[200]), .Z(n713) );
  IV U277 ( .A(B[201]), .Z(n714) );
  IV U278 ( .A(B[202]), .Z(n715) );
  IV U279 ( .A(B[203]), .Z(n716) );
  IV U280 ( .A(B[204]), .Z(n717) );
  IV U281 ( .A(B[483]), .Z(n996) );
  IV U282 ( .A(B[205]), .Z(n718) );
  IV U283 ( .A(B[206]), .Z(n719) );
  IV U284 ( .A(B[207]), .Z(n720) );
  IV U285 ( .A(B[208]), .Z(n721) );
  IV U286 ( .A(B[209]), .Z(n722) );
  IV U287 ( .A(B[210]), .Z(n723) );
  IV U288 ( .A(B[211]), .Z(n724) );
  IV U289 ( .A(B[212]), .Z(n725) );
  IV U290 ( .A(B[213]), .Z(n726) );
  IV U291 ( .A(B[214]), .Z(n727) );
  IV U292 ( .A(B[484]), .Z(n997) );
  IV U293 ( .A(B[511]), .Z(n1024) );
  IV U294 ( .A(B[215]), .Z(n728) );
  IV U295 ( .A(B[216]), .Z(n729) );
  IV U296 ( .A(B[217]), .Z(n730) );
  IV U297 ( .A(B[218]), .Z(n731) );
  IV U298 ( .A(B[219]), .Z(n732) );
  IV U299 ( .A(B[220]), .Z(n733) );
  IV U300 ( .A(B[221]), .Z(n734) );
  IV U301 ( .A(B[222]), .Z(n735) );
  IV U302 ( .A(B[223]), .Z(n736) );
  IV U303 ( .A(B[224]), .Z(n737) );
  IV U304 ( .A(B[485]), .Z(n998) );
  IV U305 ( .A(B[225]), .Z(n738) );
  IV U306 ( .A(B[226]), .Z(n739) );
  IV U307 ( .A(B[227]), .Z(n740) );
  IV U308 ( .A(B[228]), .Z(n741) );
  IV U309 ( .A(B[229]), .Z(n742) );
  IV U310 ( .A(B[230]), .Z(n743) );
  IV U311 ( .A(B[231]), .Z(n744) );
  IV U312 ( .A(B[232]), .Z(n745) );
  IV U313 ( .A(B[233]), .Z(n746) );
  IV U314 ( .A(B[234]), .Z(n747) );
  IV U315 ( .A(B[486]), .Z(n999) );
  IV U316 ( .A(B[235]), .Z(n748) );
  IV U317 ( .A(B[236]), .Z(n749) );
  IV U318 ( .A(B[237]), .Z(n750) );
  IV U319 ( .A(B[238]), .Z(n751) );
  IV U320 ( .A(B[239]), .Z(n752) );
  IV U321 ( .A(B[240]), .Z(n753) );
  IV U322 ( .A(B[241]), .Z(n754) );
  IV U323 ( .A(B[242]), .Z(n755) );
  IV U324 ( .A(B[243]), .Z(n756) );
  IV U325 ( .A(B[244]), .Z(n757) );
  IV U326 ( .A(B[487]), .Z(n1000) );
  IV U327 ( .A(B[245]), .Z(n758) );
  IV U328 ( .A(B[246]), .Z(n759) );
  IV U329 ( .A(B[247]), .Z(n760) );
  IV U330 ( .A(B[248]), .Z(n761) );
  IV U331 ( .A(B[249]), .Z(n762) );
  IV U332 ( .A(B[250]), .Z(n763) );
  IV U333 ( .A(B[251]), .Z(n764) );
  IV U334 ( .A(B[252]), .Z(n765) );
  IV U335 ( .A(B[253]), .Z(n766) );
  IV U336 ( .A(B[254]), .Z(n767) );
  IV U337 ( .A(B[488]), .Z(n1001) );
  IV U338 ( .A(B[255]), .Z(n768) );
  IV U339 ( .A(B[256]), .Z(n769) );
  IV U340 ( .A(B[257]), .Z(n770) );
  IV U341 ( .A(B[258]), .Z(n771) );
  IV U342 ( .A(B[259]), .Z(n772) );
  IV U343 ( .A(B[260]), .Z(n773) );
  IV U344 ( .A(B[261]), .Z(n774) );
  IV U345 ( .A(B[262]), .Z(n775) );
  IV U346 ( .A(B[263]), .Z(n776) );
  IV U347 ( .A(B[264]), .Z(n777) );
  IV U348 ( .A(B[489]), .Z(n1002) );
  IV U349 ( .A(B[265]), .Z(n778) );
  IV U350 ( .A(B[266]), .Z(n779) );
  IV U351 ( .A(B[267]), .Z(n780) );
  IV U352 ( .A(B[268]), .Z(n781) );
  IV U353 ( .A(B[269]), .Z(n782) );
  IV U354 ( .A(B[270]), .Z(n783) );
  IV U355 ( .A(B[271]), .Z(n784) );
  IV U356 ( .A(B[272]), .Z(n785) );
  IV U357 ( .A(B[273]), .Z(n786) );
  IV U358 ( .A(B[274]), .Z(n787) );
  IV U359 ( .A(B[490]), .Z(n1003) );
  IV U360 ( .A(B[275]), .Z(n788) );
  IV U361 ( .A(B[276]), .Z(n789) );
  IV U362 ( .A(B[277]), .Z(n790) );
  IV U363 ( .A(B[278]), .Z(n791) );
  IV U364 ( .A(B[279]), .Z(n792) );
  IV U365 ( .A(B[280]), .Z(n793) );
  IV U366 ( .A(B[281]), .Z(n794) );
  IV U367 ( .A(B[282]), .Z(n795) );
  IV U368 ( .A(B[283]), .Z(n796) );
  IV U369 ( .A(B[284]), .Z(n797) );
  IV U370 ( .A(B[491]), .Z(n1004) );
  IV U371 ( .A(B[285]), .Z(n798) );
  IV U372 ( .A(B[286]), .Z(n799) );
  IV U373 ( .A(B[287]), .Z(n800) );
  IV U374 ( .A(B[288]), .Z(n801) );
  IV U375 ( .A(B[289]), .Z(n802) );
  IV U376 ( .A(B[290]), .Z(n803) );
  IV U377 ( .A(B[291]), .Z(n804) );
  IV U378 ( .A(B[292]), .Z(n805) );
  IV U379 ( .A(B[293]), .Z(n806) );
  IV U380 ( .A(B[294]), .Z(n807) );
  IV U381 ( .A(B[492]), .Z(n1005) );
  IV U382 ( .A(B[295]), .Z(n808) );
  IV U383 ( .A(B[296]), .Z(n809) );
  IV U384 ( .A(B[297]), .Z(n810) );
  IV U385 ( .A(B[298]), .Z(n811) );
  IV U386 ( .A(B[299]), .Z(n812) );
  IV U387 ( .A(B[300]), .Z(n813) );
  IV U388 ( .A(B[301]), .Z(n814) );
  IV U389 ( .A(B[302]), .Z(n815) );
  IV U390 ( .A(B[303]), .Z(n816) );
  IV U391 ( .A(B[304]), .Z(n817) );
  IV U392 ( .A(B[493]), .Z(n1006) );
  IV U393 ( .A(B[305]), .Z(n818) );
  IV U394 ( .A(B[306]), .Z(n819) );
  IV U395 ( .A(B[307]), .Z(n820) );
  IV U396 ( .A(B[308]), .Z(n821) );
  IV U397 ( .A(B[309]), .Z(n822) );
  IV U398 ( .A(B[310]), .Z(n823) );
  IV U399 ( .A(B[311]), .Z(n824) );
  IV U400 ( .A(B[312]), .Z(n825) );
  IV U401 ( .A(B[313]), .Z(n826) );
  IV U402 ( .A(B[314]), .Z(n827) );
  IV U403 ( .A(B[494]), .Z(n1007) );
  IV U404 ( .A(B[315]), .Z(n828) );
  IV U405 ( .A(B[316]), .Z(n829) );
  IV U406 ( .A(B[317]), .Z(n830) );
  IV U407 ( .A(B[318]), .Z(n831) );
  IV U408 ( .A(B[319]), .Z(n832) );
  IV U409 ( .A(B[320]), .Z(n833) );
  IV U410 ( .A(B[321]), .Z(n834) );
  IV U411 ( .A(B[322]), .Z(n835) );
  IV U412 ( .A(B[323]), .Z(n836) );
  IV U413 ( .A(B[324]), .Z(n837) );
  IV U414 ( .A(B[495]), .Z(n1008) );
  IV U415 ( .A(B[325]), .Z(n838) );
  IV U416 ( .A(B[326]), .Z(n839) );
  IV U417 ( .A(B[327]), .Z(n840) );
  IV U418 ( .A(B[328]), .Z(n841) );
  IV U419 ( .A(B[329]), .Z(n842) );
  IV U420 ( .A(B[330]), .Z(n843) );
  IV U421 ( .A(B[331]), .Z(n844) );
  IV U422 ( .A(B[332]), .Z(n845) );
  IV U423 ( .A(B[333]), .Z(n846) );
  IV U424 ( .A(B[334]), .Z(n847) );
  IV U425 ( .A(B[496]), .Z(n1009) );
  IV U426 ( .A(B[335]), .Z(n848) );
  IV U427 ( .A(B[336]), .Z(n849) );
  IV U428 ( .A(B[337]), .Z(n850) );
  IV U429 ( .A(B[338]), .Z(n851) );
  IV U430 ( .A(B[339]), .Z(n852) );
  IV U431 ( .A(B[340]), .Z(n853) );
  IV U432 ( .A(B[341]), .Z(n854) );
  IV U433 ( .A(B[342]), .Z(n855) );
  IV U434 ( .A(B[343]), .Z(n856) );
  IV U435 ( .A(B[344]), .Z(n857) );
  IV U436 ( .A(B[497]), .Z(n1010) );
  IV U437 ( .A(B[345]), .Z(n858) );
  IV U438 ( .A(B[346]), .Z(n859) );
  IV U439 ( .A(B[347]), .Z(n860) );
  IV U440 ( .A(B[348]), .Z(n861) );
  IV U441 ( .A(B[349]), .Z(n862) );
  IV U442 ( .A(B[350]), .Z(n863) );
  IV U443 ( .A(B[351]), .Z(n864) );
  IV U444 ( .A(B[352]), .Z(n865) );
  IV U445 ( .A(B[353]), .Z(n866) );
  IV U446 ( .A(B[354]), .Z(n867) );
  IV U447 ( .A(B[498]), .Z(n1011) );
  IV U448 ( .A(B[355]), .Z(n868) );
  IV U449 ( .A(B[356]), .Z(n869) );
  IV U450 ( .A(B[357]), .Z(n870) );
  IV U451 ( .A(B[358]), .Z(n871) );
  IV U452 ( .A(B[359]), .Z(n872) );
  IV U453 ( .A(B[360]), .Z(n873) );
  IV U454 ( .A(B[361]), .Z(n874) );
  IV U455 ( .A(B[362]), .Z(n875) );
  IV U456 ( .A(B[363]), .Z(n876) );
  IV U457 ( .A(B[364]), .Z(n877) );
  IV U458 ( .A(B[499]), .Z(n1012) );
  IV U459 ( .A(B[365]), .Z(n878) );
  IV U460 ( .A(B[366]), .Z(n879) );
  IV U461 ( .A(B[367]), .Z(n880) );
  IV U462 ( .A(B[368]), .Z(n881) );
  IV U463 ( .A(B[369]), .Z(n882) );
  IV U464 ( .A(B[370]), .Z(n883) );
  IV U465 ( .A(B[371]), .Z(n884) );
  IV U466 ( .A(B[372]), .Z(n885) );
  IV U467 ( .A(B[373]), .Z(n886) );
  IV U468 ( .A(B[374]), .Z(n887) );
  IV U469 ( .A(B[500]), .Z(n1013) );
  IV U470 ( .A(B[375]), .Z(n888) );
  IV U471 ( .A(B[376]), .Z(n889) );
  IV U472 ( .A(B[377]), .Z(n890) );
  IV U473 ( .A(B[378]), .Z(n891) );
  IV U474 ( .A(B[379]), .Z(n892) );
  IV U475 ( .A(B[380]), .Z(n893) );
  IV U476 ( .A(B[381]), .Z(n894) );
  IV U477 ( .A(B[382]), .Z(n895) );
  IV U478 ( .A(B[383]), .Z(n896) );
  IV U479 ( .A(B[384]), .Z(n897) );
  IV U480 ( .A(B[501]), .Z(n1014) );
  IV U481 ( .A(B[385]), .Z(n898) );
  IV U482 ( .A(B[386]), .Z(n899) );
  IV U483 ( .A(B[387]), .Z(n900) );
  IV U484 ( .A(B[388]), .Z(n901) );
  IV U485 ( .A(B[389]), .Z(n902) );
  IV U486 ( .A(B[390]), .Z(n903) );
  IV U487 ( .A(B[391]), .Z(n904) );
  IV U488 ( .A(B[392]), .Z(n905) );
  IV U489 ( .A(B[393]), .Z(n906) );
  IV U490 ( .A(B[394]), .Z(n907) );
  IV U491 ( .A(B[502]), .Z(n1015) );
  IV U492 ( .A(B[395]), .Z(n908) );
  IV U493 ( .A(B[396]), .Z(n909) );
  IV U494 ( .A(B[397]), .Z(n910) );
  IV U495 ( .A(B[398]), .Z(n911) );
  IV U496 ( .A(B[399]), .Z(n912) );
  IV U497 ( .A(B[400]), .Z(n913) );
  IV U498 ( .A(B[401]), .Z(n914) );
  IV U499 ( .A(B[402]), .Z(n915) );
  IV U500 ( .A(B[403]), .Z(n916) );
  IV U501 ( .A(B[404]), .Z(n917) );
  IV U502 ( .A(B[503]), .Z(n1016) );
  IV U503 ( .A(B[405]), .Z(n918) );
  IV U504 ( .A(B[406]), .Z(n919) );
  IV U505 ( .A(B[407]), .Z(n920) );
  IV U506 ( .A(B[408]), .Z(n921) );
  IV U507 ( .A(B[409]), .Z(n922) );
  IV U508 ( .A(B[410]), .Z(n923) );
  IV U509 ( .A(B[411]), .Z(n924) );
  IV U510 ( .A(B[412]), .Z(n925) );
  IV U511 ( .A(B[413]), .Z(n926) );
  IV U512 ( .A(B[414]), .Z(n927) );
  IV U513 ( .A(B[504]), .Z(n1017) );
endmodule


module FA_7465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(CI), .B(A), .Z(S) );
endmodule


module FA_7466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  NANDN U1 ( .A(CI), .B(S), .Z(CO) );
  XNOR U2 ( .A(A), .B(CI), .Z(S) );
endmodule


module FA_7467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7512 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7513 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7514 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7515 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7516 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7517 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7518 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7519 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7520 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7521 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7522 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7523 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7524 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7525 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7526 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7527 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7528 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7529 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7530 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7531 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7532 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7533 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7534 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7535 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7536 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7537 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7538 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7539 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7540 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7541 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7542 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7543 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7544 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7545 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7546 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7547 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7548 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7549 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7550 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7551 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7552 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7553 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7554 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7555 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7556 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7557 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7558 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7559 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7560 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7561 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7562 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7563 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7564 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7565 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7566 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7567 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7568 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7569 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7570 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7571 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7572 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7573 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7574 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7575 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7576 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7577 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7578 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7579 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7580 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7581 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7582 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7583 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7584 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7585 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7586 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7587 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7588 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7589 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7590 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7591 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7592 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7593 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7594 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7595 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7596 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7597 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7598 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7599 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7600 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7601 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7602 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7603 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7604 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7605 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7606 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7607 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7608 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7609 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7610 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7611 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7612 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7613 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7614 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7615 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7616 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7617 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7618 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7619 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7620 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7621 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7622 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7623 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7624 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7625 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7626 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7627 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7628 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7629 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7630 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7631 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7632 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7633 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7634 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7635 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7636 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7637 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7638 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7639 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7640 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7641 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7642 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7643 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7644 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7645 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7646 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7647 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7648 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7649 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7650 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7651 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7652 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7653 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7654 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7655 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7656 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7657 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7658 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7659 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7660 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7661 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7662 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7663 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7664 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7665 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7666 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7667 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7668 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7669 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7670 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7671 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7672 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7673 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7674 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7675 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7676 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7677 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7678 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7679 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7680 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7681 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7682 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7683 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7684 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7685 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7686 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7687 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7688 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7689 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7690 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7691 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7692 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7693 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7694 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7695 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7696 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7697 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7698 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7699 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7700 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7701 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7702 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7703 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7704 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7705 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7706 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7707 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7708 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7709 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7710 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7711 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7712 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7713 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7714 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7715 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7716 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7717 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7718 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7719 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7720 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7721 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7722 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7723 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7724 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7725 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7726 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7727 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7728 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7729 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7730 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7731 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7732 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7733 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7734 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7735 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7736 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7737 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7738 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7739 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7740 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7741 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7742 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7743 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7744 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7745 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7746 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7747 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7748 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7749 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7750 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7751 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7752 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7753 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7754 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7755 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7756 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7757 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7758 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7759 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7760 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7761 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7762 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7763 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7764 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7765 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7766 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7767 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7768 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7769 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7770 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7771 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7772 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7773 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7774 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7775 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7776 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7777 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7778 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7779 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7780 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7781 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7782 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7783 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7784 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7785 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7786 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7787 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7788 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7789 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7790 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7791 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7792 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7793 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7794 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7795 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7796 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7797 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7798 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7799 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7800 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7801 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7802 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7803 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7804 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7805 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7806 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7807 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7808 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7809 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7810 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7811 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7812 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7813 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7814 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7815 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7816 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7817 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7818 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7819 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7820 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7821 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7822 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7823 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7824 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7825 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7826 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7827 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7828 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7829 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7830 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7831 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7832 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7833 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7834 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7835 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7836 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7837 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7838 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7839 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7840 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7841 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7842 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7843 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7844 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7845 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7846 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7847 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7848 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7849 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7850 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7851 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7852 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7853 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7854 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7855 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7856 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7857 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7858 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7859 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7860 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7861 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7862 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7863 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7864 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7865 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7866 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7867 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7868 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7869 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7870 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7871 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7872 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7873 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7874 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7875 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7876 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7877 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7878 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7879 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7880 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7881 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7882 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7883 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7884 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7885 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7886 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7887 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7888 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7889 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7890 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7891 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7892 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7893 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7894 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7895 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7896 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7897 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7898 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7899 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7900 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7901 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7902 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7903 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7904 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7905 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7906 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7907 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7908 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7909 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7910 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7911 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7912 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7913 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7914 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7915 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7916 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7917 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7918 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7919 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7920 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7921 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7922 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7923 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7924 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7925 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7926 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7927 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7928 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7929 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7930 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7931 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7932 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7933 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7934 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7935 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7936 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7937 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7938 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7939 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7940 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7941 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7942 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7943 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7944 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7945 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7946 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7947 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7948 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7949 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7950 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7951 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7952 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7953 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7954 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7955 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7956 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7957 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7958 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7959 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7960 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7961 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7962 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7963 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7964 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7965 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7966 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7967 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7968 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7969 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7970 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7971 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7972 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7973 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7974 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7975 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7976 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7977 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3, n4;

  XOR U1 ( .A(B), .B(n1), .Z(S) );
  XOR U2 ( .A(CI), .B(n2), .Z(CO) );
  AND U3 ( .A(n1), .B(n3), .Z(n2) );
  XNOR U4 ( .A(n4), .B(B), .Z(n3) );
  IV U5 ( .A(CI), .Z(n4) );
  XOR U6 ( .A(A), .B(CI), .Z(n1) );
endmodule


module FA_7978 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  XNOR U1 ( .A(B), .B(A), .Z(S) );
  OR U2 ( .A(B), .B(A), .Z(CO) );
endmodule


module SUB_N514_4 ( A, B, S, CO );
  input [513:0] A;
  input [513:0] B;
  output [513:0] S;
  output CO;
  wire   n2, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024;
  wire   [513:1] C;

  FA_7978 \FA_INST_0[0].FA_INST_1[0].FA_  ( .A(A[0]), .B(n2), .CI(1'b1), .S(
        S[0]), .CO(C[1]) );
  FA_7977 \FA_INST_0[0].FA_INST_1[1].FA_  ( .A(A[1]), .B(n514), .CI(C[1]), .S(
        S[1]), .CO(C[2]) );
  FA_7976 \FA_INST_0[0].FA_INST_1[2].FA_  ( .A(A[2]), .B(n515), .CI(C[2]), .S(
        S[2]), .CO(C[3]) );
  FA_7975 \FA_INST_0[0].FA_INST_1[3].FA_  ( .A(A[3]), .B(n516), .CI(C[3]), .S(
        S[3]), .CO(C[4]) );
  FA_7974 \FA_INST_0[0].FA_INST_1[4].FA_  ( .A(A[4]), .B(n517), .CI(C[4]), .S(
        S[4]), .CO(C[5]) );
  FA_7973 \FA_INST_0[0].FA_INST_1[5].FA_  ( .A(A[5]), .B(n518), .CI(C[5]), .S(
        S[5]), .CO(C[6]) );
  FA_7972 \FA_INST_0[0].FA_INST_1[6].FA_  ( .A(A[6]), .B(n519), .CI(C[6]), .S(
        S[6]), .CO(C[7]) );
  FA_7971 \FA_INST_0[0].FA_INST_1[7].FA_  ( .A(A[7]), .B(n520), .CI(C[7]), .S(
        S[7]), .CO(C[8]) );
  FA_7970 \FA_INST_0[0].FA_INST_1[8].FA_  ( .A(A[8]), .B(n521), .CI(C[8]), .S(
        S[8]), .CO(C[9]) );
  FA_7969 \FA_INST_0[0].FA_INST_1[9].FA_  ( .A(A[9]), .B(n522), .CI(C[9]), .S(
        S[9]), .CO(C[10]) );
  FA_7968 \FA_INST_0[0].FA_INST_1[10].FA_  ( .A(A[10]), .B(n523), .CI(C[10]), 
        .S(S[10]), .CO(C[11]) );
  FA_7967 \FA_INST_0[0].FA_INST_1[11].FA_  ( .A(A[11]), .B(n524), .CI(C[11]), 
        .S(S[11]), .CO(C[12]) );
  FA_7966 \FA_INST_0[0].FA_INST_1[12].FA_  ( .A(A[12]), .B(n525), .CI(C[12]), 
        .S(S[12]), .CO(C[13]) );
  FA_7965 \FA_INST_0[0].FA_INST_1[13].FA_  ( .A(A[13]), .B(n526), .CI(C[13]), 
        .S(S[13]), .CO(C[14]) );
  FA_7964 \FA_INST_0[0].FA_INST_1[14].FA_  ( .A(A[14]), .B(n527), .CI(C[14]), 
        .S(S[14]), .CO(C[15]) );
  FA_7963 \FA_INST_0[0].FA_INST_1[15].FA_  ( .A(A[15]), .B(n528), .CI(C[15]), 
        .S(S[15]), .CO(C[16]) );
  FA_7962 \FA_INST_0[0].FA_INST_1[16].FA_  ( .A(A[16]), .B(n529), .CI(C[16]), 
        .S(S[16]), .CO(C[17]) );
  FA_7961 \FA_INST_0[0].FA_INST_1[17].FA_  ( .A(A[17]), .B(n530), .CI(C[17]), 
        .S(S[17]), .CO(C[18]) );
  FA_7960 \FA_INST_0[0].FA_INST_1[18].FA_  ( .A(A[18]), .B(n531), .CI(C[18]), 
        .S(S[18]), .CO(C[19]) );
  FA_7959 \FA_INST_0[0].FA_INST_1[19].FA_  ( .A(A[19]), .B(n532), .CI(C[19]), 
        .S(S[19]), .CO(C[20]) );
  FA_7958 \FA_INST_0[0].FA_INST_1[20].FA_  ( .A(A[20]), .B(n533), .CI(C[20]), 
        .S(S[20]), .CO(C[21]) );
  FA_7957 \FA_INST_0[0].FA_INST_1[21].FA_  ( .A(A[21]), .B(n534), .CI(C[21]), 
        .S(S[21]), .CO(C[22]) );
  FA_7956 \FA_INST_0[0].FA_INST_1[22].FA_  ( .A(A[22]), .B(n535), .CI(C[22]), 
        .S(S[22]), .CO(C[23]) );
  FA_7955 \FA_INST_0[0].FA_INST_1[23].FA_  ( .A(A[23]), .B(n536), .CI(C[23]), 
        .S(S[23]), .CO(C[24]) );
  FA_7954 \FA_INST_0[0].FA_INST_1[24].FA_  ( .A(A[24]), .B(n537), .CI(C[24]), 
        .S(S[24]), .CO(C[25]) );
  FA_7953 \FA_INST_0[0].FA_INST_1[25].FA_  ( .A(A[25]), .B(n538), .CI(C[25]), 
        .S(S[25]), .CO(C[26]) );
  FA_7952 \FA_INST_0[0].FA_INST_1[26].FA_  ( .A(A[26]), .B(n539), .CI(C[26]), 
        .S(S[26]), .CO(C[27]) );
  FA_7951 \FA_INST_0[0].FA_INST_1[27].FA_  ( .A(A[27]), .B(n540), .CI(C[27]), 
        .S(S[27]), .CO(C[28]) );
  FA_7950 \FA_INST_0[0].FA_INST_1[28].FA_  ( .A(A[28]), .B(n541), .CI(C[28]), 
        .S(S[28]), .CO(C[29]) );
  FA_7949 \FA_INST_0[0].FA_INST_1[29].FA_  ( .A(A[29]), .B(n542), .CI(C[29]), 
        .S(S[29]), .CO(C[30]) );
  FA_7948 \FA_INST_0[0].FA_INST_1[30].FA_  ( .A(A[30]), .B(n543), .CI(C[30]), 
        .S(S[30]), .CO(C[31]) );
  FA_7947 \FA_INST_0[0].FA_INST_1[31].FA_  ( .A(A[31]), .B(n544), .CI(C[31]), 
        .S(S[31]), .CO(C[32]) );
  FA_7946 \FA_INST_0[0].FA_INST_1[32].FA_  ( .A(A[32]), .B(n545), .CI(C[32]), 
        .S(S[32]), .CO(C[33]) );
  FA_7945 \FA_INST_0[0].FA_INST_1[33].FA_  ( .A(A[33]), .B(n546), .CI(C[33]), 
        .S(S[33]), .CO(C[34]) );
  FA_7944 \FA_INST_0[0].FA_INST_1[34].FA_  ( .A(A[34]), .B(n547), .CI(C[34]), 
        .S(S[34]), .CO(C[35]) );
  FA_7943 \FA_INST_0[0].FA_INST_1[35].FA_  ( .A(A[35]), .B(n548), .CI(C[35]), 
        .S(S[35]), .CO(C[36]) );
  FA_7942 \FA_INST_0[0].FA_INST_1[36].FA_  ( .A(A[36]), .B(n549), .CI(C[36]), 
        .S(S[36]), .CO(C[37]) );
  FA_7941 \FA_INST_0[0].FA_INST_1[37].FA_  ( .A(A[37]), .B(n550), .CI(C[37]), 
        .S(S[37]), .CO(C[38]) );
  FA_7940 \FA_INST_0[0].FA_INST_1[38].FA_  ( .A(A[38]), .B(n551), .CI(C[38]), 
        .S(S[38]), .CO(C[39]) );
  FA_7939 \FA_INST_0[0].FA_INST_1[39].FA_  ( .A(A[39]), .B(n552), .CI(C[39]), 
        .S(S[39]), .CO(C[40]) );
  FA_7938 \FA_INST_0[0].FA_INST_1[40].FA_  ( .A(A[40]), .B(n553), .CI(C[40]), 
        .S(S[40]), .CO(C[41]) );
  FA_7937 \FA_INST_0[0].FA_INST_1[41].FA_  ( .A(A[41]), .B(n554), .CI(C[41]), 
        .S(S[41]), .CO(C[42]) );
  FA_7936 \FA_INST_0[0].FA_INST_1[42].FA_  ( .A(A[42]), .B(n555), .CI(C[42]), 
        .S(S[42]), .CO(C[43]) );
  FA_7935 \FA_INST_0[0].FA_INST_1[43].FA_  ( .A(A[43]), .B(n556), .CI(C[43]), 
        .S(S[43]), .CO(C[44]) );
  FA_7934 \FA_INST_0[0].FA_INST_1[44].FA_  ( .A(A[44]), .B(n557), .CI(C[44]), 
        .S(S[44]), .CO(C[45]) );
  FA_7933 \FA_INST_0[0].FA_INST_1[45].FA_  ( .A(A[45]), .B(n558), .CI(C[45]), 
        .S(S[45]), .CO(C[46]) );
  FA_7932 \FA_INST_0[0].FA_INST_1[46].FA_  ( .A(A[46]), .B(n559), .CI(C[46]), 
        .S(S[46]), .CO(C[47]) );
  FA_7931 \FA_INST_0[0].FA_INST_1[47].FA_  ( .A(A[47]), .B(n560), .CI(C[47]), 
        .S(S[47]), .CO(C[48]) );
  FA_7930 \FA_INST_0[0].FA_INST_1[48].FA_  ( .A(A[48]), .B(n561), .CI(C[48]), 
        .S(S[48]), .CO(C[49]) );
  FA_7929 \FA_INST_0[0].FA_INST_1[49].FA_  ( .A(A[49]), .B(n562), .CI(C[49]), 
        .S(S[49]), .CO(C[50]) );
  FA_7928 \FA_INST_0[0].FA_INST_1[50].FA_  ( .A(A[50]), .B(n563), .CI(C[50]), 
        .S(S[50]), .CO(C[51]) );
  FA_7927 \FA_INST_0[0].FA_INST_1[51].FA_  ( .A(A[51]), .B(n564), .CI(C[51]), 
        .S(S[51]), .CO(C[52]) );
  FA_7926 \FA_INST_0[0].FA_INST_1[52].FA_  ( .A(A[52]), .B(n565), .CI(C[52]), 
        .S(S[52]), .CO(C[53]) );
  FA_7925 \FA_INST_0[0].FA_INST_1[53].FA_  ( .A(A[53]), .B(n566), .CI(C[53]), 
        .S(S[53]), .CO(C[54]) );
  FA_7924 \FA_INST_0[0].FA_INST_1[54].FA_  ( .A(A[54]), .B(n567), .CI(C[54]), 
        .S(S[54]), .CO(C[55]) );
  FA_7923 \FA_INST_0[0].FA_INST_1[55].FA_  ( .A(A[55]), .B(n568), .CI(C[55]), 
        .S(S[55]), .CO(C[56]) );
  FA_7922 \FA_INST_0[0].FA_INST_1[56].FA_  ( .A(A[56]), .B(n569), .CI(C[56]), 
        .S(S[56]), .CO(C[57]) );
  FA_7921 \FA_INST_0[0].FA_INST_1[57].FA_  ( .A(A[57]), .B(n570), .CI(C[57]), 
        .S(S[57]), .CO(C[58]) );
  FA_7920 \FA_INST_0[0].FA_INST_1[58].FA_  ( .A(A[58]), .B(n571), .CI(C[58]), 
        .S(S[58]), .CO(C[59]) );
  FA_7919 \FA_INST_0[0].FA_INST_1[59].FA_  ( .A(A[59]), .B(n572), .CI(C[59]), 
        .S(S[59]), .CO(C[60]) );
  FA_7918 \FA_INST_0[0].FA_INST_1[60].FA_  ( .A(A[60]), .B(n573), .CI(C[60]), 
        .S(S[60]), .CO(C[61]) );
  FA_7917 \FA_INST_0[0].FA_INST_1[61].FA_  ( .A(A[61]), .B(n574), .CI(C[61]), 
        .S(S[61]), .CO(C[62]) );
  FA_7916 \FA_INST_0[0].FA_INST_1[62].FA_  ( .A(A[62]), .B(n575), .CI(C[62]), 
        .S(S[62]), .CO(C[63]) );
  FA_7915 \FA_INST_0[0].FA_INST_1[63].FA_  ( .A(A[63]), .B(n576), .CI(C[63]), 
        .S(S[63]), .CO(C[64]) );
  FA_7914 \FA_INST_0[0].FA_INST_1[64].FA_  ( .A(A[64]), .B(n577), .CI(C[64]), 
        .S(S[64]), .CO(C[65]) );
  FA_7913 \FA_INST_0[0].FA_INST_1[65].FA_  ( .A(A[65]), .B(n578), .CI(C[65]), 
        .S(S[65]), .CO(C[66]) );
  FA_7912 \FA_INST_0[0].FA_INST_1[66].FA_  ( .A(A[66]), .B(n579), .CI(C[66]), 
        .S(S[66]), .CO(C[67]) );
  FA_7911 \FA_INST_0[0].FA_INST_1[67].FA_  ( .A(A[67]), .B(n580), .CI(C[67]), 
        .S(S[67]), .CO(C[68]) );
  FA_7910 \FA_INST_0[0].FA_INST_1[68].FA_  ( .A(A[68]), .B(n581), .CI(C[68]), 
        .S(S[68]), .CO(C[69]) );
  FA_7909 \FA_INST_0[0].FA_INST_1[69].FA_  ( .A(A[69]), .B(n582), .CI(C[69]), 
        .S(S[69]), .CO(C[70]) );
  FA_7908 \FA_INST_0[0].FA_INST_1[70].FA_  ( .A(A[70]), .B(n583), .CI(C[70]), 
        .S(S[70]), .CO(C[71]) );
  FA_7907 \FA_INST_0[0].FA_INST_1[71].FA_  ( .A(A[71]), .B(n584), .CI(C[71]), 
        .S(S[71]), .CO(C[72]) );
  FA_7906 \FA_INST_0[0].FA_INST_1[72].FA_  ( .A(A[72]), .B(n585), .CI(C[72]), 
        .S(S[72]), .CO(C[73]) );
  FA_7905 \FA_INST_0[0].FA_INST_1[73].FA_  ( .A(A[73]), .B(n586), .CI(C[73]), 
        .S(S[73]), .CO(C[74]) );
  FA_7904 \FA_INST_0[0].FA_INST_1[74].FA_  ( .A(A[74]), .B(n587), .CI(C[74]), 
        .S(S[74]), .CO(C[75]) );
  FA_7903 \FA_INST_0[0].FA_INST_1[75].FA_  ( .A(A[75]), .B(n588), .CI(C[75]), 
        .S(S[75]), .CO(C[76]) );
  FA_7902 \FA_INST_0[0].FA_INST_1[76].FA_  ( .A(A[76]), .B(n589), .CI(C[76]), 
        .S(S[76]), .CO(C[77]) );
  FA_7901 \FA_INST_0[0].FA_INST_1[77].FA_  ( .A(A[77]), .B(n590), .CI(C[77]), 
        .S(S[77]), .CO(C[78]) );
  FA_7900 \FA_INST_0[0].FA_INST_1[78].FA_  ( .A(A[78]), .B(n591), .CI(C[78]), 
        .S(S[78]), .CO(C[79]) );
  FA_7899 \FA_INST_0[0].FA_INST_1[79].FA_  ( .A(A[79]), .B(n592), .CI(C[79]), 
        .S(S[79]), .CO(C[80]) );
  FA_7898 \FA_INST_0[0].FA_INST_1[80].FA_  ( .A(A[80]), .B(n593), .CI(C[80]), 
        .S(S[80]), .CO(C[81]) );
  FA_7897 \FA_INST_0[0].FA_INST_1[81].FA_  ( .A(A[81]), .B(n594), .CI(C[81]), 
        .S(S[81]), .CO(C[82]) );
  FA_7896 \FA_INST_0[0].FA_INST_1[82].FA_  ( .A(A[82]), .B(n595), .CI(C[82]), 
        .S(S[82]), .CO(C[83]) );
  FA_7895 \FA_INST_0[0].FA_INST_1[83].FA_  ( .A(A[83]), .B(n596), .CI(C[83]), 
        .S(S[83]), .CO(C[84]) );
  FA_7894 \FA_INST_0[0].FA_INST_1[84].FA_  ( .A(A[84]), .B(n597), .CI(C[84]), 
        .S(S[84]), .CO(C[85]) );
  FA_7893 \FA_INST_0[0].FA_INST_1[85].FA_  ( .A(A[85]), .B(n598), .CI(C[85]), 
        .S(S[85]), .CO(C[86]) );
  FA_7892 \FA_INST_0[0].FA_INST_1[86].FA_  ( .A(A[86]), .B(n599), .CI(C[86]), 
        .S(S[86]), .CO(C[87]) );
  FA_7891 \FA_INST_0[0].FA_INST_1[87].FA_  ( .A(A[87]), .B(n600), .CI(C[87]), 
        .S(S[87]), .CO(C[88]) );
  FA_7890 \FA_INST_0[0].FA_INST_1[88].FA_  ( .A(A[88]), .B(n601), .CI(C[88]), 
        .S(S[88]), .CO(C[89]) );
  FA_7889 \FA_INST_0[0].FA_INST_1[89].FA_  ( .A(A[89]), .B(n602), .CI(C[89]), 
        .S(S[89]), .CO(C[90]) );
  FA_7888 \FA_INST_0[0].FA_INST_1[90].FA_  ( .A(A[90]), .B(n603), .CI(C[90]), 
        .S(S[90]), .CO(C[91]) );
  FA_7887 \FA_INST_0[0].FA_INST_1[91].FA_  ( .A(A[91]), .B(n604), .CI(C[91]), 
        .S(S[91]), .CO(C[92]) );
  FA_7886 \FA_INST_0[0].FA_INST_1[92].FA_  ( .A(A[92]), .B(n605), .CI(C[92]), 
        .S(S[92]), .CO(C[93]) );
  FA_7885 \FA_INST_0[0].FA_INST_1[93].FA_  ( .A(A[93]), .B(n606), .CI(C[93]), 
        .S(S[93]), .CO(C[94]) );
  FA_7884 \FA_INST_0[0].FA_INST_1[94].FA_  ( .A(A[94]), .B(n607), .CI(C[94]), 
        .S(S[94]), .CO(C[95]) );
  FA_7883 \FA_INST_0[0].FA_INST_1[95].FA_  ( .A(A[95]), .B(n608), .CI(C[95]), 
        .S(S[95]), .CO(C[96]) );
  FA_7882 \FA_INST_0[0].FA_INST_1[96].FA_  ( .A(A[96]), .B(n609), .CI(C[96]), 
        .S(S[96]), .CO(C[97]) );
  FA_7881 \FA_INST_0[0].FA_INST_1[97].FA_  ( .A(A[97]), .B(n610), .CI(C[97]), 
        .S(S[97]), .CO(C[98]) );
  FA_7880 \FA_INST_0[0].FA_INST_1[98].FA_  ( .A(A[98]), .B(n611), .CI(C[98]), 
        .S(S[98]), .CO(C[99]) );
  FA_7879 \FA_INST_0[0].FA_INST_1[99].FA_  ( .A(A[99]), .B(n612), .CI(C[99]), 
        .S(S[99]), .CO(C[100]) );
  FA_7878 \FA_INST_0[0].FA_INST_1[100].FA_  ( .A(A[100]), .B(n613), .CI(C[100]), .S(S[100]), .CO(C[101]) );
  FA_7877 \FA_INST_0[0].FA_INST_1[101].FA_  ( .A(A[101]), .B(n614), .CI(C[101]), .S(S[101]), .CO(C[102]) );
  FA_7876 \FA_INST_0[0].FA_INST_1[102].FA_  ( .A(A[102]), .B(n615), .CI(C[102]), .S(S[102]), .CO(C[103]) );
  FA_7875 \FA_INST_0[0].FA_INST_1[103].FA_  ( .A(A[103]), .B(n616), .CI(C[103]), .S(S[103]), .CO(C[104]) );
  FA_7874 \FA_INST_0[0].FA_INST_1[104].FA_  ( .A(A[104]), .B(n617), .CI(C[104]), .S(S[104]), .CO(C[105]) );
  FA_7873 \FA_INST_0[0].FA_INST_1[105].FA_  ( .A(A[105]), .B(n618), .CI(C[105]), .S(S[105]), .CO(C[106]) );
  FA_7872 \FA_INST_0[0].FA_INST_1[106].FA_  ( .A(A[106]), .B(n619), .CI(C[106]), .S(S[106]), .CO(C[107]) );
  FA_7871 \FA_INST_0[0].FA_INST_1[107].FA_  ( .A(A[107]), .B(n620), .CI(C[107]), .S(S[107]), .CO(C[108]) );
  FA_7870 \FA_INST_0[0].FA_INST_1[108].FA_  ( .A(A[108]), .B(n621), .CI(C[108]), .S(S[108]), .CO(C[109]) );
  FA_7869 \FA_INST_0[0].FA_INST_1[109].FA_  ( .A(A[109]), .B(n622), .CI(C[109]), .S(S[109]), .CO(C[110]) );
  FA_7868 \FA_INST_0[0].FA_INST_1[110].FA_  ( .A(A[110]), .B(n623), .CI(C[110]), .S(S[110]), .CO(C[111]) );
  FA_7867 \FA_INST_0[0].FA_INST_1[111].FA_  ( .A(A[111]), .B(n624), .CI(C[111]), .S(S[111]), .CO(C[112]) );
  FA_7866 \FA_INST_0[0].FA_INST_1[112].FA_  ( .A(A[112]), .B(n625), .CI(C[112]), .S(S[112]), .CO(C[113]) );
  FA_7865 \FA_INST_0[0].FA_INST_1[113].FA_  ( .A(A[113]), .B(n626), .CI(C[113]), .S(S[113]), .CO(C[114]) );
  FA_7864 \FA_INST_0[0].FA_INST_1[114].FA_  ( .A(A[114]), .B(n627), .CI(C[114]), .S(S[114]), .CO(C[115]) );
  FA_7863 \FA_INST_0[0].FA_INST_1[115].FA_  ( .A(A[115]), .B(n628), .CI(C[115]), .S(S[115]), .CO(C[116]) );
  FA_7862 \FA_INST_0[0].FA_INST_1[116].FA_  ( .A(A[116]), .B(n629), .CI(C[116]), .S(S[116]), .CO(C[117]) );
  FA_7861 \FA_INST_0[0].FA_INST_1[117].FA_  ( .A(A[117]), .B(n630), .CI(C[117]), .S(S[117]), .CO(C[118]) );
  FA_7860 \FA_INST_0[0].FA_INST_1[118].FA_  ( .A(A[118]), .B(n631), .CI(C[118]), .S(S[118]), .CO(C[119]) );
  FA_7859 \FA_INST_0[0].FA_INST_1[119].FA_  ( .A(A[119]), .B(n632), .CI(C[119]), .S(S[119]), .CO(C[120]) );
  FA_7858 \FA_INST_0[0].FA_INST_1[120].FA_  ( .A(A[120]), .B(n633), .CI(C[120]), .S(S[120]), .CO(C[121]) );
  FA_7857 \FA_INST_0[0].FA_INST_1[121].FA_  ( .A(A[121]), .B(n634), .CI(C[121]), .S(S[121]), .CO(C[122]) );
  FA_7856 \FA_INST_0[0].FA_INST_1[122].FA_  ( .A(A[122]), .B(n635), .CI(C[122]), .S(S[122]), .CO(C[123]) );
  FA_7855 \FA_INST_0[0].FA_INST_1[123].FA_  ( .A(A[123]), .B(n636), .CI(C[123]), .S(S[123]), .CO(C[124]) );
  FA_7854 \FA_INST_0[0].FA_INST_1[124].FA_  ( .A(A[124]), .B(n637), .CI(C[124]), .S(S[124]), .CO(C[125]) );
  FA_7853 \FA_INST_0[0].FA_INST_1[125].FA_  ( .A(A[125]), .B(n638), .CI(C[125]), .S(S[125]), .CO(C[126]) );
  FA_7852 \FA_INST_0[0].FA_INST_1[126].FA_  ( .A(A[126]), .B(n639), .CI(C[126]), .S(S[126]), .CO(C[127]) );
  FA_7851 \FA_INST_0[0].FA_INST_1[127].FA_  ( .A(A[127]), .B(n640), .CI(C[127]), .S(S[127]), .CO(C[128]) );
  FA_7850 \FA_INST_0[0].FA_INST_1[128].FA_  ( .A(A[128]), .B(n641), .CI(C[128]), .S(S[128]), .CO(C[129]) );
  FA_7849 \FA_INST_0[0].FA_INST_1[129].FA_  ( .A(A[129]), .B(n642), .CI(C[129]), .S(S[129]), .CO(C[130]) );
  FA_7848 \FA_INST_0[0].FA_INST_1[130].FA_  ( .A(A[130]), .B(n643), .CI(C[130]), .S(S[130]), .CO(C[131]) );
  FA_7847 \FA_INST_0[0].FA_INST_1[131].FA_  ( .A(A[131]), .B(n644), .CI(C[131]), .S(S[131]), .CO(C[132]) );
  FA_7846 \FA_INST_0[0].FA_INST_1[132].FA_  ( .A(A[132]), .B(n645), .CI(C[132]), .S(S[132]), .CO(C[133]) );
  FA_7845 \FA_INST_0[0].FA_INST_1[133].FA_  ( .A(A[133]), .B(n646), .CI(C[133]), .S(S[133]), .CO(C[134]) );
  FA_7844 \FA_INST_0[0].FA_INST_1[134].FA_  ( .A(A[134]), .B(n647), .CI(C[134]), .S(S[134]), .CO(C[135]) );
  FA_7843 \FA_INST_0[0].FA_INST_1[135].FA_  ( .A(A[135]), .B(n648), .CI(C[135]), .S(S[135]), .CO(C[136]) );
  FA_7842 \FA_INST_0[0].FA_INST_1[136].FA_  ( .A(A[136]), .B(n649), .CI(C[136]), .S(S[136]), .CO(C[137]) );
  FA_7841 \FA_INST_0[0].FA_INST_1[137].FA_  ( .A(A[137]), .B(n650), .CI(C[137]), .S(S[137]), .CO(C[138]) );
  FA_7840 \FA_INST_0[0].FA_INST_1[138].FA_  ( .A(A[138]), .B(n651), .CI(C[138]), .S(S[138]), .CO(C[139]) );
  FA_7839 \FA_INST_0[0].FA_INST_1[139].FA_  ( .A(A[139]), .B(n652), .CI(C[139]), .S(S[139]), .CO(C[140]) );
  FA_7838 \FA_INST_0[0].FA_INST_1[140].FA_  ( .A(A[140]), .B(n653), .CI(C[140]), .S(S[140]), .CO(C[141]) );
  FA_7837 \FA_INST_0[0].FA_INST_1[141].FA_  ( .A(A[141]), .B(n654), .CI(C[141]), .S(S[141]), .CO(C[142]) );
  FA_7836 \FA_INST_0[0].FA_INST_1[142].FA_  ( .A(A[142]), .B(n655), .CI(C[142]), .S(S[142]), .CO(C[143]) );
  FA_7835 \FA_INST_0[0].FA_INST_1[143].FA_  ( .A(A[143]), .B(n656), .CI(C[143]), .S(S[143]), .CO(C[144]) );
  FA_7834 \FA_INST_0[0].FA_INST_1[144].FA_  ( .A(A[144]), .B(n657), .CI(C[144]), .S(S[144]), .CO(C[145]) );
  FA_7833 \FA_INST_0[0].FA_INST_1[145].FA_  ( .A(A[145]), .B(n658), .CI(C[145]), .S(S[145]), .CO(C[146]) );
  FA_7832 \FA_INST_0[0].FA_INST_1[146].FA_  ( .A(A[146]), .B(n659), .CI(C[146]), .S(S[146]), .CO(C[147]) );
  FA_7831 \FA_INST_0[0].FA_INST_1[147].FA_  ( .A(A[147]), .B(n660), .CI(C[147]), .S(S[147]), .CO(C[148]) );
  FA_7830 \FA_INST_0[0].FA_INST_1[148].FA_  ( .A(A[148]), .B(n661), .CI(C[148]), .S(S[148]), .CO(C[149]) );
  FA_7829 \FA_INST_0[0].FA_INST_1[149].FA_  ( .A(A[149]), .B(n662), .CI(C[149]), .S(S[149]), .CO(C[150]) );
  FA_7828 \FA_INST_0[0].FA_INST_1[150].FA_  ( .A(A[150]), .B(n663), .CI(C[150]), .S(S[150]), .CO(C[151]) );
  FA_7827 \FA_INST_0[0].FA_INST_1[151].FA_  ( .A(A[151]), .B(n664), .CI(C[151]), .S(S[151]), .CO(C[152]) );
  FA_7826 \FA_INST_0[0].FA_INST_1[152].FA_  ( .A(A[152]), .B(n665), .CI(C[152]), .S(S[152]), .CO(C[153]) );
  FA_7825 \FA_INST_0[0].FA_INST_1[153].FA_  ( .A(A[153]), .B(n666), .CI(C[153]), .S(S[153]), .CO(C[154]) );
  FA_7824 \FA_INST_0[0].FA_INST_1[154].FA_  ( .A(A[154]), .B(n667), .CI(C[154]), .S(S[154]), .CO(C[155]) );
  FA_7823 \FA_INST_0[0].FA_INST_1[155].FA_  ( .A(A[155]), .B(n668), .CI(C[155]), .S(S[155]), .CO(C[156]) );
  FA_7822 \FA_INST_0[0].FA_INST_1[156].FA_  ( .A(A[156]), .B(n669), .CI(C[156]), .S(S[156]), .CO(C[157]) );
  FA_7821 \FA_INST_0[0].FA_INST_1[157].FA_  ( .A(A[157]), .B(n670), .CI(C[157]), .S(S[157]), .CO(C[158]) );
  FA_7820 \FA_INST_0[0].FA_INST_1[158].FA_  ( .A(A[158]), .B(n671), .CI(C[158]), .S(S[158]), .CO(C[159]) );
  FA_7819 \FA_INST_0[0].FA_INST_1[159].FA_  ( .A(A[159]), .B(n672), .CI(C[159]), .S(S[159]), .CO(C[160]) );
  FA_7818 \FA_INST_0[0].FA_INST_1[160].FA_  ( .A(A[160]), .B(n673), .CI(C[160]), .S(S[160]), .CO(C[161]) );
  FA_7817 \FA_INST_0[0].FA_INST_1[161].FA_  ( .A(A[161]), .B(n674), .CI(C[161]), .S(S[161]), .CO(C[162]) );
  FA_7816 \FA_INST_0[0].FA_INST_1[162].FA_  ( .A(A[162]), .B(n675), .CI(C[162]), .S(S[162]), .CO(C[163]) );
  FA_7815 \FA_INST_0[0].FA_INST_1[163].FA_  ( .A(A[163]), .B(n676), .CI(C[163]), .S(S[163]), .CO(C[164]) );
  FA_7814 \FA_INST_0[0].FA_INST_1[164].FA_  ( .A(A[164]), .B(n677), .CI(C[164]), .S(S[164]), .CO(C[165]) );
  FA_7813 \FA_INST_0[0].FA_INST_1[165].FA_  ( .A(A[165]), .B(n678), .CI(C[165]), .S(S[165]), .CO(C[166]) );
  FA_7812 \FA_INST_0[0].FA_INST_1[166].FA_  ( .A(A[166]), .B(n679), .CI(C[166]), .S(S[166]), .CO(C[167]) );
  FA_7811 \FA_INST_0[0].FA_INST_1[167].FA_  ( .A(A[167]), .B(n680), .CI(C[167]), .S(S[167]), .CO(C[168]) );
  FA_7810 \FA_INST_0[0].FA_INST_1[168].FA_  ( .A(A[168]), .B(n681), .CI(C[168]), .S(S[168]), .CO(C[169]) );
  FA_7809 \FA_INST_0[0].FA_INST_1[169].FA_  ( .A(A[169]), .B(n682), .CI(C[169]), .S(S[169]), .CO(C[170]) );
  FA_7808 \FA_INST_0[0].FA_INST_1[170].FA_  ( .A(A[170]), .B(n683), .CI(C[170]), .S(S[170]), .CO(C[171]) );
  FA_7807 \FA_INST_0[0].FA_INST_1[171].FA_  ( .A(A[171]), .B(n684), .CI(C[171]), .S(S[171]), .CO(C[172]) );
  FA_7806 \FA_INST_0[0].FA_INST_1[172].FA_  ( .A(A[172]), .B(n685), .CI(C[172]), .S(S[172]), .CO(C[173]) );
  FA_7805 \FA_INST_0[0].FA_INST_1[173].FA_  ( .A(A[173]), .B(n686), .CI(C[173]), .S(S[173]), .CO(C[174]) );
  FA_7804 \FA_INST_0[0].FA_INST_1[174].FA_  ( .A(A[174]), .B(n687), .CI(C[174]), .S(S[174]), .CO(C[175]) );
  FA_7803 \FA_INST_0[0].FA_INST_1[175].FA_  ( .A(A[175]), .B(n688), .CI(C[175]), .S(S[175]), .CO(C[176]) );
  FA_7802 \FA_INST_0[0].FA_INST_1[176].FA_  ( .A(A[176]), .B(n689), .CI(C[176]), .S(S[176]), .CO(C[177]) );
  FA_7801 \FA_INST_0[0].FA_INST_1[177].FA_  ( .A(A[177]), .B(n690), .CI(C[177]), .S(S[177]), .CO(C[178]) );
  FA_7800 \FA_INST_0[0].FA_INST_1[178].FA_  ( .A(A[178]), .B(n691), .CI(C[178]), .S(S[178]), .CO(C[179]) );
  FA_7799 \FA_INST_0[0].FA_INST_1[179].FA_  ( .A(A[179]), .B(n692), .CI(C[179]), .S(S[179]), .CO(C[180]) );
  FA_7798 \FA_INST_0[0].FA_INST_1[180].FA_  ( .A(A[180]), .B(n693), .CI(C[180]), .S(S[180]), .CO(C[181]) );
  FA_7797 \FA_INST_0[0].FA_INST_1[181].FA_  ( .A(A[181]), .B(n694), .CI(C[181]), .S(S[181]), .CO(C[182]) );
  FA_7796 \FA_INST_0[0].FA_INST_1[182].FA_  ( .A(A[182]), .B(n695), .CI(C[182]), .S(S[182]), .CO(C[183]) );
  FA_7795 \FA_INST_0[0].FA_INST_1[183].FA_  ( .A(A[183]), .B(n696), .CI(C[183]), .S(S[183]), .CO(C[184]) );
  FA_7794 \FA_INST_0[0].FA_INST_1[184].FA_  ( .A(A[184]), .B(n697), .CI(C[184]), .S(S[184]), .CO(C[185]) );
  FA_7793 \FA_INST_0[0].FA_INST_1[185].FA_  ( .A(A[185]), .B(n698), .CI(C[185]), .S(S[185]), .CO(C[186]) );
  FA_7792 \FA_INST_0[0].FA_INST_1[186].FA_  ( .A(A[186]), .B(n699), .CI(C[186]), .S(S[186]), .CO(C[187]) );
  FA_7791 \FA_INST_0[0].FA_INST_1[187].FA_  ( .A(A[187]), .B(n700), .CI(C[187]), .S(S[187]), .CO(C[188]) );
  FA_7790 \FA_INST_0[0].FA_INST_1[188].FA_  ( .A(A[188]), .B(n701), .CI(C[188]), .S(S[188]), .CO(C[189]) );
  FA_7789 \FA_INST_0[0].FA_INST_1[189].FA_  ( .A(A[189]), .B(n702), .CI(C[189]), .S(S[189]), .CO(C[190]) );
  FA_7788 \FA_INST_0[0].FA_INST_1[190].FA_  ( .A(A[190]), .B(n703), .CI(C[190]), .S(S[190]), .CO(C[191]) );
  FA_7787 \FA_INST_0[0].FA_INST_1[191].FA_  ( .A(A[191]), .B(n704), .CI(C[191]), .S(S[191]), .CO(C[192]) );
  FA_7786 \FA_INST_0[0].FA_INST_1[192].FA_  ( .A(A[192]), .B(n705), .CI(C[192]), .S(S[192]), .CO(C[193]) );
  FA_7785 \FA_INST_0[0].FA_INST_1[193].FA_  ( .A(A[193]), .B(n706), .CI(C[193]), .S(S[193]), .CO(C[194]) );
  FA_7784 \FA_INST_0[0].FA_INST_1[194].FA_  ( .A(A[194]), .B(n707), .CI(C[194]), .S(S[194]), .CO(C[195]) );
  FA_7783 \FA_INST_0[0].FA_INST_1[195].FA_  ( .A(A[195]), .B(n708), .CI(C[195]), .S(S[195]), .CO(C[196]) );
  FA_7782 \FA_INST_0[0].FA_INST_1[196].FA_  ( .A(A[196]), .B(n709), .CI(C[196]), .S(S[196]), .CO(C[197]) );
  FA_7781 \FA_INST_0[0].FA_INST_1[197].FA_  ( .A(A[197]), .B(n710), .CI(C[197]), .S(S[197]), .CO(C[198]) );
  FA_7780 \FA_INST_0[0].FA_INST_1[198].FA_  ( .A(A[198]), .B(n711), .CI(C[198]), .S(S[198]), .CO(C[199]) );
  FA_7779 \FA_INST_0[0].FA_INST_1[199].FA_  ( .A(A[199]), .B(n712), .CI(C[199]), .S(S[199]), .CO(C[200]) );
  FA_7778 \FA_INST_0[0].FA_INST_1[200].FA_  ( .A(A[200]), .B(n713), .CI(C[200]), .S(S[200]), .CO(C[201]) );
  FA_7777 \FA_INST_0[0].FA_INST_1[201].FA_  ( .A(A[201]), .B(n714), .CI(C[201]), .S(S[201]), .CO(C[202]) );
  FA_7776 \FA_INST_0[0].FA_INST_1[202].FA_  ( .A(A[202]), .B(n715), .CI(C[202]), .S(S[202]), .CO(C[203]) );
  FA_7775 \FA_INST_0[0].FA_INST_1[203].FA_  ( .A(A[203]), .B(n716), .CI(C[203]), .S(S[203]), .CO(C[204]) );
  FA_7774 \FA_INST_0[0].FA_INST_1[204].FA_  ( .A(A[204]), .B(n717), .CI(C[204]), .S(S[204]), .CO(C[205]) );
  FA_7773 \FA_INST_0[0].FA_INST_1[205].FA_  ( .A(A[205]), .B(n718), .CI(C[205]), .S(S[205]), .CO(C[206]) );
  FA_7772 \FA_INST_0[0].FA_INST_1[206].FA_  ( .A(A[206]), .B(n719), .CI(C[206]), .S(S[206]), .CO(C[207]) );
  FA_7771 \FA_INST_0[0].FA_INST_1[207].FA_  ( .A(A[207]), .B(n720), .CI(C[207]), .S(S[207]), .CO(C[208]) );
  FA_7770 \FA_INST_0[0].FA_INST_1[208].FA_  ( .A(A[208]), .B(n721), .CI(C[208]), .S(S[208]), .CO(C[209]) );
  FA_7769 \FA_INST_0[0].FA_INST_1[209].FA_  ( .A(A[209]), .B(n722), .CI(C[209]), .S(S[209]), .CO(C[210]) );
  FA_7768 \FA_INST_0[0].FA_INST_1[210].FA_  ( .A(A[210]), .B(n723), .CI(C[210]), .S(S[210]), .CO(C[211]) );
  FA_7767 \FA_INST_0[0].FA_INST_1[211].FA_  ( .A(A[211]), .B(n724), .CI(C[211]), .S(S[211]), .CO(C[212]) );
  FA_7766 \FA_INST_0[0].FA_INST_1[212].FA_  ( .A(A[212]), .B(n725), .CI(C[212]), .S(S[212]), .CO(C[213]) );
  FA_7765 \FA_INST_0[0].FA_INST_1[213].FA_  ( .A(A[213]), .B(n726), .CI(C[213]), .S(S[213]), .CO(C[214]) );
  FA_7764 \FA_INST_0[0].FA_INST_1[214].FA_  ( .A(A[214]), .B(n727), .CI(C[214]), .S(S[214]), .CO(C[215]) );
  FA_7763 \FA_INST_0[0].FA_INST_1[215].FA_  ( .A(A[215]), .B(n728), .CI(C[215]), .S(S[215]), .CO(C[216]) );
  FA_7762 \FA_INST_0[0].FA_INST_1[216].FA_  ( .A(A[216]), .B(n729), .CI(C[216]), .S(S[216]), .CO(C[217]) );
  FA_7761 \FA_INST_0[0].FA_INST_1[217].FA_  ( .A(A[217]), .B(n730), .CI(C[217]), .S(S[217]), .CO(C[218]) );
  FA_7760 \FA_INST_0[0].FA_INST_1[218].FA_  ( .A(A[218]), .B(n731), .CI(C[218]), .S(S[218]), .CO(C[219]) );
  FA_7759 \FA_INST_0[0].FA_INST_1[219].FA_  ( .A(A[219]), .B(n732), .CI(C[219]), .S(S[219]), .CO(C[220]) );
  FA_7758 \FA_INST_0[0].FA_INST_1[220].FA_  ( .A(A[220]), .B(n733), .CI(C[220]), .S(S[220]), .CO(C[221]) );
  FA_7757 \FA_INST_0[0].FA_INST_1[221].FA_  ( .A(A[221]), .B(n734), .CI(C[221]), .S(S[221]), .CO(C[222]) );
  FA_7756 \FA_INST_0[0].FA_INST_1[222].FA_  ( .A(A[222]), .B(n735), .CI(C[222]), .S(S[222]), .CO(C[223]) );
  FA_7755 \FA_INST_0[0].FA_INST_1[223].FA_  ( .A(A[223]), .B(n736), .CI(C[223]), .S(S[223]), .CO(C[224]) );
  FA_7754 \FA_INST_0[0].FA_INST_1[224].FA_  ( .A(A[224]), .B(n737), .CI(C[224]), .S(S[224]), .CO(C[225]) );
  FA_7753 \FA_INST_0[0].FA_INST_1[225].FA_  ( .A(A[225]), .B(n738), .CI(C[225]), .S(S[225]), .CO(C[226]) );
  FA_7752 \FA_INST_0[0].FA_INST_1[226].FA_  ( .A(A[226]), .B(n739), .CI(C[226]), .S(S[226]), .CO(C[227]) );
  FA_7751 \FA_INST_0[0].FA_INST_1[227].FA_  ( .A(A[227]), .B(n740), .CI(C[227]), .S(S[227]), .CO(C[228]) );
  FA_7750 \FA_INST_0[0].FA_INST_1[228].FA_  ( .A(A[228]), .B(n741), .CI(C[228]), .S(S[228]), .CO(C[229]) );
  FA_7749 \FA_INST_0[0].FA_INST_1[229].FA_  ( .A(A[229]), .B(n742), .CI(C[229]), .S(S[229]), .CO(C[230]) );
  FA_7748 \FA_INST_0[0].FA_INST_1[230].FA_  ( .A(A[230]), .B(n743), .CI(C[230]), .S(S[230]), .CO(C[231]) );
  FA_7747 \FA_INST_0[0].FA_INST_1[231].FA_  ( .A(A[231]), .B(n744), .CI(C[231]), .S(S[231]), .CO(C[232]) );
  FA_7746 \FA_INST_0[0].FA_INST_1[232].FA_  ( .A(A[232]), .B(n745), .CI(C[232]), .S(S[232]), .CO(C[233]) );
  FA_7745 \FA_INST_0[0].FA_INST_1[233].FA_  ( .A(A[233]), .B(n746), .CI(C[233]), .S(S[233]), .CO(C[234]) );
  FA_7744 \FA_INST_0[0].FA_INST_1[234].FA_  ( .A(A[234]), .B(n747), .CI(C[234]), .S(S[234]), .CO(C[235]) );
  FA_7743 \FA_INST_0[0].FA_INST_1[235].FA_  ( .A(A[235]), .B(n748), .CI(C[235]), .S(S[235]), .CO(C[236]) );
  FA_7742 \FA_INST_0[0].FA_INST_1[236].FA_  ( .A(A[236]), .B(n749), .CI(C[236]), .S(S[236]), .CO(C[237]) );
  FA_7741 \FA_INST_0[0].FA_INST_1[237].FA_  ( .A(A[237]), .B(n750), .CI(C[237]), .S(S[237]), .CO(C[238]) );
  FA_7740 \FA_INST_0[0].FA_INST_1[238].FA_  ( .A(A[238]), .B(n751), .CI(C[238]), .S(S[238]), .CO(C[239]) );
  FA_7739 \FA_INST_0[0].FA_INST_1[239].FA_  ( .A(A[239]), .B(n752), .CI(C[239]), .S(S[239]), .CO(C[240]) );
  FA_7738 \FA_INST_0[0].FA_INST_1[240].FA_  ( .A(A[240]), .B(n753), .CI(C[240]), .S(S[240]), .CO(C[241]) );
  FA_7737 \FA_INST_0[0].FA_INST_1[241].FA_  ( .A(A[241]), .B(n754), .CI(C[241]), .S(S[241]), .CO(C[242]) );
  FA_7736 \FA_INST_0[0].FA_INST_1[242].FA_  ( .A(A[242]), .B(n755), .CI(C[242]), .S(S[242]), .CO(C[243]) );
  FA_7735 \FA_INST_0[0].FA_INST_1[243].FA_  ( .A(A[243]), .B(n756), .CI(C[243]), .S(S[243]), .CO(C[244]) );
  FA_7734 \FA_INST_0[0].FA_INST_1[244].FA_  ( .A(A[244]), .B(n757), .CI(C[244]), .S(S[244]), .CO(C[245]) );
  FA_7733 \FA_INST_0[0].FA_INST_1[245].FA_  ( .A(A[245]), .B(n758), .CI(C[245]), .S(S[245]), .CO(C[246]) );
  FA_7732 \FA_INST_0[0].FA_INST_1[246].FA_  ( .A(A[246]), .B(n759), .CI(C[246]), .S(S[246]), .CO(C[247]) );
  FA_7731 \FA_INST_0[0].FA_INST_1[247].FA_  ( .A(A[247]), .B(n760), .CI(C[247]), .S(S[247]), .CO(C[248]) );
  FA_7730 \FA_INST_0[0].FA_INST_1[248].FA_  ( .A(A[248]), .B(n761), .CI(C[248]), .S(S[248]), .CO(C[249]) );
  FA_7729 \FA_INST_0[0].FA_INST_1[249].FA_  ( .A(A[249]), .B(n762), .CI(C[249]), .S(S[249]), .CO(C[250]) );
  FA_7728 \FA_INST_0[0].FA_INST_1[250].FA_  ( .A(A[250]), .B(n763), .CI(C[250]), .S(S[250]), .CO(C[251]) );
  FA_7727 \FA_INST_0[0].FA_INST_1[251].FA_  ( .A(A[251]), .B(n764), .CI(C[251]), .S(S[251]), .CO(C[252]) );
  FA_7726 \FA_INST_0[0].FA_INST_1[252].FA_  ( .A(A[252]), .B(n765), .CI(C[252]), .S(S[252]), .CO(C[253]) );
  FA_7725 \FA_INST_0[0].FA_INST_1[253].FA_  ( .A(A[253]), .B(n766), .CI(C[253]), .S(S[253]), .CO(C[254]) );
  FA_7724 \FA_INST_0[0].FA_INST_1[254].FA_  ( .A(A[254]), .B(n767), .CI(C[254]), .S(S[254]), .CO(C[255]) );
  FA_7723 \FA_INST_0[0].FA_INST_1[255].FA_  ( .A(A[255]), .B(n768), .CI(C[255]), .S(S[255]), .CO(C[256]) );
  FA_7722 \FA_INST_0[0].FA_INST_1[256].FA_  ( .A(A[256]), .B(n769), .CI(C[256]), .S(S[256]), .CO(C[257]) );
  FA_7721 \FA_INST_0[0].FA_INST_1[257].FA_  ( .A(A[257]), .B(n770), .CI(C[257]), .S(S[257]), .CO(C[258]) );
  FA_7720 \FA_INST_0[0].FA_INST_1[258].FA_  ( .A(A[258]), .B(n771), .CI(C[258]), .S(S[258]), .CO(C[259]) );
  FA_7719 \FA_INST_0[0].FA_INST_1[259].FA_  ( .A(A[259]), .B(n772), .CI(C[259]), .S(S[259]), .CO(C[260]) );
  FA_7718 \FA_INST_0[0].FA_INST_1[260].FA_  ( .A(A[260]), .B(n773), .CI(C[260]), .S(S[260]), .CO(C[261]) );
  FA_7717 \FA_INST_0[0].FA_INST_1[261].FA_  ( .A(A[261]), .B(n774), .CI(C[261]), .S(S[261]), .CO(C[262]) );
  FA_7716 \FA_INST_0[0].FA_INST_1[262].FA_  ( .A(A[262]), .B(n775), .CI(C[262]), .S(S[262]), .CO(C[263]) );
  FA_7715 \FA_INST_0[0].FA_INST_1[263].FA_  ( .A(A[263]), .B(n776), .CI(C[263]), .S(S[263]), .CO(C[264]) );
  FA_7714 \FA_INST_0[0].FA_INST_1[264].FA_  ( .A(A[264]), .B(n777), .CI(C[264]), .S(S[264]), .CO(C[265]) );
  FA_7713 \FA_INST_0[0].FA_INST_1[265].FA_  ( .A(A[265]), .B(n778), .CI(C[265]), .S(S[265]), .CO(C[266]) );
  FA_7712 \FA_INST_0[0].FA_INST_1[266].FA_  ( .A(A[266]), .B(n779), .CI(C[266]), .S(S[266]), .CO(C[267]) );
  FA_7711 \FA_INST_0[0].FA_INST_1[267].FA_  ( .A(A[267]), .B(n780), .CI(C[267]), .S(S[267]), .CO(C[268]) );
  FA_7710 \FA_INST_0[0].FA_INST_1[268].FA_  ( .A(A[268]), .B(n781), .CI(C[268]), .S(S[268]), .CO(C[269]) );
  FA_7709 \FA_INST_0[0].FA_INST_1[269].FA_  ( .A(A[269]), .B(n782), .CI(C[269]), .S(S[269]), .CO(C[270]) );
  FA_7708 \FA_INST_0[0].FA_INST_1[270].FA_  ( .A(A[270]), .B(n783), .CI(C[270]), .S(S[270]), .CO(C[271]) );
  FA_7707 \FA_INST_0[0].FA_INST_1[271].FA_  ( .A(A[271]), .B(n784), .CI(C[271]), .S(S[271]), .CO(C[272]) );
  FA_7706 \FA_INST_0[0].FA_INST_1[272].FA_  ( .A(A[272]), .B(n785), .CI(C[272]), .S(S[272]), .CO(C[273]) );
  FA_7705 \FA_INST_0[0].FA_INST_1[273].FA_  ( .A(A[273]), .B(n786), .CI(C[273]), .S(S[273]), .CO(C[274]) );
  FA_7704 \FA_INST_0[0].FA_INST_1[274].FA_  ( .A(A[274]), .B(n787), .CI(C[274]), .S(S[274]), .CO(C[275]) );
  FA_7703 \FA_INST_0[0].FA_INST_1[275].FA_  ( .A(A[275]), .B(n788), .CI(C[275]), .S(S[275]), .CO(C[276]) );
  FA_7702 \FA_INST_0[0].FA_INST_1[276].FA_  ( .A(A[276]), .B(n789), .CI(C[276]), .S(S[276]), .CO(C[277]) );
  FA_7701 \FA_INST_0[0].FA_INST_1[277].FA_  ( .A(A[277]), .B(n790), .CI(C[277]), .S(S[277]), .CO(C[278]) );
  FA_7700 \FA_INST_0[0].FA_INST_1[278].FA_  ( .A(A[278]), .B(n791), .CI(C[278]), .S(S[278]), .CO(C[279]) );
  FA_7699 \FA_INST_0[0].FA_INST_1[279].FA_  ( .A(A[279]), .B(n792), .CI(C[279]), .S(S[279]), .CO(C[280]) );
  FA_7698 \FA_INST_0[0].FA_INST_1[280].FA_  ( .A(A[280]), .B(n793), .CI(C[280]), .S(S[280]), .CO(C[281]) );
  FA_7697 \FA_INST_0[0].FA_INST_1[281].FA_  ( .A(A[281]), .B(n794), .CI(C[281]), .S(S[281]), .CO(C[282]) );
  FA_7696 \FA_INST_0[0].FA_INST_1[282].FA_  ( .A(A[282]), .B(n795), .CI(C[282]), .S(S[282]), .CO(C[283]) );
  FA_7695 \FA_INST_0[0].FA_INST_1[283].FA_  ( .A(A[283]), .B(n796), .CI(C[283]), .S(S[283]), .CO(C[284]) );
  FA_7694 \FA_INST_0[0].FA_INST_1[284].FA_  ( .A(A[284]), .B(n797), .CI(C[284]), .S(S[284]), .CO(C[285]) );
  FA_7693 \FA_INST_0[0].FA_INST_1[285].FA_  ( .A(A[285]), .B(n798), .CI(C[285]), .S(S[285]), .CO(C[286]) );
  FA_7692 \FA_INST_0[0].FA_INST_1[286].FA_  ( .A(A[286]), .B(n799), .CI(C[286]), .S(S[286]), .CO(C[287]) );
  FA_7691 \FA_INST_0[0].FA_INST_1[287].FA_  ( .A(A[287]), .B(n800), .CI(C[287]), .S(S[287]), .CO(C[288]) );
  FA_7690 \FA_INST_0[0].FA_INST_1[288].FA_  ( .A(A[288]), .B(n801), .CI(C[288]), .S(S[288]), .CO(C[289]) );
  FA_7689 \FA_INST_0[0].FA_INST_1[289].FA_  ( .A(A[289]), .B(n802), .CI(C[289]), .S(S[289]), .CO(C[290]) );
  FA_7688 \FA_INST_0[0].FA_INST_1[290].FA_  ( .A(A[290]), .B(n803), .CI(C[290]), .S(S[290]), .CO(C[291]) );
  FA_7687 \FA_INST_0[0].FA_INST_1[291].FA_  ( .A(A[291]), .B(n804), .CI(C[291]), .S(S[291]), .CO(C[292]) );
  FA_7686 \FA_INST_0[0].FA_INST_1[292].FA_  ( .A(A[292]), .B(n805), .CI(C[292]), .S(S[292]), .CO(C[293]) );
  FA_7685 \FA_INST_0[0].FA_INST_1[293].FA_  ( .A(A[293]), .B(n806), .CI(C[293]), .S(S[293]), .CO(C[294]) );
  FA_7684 \FA_INST_0[0].FA_INST_1[294].FA_  ( .A(A[294]), .B(n807), .CI(C[294]), .S(S[294]), .CO(C[295]) );
  FA_7683 \FA_INST_0[0].FA_INST_1[295].FA_  ( .A(A[295]), .B(n808), .CI(C[295]), .S(S[295]), .CO(C[296]) );
  FA_7682 \FA_INST_0[0].FA_INST_1[296].FA_  ( .A(A[296]), .B(n809), .CI(C[296]), .S(S[296]), .CO(C[297]) );
  FA_7681 \FA_INST_0[0].FA_INST_1[297].FA_  ( .A(A[297]), .B(n810), .CI(C[297]), .S(S[297]), .CO(C[298]) );
  FA_7680 \FA_INST_0[0].FA_INST_1[298].FA_  ( .A(A[298]), .B(n811), .CI(C[298]), .S(S[298]), .CO(C[299]) );
  FA_7679 \FA_INST_0[0].FA_INST_1[299].FA_  ( .A(A[299]), .B(n812), .CI(C[299]), .S(S[299]), .CO(C[300]) );
  FA_7678 \FA_INST_0[0].FA_INST_1[300].FA_  ( .A(A[300]), .B(n813), .CI(C[300]), .S(S[300]), .CO(C[301]) );
  FA_7677 \FA_INST_0[0].FA_INST_1[301].FA_  ( .A(A[301]), .B(n814), .CI(C[301]), .S(S[301]), .CO(C[302]) );
  FA_7676 \FA_INST_0[0].FA_INST_1[302].FA_  ( .A(A[302]), .B(n815), .CI(C[302]), .S(S[302]), .CO(C[303]) );
  FA_7675 \FA_INST_0[0].FA_INST_1[303].FA_  ( .A(A[303]), .B(n816), .CI(C[303]), .S(S[303]), .CO(C[304]) );
  FA_7674 \FA_INST_0[0].FA_INST_1[304].FA_  ( .A(A[304]), .B(n817), .CI(C[304]), .S(S[304]), .CO(C[305]) );
  FA_7673 \FA_INST_0[0].FA_INST_1[305].FA_  ( .A(A[305]), .B(n818), .CI(C[305]), .S(S[305]), .CO(C[306]) );
  FA_7672 \FA_INST_0[0].FA_INST_1[306].FA_  ( .A(A[306]), .B(n819), .CI(C[306]), .S(S[306]), .CO(C[307]) );
  FA_7671 \FA_INST_0[0].FA_INST_1[307].FA_  ( .A(A[307]), .B(n820), .CI(C[307]), .S(S[307]), .CO(C[308]) );
  FA_7670 \FA_INST_0[0].FA_INST_1[308].FA_  ( .A(A[308]), .B(n821), .CI(C[308]), .S(S[308]), .CO(C[309]) );
  FA_7669 \FA_INST_0[0].FA_INST_1[309].FA_  ( .A(A[309]), .B(n822), .CI(C[309]), .S(S[309]), .CO(C[310]) );
  FA_7668 \FA_INST_0[0].FA_INST_1[310].FA_  ( .A(A[310]), .B(n823), .CI(C[310]), .S(S[310]), .CO(C[311]) );
  FA_7667 \FA_INST_0[0].FA_INST_1[311].FA_  ( .A(A[311]), .B(n824), .CI(C[311]), .S(S[311]), .CO(C[312]) );
  FA_7666 \FA_INST_0[0].FA_INST_1[312].FA_  ( .A(A[312]), .B(n825), .CI(C[312]), .S(S[312]), .CO(C[313]) );
  FA_7665 \FA_INST_0[0].FA_INST_1[313].FA_  ( .A(A[313]), .B(n826), .CI(C[313]), .S(S[313]), .CO(C[314]) );
  FA_7664 \FA_INST_0[0].FA_INST_1[314].FA_  ( .A(A[314]), .B(n827), .CI(C[314]), .S(S[314]), .CO(C[315]) );
  FA_7663 \FA_INST_0[0].FA_INST_1[315].FA_  ( .A(A[315]), .B(n828), .CI(C[315]), .S(S[315]), .CO(C[316]) );
  FA_7662 \FA_INST_0[0].FA_INST_1[316].FA_  ( .A(A[316]), .B(n829), .CI(C[316]), .S(S[316]), .CO(C[317]) );
  FA_7661 \FA_INST_0[0].FA_INST_1[317].FA_  ( .A(A[317]), .B(n830), .CI(C[317]), .S(S[317]), .CO(C[318]) );
  FA_7660 \FA_INST_0[0].FA_INST_1[318].FA_  ( .A(A[318]), .B(n831), .CI(C[318]), .S(S[318]), .CO(C[319]) );
  FA_7659 \FA_INST_0[0].FA_INST_1[319].FA_  ( .A(A[319]), .B(n832), .CI(C[319]), .S(S[319]), .CO(C[320]) );
  FA_7658 \FA_INST_0[0].FA_INST_1[320].FA_  ( .A(A[320]), .B(n833), .CI(C[320]), .S(S[320]), .CO(C[321]) );
  FA_7657 \FA_INST_0[0].FA_INST_1[321].FA_  ( .A(A[321]), .B(n834), .CI(C[321]), .S(S[321]), .CO(C[322]) );
  FA_7656 \FA_INST_0[0].FA_INST_1[322].FA_  ( .A(A[322]), .B(n835), .CI(C[322]), .S(S[322]), .CO(C[323]) );
  FA_7655 \FA_INST_0[0].FA_INST_1[323].FA_  ( .A(A[323]), .B(n836), .CI(C[323]), .S(S[323]), .CO(C[324]) );
  FA_7654 \FA_INST_0[0].FA_INST_1[324].FA_  ( .A(A[324]), .B(n837), .CI(C[324]), .S(S[324]), .CO(C[325]) );
  FA_7653 \FA_INST_0[0].FA_INST_1[325].FA_  ( .A(A[325]), .B(n838), .CI(C[325]), .S(S[325]), .CO(C[326]) );
  FA_7652 \FA_INST_0[0].FA_INST_1[326].FA_  ( .A(A[326]), .B(n839), .CI(C[326]), .S(S[326]), .CO(C[327]) );
  FA_7651 \FA_INST_0[0].FA_INST_1[327].FA_  ( .A(A[327]), .B(n840), .CI(C[327]), .S(S[327]), .CO(C[328]) );
  FA_7650 \FA_INST_0[0].FA_INST_1[328].FA_  ( .A(A[328]), .B(n841), .CI(C[328]), .S(S[328]), .CO(C[329]) );
  FA_7649 \FA_INST_0[0].FA_INST_1[329].FA_  ( .A(A[329]), .B(n842), .CI(C[329]), .S(S[329]), .CO(C[330]) );
  FA_7648 \FA_INST_0[0].FA_INST_1[330].FA_  ( .A(A[330]), .B(n843), .CI(C[330]), .S(S[330]), .CO(C[331]) );
  FA_7647 \FA_INST_0[0].FA_INST_1[331].FA_  ( .A(A[331]), .B(n844), .CI(C[331]), .S(S[331]), .CO(C[332]) );
  FA_7646 \FA_INST_0[0].FA_INST_1[332].FA_  ( .A(A[332]), .B(n845), .CI(C[332]), .S(S[332]), .CO(C[333]) );
  FA_7645 \FA_INST_0[0].FA_INST_1[333].FA_  ( .A(A[333]), .B(n846), .CI(C[333]), .S(S[333]), .CO(C[334]) );
  FA_7644 \FA_INST_0[0].FA_INST_1[334].FA_  ( .A(A[334]), .B(n847), .CI(C[334]), .S(S[334]), .CO(C[335]) );
  FA_7643 \FA_INST_0[0].FA_INST_1[335].FA_  ( .A(A[335]), .B(n848), .CI(C[335]), .S(S[335]), .CO(C[336]) );
  FA_7642 \FA_INST_0[0].FA_INST_1[336].FA_  ( .A(A[336]), .B(n849), .CI(C[336]), .S(S[336]), .CO(C[337]) );
  FA_7641 \FA_INST_0[0].FA_INST_1[337].FA_  ( .A(A[337]), .B(n850), .CI(C[337]), .S(S[337]), .CO(C[338]) );
  FA_7640 \FA_INST_0[0].FA_INST_1[338].FA_  ( .A(A[338]), .B(n851), .CI(C[338]), .S(S[338]), .CO(C[339]) );
  FA_7639 \FA_INST_0[0].FA_INST_1[339].FA_  ( .A(A[339]), .B(n852), .CI(C[339]), .S(S[339]), .CO(C[340]) );
  FA_7638 \FA_INST_0[0].FA_INST_1[340].FA_  ( .A(A[340]), .B(n853), .CI(C[340]), .S(S[340]), .CO(C[341]) );
  FA_7637 \FA_INST_0[0].FA_INST_1[341].FA_  ( .A(A[341]), .B(n854), .CI(C[341]), .S(S[341]), .CO(C[342]) );
  FA_7636 \FA_INST_0[0].FA_INST_1[342].FA_  ( .A(A[342]), .B(n855), .CI(C[342]), .S(S[342]), .CO(C[343]) );
  FA_7635 \FA_INST_0[0].FA_INST_1[343].FA_  ( .A(A[343]), .B(n856), .CI(C[343]), .S(S[343]), .CO(C[344]) );
  FA_7634 \FA_INST_0[0].FA_INST_1[344].FA_  ( .A(A[344]), .B(n857), .CI(C[344]), .S(S[344]), .CO(C[345]) );
  FA_7633 \FA_INST_0[0].FA_INST_1[345].FA_  ( .A(A[345]), .B(n858), .CI(C[345]), .S(S[345]), .CO(C[346]) );
  FA_7632 \FA_INST_0[0].FA_INST_1[346].FA_  ( .A(A[346]), .B(n859), .CI(C[346]), .S(S[346]), .CO(C[347]) );
  FA_7631 \FA_INST_0[0].FA_INST_1[347].FA_  ( .A(A[347]), .B(n860), .CI(C[347]), .S(S[347]), .CO(C[348]) );
  FA_7630 \FA_INST_0[0].FA_INST_1[348].FA_  ( .A(A[348]), .B(n861), .CI(C[348]), .S(S[348]), .CO(C[349]) );
  FA_7629 \FA_INST_0[0].FA_INST_1[349].FA_  ( .A(A[349]), .B(n862), .CI(C[349]), .S(S[349]), .CO(C[350]) );
  FA_7628 \FA_INST_0[0].FA_INST_1[350].FA_  ( .A(A[350]), .B(n863), .CI(C[350]), .S(S[350]), .CO(C[351]) );
  FA_7627 \FA_INST_0[0].FA_INST_1[351].FA_  ( .A(A[351]), .B(n864), .CI(C[351]), .S(S[351]), .CO(C[352]) );
  FA_7626 \FA_INST_0[0].FA_INST_1[352].FA_  ( .A(A[352]), .B(n865), .CI(C[352]), .S(S[352]), .CO(C[353]) );
  FA_7625 \FA_INST_0[0].FA_INST_1[353].FA_  ( .A(A[353]), .B(n866), .CI(C[353]), .S(S[353]), .CO(C[354]) );
  FA_7624 \FA_INST_0[0].FA_INST_1[354].FA_  ( .A(A[354]), .B(n867), .CI(C[354]), .S(S[354]), .CO(C[355]) );
  FA_7623 \FA_INST_0[0].FA_INST_1[355].FA_  ( .A(A[355]), .B(n868), .CI(C[355]), .S(S[355]), .CO(C[356]) );
  FA_7622 \FA_INST_0[0].FA_INST_1[356].FA_  ( .A(A[356]), .B(n869), .CI(C[356]), .S(S[356]), .CO(C[357]) );
  FA_7621 \FA_INST_0[0].FA_INST_1[357].FA_  ( .A(A[357]), .B(n870), .CI(C[357]), .S(S[357]), .CO(C[358]) );
  FA_7620 \FA_INST_0[0].FA_INST_1[358].FA_  ( .A(A[358]), .B(n871), .CI(C[358]), .S(S[358]), .CO(C[359]) );
  FA_7619 \FA_INST_0[0].FA_INST_1[359].FA_  ( .A(A[359]), .B(n872), .CI(C[359]), .S(S[359]), .CO(C[360]) );
  FA_7618 \FA_INST_0[0].FA_INST_1[360].FA_  ( .A(A[360]), .B(n873), .CI(C[360]), .S(S[360]), .CO(C[361]) );
  FA_7617 \FA_INST_0[0].FA_INST_1[361].FA_  ( .A(A[361]), .B(n874), .CI(C[361]), .S(S[361]), .CO(C[362]) );
  FA_7616 \FA_INST_0[0].FA_INST_1[362].FA_  ( .A(A[362]), .B(n875), .CI(C[362]), .S(S[362]), .CO(C[363]) );
  FA_7615 \FA_INST_0[0].FA_INST_1[363].FA_  ( .A(A[363]), .B(n876), .CI(C[363]), .S(S[363]), .CO(C[364]) );
  FA_7614 \FA_INST_0[0].FA_INST_1[364].FA_  ( .A(A[364]), .B(n877), .CI(C[364]), .S(S[364]), .CO(C[365]) );
  FA_7613 \FA_INST_0[0].FA_INST_1[365].FA_  ( .A(A[365]), .B(n878), .CI(C[365]), .S(S[365]), .CO(C[366]) );
  FA_7612 \FA_INST_0[0].FA_INST_1[366].FA_  ( .A(A[366]), .B(n879), .CI(C[366]), .S(S[366]), .CO(C[367]) );
  FA_7611 \FA_INST_0[0].FA_INST_1[367].FA_  ( .A(A[367]), .B(n880), .CI(C[367]), .S(S[367]), .CO(C[368]) );
  FA_7610 \FA_INST_0[0].FA_INST_1[368].FA_  ( .A(A[368]), .B(n881), .CI(C[368]), .S(S[368]), .CO(C[369]) );
  FA_7609 \FA_INST_0[0].FA_INST_1[369].FA_  ( .A(A[369]), .B(n882), .CI(C[369]), .S(S[369]), .CO(C[370]) );
  FA_7608 \FA_INST_0[0].FA_INST_1[370].FA_  ( .A(A[370]), .B(n883), .CI(C[370]), .S(S[370]), .CO(C[371]) );
  FA_7607 \FA_INST_0[0].FA_INST_1[371].FA_  ( .A(A[371]), .B(n884), .CI(C[371]), .S(S[371]), .CO(C[372]) );
  FA_7606 \FA_INST_0[0].FA_INST_1[372].FA_  ( .A(A[372]), .B(n885), .CI(C[372]), .S(S[372]), .CO(C[373]) );
  FA_7605 \FA_INST_0[0].FA_INST_1[373].FA_  ( .A(A[373]), .B(n886), .CI(C[373]), .S(S[373]), .CO(C[374]) );
  FA_7604 \FA_INST_0[0].FA_INST_1[374].FA_  ( .A(A[374]), .B(n887), .CI(C[374]), .S(S[374]), .CO(C[375]) );
  FA_7603 \FA_INST_0[0].FA_INST_1[375].FA_  ( .A(A[375]), .B(n888), .CI(C[375]), .S(S[375]), .CO(C[376]) );
  FA_7602 \FA_INST_0[0].FA_INST_1[376].FA_  ( .A(A[376]), .B(n889), .CI(C[376]), .S(S[376]), .CO(C[377]) );
  FA_7601 \FA_INST_0[0].FA_INST_1[377].FA_  ( .A(A[377]), .B(n890), .CI(C[377]), .S(S[377]), .CO(C[378]) );
  FA_7600 \FA_INST_0[0].FA_INST_1[378].FA_  ( .A(A[378]), .B(n891), .CI(C[378]), .S(S[378]), .CO(C[379]) );
  FA_7599 \FA_INST_0[0].FA_INST_1[379].FA_  ( .A(A[379]), .B(n892), .CI(C[379]), .S(S[379]), .CO(C[380]) );
  FA_7598 \FA_INST_0[0].FA_INST_1[380].FA_  ( .A(A[380]), .B(n893), .CI(C[380]), .S(S[380]), .CO(C[381]) );
  FA_7597 \FA_INST_0[0].FA_INST_1[381].FA_  ( .A(A[381]), .B(n894), .CI(C[381]), .S(S[381]), .CO(C[382]) );
  FA_7596 \FA_INST_0[0].FA_INST_1[382].FA_  ( .A(A[382]), .B(n895), .CI(C[382]), .S(S[382]), .CO(C[383]) );
  FA_7595 \FA_INST_0[0].FA_INST_1[383].FA_  ( .A(A[383]), .B(n896), .CI(C[383]), .S(S[383]), .CO(C[384]) );
  FA_7594 \FA_INST_0[0].FA_INST_1[384].FA_  ( .A(A[384]), .B(n897), .CI(C[384]), .S(S[384]), .CO(C[385]) );
  FA_7593 \FA_INST_0[0].FA_INST_1[385].FA_  ( .A(A[385]), .B(n898), .CI(C[385]), .S(S[385]), .CO(C[386]) );
  FA_7592 \FA_INST_0[0].FA_INST_1[386].FA_  ( .A(A[386]), .B(n899), .CI(C[386]), .S(S[386]), .CO(C[387]) );
  FA_7591 \FA_INST_0[0].FA_INST_1[387].FA_  ( .A(A[387]), .B(n900), .CI(C[387]), .S(S[387]), .CO(C[388]) );
  FA_7590 \FA_INST_0[0].FA_INST_1[388].FA_  ( .A(A[388]), .B(n901), .CI(C[388]), .S(S[388]), .CO(C[389]) );
  FA_7589 \FA_INST_0[0].FA_INST_1[389].FA_  ( .A(A[389]), .B(n902), .CI(C[389]), .S(S[389]), .CO(C[390]) );
  FA_7588 \FA_INST_0[0].FA_INST_1[390].FA_  ( .A(A[390]), .B(n903), .CI(C[390]), .S(S[390]), .CO(C[391]) );
  FA_7587 \FA_INST_0[0].FA_INST_1[391].FA_  ( .A(A[391]), .B(n904), .CI(C[391]), .S(S[391]), .CO(C[392]) );
  FA_7586 \FA_INST_0[0].FA_INST_1[392].FA_  ( .A(A[392]), .B(n905), .CI(C[392]), .S(S[392]), .CO(C[393]) );
  FA_7585 \FA_INST_0[0].FA_INST_1[393].FA_  ( .A(A[393]), .B(n906), .CI(C[393]), .S(S[393]), .CO(C[394]) );
  FA_7584 \FA_INST_0[0].FA_INST_1[394].FA_  ( .A(A[394]), .B(n907), .CI(C[394]), .S(S[394]), .CO(C[395]) );
  FA_7583 \FA_INST_0[0].FA_INST_1[395].FA_  ( .A(A[395]), .B(n908), .CI(C[395]), .S(S[395]), .CO(C[396]) );
  FA_7582 \FA_INST_0[0].FA_INST_1[396].FA_  ( .A(A[396]), .B(n909), .CI(C[396]), .S(S[396]), .CO(C[397]) );
  FA_7581 \FA_INST_0[0].FA_INST_1[397].FA_  ( .A(A[397]), .B(n910), .CI(C[397]), .S(S[397]), .CO(C[398]) );
  FA_7580 \FA_INST_0[0].FA_INST_1[398].FA_  ( .A(A[398]), .B(n911), .CI(C[398]), .S(S[398]), .CO(C[399]) );
  FA_7579 \FA_INST_0[0].FA_INST_1[399].FA_  ( .A(A[399]), .B(n912), .CI(C[399]), .S(S[399]), .CO(C[400]) );
  FA_7578 \FA_INST_0[0].FA_INST_1[400].FA_  ( .A(A[400]), .B(n913), .CI(C[400]), .S(S[400]), .CO(C[401]) );
  FA_7577 \FA_INST_0[0].FA_INST_1[401].FA_  ( .A(A[401]), .B(n914), .CI(C[401]), .S(S[401]), .CO(C[402]) );
  FA_7576 \FA_INST_0[0].FA_INST_1[402].FA_  ( .A(A[402]), .B(n915), .CI(C[402]), .S(S[402]), .CO(C[403]) );
  FA_7575 \FA_INST_0[0].FA_INST_1[403].FA_  ( .A(A[403]), .B(n916), .CI(C[403]), .S(S[403]), .CO(C[404]) );
  FA_7574 \FA_INST_0[0].FA_INST_1[404].FA_  ( .A(A[404]), .B(n917), .CI(C[404]), .S(S[404]), .CO(C[405]) );
  FA_7573 \FA_INST_0[0].FA_INST_1[405].FA_  ( .A(A[405]), .B(n918), .CI(C[405]), .S(S[405]), .CO(C[406]) );
  FA_7572 \FA_INST_0[0].FA_INST_1[406].FA_  ( .A(A[406]), .B(n919), .CI(C[406]), .S(S[406]), .CO(C[407]) );
  FA_7571 \FA_INST_0[0].FA_INST_1[407].FA_  ( .A(A[407]), .B(n920), .CI(C[407]), .S(S[407]), .CO(C[408]) );
  FA_7570 \FA_INST_0[0].FA_INST_1[408].FA_  ( .A(A[408]), .B(n921), .CI(C[408]), .S(S[408]), .CO(C[409]) );
  FA_7569 \FA_INST_0[0].FA_INST_1[409].FA_  ( .A(A[409]), .B(n922), .CI(C[409]), .S(S[409]), .CO(C[410]) );
  FA_7568 \FA_INST_0[0].FA_INST_1[410].FA_  ( .A(A[410]), .B(n923), .CI(C[410]), .S(S[410]), .CO(C[411]) );
  FA_7567 \FA_INST_0[0].FA_INST_1[411].FA_  ( .A(A[411]), .B(n924), .CI(C[411]), .S(S[411]), .CO(C[412]) );
  FA_7566 \FA_INST_0[0].FA_INST_1[412].FA_  ( .A(A[412]), .B(n925), .CI(C[412]), .S(S[412]), .CO(C[413]) );
  FA_7565 \FA_INST_0[0].FA_INST_1[413].FA_  ( .A(A[413]), .B(n926), .CI(C[413]), .S(S[413]), .CO(C[414]) );
  FA_7564 \FA_INST_0[0].FA_INST_1[414].FA_  ( .A(A[414]), .B(n927), .CI(C[414]), .S(S[414]), .CO(C[415]) );
  FA_7563 \FA_INST_0[0].FA_INST_1[415].FA_  ( .A(A[415]), .B(n928), .CI(C[415]), .S(S[415]), .CO(C[416]) );
  FA_7562 \FA_INST_0[0].FA_INST_1[416].FA_  ( .A(A[416]), .B(n929), .CI(C[416]), .S(S[416]), .CO(C[417]) );
  FA_7561 \FA_INST_0[0].FA_INST_1[417].FA_  ( .A(A[417]), .B(n930), .CI(C[417]), .S(S[417]), .CO(C[418]) );
  FA_7560 \FA_INST_0[0].FA_INST_1[418].FA_  ( .A(A[418]), .B(n931), .CI(C[418]), .S(S[418]), .CO(C[419]) );
  FA_7559 \FA_INST_0[0].FA_INST_1[419].FA_  ( .A(A[419]), .B(n932), .CI(C[419]), .S(S[419]), .CO(C[420]) );
  FA_7558 \FA_INST_0[0].FA_INST_1[420].FA_  ( .A(A[420]), .B(n933), .CI(C[420]), .S(S[420]), .CO(C[421]) );
  FA_7557 \FA_INST_0[0].FA_INST_1[421].FA_  ( .A(A[421]), .B(n934), .CI(C[421]), .S(S[421]), .CO(C[422]) );
  FA_7556 \FA_INST_0[0].FA_INST_1[422].FA_  ( .A(A[422]), .B(n935), .CI(C[422]), .S(S[422]), .CO(C[423]) );
  FA_7555 \FA_INST_0[0].FA_INST_1[423].FA_  ( .A(A[423]), .B(n936), .CI(C[423]), .S(S[423]), .CO(C[424]) );
  FA_7554 \FA_INST_0[0].FA_INST_1[424].FA_  ( .A(A[424]), .B(n937), .CI(C[424]), .S(S[424]), .CO(C[425]) );
  FA_7553 \FA_INST_0[0].FA_INST_1[425].FA_  ( .A(A[425]), .B(n938), .CI(C[425]), .S(S[425]), .CO(C[426]) );
  FA_7552 \FA_INST_0[0].FA_INST_1[426].FA_  ( .A(A[426]), .B(n939), .CI(C[426]), .S(S[426]), .CO(C[427]) );
  FA_7551 \FA_INST_0[0].FA_INST_1[427].FA_  ( .A(A[427]), .B(n940), .CI(C[427]), .S(S[427]), .CO(C[428]) );
  FA_7550 \FA_INST_0[0].FA_INST_1[428].FA_  ( .A(A[428]), .B(n941), .CI(C[428]), .S(S[428]), .CO(C[429]) );
  FA_7549 \FA_INST_0[0].FA_INST_1[429].FA_  ( .A(A[429]), .B(n942), .CI(C[429]), .S(S[429]), .CO(C[430]) );
  FA_7548 \FA_INST_0[0].FA_INST_1[430].FA_  ( .A(A[430]), .B(n943), .CI(C[430]), .S(S[430]), .CO(C[431]) );
  FA_7547 \FA_INST_0[0].FA_INST_1[431].FA_  ( .A(A[431]), .B(n944), .CI(C[431]), .S(S[431]), .CO(C[432]) );
  FA_7546 \FA_INST_0[0].FA_INST_1[432].FA_  ( .A(A[432]), .B(n945), .CI(C[432]), .S(S[432]), .CO(C[433]) );
  FA_7545 \FA_INST_0[0].FA_INST_1[433].FA_  ( .A(A[433]), .B(n946), .CI(C[433]), .S(S[433]), .CO(C[434]) );
  FA_7544 \FA_INST_0[0].FA_INST_1[434].FA_  ( .A(A[434]), .B(n947), .CI(C[434]), .S(S[434]), .CO(C[435]) );
  FA_7543 \FA_INST_0[0].FA_INST_1[435].FA_  ( .A(A[435]), .B(n948), .CI(C[435]), .S(S[435]), .CO(C[436]) );
  FA_7542 \FA_INST_0[0].FA_INST_1[436].FA_  ( .A(A[436]), .B(n949), .CI(C[436]), .S(S[436]), .CO(C[437]) );
  FA_7541 \FA_INST_0[0].FA_INST_1[437].FA_  ( .A(A[437]), .B(n950), .CI(C[437]), .S(S[437]), .CO(C[438]) );
  FA_7540 \FA_INST_0[0].FA_INST_1[438].FA_  ( .A(A[438]), .B(n951), .CI(C[438]), .S(S[438]), .CO(C[439]) );
  FA_7539 \FA_INST_0[0].FA_INST_1[439].FA_  ( .A(A[439]), .B(n952), .CI(C[439]), .S(S[439]), .CO(C[440]) );
  FA_7538 \FA_INST_0[0].FA_INST_1[440].FA_  ( .A(A[440]), .B(n953), .CI(C[440]), .S(S[440]), .CO(C[441]) );
  FA_7537 \FA_INST_0[0].FA_INST_1[441].FA_  ( .A(A[441]), .B(n954), .CI(C[441]), .S(S[441]), .CO(C[442]) );
  FA_7536 \FA_INST_0[0].FA_INST_1[442].FA_  ( .A(A[442]), .B(n955), .CI(C[442]), .S(S[442]), .CO(C[443]) );
  FA_7535 \FA_INST_0[0].FA_INST_1[443].FA_  ( .A(A[443]), .B(n956), .CI(C[443]), .S(S[443]), .CO(C[444]) );
  FA_7534 \FA_INST_0[0].FA_INST_1[444].FA_  ( .A(A[444]), .B(n957), .CI(C[444]), .S(S[444]), .CO(C[445]) );
  FA_7533 \FA_INST_0[0].FA_INST_1[445].FA_  ( .A(A[445]), .B(n958), .CI(C[445]), .S(S[445]), .CO(C[446]) );
  FA_7532 \FA_INST_0[0].FA_INST_1[446].FA_  ( .A(A[446]), .B(n959), .CI(C[446]), .S(S[446]), .CO(C[447]) );
  FA_7531 \FA_INST_0[0].FA_INST_1[447].FA_  ( .A(A[447]), .B(n960), .CI(C[447]), .S(S[447]), .CO(C[448]) );
  FA_7530 \FA_INST_0[0].FA_INST_1[448].FA_  ( .A(A[448]), .B(n961), .CI(C[448]), .S(S[448]), .CO(C[449]) );
  FA_7529 \FA_INST_0[0].FA_INST_1[449].FA_  ( .A(A[449]), .B(n962), .CI(C[449]), .S(S[449]), .CO(C[450]) );
  FA_7528 \FA_INST_0[0].FA_INST_1[450].FA_  ( .A(A[450]), .B(n963), .CI(C[450]), .S(S[450]), .CO(C[451]) );
  FA_7527 \FA_INST_0[0].FA_INST_1[451].FA_  ( .A(A[451]), .B(n964), .CI(C[451]), .S(S[451]), .CO(C[452]) );
  FA_7526 \FA_INST_0[0].FA_INST_1[452].FA_  ( .A(A[452]), .B(n965), .CI(C[452]), .S(S[452]), .CO(C[453]) );
  FA_7525 \FA_INST_0[0].FA_INST_1[453].FA_  ( .A(A[453]), .B(n966), .CI(C[453]), .S(S[453]), .CO(C[454]) );
  FA_7524 \FA_INST_0[0].FA_INST_1[454].FA_  ( .A(A[454]), .B(n967), .CI(C[454]), .S(S[454]), .CO(C[455]) );
  FA_7523 \FA_INST_0[0].FA_INST_1[455].FA_  ( .A(A[455]), .B(n968), .CI(C[455]), .S(S[455]), .CO(C[456]) );
  FA_7522 \FA_INST_0[0].FA_INST_1[456].FA_  ( .A(A[456]), .B(n969), .CI(C[456]), .S(S[456]), .CO(C[457]) );
  FA_7521 \FA_INST_0[0].FA_INST_1[457].FA_  ( .A(A[457]), .B(n970), .CI(C[457]), .S(S[457]), .CO(C[458]) );
  FA_7520 \FA_INST_0[0].FA_INST_1[458].FA_  ( .A(A[458]), .B(n971), .CI(C[458]), .S(S[458]), .CO(C[459]) );
  FA_7519 \FA_INST_0[0].FA_INST_1[459].FA_  ( .A(A[459]), .B(n972), .CI(C[459]), .S(S[459]), .CO(C[460]) );
  FA_7518 \FA_INST_0[0].FA_INST_1[460].FA_  ( .A(A[460]), .B(n973), .CI(C[460]), .S(S[460]), .CO(C[461]) );
  FA_7517 \FA_INST_0[0].FA_INST_1[461].FA_  ( .A(A[461]), .B(n974), .CI(C[461]), .S(S[461]), .CO(C[462]) );
  FA_7516 \FA_INST_0[0].FA_INST_1[462].FA_  ( .A(A[462]), .B(n975), .CI(C[462]), .S(S[462]), .CO(C[463]) );
  FA_7515 \FA_INST_0[0].FA_INST_1[463].FA_  ( .A(A[463]), .B(n976), .CI(C[463]), .S(S[463]), .CO(C[464]) );
  FA_7514 \FA_INST_0[0].FA_INST_1[464].FA_  ( .A(A[464]), .B(n977), .CI(C[464]), .S(S[464]), .CO(C[465]) );
  FA_7513 \FA_INST_0[0].FA_INST_1[465].FA_  ( .A(A[465]), .B(n978), .CI(C[465]), .S(S[465]), .CO(C[466]) );
  FA_7512 \FA_INST_0[0].FA_INST_1[466].FA_  ( .A(A[466]), .B(n979), .CI(C[466]), .S(S[466]), .CO(C[467]) );
  FA_7511 \FA_INST_0[0].FA_INST_1[467].FA_  ( .A(A[467]), .B(n980), .CI(C[467]), .S(S[467]), .CO(C[468]) );
  FA_7510 \FA_INST_0[0].FA_INST_1[468].FA_  ( .A(A[468]), .B(n981), .CI(C[468]), .S(S[468]), .CO(C[469]) );
  FA_7509 \FA_INST_0[0].FA_INST_1[469].FA_  ( .A(A[469]), .B(n982), .CI(C[469]), .S(S[469]), .CO(C[470]) );
  FA_7508 \FA_INST_0[0].FA_INST_1[470].FA_  ( .A(A[470]), .B(n983), .CI(C[470]), .S(S[470]), .CO(C[471]) );
  FA_7507 \FA_INST_0[0].FA_INST_1[471].FA_  ( .A(A[471]), .B(n984), .CI(C[471]), .S(S[471]), .CO(C[472]) );
  FA_7506 \FA_INST_0[0].FA_INST_1[472].FA_  ( .A(A[472]), .B(n985), .CI(C[472]), .S(S[472]), .CO(C[473]) );
  FA_7505 \FA_INST_0[0].FA_INST_1[473].FA_  ( .A(A[473]), .B(n986), .CI(C[473]), .S(S[473]), .CO(C[474]) );
  FA_7504 \FA_INST_0[0].FA_INST_1[474].FA_  ( .A(A[474]), .B(n987), .CI(C[474]), .S(S[474]), .CO(C[475]) );
  FA_7503 \FA_INST_0[0].FA_INST_1[475].FA_  ( .A(A[475]), .B(n988), .CI(C[475]), .S(S[475]), .CO(C[476]) );
  FA_7502 \FA_INST_0[0].FA_INST_1[476].FA_  ( .A(A[476]), .B(n989), .CI(C[476]), .S(S[476]), .CO(C[477]) );
  FA_7501 \FA_INST_0[0].FA_INST_1[477].FA_  ( .A(A[477]), .B(n990), .CI(C[477]), .S(S[477]), .CO(C[478]) );
  FA_7500 \FA_INST_0[0].FA_INST_1[478].FA_  ( .A(A[478]), .B(n991), .CI(C[478]), .S(S[478]), .CO(C[479]) );
  FA_7499 \FA_INST_0[0].FA_INST_1[479].FA_  ( .A(A[479]), .B(n992), .CI(C[479]), .S(S[479]), .CO(C[480]) );
  FA_7498 \FA_INST_0[0].FA_INST_1[480].FA_  ( .A(A[480]), .B(n993), .CI(C[480]), .S(S[480]), .CO(C[481]) );
  FA_7497 \FA_INST_0[0].FA_INST_1[481].FA_  ( .A(A[481]), .B(n994), .CI(C[481]), .S(S[481]), .CO(C[482]) );
  FA_7496 \FA_INST_0[0].FA_INST_1[482].FA_  ( .A(A[482]), .B(n995), .CI(C[482]), .S(S[482]), .CO(C[483]) );
  FA_7495 \FA_INST_0[0].FA_INST_1[483].FA_  ( .A(A[483]), .B(n996), .CI(C[483]), .S(S[483]), .CO(C[484]) );
  FA_7494 \FA_INST_0[0].FA_INST_1[484].FA_  ( .A(A[484]), .B(n997), .CI(C[484]), .S(S[484]), .CO(C[485]) );
  FA_7493 \FA_INST_0[0].FA_INST_1[485].FA_  ( .A(A[485]), .B(n998), .CI(C[485]), .S(S[485]), .CO(C[486]) );
  FA_7492 \FA_INST_0[0].FA_INST_1[486].FA_  ( .A(A[486]), .B(n999), .CI(C[486]), .S(S[486]), .CO(C[487]) );
  FA_7491 \FA_INST_0[0].FA_INST_1[487].FA_  ( .A(A[487]), .B(n1000), .CI(
        C[487]), .S(S[487]), .CO(C[488]) );
  FA_7490 \FA_INST_0[0].FA_INST_1[488].FA_  ( .A(A[488]), .B(n1001), .CI(
        C[488]), .S(S[488]), .CO(C[489]) );
  FA_7489 \FA_INST_0[0].FA_INST_1[489].FA_  ( .A(A[489]), .B(n1002), .CI(
        C[489]), .S(S[489]), .CO(C[490]) );
  FA_7488 \FA_INST_0[0].FA_INST_1[490].FA_  ( .A(A[490]), .B(n1003), .CI(
        C[490]), .S(S[490]), .CO(C[491]) );
  FA_7487 \FA_INST_0[0].FA_INST_1[491].FA_  ( .A(A[491]), .B(n1004), .CI(
        C[491]), .S(S[491]), .CO(C[492]) );
  FA_7486 \FA_INST_0[0].FA_INST_1[492].FA_  ( .A(A[492]), .B(n1005), .CI(
        C[492]), .S(S[492]), .CO(C[493]) );
  FA_7485 \FA_INST_0[0].FA_INST_1[493].FA_  ( .A(A[493]), .B(n1006), .CI(
        C[493]), .S(S[493]), .CO(C[494]) );
  FA_7484 \FA_INST_0[0].FA_INST_1[494].FA_  ( .A(A[494]), .B(n1007), .CI(
        C[494]), .S(S[494]), .CO(C[495]) );
  FA_7483 \FA_INST_0[0].FA_INST_1[495].FA_  ( .A(A[495]), .B(n1008), .CI(
        C[495]), .S(S[495]), .CO(C[496]) );
  FA_7482 \FA_INST_0[0].FA_INST_1[496].FA_  ( .A(A[496]), .B(n1009), .CI(
        C[496]), .S(S[496]), .CO(C[497]) );
  FA_7481 \FA_INST_0[0].FA_INST_1[497].FA_  ( .A(A[497]), .B(n1010), .CI(
        C[497]), .S(S[497]), .CO(C[498]) );
  FA_7480 \FA_INST_0[0].FA_INST_1[498].FA_  ( .A(A[498]), .B(n1011), .CI(
        C[498]), .S(S[498]), .CO(C[499]) );
  FA_7479 \FA_INST_0[0].FA_INST_1[499].FA_  ( .A(A[499]), .B(n1012), .CI(
        C[499]), .S(S[499]), .CO(C[500]) );
  FA_7478 \FA_INST_0[0].FA_INST_1[500].FA_  ( .A(A[500]), .B(n1013), .CI(
        C[500]), .S(S[500]), .CO(C[501]) );
  FA_7477 \FA_INST_0[0].FA_INST_1[501].FA_  ( .A(A[501]), .B(n1014), .CI(
        C[501]), .S(S[501]), .CO(C[502]) );
  FA_7476 \FA_INST_0[0].FA_INST_1[502].FA_  ( .A(A[502]), .B(n1015), .CI(
        C[502]), .S(S[502]), .CO(C[503]) );
  FA_7475 \FA_INST_0[0].FA_INST_1[503].FA_  ( .A(A[503]), .B(n1016), .CI(
        C[503]), .S(S[503]), .CO(C[504]) );
  FA_7474 \FA_INST_0[0].FA_INST_1[504].FA_  ( .A(A[504]), .B(n1017), .CI(
        C[504]), .S(S[504]), .CO(C[505]) );
  FA_7473 \FA_INST_0[0].FA_INST_1[505].FA_  ( .A(A[505]), .B(n1018), .CI(
        C[505]), .S(S[505]), .CO(C[506]) );
  FA_7472 \FA_INST_0[0].FA_INST_1[506].FA_  ( .A(A[506]), .B(n1019), .CI(
        C[506]), .S(S[506]), .CO(C[507]) );
  FA_7471 \FA_INST_0[0].FA_INST_1[507].FA_  ( .A(A[507]), .B(n1020), .CI(
        C[507]), .S(S[507]), .CO(C[508]) );
  FA_7470 \FA_INST_0[0].FA_INST_1[508].FA_  ( .A(A[508]), .B(n1021), .CI(
        C[508]), .S(S[508]), .CO(C[509]) );
  FA_7469 \FA_INST_0[0].FA_INST_1[509].FA_  ( .A(A[509]), .B(n1022), .CI(
        C[509]), .S(S[509]), .CO(C[510]) );
  FA_7468 \FA_INST_0[0].FA_INST_1[510].FA_  ( .A(A[510]), .B(n1023), .CI(
        C[510]), .S(S[510]), .CO(C[511]) );
  FA_7467 \FA_INST_0[0].FA_INST_1[511].FA_  ( .A(A[511]), .B(n1024), .CI(
        C[511]), .S(S[511]), .CO(C[512]) );
  FA_7466 \FA_INST_1[512].FA_  ( .A(A[512]), .B(1'b1), .CI(C[512]), .S(S[512]), 
        .CO(C[513]) );
  FA_7465 \FA_INST_1[513].FA_  ( .A(A[513]), .B(1'b1), .CI(C[513]), .S(S[513])
         );
  IV U2 ( .A(B[415]), .Z(n928) );
  IV U3 ( .A(B[416]), .Z(n929) );
  IV U4 ( .A(B[417]), .Z(n930) );
  IV U5 ( .A(B[418]), .Z(n931) );
  IV U6 ( .A(B[419]), .Z(n932) );
  IV U7 ( .A(B[420]), .Z(n933) );
  IV U8 ( .A(B[421]), .Z(n934) );
  IV U9 ( .A(B[422]), .Z(n935) );
  IV U10 ( .A(B[423]), .Z(n936) );
  IV U11 ( .A(B[424]), .Z(n937) );
  IV U12 ( .A(B[505]), .Z(n1018) );
  IV U13 ( .A(B[425]), .Z(n938) );
  IV U14 ( .A(B[426]), .Z(n939) );
  IV U15 ( .A(B[427]), .Z(n940) );
  IV U16 ( .A(B[428]), .Z(n941) );
  IV U17 ( .A(B[429]), .Z(n942) );
  IV U18 ( .A(B[430]), .Z(n943) );
  IV U19 ( .A(B[431]), .Z(n944) );
  IV U20 ( .A(B[432]), .Z(n945) );
  IV U21 ( .A(B[433]), .Z(n946) );
  IV U22 ( .A(B[434]), .Z(n947) );
  IV U23 ( .A(B[506]), .Z(n1019) );
  IV U24 ( .A(B[435]), .Z(n948) );
  IV U25 ( .A(B[436]), .Z(n949) );
  IV U26 ( .A(B[437]), .Z(n950) );
  IV U27 ( .A(B[438]), .Z(n951) );
  IV U28 ( .A(B[439]), .Z(n952) );
  IV U29 ( .A(B[440]), .Z(n953) );
  IV U30 ( .A(B[441]), .Z(n954) );
  IV U31 ( .A(B[442]), .Z(n955) );
  IV U32 ( .A(B[443]), .Z(n956) );
  IV U33 ( .A(B[444]), .Z(n957) );
  IV U34 ( .A(B[507]), .Z(n1020) );
  IV U35 ( .A(B[445]), .Z(n958) );
  IV U36 ( .A(B[446]), .Z(n959) );
  IV U37 ( .A(B[447]), .Z(n960) );
  IV U38 ( .A(B[448]), .Z(n961) );
  IV U39 ( .A(B[449]), .Z(n962) );
  IV U40 ( .A(B[450]), .Z(n963) );
  IV U41 ( .A(B[451]), .Z(n964) );
  IV U42 ( .A(B[452]), .Z(n965) );
  IV U43 ( .A(B[453]), .Z(n966) );
  IV U44 ( .A(B[454]), .Z(n967) );
  IV U45 ( .A(B[508]), .Z(n1021) );
  IV U46 ( .A(B[455]), .Z(n968) );
  IV U47 ( .A(B[456]), .Z(n969) );
  IV U48 ( .A(B[457]), .Z(n970) );
  IV U49 ( .A(B[458]), .Z(n971) );
  IV U50 ( .A(B[459]), .Z(n972) );
  IV U51 ( .A(B[460]), .Z(n973) );
  IV U52 ( .A(B[461]), .Z(n974) );
  IV U53 ( .A(B[462]), .Z(n975) );
  IV U54 ( .A(B[0]), .Z(n2) );
  IV U55 ( .A(B[1]), .Z(n514) );
  IV U56 ( .A(B[2]), .Z(n515) );
  IV U57 ( .A(B[3]), .Z(n516) );
  IV U58 ( .A(B[4]), .Z(n517) );
  IV U59 ( .A(B[463]), .Z(n976) );
  IV U60 ( .A(B[5]), .Z(n518) );
  IV U61 ( .A(B[6]), .Z(n519) );
  IV U62 ( .A(B[7]), .Z(n520) );
  IV U63 ( .A(B[8]), .Z(n521) );
  IV U64 ( .A(B[9]), .Z(n522) );
  IV U65 ( .A(B[10]), .Z(n523) );
  IV U66 ( .A(B[11]), .Z(n524) );
  IV U67 ( .A(B[12]), .Z(n525) );
  IV U68 ( .A(B[13]), .Z(n526) );
  IV U69 ( .A(B[14]), .Z(n527) );
  IV U70 ( .A(B[464]), .Z(n977) );
  IV U71 ( .A(B[509]), .Z(n1022) );
  IV U72 ( .A(B[15]), .Z(n528) );
  IV U73 ( .A(B[16]), .Z(n529) );
  IV U74 ( .A(B[17]), .Z(n530) );
  IV U75 ( .A(B[18]), .Z(n531) );
  IV U76 ( .A(B[19]), .Z(n532) );
  IV U77 ( .A(B[20]), .Z(n533) );
  IV U78 ( .A(B[21]), .Z(n534) );
  IV U79 ( .A(B[22]), .Z(n535) );
  IV U80 ( .A(B[23]), .Z(n536) );
  IV U81 ( .A(B[24]), .Z(n537) );
  IV U82 ( .A(B[465]), .Z(n978) );
  IV U83 ( .A(B[25]), .Z(n538) );
  IV U84 ( .A(B[26]), .Z(n539) );
  IV U85 ( .A(B[27]), .Z(n540) );
  IV U86 ( .A(B[28]), .Z(n541) );
  IV U87 ( .A(B[29]), .Z(n542) );
  IV U88 ( .A(B[30]), .Z(n543) );
  IV U89 ( .A(B[31]), .Z(n544) );
  IV U90 ( .A(B[32]), .Z(n545) );
  IV U91 ( .A(B[33]), .Z(n546) );
  IV U92 ( .A(B[34]), .Z(n547) );
  IV U93 ( .A(B[466]), .Z(n979) );
  IV U94 ( .A(B[35]), .Z(n548) );
  IV U95 ( .A(B[36]), .Z(n549) );
  IV U96 ( .A(B[37]), .Z(n550) );
  IV U97 ( .A(B[38]), .Z(n551) );
  IV U98 ( .A(B[39]), .Z(n552) );
  IV U99 ( .A(B[40]), .Z(n553) );
  IV U100 ( .A(B[41]), .Z(n554) );
  IV U101 ( .A(B[42]), .Z(n555) );
  IV U102 ( .A(B[43]), .Z(n556) );
  IV U103 ( .A(B[44]), .Z(n557) );
  IV U104 ( .A(B[467]), .Z(n980) );
  IV U105 ( .A(B[45]), .Z(n558) );
  IV U106 ( .A(B[46]), .Z(n559) );
  IV U107 ( .A(B[47]), .Z(n560) );
  IV U108 ( .A(B[48]), .Z(n561) );
  IV U109 ( .A(B[49]), .Z(n562) );
  IV U110 ( .A(B[50]), .Z(n563) );
  IV U111 ( .A(B[51]), .Z(n564) );
  IV U112 ( .A(B[52]), .Z(n565) );
  IV U113 ( .A(B[53]), .Z(n566) );
  IV U114 ( .A(B[54]), .Z(n567) );
  IV U115 ( .A(B[468]), .Z(n981) );
  IV U116 ( .A(B[55]), .Z(n568) );
  IV U117 ( .A(B[56]), .Z(n569) );
  IV U118 ( .A(B[57]), .Z(n570) );
  IV U119 ( .A(B[58]), .Z(n571) );
  IV U120 ( .A(B[59]), .Z(n572) );
  IV U121 ( .A(B[60]), .Z(n573) );
  IV U122 ( .A(B[61]), .Z(n574) );
  IV U123 ( .A(B[62]), .Z(n575) );
  IV U124 ( .A(B[63]), .Z(n576) );
  IV U125 ( .A(B[64]), .Z(n577) );
  IV U126 ( .A(B[469]), .Z(n982) );
  IV U127 ( .A(B[65]), .Z(n578) );
  IV U128 ( .A(B[66]), .Z(n579) );
  IV U129 ( .A(B[67]), .Z(n580) );
  IV U130 ( .A(B[68]), .Z(n581) );
  IV U131 ( .A(B[69]), .Z(n582) );
  IV U132 ( .A(B[70]), .Z(n583) );
  IV U133 ( .A(B[71]), .Z(n584) );
  IV U134 ( .A(B[72]), .Z(n585) );
  IV U135 ( .A(B[73]), .Z(n586) );
  IV U136 ( .A(B[74]), .Z(n587) );
  IV U137 ( .A(B[470]), .Z(n983) );
  IV U138 ( .A(B[75]), .Z(n588) );
  IV U139 ( .A(B[76]), .Z(n589) );
  IV U140 ( .A(B[77]), .Z(n590) );
  IV U141 ( .A(B[78]), .Z(n591) );
  IV U142 ( .A(B[79]), .Z(n592) );
  IV U143 ( .A(B[80]), .Z(n593) );
  IV U144 ( .A(B[81]), .Z(n594) );
  IV U145 ( .A(B[82]), .Z(n595) );
  IV U146 ( .A(B[83]), .Z(n596) );
  IV U147 ( .A(B[84]), .Z(n597) );
  IV U148 ( .A(B[471]), .Z(n984) );
  IV U149 ( .A(B[85]), .Z(n598) );
  IV U150 ( .A(B[86]), .Z(n599) );
  IV U151 ( .A(B[87]), .Z(n600) );
  IV U152 ( .A(B[88]), .Z(n601) );
  IV U153 ( .A(B[89]), .Z(n602) );
  IV U154 ( .A(B[90]), .Z(n603) );
  IV U155 ( .A(B[91]), .Z(n604) );
  IV U156 ( .A(B[92]), .Z(n605) );
  IV U157 ( .A(B[93]), .Z(n606) );
  IV U158 ( .A(B[94]), .Z(n607) );
  IV U159 ( .A(B[472]), .Z(n985) );
  IV U160 ( .A(B[95]), .Z(n608) );
  IV U161 ( .A(B[96]), .Z(n609) );
  IV U162 ( .A(B[97]), .Z(n610) );
  IV U163 ( .A(B[98]), .Z(n611) );
  IV U164 ( .A(B[99]), .Z(n612) );
  IV U165 ( .A(B[100]), .Z(n613) );
  IV U166 ( .A(B[101]), .Z(n614) );
  IV U167 ( .A(B[102]), .Z(n615) );
  IV U168 ( .A(B[103]), .Z(n616) );
  IV U169 ( .A(B[104]), .Z(n617) );
  IV U170 ( .A(B[473]), .Z(n986) );
  IV U171 ( .A(B[105]), .Z(n618) );
  IV U172 ( .A(B[106]), .Z(n619) );
  IV U173 ( .A(B[107]), .Z(n620) );
  IV U174 ( .A(B[108]), .Z(n621) );
  IV U175 ( .A(B[109]), .Z(n622) );
  IV U176 ( .A(B[110]), .Z(n623) );
  IV U177 ( .A(B[111]), .Z(n624) );
  IV U178 ( .A(B[112]), .Z(n625) );
  IV U179 ( .A(B[113]), .Z(n626) );
  IV U180 ( .A(B[114]), .Z(n627) );
  IV U181 ( .A(B[474]), .Z(n987) );
  IV U182 ( .A(B[510]), .Z(n1023) );
  IV U183 ( .A(B[115]), .Z(n628) );
  IV U184 ( .A(B[116]), .Z(n629) );
  IV U185 ( .A(B[117]), .Z(n630) );
  IV U186 ( .A(B[118]), .Z(n631) );
  IV U187 ( .A(B[119]), .Z(n632) );
  IV U188 ( .A(B[120]), .Z(n633) );
  IV U189 ( .A(B[121]), .Z(n634) );
  IV U190 ( .A(B[122]), .Z(n635) );
  IV U191 ( .A(B[123]), .Z(n636) );
  IV U192 ( .A(B[124]), .Z(n637) );
  IV U193 ( .A(B[475]), .Z(n988) );
  IV U194 ( .A(B[125]), .Z(n638) );
  IV U195 ( .A(B[126]), .Z(n639) );
  IV U196 ( .A(B[127]), .Z(n640) );
  IV U197 ( .A(B[128]), .Z(n641) );
  IV U198 ( .A(B[129]), .Z(n642) );
  IV U199 ( .A(B[130]), .Z(n643) );
  IV U200 ( .A(B[131]), .Z(n644) );
  IV U201 ( .A(B[132]), .Z(n645) );
  IV U202 ( .A(B[133]), .Z(n646) );
  IV U203 ( .A(B[134]), .Z(n647) );
  IV U204 ( .A(B[476]), .Z(n989) );
  IV U205 ( .A(B[135]), .Z(n648) );
  IV U206 ( .A(B[136]), .Z(n649) );
  IV U207 ( .A(B[137]), .Z(n650) );
  IV U208 ( .A(B[138]), .Z(n651) );
  IV U209 ( .A(B[139]), .Z(n652) );
  IV U210 ( .A(B[140]), .Z(n653) );
  IV U211 ( .A(B[141]), .Z(n654) );
  IV U212 ( .A(B[142]), .Z(n655) );
  IV U213 ( .A(B[143]), .Z(n656) );
  IV U214 ( .A(B[144]), .Z(n657) );
  IV U215 ( .A(B[477]), .Z(n990) );
  IV U216 ( .A(B[145]), .Z(n658) );
  IV U217 ( .A(B[146]), .Z(n659) );
  IV U218 ( .A(B[147]), .Z(n660) );
  IV U219 ( .A(B[148]), .Z(n661) );
  IV U220 ( .A(B[149]), .Z(n662) );
  IV U221 ( .A(B[150]), .Z(n663) );
  IV U222 ( .A(B[151]), .Z(n664) );
  IV U223 ( .A(B[152]), .Z(n665) );
  IV U224 ( .A(B[153]), .Z(n666) );
  IV U225 ( .A(B[154]), .Z(n667) );
  IV U226 ( .A(B[478]), .Z(n991) );
  IV U227 ( .A(B[155]), .Z(n668) );
  IV U228 ( .A(B[156]), .Z(n669) );
  IV U229 ( .A(B[157]), .Z(n670) );
  IV U230 ( .A(B[158]), .Z(n671) );
  IV U231 ( .A(B[159]), .Z(n672) );
  IV U232 ( .A(B[160]), .Z(n673) );
  IV U233 ( .A(B[161]), .Z(n674) );
  IV U234 ( .A(B[162]), .Z(n675) );
  IV U235 ( .A(B[163]), .Z(n676) );
  IV U236 ( .A(B[164]), .Z(n677) );
  IV U237 ( .A(B[479]), .Z(n992) );
  IV U238 ( .A(B[165]), .Z(n678) );
  IV U239 ( .A(B[166]), .Z(n679) );
  IV U240 ( .A(B[167]), .Z(n680) );
  IV U241 ( .A(B[168]), .Z(n681) );
  IV U242 ( .A(B[169]), .Z(n682) );
  IV U243 ( .A(B[170]), .Z(n683) );
  IV U244 ( .A(B[171]), .Z(n684) );
  IV U245 ( .A(B[172]), .Z(n685) );
  IV U246 ( .A(B[173]), .Z(n686) );
  IV U247 ( .A(B[174]), .Z(n687) );
  IV U248 ( .A(B[480]), .Z(n993) );
  IV U249 ( .A(B[175]), .Z(n688) );
  IV U250 ( .A(B[176]), .Z(n689) );
  IV U251 ( .A(B[177]), .Z(n690) );
  IV U252 ( .A(B[178]), .Z(n691) );
  IV U253 ( .A(B[179]), .Z(n692) );
  IV U254 ( .A(B[180]), .Z(n693) );
  IV U255 ( .A(B[181]), .Z(n694) );
  IV U256 ( .A(B[182]), .Z(n695) );
  IV U257 ( .A(B[183]), .Z(n696) );
  IV U258 ( .A(B[184]), .Z(n697) );
  IV U259 ( .A(B[481]), .Z(n994) );
  IV U260 ( .A(B[185]), .Z(n698) );
  IV U261 ( .A(B[186]), .Z(n699) );
  IV U262 ( .A(B[187]), .Z(n700) );
  IV U263 ( .A(B[188]), .Z(n701) );
  IV U264 ( .A(B[189]), .Z(n702) );
  IV U265 ( .A(B[190]), .Z(n703) );
  IV U266 ( .A(B[191]), .Z(n704) );
  IV U267 ( .A(B[192]), .Z(n705) );
  IV U268 ( .A(B[193]), .Z(n706) );
  IV U269 ( .A(B[194]), .Z(n707) );
  IV U270 ( .A(B[482]), .Z(n995) );
  IV U271 ( .A(B[195]), .Z(n708) );
  IV U272 ( .A(B[196]), .Z(n709) );
  IV U273 ( .A(B[197]), .Z(n710) );
  IV U274 ( .A(B[198]), .Z(n711) );
  IV U275 ( .A(B[199]), .Z(n712) );
  IV U276 ( .A(B[200]), .Z(n713) );
  IV U277 ( .A(B[201]), .Z(n714) );
  IV U278 ( .A(B[202]), .Z(n715) );
  IV U279 ( .A(B[203]), .Z(n716) );
  IV U280 ( .A(B[204]), .Z(n717) );
  IV U281 ( .A(B[483]), .Z(n996) );
  IV U282 ( .A(B[205]), .Z(n718) );
  IV U283 ( .A(B[206]), .Z(n719) );
  IV U284 ( .A(B[207]), .Z(n720) );
  IV U285 ( .A(B[208]), .Z(n721) );
  IV U286 ( .A(B[209]), .Z(n722) );
  IV U287 ( .A(B[210]), .Z(n723) );
  IV U288 ( .A(B[211]), .Z(n724) );
  IV U289 ( .A(B[212]), .Z(n725) );
  IV U290 ( .A(B[213]), .Z(n726) );
  IV U291 ( .A(B[214]), .Z(n727) );
  IV U292 ( .A(B[484]), .Z(n997) );
  IV U293 ( .A(B[511]), .Z(n1024) );
  IV U294 ( .A(B[215]), .Z(n728) );
  IV U295 ( .A(B[216]), .Z(n729) );
  IV U296 ( .A(B[217]), .Z(n730) );
  IV U297 ( .A(B[218]), .Z(n731) );
  IV U298 ( .A(B[219]), .Z(n732) );
  IV U299 ( .A(B[220]), .Z(n733) );
  IV U300 ( .A(B[221]), .Z(n734) );
  IV U301 ( .A(B[222]), .Z(n735) );
  IV U302 ( .A(B[223]), .Z(n736) );
  IV U303 ( .A(B[224]), .Z(n737) );
  IV U304 ( .A(B[485]), .Z(n998) );
  IV U305 ( .A(B[225]), .Z(n738) );
  IV U306 ( .A(B[226]), .Z(n739) );
  IV U307 ( .A(B[227]), .Z(n740) );
  IV U308 ( .A(B[228]), .Z(n741) );
  IV U309 ( .A(B[229]), .Z(n742) );
  IV U310 ( .A(B[230]), .Z(n743) );
  IV U311 ( .A(B[231]), .Z(n744) );
  IV U312 ( .A(B[232]), .Z(n745) );
  IV U313 ( .A(B[233]), .Z(n746) );
  IV U314 ( .A(B[234]), .Z(n747) );
  IV U315 ( .A(B[486]), .Z(n999) );
  IV U316 ( .A(B[235]), .Z(n748) );
  IV U317 ( .A(B[236]), .Z(n749) );
  IV U318 ( .A(B[237]), .Z(n750) );
  IV U319 ( .A(B[238]), .Z(n751) );
  IV U320 ( .A(B[239]), .Z(n752) );
  IV U321 ( .A(B[240]), .Z(n753) );
  IV U322 ( .A(B[241]), .Z(n754) );
  IV U323 ( .A(B[242]), .Z(n755) );
  IV U324 ( .A(B[243]), .Z(n756) );
  IV U325 ( .A(B[244]), .Z(n757) );
  IV U326 ( .A(B[487]), .Z(n1000) );
  IV U327 ( .A(B[245]), .Z(n758) );
  IV U328 ( .A(B[246]), .Z(n759) );
  IV U329 ( .A(B[247]), .Z(n760) );
  IV U330 ( .A(B[248]), .Z(n761) );
  IV U331 ( .A(B[249]), .Z(n762) );
  IV U332 ( .A(B[250]), .Z(n763) );
  IV U333 ( .A(B[251]), .Z(n764) );
  IV U334 ( .A(B[252]), .Z(n765) );
  IV U335 ( .A(B[253]), .Z(n766) );
  IV U336 ( .A(B[254]), .Z(n767) );
  IV U337 ( .A(B[488]), .Z(n1001) );
  IV U338 ( .A(B[255]), .Z(n768) );
  IV U339 ( .A(B[256]), .Z(n769) );
  IV U340 ( .A(B[257]), .Z(n770) );
  IV U341 ( .A(B[258]), .Z(n771) );
  IV U342 ( .A(B[259]), .Z(n772) );
  IV U343 ( .A(B[260]), .Z(n773) );
  IV U344 ( .A(B[261]), .Z(n774) );
  IV U345 ( .A(B[262]), .Z(n775) );
  IV U346 ( .A(B[263]), .Z(n776) );
  IV U347 ( .A(B[264]), .Z(n777) );
  IV U348 ( .A(B[489]), .Z(n1002) );
  IV U349 ( .A(B[265]), .Z(n778) );
  IV U350 ( .A(B[266]), .Z(n779) );
  IV U351 ( .A(B[267]), .Z(n780) );
  IV U352 ( .A(B[268]), .Z(n781) );
  IV U353 ( .A(B[269]), .Z(n782) );
  IV U354 ( .A(B[270]), .Z(n783) );
  IV U355 ( .A(B[271]), .Z(n784) );
  IV U356 ( .A(B[272]), .Z(n785) );
  IV U357 ( .A(B[273]), .Z(n786) );
  IV U358 ( .A(B[274]), .Z(n787) );
  IV U359 ( .A(B[490]), .Z(n1003) );
  IV U360 ( .A(B[275]), .Z(n788) );
  IV U361 ( .A(B[276]), .Z(n789) );
  IV U362 ( .A(B[277]), .Z(n790) );
  IV U363 ( .A(B[278]), .Z(n791) );
  IV U364 ( .A(B[279]), .Z(n792) );
  IV U365 ( .A(B[280]), .Z(n793) );
  IV U366 ( .A(B[281]), .Z(n794) );
  IV U367 ( .A(B[282]), .Z(n795) );
  IV U368 ( .A(B[283]), .Z(n796) );
  IV U369 ( .A(B[284]), .Z(n797) );
  IV U370 ( .A(B[491]), .Z(n1004) );
  IV U371 ( .A(B[285]), .Z(n798) );
  IV U372 ( .A(B[286]), .Z(n799) );
  IV U373 ( .A(B[287]), .Z(n800) );
  IV U374 ( .A(B[288]), .Z(n801) );
  IV U375 ( .A(B[289]), .Z(n802) );
  IV U376 ( .A(B[290]), .Z(n803) );
  IV U377 ( .A(B[291]), .Z(n804) );
  IV U378 ( .A(B[292]), .Z(n805) );
  IV U379 ( .A(B[293]), .Z(n806) );
  IV U380 ( .A(B[294]), .Z(n807) );
  IV U381 ( .A(B[492]), .Z(n1005) );
  IV U382 ( .A(B[295]), .Z(n808) );
  IV U383 ( .A(B[296]), .Z(n809) );
  IV U384 ( .A(B[297]), .Z(n810) );
  IV U385 ( .A(B[298]), .Z(n811) );
  IV U386 ( .A(B[299]), .Z(n812) );
  IV U387 ( .A(B[300]), .Z(n813) );
  IV U388 ( .A(B[301]), .Z(n814) );
  IV U389 ( .A(B[302]), .Z(n815) );
  IV U390 ( .A(B[303]), .Z(n816) );
  IV U391 ( .A(B[304]), .Z(n817) );
  IV U392 ( .A(B[493]), .Z(n1006) );
  IV U393 ( .A(B[305]), .Z(n818) );
  IV U394 ( .A(B[306]), .Z(n819) );
  IV U395 ( .A(B[307]), .Z(n820) );
  IV U396 ( .A(B[308]), .Z(n821) );
  IV U397 ( .A(B[309]), .Z(n822) );
  IV U398 ( .A(B[310]), .Z(n823) );
  IV U399 ( .A(B[311]), .Z(n824) );
  IV U400 ( .A(B[312]), .Z(n825) );
  IV U401 ( .A(B[313]), .Z(n826) );
  IV U402 ( .A(B[314]), .Z(n827) );
  IV U403 ( .A(B[494]), .Z(n1007) );
  IV U404 ( .A(B[315]), .Z(n828) );
  IV U405 ( .A(B[316]), .Z(n829) );
  IV U406 ( .A(B[317]), .Z(n830) );
  IV U407 ( .A(B[318]), .Z(n831) );
  IV U408 ( .A(B[319]), .Z(n832) );
  IV U409 ( .A(B[320]), .Z(n833) );
  IV U410 ( .A(B[321]), .Z(n834) );
  IV U411 ( .A(B[322]), .Z(n835) );
  IV U412 ( .A(B[323]), .Z(n836) );
  IV U413 ( .A(B[324]), .Z(n837) );
  IV U414 ( .A(B[495]), .Z(n1008) );
  IV U415 ( .A(B[325]), .Z(n838) );
  IV U416 ( .A(B[326]), .Z(n839) );
  IV U417 ( .A(B[327]), .Z(n840) );
  IV U418 ( .A(B[328]), .Z(n841) );
  IV U419 ( .A(B[329]), .Z(n842) );
  IV U420 ( .A(B[330]), .Z(n843) );
  IV U421 ( .A(B[331]), .Z(n844) );
  IV U422 ( .A(B[332]), .Z(n845) );
  IV U423 ( .A(B[333]), .Z(n846) );
  IV U424 ( .A(B[334]), .Z(n847) );
  IV U425 ( .A(B[496]), .Z(n1009) );
  IV U426 ( .A(B[335]), .Z(n848) );
  IV U427 ( .A(B[336]), .Z(n849) );
  IV U428 ( .A(B[337]), .Z(n850) );
  IV U429 ( .A(B[338]), .Z(n851) );
  IV U430 ( .A(B[339]), .Z(n852) );
  IV U431 ( .A(B[340]), .Z(n853) );
  IV U432 ( .A(B[341]), .Z(n854) );
  IV U433 ( .A(B[342]), .Z(n855) );
  IV U434 ( .A(B[343]), .Z(n856) );
  IV U435 ( .A(B[344]), .Z(n857) );
  IV U436 ( .A(B[497]), .Z(n1010) );
  IV U437 ( .A(B[345]), .Z(n858) );
  IV U438 ( .A(B[346]), .Z(n859) );
  IV U439 ( .A(B[347]), .Z(n860) );
  IV U440 ( .A(B[348]), .Z(n861) );
  IV U441 ( .A(B[349]), .Z(n862) );
  IV U442 ( .A(B[350]), .Z(n863) );
  IV U443 ( .A(B[351]), .Z(n864) );
  IV U444 ( .A(B[352]), .Z(n865) );
  IV U445 ( .A(B[353]), .Z(n866) );
  IV U446 ( .A(B[354]), .Z(n867) );
  IV U447 ( .A(B[498]), .Z(n1011) );
  IV U448 ( .A(B[355]), .Z(n868) );
  IV U449 ( .A(B[356]), .Z(n869) );
  IV U450 ( .A(B[357]), .Z(n870) );
  IV U451 ( .A(B[358]), .Z(n871) );
  IV U452 ( .A(B[359]), .Z(n872) );
  IV U453 ( .A(B[360]), .Z(n873) );
  IV U454 ( .A(B[361]), .Z(n874) );
  IV U455 ( .A(B[362]), .Z(n875) );
  IV U456 ( .A(B[363]), .Z(n876) );
  IV U457 ( .A(B[364]), .Z(n877) );
  IV U458 ( .A(B[499]), .Z(n1012) );
  IV U459 ( .A(B[365]), .Z(n878) );
  IV U460 ( .A(B[366]), .Z(n879) );
  IV U461 ( .A(B[367]), .Z(n880) );
  IV U462 ( .A(B[368]), .Z(n881) );
  IV U463 ( .A(B[369]), .Z(n882) );
  IV U464 ( .A(B[370]), .Z(n883) );
  IV U465 ( .A(B[371]), .Z(n884) );
  IV U466 ( .A(B[372]), .Z(n885) );
  IV U467 ( .A(B[373]), .Z(n886) );
  IV U468 ( .A(B[374]), .Z(n887) );
  IV U469 ( .A(B[500]), .Z(n1013) );
  IV U470 ( .A(B[375]), .Z(n888) );
  IV U471 ( .A(B[376]), .Z(n889) );
  IV U472 ( .A(B[377]), .Z(n890) );
  IV U473 ( .A(B[378]), .Z(n891) );
  IV U474 ( .A(B[379]), .Z(n892) );
  IV U475 ( .A(B[380]), .Z(n893) );
  IV U476 ( .A(B[381]), .Z(n894) );
  IV U477 ( .A(B[382]), .Z(n895) );
  IV U478 ( .A(B[383]), .Z(n896) );
  IV U479 ( .A(B[384]), .Z(n897) );
  IV U480 ( .A(B[501]), .Z(n1014) );
  IV U481 ( .A(B[385]), .Z(n898) );
  IV U482 ( .A(B[386]), .Z(n899) );
  IV U483 ( .A(B[387]), .Z(n900) );
  IV U484 ( .A(B[388]), .Z(n901) );
  IV U485 ( .A(B[389]), .Z(n902) );
  IV U486 ( .A(B[390]), .Z(n903) );
  IV U487 ( .A(B[391]), .Z(n904) );
  IV U488 ( .A(B[392]), .Z(n905) );
  IV U489 ( .A(B[393]), .Z(n906) );
  IV U490 ( .A(B[394]), .Z(n907) );
  IV U491 ( .A(B[502]), .Z(n1015) );
  IV U492 ( .A(B[395]), .Z(n908) );
  IV U493 ( .A(B[396]), .Z(n909) );
  IV U494 ( .A(B[397]), .Z(n910) );
  IV U495 ( .A(B[398]), .Z(n911) );
  IV U496 ( .A(B[399]), .Z(n912) );
  IV U497 ( .A(B[400]), .Z(n913) );
  IV U498 ( .A(B[401]), .Z(n914) );
  IV U499 ( .A(B[402]), .Z(n915) );
  IV U500 ( .A(B[403]), .Z(n916) );
  IV U501 ( .A(B[404]), .Z(n917) );
  IV U502 ( .A(B[503]), .Z(n1016) );
  IV U503 ( .A(B[405]), .Z(n918) );
  IV U504 ( .A(B[406]), .Z(n919) );
  IV U505 ( .A(B[407]), .Z(n920) );
  IV U506 ( .A(B[408]), .Z(n921) );
  IV U507 ( .A(B[409]), .Z(n922) );
  IV U508 ( .A(B[410]), .Z(n923) );
  IV U509 ( .A(B[411]), .Z(n924) );
  IV U510 ( .A(B[412]), .Z(n925) );
  IV U511 ( .A(B[413]), .Z(n926) );
  IV U512 ( .A(B[414]), .Z(n927) );
  IV U513 ( .A(B[504]), .Z(n1017) );
endmodule


module modmult_step_N512_1_1 ( xregN_1, y, n, zin, zout );
  input [511:0] y;
  input [511:0] n;
  input [513:0] zin;
  output [513:0] zout;
  input xregN_1;
  wire   c1, c2, n4;
  wire   [513:0] w1;
  wire   [513:0] w2;
  wire   [513:0] w3;
  wire   [513:0] z2;
  wire   [513:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6;

  MUX_N514_6 MUX_1 ( .A({1'b0, 1'b0, y}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(xregN_1), .O({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, w1[511:0]}) );
  MUX_N514_5 MUX_2 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(c1), .O({SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, w2[511:0]}) );
  MUX_N514_4 MUX_3 ( .A({1'b0, 1'b0, n}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .S(n4), .O({SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, w3[511:0]}) );
  ADD_N514_1_1 ADD_1 ( .A({zin[512:0], 1'b0}), .B({1'b0, 1'b0, w1[511:0]}), 
        .CI(1'b0), .S(z2) );
  COMP_N514_4 COMP_1 ( .A(z2), .B({1'b0, 1'b0, n}), .O(c1) );
  SUB_N514_4 SUB_1 ( .A(z2), .B({1'b0, 1'b0, w2[511:0]}), .S(z3) );
  COMP_N514_3 COMP_2 ( .A({1'b0, 1'b0, n}), .B(z3), .O(c2) );
  SUB_N514_3 SUB_2 ( .A({1'b0, z3[512:0]}), .B({1'b0, 1'b0, w3[511:0]}), .S({
        SYNOPSYS_UNCONNECTED__6, zout[512:0]}) );
  IV U2 ( .A(c2), .Z(n4) );
endmodule


module modmult_N512_CC256 ( clk, rst, start, x, y, n, o );
  input [511:0] x;
  input [511:0] y;
  input [511:0] n;
  output [511:0] o;
  input clk, rst, start;
  wire   \zout[1][512] , \zin[1][512] , \zin[1][511] , \zin[1][510] ,
         \zin[1][509] , \zin[1][508] , \zin[1][507] , \zin[1][506] ,
         \zin[1][505] , \zin[1][504] , \zin[1][503] , \zin[1][502] ,
         \zin[1][501] , \zin[1][500] , \zin[1][499] , \zin[1][498] ,
         \zin[1][497] , \zin[1][496] , \zin[1][495] , \zin[1][494] ,
         \zin[1][493] , \zin[1][492] , \zin[1][491] , \zin[1][490] ,
         \zin[1][489] , \zin[1][488] , \zin[1][487] , \zin[1][486] ,
         \zin[1][485] , \zin[1][484] , \zin[1][483] , \zin[1][482] ,
         \zin[1][481] , \zin[1][480] , \zin[1][479] , \zin[1][478] ,
         \zin[1][477] , \zin[1][476] , \zin[1][475] , \zin[1][474] ,
         \zin[1][473] , \zin[1][472] , \zin[1][471] , \zin[1][470] ,
         \zin[1][469] , \zin[1][468] , \zin[1][467] , \zin[1][466] ,
         \zin[1][465] , \zin[1][464] , \zin[1][463] , \zin[1][462] ,
         \zin[1][461] , \zin[1][460] , \zin[1][459] , \zin[1][458] ,
         \zin[1][457] , \zin[1][456] , \zin[1][455] , \zin[1][454] ,
         \zin[1][453] , \zin[1][452] , \zin[1][451] , \zin[1][450] ,
         \zin[1][449] , \zin[1][448] , \zin[1][447] , \zin[1][446] ,
         \zin[1][445] , \zin[1][444] , \zin[1][443] , \zin[1][442] ,
         \zin[1][441] , \zin[1][440] , \zin[1][439] , \zin[1][438] ,
         \zin[1][437] , \zin[1][436] , \zin[1][435] , \zin[1][434] ,
         \zin[1][433] , \zin[1][432] , \zin[1][431] , \zin[1][430] ,
         \zin[1][429] , \zin[1][428] , \zin[1][427] , \zin[1][426] ,
         \zin[1][425] , \zin[1][424] , \zin[1][423] , \zin[1][422] ,
         \zin[1][421] , \zin[1][420] , \zin[1][419] , \zin[1][418] ,
         \zin[1][417] , \zin[1][416] , \zin[1][415] , \zin[1][414] ,
         \zin[1][413] , \zin[1][412] , \zin[1][411] , \zin[1][410] ,
         \zin[1][409] , \zin[1][408] , \zin[1][407] , \zin[1][406] ,
         \zin[1][405] , \zin[1][404] , \zin[1][403] , \zin[1][402] ,
         \zin[1][401] , \zin[1][400] , \zin[1][399] , \zin[1][398] ,
         \zin[1][397] , \zin[1][396] , \zin[1][395] , \zin[1][394] ,
         \zin[1][393] , \zin[1][392] , \zin[1][391] , \zin[1][390] ,
         \zin[1][389] , \zin[1][388] , \zin[1][387] , \zin[1][386] ,
         \zin[1][385] , \zin[1][384] , \zin[1][383] , \zin[1][382] ,
         \zin[1][381] , \zin[1][380] , \zin[1][379] , \zin[1][378] ,
         \zin[1][377] , \zin[1][376] , \zin[1][375] , \zin[1][374] ,
         \zin[1][373] , \zin[1][372] , \zin[1][371] , \zin[1][370] ,
         \zin[1][369] , \zin[1][368] , \zin[1][367] , \zin[1][366] ,
         \zin[1][365] , \zin[1][364] , \zin[1][363] , \zin[1][362] ,
         \zin[1][361] , \zin[1][360] , \zin[1][359] , \zin[1][358] ,
         \zin[1][357] , \zin[1][356] , \zin[1][355] , \zin[1][354] ,
         \zin[1][353] , \zin[1][352] , \zin[1][351] , \zin[1][350] ,
         \zin[1][349] , \zin[1][348] , \zin[1][347] , \zin[1][346] ,
         \zin[1][345] , \zin[1][344] , \zin[1][343] , \zin[1][342] ,
         \zin[1][341] , \zin[1][340] , \zin[1][339] , \zin[1][338] ,
         \zin[1][337] , \zin[1][336] , \zin[1][335] , \zin[1][334] ,
         \zin[1][333] , \zin[1][332] , \zin[1][331] , \zin[1][330] ,
         \zin[1][329] , \zin[1][328] , \zin[1][327] , \zin[1][326] ,
         \zin[1][325] , \zin[1][324] , \zin[1][323] , \zin[1][322] ,
         \zin[1][321] , \zin[1][320] , \zin[1][319] , \zin[1][318] ,
         \zin[1][317] , \zin[1][316] , \zin[1][315] , \zin[1][314] ,
         \zin[1][313] , \zin[1][312] , \zin[1][311] , \zin[1][310] ,
         \zin[1][309] , \zin[1][308] , \zin[1][307] , \zin[1][306] ,
         \zin[1][305] , \zin[1][304] , \zin[1][303] , \zin[1][302] ,
         \zin[1][301] , \zin[1][300] , \zin[1][299] , \zin[1][298] ,
         \zin[1][297] , \zin[1][296] , \zin[1][295] , \zin[1][294] ,
         \zin[1][293] , \zin[1][292] , \zin[1][291] , \zin[1][290] ,
         \zin[1][289] , \zin[1][288] , \zin[1][287] , \zin[1][286] ,
         \zin[1][285] , \zin[1][284] , \zin[1][283] , \zin[1][282] ,
         \zin[1][281] , \zin[1][280] , \zin[1][279] , \zin[1][278] ,
         \zin[1][277] , \zin[1][276] , \zin[1][275] , \zin[1][274] ,
         \zin[1][273] , \zin[1][272] , \zin[1][271] , \zin[1][270] ,
         \zin[1][269] , \zin[1][268] , \zin[1][267] , \zin[1][266] ,
         \zin[1][265] , \zin[1][264] , \zin[1][263] , \zin[1][262] ,
         \zin[1][261] , \zin[1][260] , \zin[1][259] , \zin[1][258] ,
         \zin[1][257] , \zin[1][256] , \zin[1][255] , \zin[1][254] ,
         \zin[1][253] , \zin[1][252] , \zin[1][251] , \zin[1][250] ,
         \zin[1][249] , \zin[1][248] , \zin[1][247] , \zin[1][246] ,
         \zin[1][245] , \zin[1][244] , \zin[1][243] , \zin[1][242] ,
         \zin[1][241] , \zin[1][240] , \zin[1][239] , \zin[1][238] ,
         \zin[1][237] , \zin[1][236] , \zin[1][235] , \zin[1][234] ,
         \zin[1][233] , \zin[1][232] , \zin[1][231] , \zin[1][230] ,
         \zin[1][229] , \zin[1][228] , \zin[1][227] , \zin[1][226] ,
         \zin[1][225] , \zin[1][224] , \zin[1][223] , \zin[1][222] ,
         \zin[1][221] , \zin[1][220] , \zin[1][219] , \zin[1][218] ,
         \zin[1][217] , \zin[1][216] , \zin[1][215] , \zin[1][214] ,
         \zin[1][213] , \zin[1][212] , \zin[1][211] , \zin[1][210] ,
         \zin[1][209] , \zin[1][208] , \zin[1][207] , \zin[1][206] ,
         \zin[1][205] , \zin[1][204] , \zin[1][203] , \zin[1][202] ,
         \zin[1][201] , \zin[1][200] , \zin[1][199] , \zin[1][198] ,
         \zin[1][197] , \zin[1][196] , \zin[1][195] , \zin[1][194] ,
         \zin[1][193] , \zin[1][192] , \zin[1][191] , \zin[1][190] ,
         \zin[1][189] , \zin[1][188] , \zin[1][187] , \zin[1][186] ,
         \zin[1][185] , \zin[1][184] , \zin[1][183] , \zin[1][182] ,
         \zin[1][181] , \zin[1][180] , \zin[1][179] , \zin[1][178] ,
         \zin[1][177] , \zin[1][176] , \zin[1][175] , \zin[1][174] ,
         \zin[1][173] , \zin[1][172] , \zin[1][171] , \zin[1][170] ,
         \zin[1][169] , \zin[1][168] , \zin[1][167] , \zin[1][166] ,
         \zin[1][165] , \zin[1][164] , \zin[1][163] , \zin[1][162] ,
         \zin[1][161] , \zin[1][160] , \zin[1][159] , \zin[1][158] ,
         \zin[1][157] , \zin[1][156] , \zin[1][155] , \zin[1][154] ,
         \zin[1][153] , \zin[1][152] , \zin[1][151] , \zin[1][150] ,
         \zin[1][149] , \zin[1][148] , \zin[1][147] , \zin[1][146] ,
         \zin[1][145] , \zin[1][144] , \zin[1][143] , \zin[1][142] ,
         \zin[1][141] , \zin[1][140] , \zin[1][139] , \zin[1][138] ,
         \zin[1][137] , \zin[1][136] , \zin[1][135] , \zin[1][134] ,
         \zin[1][133] , \zin[1][132] , \zin[1][131] , \zin[1][130] ,
         \zin[1][129] , \zin[1][128] , \zin[1][127] , \zin[1][126] ,
         \zin[1][125] , \zin[1][124] , \zin[1][123] , \zin[1][122] ,
         \zin[1][121] , \zin[1][120] , \zin[1][119] , \zin[1][118] ,
         \zin[1][117] , \zin[1][116] , \zin[1][115] , \zin[1][114] ,
         \zin[1][113] , \zin[1][112] , \zin[1][111] , \zin[1][110] ,
         \zin[1][109] , \zin[1][108] , \zin[1][107] , \zin[1][106] ,
         \zin[1][105] , \zin[1][104] , \zin[1][103] , \zin[1][102] ,
         \zin[1][101] , \zin[1][100] , \zin[1][99] , \zin[1][98] ,
         \zin[1][97] , \zin[1][96] , \zin[1][95] , \zin[1][94] , \zin[1][93] ,
         \zin[1][92] , \zin[1][91] , \zin[1][90] , \zin[1][89] , \zin[1][88] ,
         \zin[1][87] , \zin[1][86] , \zin[1][85] , \zin[1][84] , \zin[1][83] ,
         \zin[1][82] , \zin[1][81] , \zin[1][80] , \zin[1][79] , \zin[1][78] ,
         \zin[1][77] , \zin[1][76] , \zin[1][75] , \zin[1][74] , \zin[1][73] ,
         \zin[1][72] , \zin[1][71] , \zin[1][70] , \zin[1][69] , \zin[1][68] ,
         \zin[1][67] , \zin[1][66] , \zin[1][65] , \zin[1][64] , \zin[1][63] ,
         \zin[1][62] , \zin[1][61] , \zin[1][60] , \zin[1][59] , \zin[1][58] ,
         \zin[1][57] , \zin[1][56] , \zin[1][55] , \zin[1][54] , \zin[1][53] ,
         \zin[1][52] , \zin[1][51] , \zin[1][50] , \zin[1][49] , \zin[1][48] ,
         \zin[1][47] , \zin[1][46] , \zin[1][45] , \zin[1][44] , \zin[1][43] ,
         \zin[1][42] , \zin[1][41] , \zin[1][40] , \zin[1][39] , \zin[1][38] ,
         \zin[1][37] , \zin[1][36] , \zin[1][35] , \zin[1][34] , \zin[1][33] ,
         \zin[1][32] , \zin[1][31] , \zin[1][30] , \zin[1][29] , \zin[1][28] ,
         \zin[1][27] , \zin[1][26] , \zin[1][25] , \zin[1][24] , \zin[1][23] ,
         \zin[1][22] , \zin[1][21] , \zin[1][20] , \zin[1][19] , \zin[1][18] ,
         \zin[1][17] , \zin[1][16] , \zin[1][15] , \zin[1][14] , \zin[1][13] ,
         \zin[1][12] , \zin[1][11] , \zin[1][10] , \zin[1][9] , \zin[1][8] ,
         \zin[1][7] , \zin[1][6] , \zin[1][5] , \zin[1][4] , \zin[1][3] ,
         \zin[1][2] , \zin[1][1] , \zin[1][0] , \zin[0][512] , \zin[0][511] ,
         \zin[0][510] , \zin[0][509] , \zin[0][508] , \zin[0][507] ,
         \zin[0][506] , \zin[0][505] , \zin[0][504] , \zin[0][503] ,
         \zin[0][502] , \zin[0][501] , \zin[0][500] , \zin[0][499] ,
         \zin[0][498] , \zin[0][497] , \zin[0][496] , \zin[0][495] ,
         \zin[0][494] , \zin[0][493] , \zin[0][492] , \zin[0][491] ,
         \zin[0][490] , \zin[0][489] , \zin[0][488] , \zin[0][487] ,
         \zin[0][486] , \zin[0][485] , \zin[0][484] , \zin[0][483] ,
         \zin[0][482] , \zin[0][481] , \zin[0][480] , \zin[0][479] ,
         \zin[0][478] , \zin[0][477] , \zin[0][476] , \zin[0][475] ,
         \zin[0][474] , \zin[0][473] , \zin[0][472] , \zin[0][471] ,
         \zin[0][470] , \zin[0][469] , \zin[0][468] , \zin[0][467] ,
         \zin[0][466] , \zin[0][465] , \zin[0][464] , \zin[0][463] ,
         \zin[0][462] , \zin[0][461] , \zin[0][460] , \zin[0][459] ,
         \zin[0][458] , \zin[0][457] , \zin[0][456] , \zin[0][455] ,
         \zin[0][454] , \zin[0][453] , \zin[0][452] , \zin[0][451] ,
         \zin[0][450] , \zin[0][449] , \zin[0][448] , \zin[0][447] ,
         \zin[0][446] , \zin[0][445] , \zin[0][444] , \zin[0][443] ,
         \zin[0][442] , \zin[0][441] , \zin[0][440] , \zin[0][439] ,
         \zin[0][438] , \zin[0][437] , \zin[0][436] , \zin[0][435] ,
         \zin[0][434] , \zin[0][433] , \zin[0][432] , \zin[0][431] ,
         \zin[0][430] , \zin[0][429] , \zin[0][428] , \zin[0][427] ,
         \zin[0][426] , \zin[0][425] , \zin[0][424] , \zin[0][423] ,
         \zin[0][422] , \zin[0][421] , \zin[0][420] , \zin[0][419] ,
         \zin[0][418] , \zin[0][417] , \zin[0][416] , \zin[0][415] ,
         \zin[0][414] , \zin[0][413] , \zin[0][412] , \zin[0][411] ,
         \zin[0][410] , \zin[0][409] , \zin[0][408] , \zin[0][407] ,
         \zin[0][406] , \zin[0][405] , \zin[0][404] , \zin[0][403] ,
         \zin[0][402] , \zin[0][401] , \zin[0][400] , \zin[0][399] ,
         \zin[0][398] , \zin[0][397] , \zin[0][396] , \zin[0][395] ,
         \zin[0][394] , \zin[0][393] , \zin[0][392] , \zin[0][391] ,
         \zin[0][390] , \zin[0][389] , \zin[0][388] , \zin[0][387] ,
         \zin[0][386] , \zin[0][385] , \zin[0][384] , \zin[0][383] ,
         \zin[0][382] , \zin[0][381] , \zin[0][380] , \zin[0][379] ,
         \zin[0][378] , \zin[0][377] , \zin[0][376] , \zin[0][375] ,
         \zin[0][374] , \zin[0][373] , \zin[0][372] , \zin[0][371] ,
         \zin[0][370] , \zin[0][369] , \zin[0][368] , \zin[0][367] ,
         \zin[0][366] , \zin[0][365] , \zin[0][364] , \zin[0][363] ,
         \zin[0][362] , \zin[0][361] , \zin[0][360] , \zin[0][359] ,
         \zin[0][358] , \zin[0][357] , \zin[0][356] , \zin[0][355] ,
         \zin[0][354] , \zin[0][353] , \zin[0][352] , \zin[0][351] ,
         \zin[0][350] , \zin[0][349] , \zin[0][348] , \zin[0][347] ,
         \zin[0][346] , \zin[0][345] , \zin[0][344] , \zin[0][343] ,
         \zin[0][342] , \zin[0][341] , \zin[0][340] , \zin[0][339] ,
         \zin[0][338] , \zin[0][337] , \zin[0][336] , \zin[0][335] ,
         \zin[0][334] , \zin[0][333] , \zin[0][332] , \zin[0][331] ,
         \zin[0][330] , \zin[0][329] , \zin[0][328] , \zin[0][327] ,
         \zin[0][326] , \zin[0][325] , \zin[0][324] , \zin[0][323] ,
         \zin[0][322] , \zin[0][321] , \zin[0][320] , \zin[0][319] ,
         \zin[0][318] , \zin[0][317] , \zin[0][316] , \zin[0][315] ,
         \zin[0][314] , \zin[0][313] , \zin[0][312] , \zin[0][311] ,
         \zin[0][310] , \zin[0][309] , \zin[0][308] , \zin[0][307] ,
         \zin[0][306] , \zin[0][305] , \zin[0][304] , \zin[0][303] ,
         \zin[0][302] , \zin[0][301] , \zin[0][300] , \zin[0][299] ,
         \zin[0][298] , \zin[0][297] , \zin[0][296] , \zin[0][295] ,
         \zin[0][294] , \zin[0][293] , \zin[0][292] , \zin[0][291] ,
         \zin[0][290] , \zin[0][289] , \zin[0][288] , \zin[0][287] ,
         \zin[0][286] , \zin[0][285] , \zin[0][284] , \zin[0][283] ,
         \zin[0][282] , \zin[0][281] , \zin[0][280] , \zin[0][279] ,
         \zin[0][278] , \zin[0][277] , \zin[0][276] , \zin[0][275] ,
         \zin[0][274] , \zin[0][273] , \zin[0][272] , \zin[0][271] ,
         \zin[0][270] , \zin[0][269] , \zin[0][268] , \zin[0][267] ,
         \zin[0][266] , \zin[0][265] , \zin[0][264] , \zin[0][263] ,
         \zin[0][262] , \zin[0][261] , \zin[0][260] , \zin[0][259] ,
         \zin[0][258] , \zin[0][257] , \zin[0][256] , \zin[0][255] ,
         \zin[0][254] , \zin[0][253] , \zin[0][252] , \zin[0][251] ,
         \zin[0][250] , \zin[0][249] , \zin[0][248] , \zin[0][247] ,
         \zin[0][246] , \zin[0][245] , \zin[0][244] , \zin[0][243] ,
         \zin[0][242] , \zin[0][241] , \zin[0][240] , \zin[0][239] ,
         \zin[0][238] , \zin[0][237] , \zin[0][236] , \zin[0][235] ,
         \zin[0][234] , \zin[0][233] , \zin[0][232] , \zin[0][231] ,
         \zin[0][230] , \zin[0][229] , \zin[0][228] , \zin[0][227] ,
         \zin[0][226] , \zin[0][225] , \zin[0][224] , \zin[0][223] ,
         \zin[0][222] , \zin[0][221] , \zin[0][220] , \zin[0][219] ,
         \zin[0][218] , \zin[0][217] , \zin[0][216] , \zin[0][215] ,
         \zin[0][214] , \zin[0][213] , \zin[0][212] , \zin[0][211] ,
         \zin[0][210] , \zin[0][209] , \zin[0][208] , \zin[0][207] ,
         \zin[0][206] , \zin[0][205] , \zin[0][204] , \zin[0][203] ,
         \zin[0][202] , \zin[0][201] , \zin[0][200] , \zin[0][199] ,
         \zin[0][198] , \zin[0][197] , \zin[0][196] , \zin[0][195] ,
         \zin[0][194] , \zin[0][193] , \zin[0][192] , \zin[0][191] ,
         \zin[0][190] , \zin[0][189] , \zin[0][188] , \zin[0][187] ,
         \zin[0][186] , \zin[0][185] , \zin[0][184] , \zin[0][183] ,
         \zin[0][182] , \zin[0][181] , \zin[0][180] , \zin[0][179] ,
         \zin[0][178] , \zin[0][177] , \zin[0][176] , \zin[0][175] ,
         \zin[0][174] , \zin[0][173] , \zin[0][172] , \zin[0][171] ,
         \zin[0][170] , \zin[0][169] , \zin[0][168] , \zin[0][167] ,
         \zin[0][166] , \zin[0][165] , \zin[0][164] , \zin[0][163] ,
         \zin[0][162] , \zin[0][161] , \zin[0][160] , \zin[0][159] ,
         \zin[0][158] , \zin[0][157] , \zin[0][156] , \zin[0][155] ,
         \zin[0][154] , \zin[0][153] , \zin[0][152] , \zin[0][151] ,
         \zin[0][150] , \zin[0][149] , \zin[0][148] , \zin[0][147] ,
         \zin[0][146] , \zin[0][145] , \zin[0][144] , \zin[0][143] ,
         \zin[0][142] , \zin[0][141] , \zin[0][140] , \zin[0][139] ,
         \zin[0][138] , \zin[0][137] , \zin[0][136] , \zin[0][135] ,
         \zin[0][134] , \zin[0][133] , \zin[0][132] , \zin[0][131] ,
         \zin[0][130] , \zin[0][129] , \zin[0][128] , \zin[0][127] ,
         \zin[0][126] , \zin[0][125] , \zin[0][124] , \zin[0][123] ,
         \zin[0][122] , \zin[0][121] , \zin[0][120] , \zin[0][119] ,
         \zin[0][118] , \zin[0][117] , \zin[0][116] , \zin[0][115] ,
         \zin[0][114] , \zin[0][113] , \zin[0][112] , \zin[0][111] ,
         \zin[0][110] , \zin[0][109] , \zin[0][108] , \zin[0][107] ,
         \zin[0][106] , \zin[0][105] , \zin[0][104] , \zin[0][103] ,
         \zin[0][102] , \zin[0][101] , \zin[0][100] , \zin[0][99] ,
         \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] ,
         \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] ,
         \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] ,
         \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] ,
         \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] ,
         \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] ,
         \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] ,
         \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] ,
         \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] ,
         \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] ,
         \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] ,
         \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] ,
         \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] ,
         \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] ,
         \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] ,
         \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] ,
         \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] ,
         \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] ,
         \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] ,
         \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] ;
  wire   [511:0] xin;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1;

  modmult_step_N512_1_0 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[511]), 
        .y(y), .n(n), .zin({1'b0, \zin[0][512] , \zin[0][511] , \zin[0][510] , 
        \zin[0][509] , \zin[0][508] , \zin[0][507] , \zin[0][506] , 
        \zin[0][505] , \zin[0][504] , \zin[0][503] , \zin[0][502] , 
        \zin[0][501] , \zin[0][500] , \zin[0][499] , \zin[0][498] , 
        \zin[0][497] , \zin[0][496] , \zin[0][495] , \zin[0][494] , 
        \zin[0][493] , \zin[0][492] , \zin[0][491] , \zin[0][490] , 
        \zin[0][489] , \zin[0][488] , \zin[0][487] , \zin[0][486] , 
        \zin[0][485] , \zin[0][484] , \zin[0][483] , \zin[0][482] , 
        \zin[0][481] , \zin[0][480] , \zin[0][479] , \zin[0][478] , 
        \zin[0][477] , \zin[0][476] , \zin[0][475] , \zin[0][474] , 
        \zin[0][473] , \zin[0][472] , \zin[0][471] , \zin[0][470] , 
        \zin[0][469] , \zin[0][468] , \zin[0][467] , \zin[0][466] , 
        \zin[0][465] , \zin[0][464] , \zin[0][463] , \zin[0][462] , 
        \zin[0][461] , \zin[0][460] , \zin[0][459] , \zin[0][458] , 
        \zin[0][457] , \zin[0][456] , \zin[0][455] , \zin[0][454] , 
        \zin[0][453] , \zin[0][452] , \zin[0][451] , \zin[0][450] , 
        \zin[0][449] , \zin[0][448] , \zin[0][447] , \zin[0][446] , 
        \zin[0][445] , \zin[0][444] , \zin[0][443] , \zin[0][442] , 
        \zin[0][441] , \zin[0][440] , \zin[0][439] , \zin[0][438] , 
        \zin[0][437] , \zin[0][436] , \zin[0][435] , \zin[0][434] , 
        \zin[0][433] , \zin[0][432] , \zin[0][431] , \zin[0][430] , 
        \zin[0][429] , \zin[0][428] , \zin[0][427] , \zin[0][426] , 
        \zin[0][425] , \zin[0][424] , \zin[0][423] , \zin[0][422] , 
        \zin[0][421] , \zin[0][420] , \zin[0][419] , \zin[0][418] , 
        \zin[0][417] , \zin[0][416] , \zin[0][415] , \zin[0][414] , 
        \zin[0][413] , \zin[0][412] , \zin[0][411] , \zin[0][410] , 
        \zin[0][409] , \zin[0][408] , \zin[0][407] , \zin[0][406] , 
        \zin[0][405] , \zin[0][404] , \zin[0][403] , \zin[0][402] , 
        \zin[0][401] , \zin[0][400] , \zin[0][399] , \zin[0][398] , 
        \zin[0][397] , \zin[0][396] , \zin[0][395] , \zin[0][394] , 
        \zin[0][393] , \zin[0][392] , \zin[0][391] , \zin[0][390] , 
        \zin[0][389] , \zin[0][388] , \zin[0][387] , \zin[0][386] , 
        \zin[0][385] , \zin[0][384] , \zin[0][383] , \zin[0][382] , 
        \zin[0][381] , \zin[0][380] , \zin[0][379] , \zin[0][378] , 
        \zin[0][377] , \zin[0][376] , \zin[0][375] , \zin[0][374] , 
        \zin[0][373] , \zin[0][372] , \zin[0][371] , \zin[0][370] , 
        \zin[0][369] , \zin[0][368] , \zin[0][367] , \zin[0][366] , 
        \zin[0][365] , \zin[0][364] , \zin[0][363] , \zin[0][362] , 
        \zin[0][361] , \zin[0][360] , \zin[0][359] , \zin[0][358] , 
        \zin[0][357] , \zin[0][356] , \zin[0][355] , \zin[0][354] , 
        \zin[0][353] , \zin[0][352] , \zin[0][351] , \zin[0][350] , 
        \zin[0][349] , \zin[0][348] , \zin[0][347] , \zin[0][346] , 
        \zin[0][345] , \zin[0][344] , \zin[0][343] , \zin[0][342] , 
        \zin[0][341] , \zin[0][340] , \zin[0][339] , \zin[0][338] , 
        \zin[0][337] , \zin[0][336] , \zin[0][335] , \zin[0][334] , 
        \zin[0][333] , \zin[0][332] , \zin[0][331] , \zin[0][330] , 
        \zin[0][329] , \zin[0][328] , \zin[0][327] , \zin[0][326] , 
        \zin[0][325] , \zin[0][324] , \zin[0][323] , \zin[0][322] , 
        \zin[0][321] , \zin[0][320] , \zin[0][319] , \zin[0][318] , 
        \zin[0][317] , \zin[0][316] , \zin[0][315] , \zin[0][314] , 
        \zin[0][313] , \zin[0][312] , \zin[0][311] , \zin[0][310] , 
        \zin[0][309] , \zin[0][308] , \zin[0][307] , \zin[0][306] , 
        \zin[0][305] , \zin[0][304] , \zin[0][303] , \zin[0][302] , 
        \zin[0][301] , \zin[0][300] , \zin[0][299] , \zin[0][298] , 
        \zin[0][297] , \zin[0][296] , \zin[0][295] , \zin[0][294] , 
        \zin[0][293] , \zin[0][292] , \zin[0][291] , \zin[0][290] , 
        \zin[0][289] , \zin[0][288] , \zin[0][287] , \zin[0][286] , 
        \zin[0][285] , \zin[0][284] , \zin[0][283] , \zin[0][282] , 
        \zin[0][281] , \zin[0][280] , \zin[0][279] , \zin[0][278] , 
        \zin[0][277] , \zin[0][276] , \zin[0][275] , \zin[0][274] , 
        \zin[0][273] , \zin[0][272] , \zin[0][271] , \zin[0][270] , 
        \zin[0][269] , \zin[0][268] , \zin[0][267] , \zin[0][266] , 
        \zin[0][265] , \zin[0][264] , \zin[0][263] , \zin[0][262] , 
        \zin[0][261] , \zin[0][260] , \zin[0][259] , \zin[0][258] , 
        \zin[0][257] , \zin[0][256] , \zin[0][255] , \zin[0][254] , 
        \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] , 
        \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] , 
        \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] , 
        \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] , 
        \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] , 
        \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] , 
        \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] , 
        \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] , 
        \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] , 
        \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] , 
        \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] , 
        \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] , 
        \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] , 
        \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] , 
        \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] , 
        \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] , 
        \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] , 
        \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] , 
        \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] , 
        \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] , 
        \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] , 
        \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] , 
        \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] , 
        \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] , 
        \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] , 
        \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] , 
        \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] , 
        \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] , 
        \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] , 
        \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] , 
        \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] , 
        \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] , 
        \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] , 
        \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] , 
        \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] , 
        \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] , 
        \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] , 
        \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] , 
        \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] , \zin[0][97] , 
        \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] , \zin[0][92] , 
        \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] , \zin[0][87] , 
        \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] , \zin[0][82] , 
        \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] , \zin[0][77] , 
        \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] , \zin[0][72] , 
        \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] , \zin[0][67] , 
        \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] , \zin[0][62] , 
        \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] , \zin[0][57] , 
        \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] , \zin[0][52] , 
        \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] , \zin[0][47] , 
        \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] , \zin[0][42] , 
        \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] , \zin[0][37] , 
        \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] , \zin[0][32] , 
        \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] , \zin[0][27] , 
        \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] , \zin[0][22] , 
        \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] , \zin[0][17] , 
        \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] , \zin[0][12] , 
        \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] , \zin[0][7] , 
        \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] , \zin[0][2] , 
        \zin[0][1] , \zin[0][0] }), .zout({SYNOPSYS_UNCONNECTED__0, 
        \zin[1][512] , \zin[1][511] , \zin[1][510] , \zin[1][509] , 
        \zin[1][508] , \zin[1][507] , \zin[1][506] , \zin[1][505] , 
        \zin[1][504] , \zin[1][503] , \zin[1][502] , \zin[1][501] , 
        \zin[1][500] , \zin[1][499] , \zin[1][498] , \zin[1][497] , 
        \zin[1][496] , \zin[1][495] , \zin[1][494] , \zin[1][493] , 
        \zin[1][492] , \zin[1][491] , \zin[1][490] , \zin[1][489] , 
        \zin[1][488] , \zin[1][487] , \zin[1][486] , \zin[1][485] , 
        \zin[1][484] , \zin[1][483] , \zin[1][482] , \zin[1][481] , 
        \zin[1][480] , \zin[1][479] , \zin[1][478] , \zin[1][477] , 
        \zin[1][476] , \zin[1][475] , \zin[1][474] , \zin[1][473] , 
        \zin[1][472] , \zin[1][471] , \zin[1][470] , \zin[1][469] , 
        \zin[1][468] , \zin[1][467] , \zin[1][466] , \zin[1][465] , 
        \zin[1][464] , \zin[1][463] , \zin[1][462] , \zin[1][461] , 
        \zin[1][460] , \zin[1][459] , \zin[1][458] , \zin[1][457] , 
        \zin[1][456] , \zin[1][455] , \zin[1][454] , \zin[1][453] , 
        \zin[1][452] , \zin[1][451] , \zin[1][450] , \zin[1][449] , 
        \zin[1][448] , \zin[1][447] , \zin[1][446] , \zin[1][445] , 
        \zin[1][444] , \zin[1][443] , \zin[1][442] , \zin[1][441] , 
        \zin[1][440] , \zin[1][439] , \zin[1][438] , \zin[1][437] , 
        \zin[1][436] , \zin[1][435] , \zin[1][434] , \zin[1][433] , 
        \zin[1][432] , \zin[1][431] , \zin[1][430] , \zin[1][429] , 
        \zin[1][428] , \zin[1][427] , \zin[1][426] , \zin[1][425] , 
        \zin[1][424] , \zin[1][423] , \zin[1][422] , \zin[1][421] , 
        \zin[1][420] , \zin[1][419] , \zin[1][418] , \zin[1][417] , 
        \zin[1][416] , \zin[1][415] , \zin[1][414] , \zin[1][413] , 
        \zin[1][412] , \zin[1][411] , \zin[1][410] , \zin[1][409] , 
        \zin[1][408] , \zin[1][407] , \zin[1][406] , \zin[1][405] , 
        \zin[1][404] , \zin[1][403] , \zin[1][402] , \zin[1][401] , 
        \zin[1][400] , \zin[1][399] , \zin[1][398] , \zin[1][397] , 
        \zin[1][396] , \zin[1][395] , \zin[1][394] , \zin[1][393] , 
        \zin[1][392] , \zin[1][391] , \zin[1][390] , \zin[1][389] , 
        \zin[1][388] , \zin[1][387] , \zin[1][386] , \zin[1][385] , 
        \zin[1][384] , \zin[1][383] , \zin[1][382] , \zin[1][381] , 
        \zin[1][380] , \zin[1][379] , \zin[1][378] , \zin[1][377] , 
        \zin[1][376] , \zin[1][375] , \zin[1][374] , \zin[1][373] , 
        \zin[1][372] , \zin[1][371] , \zin[1][370] , \zin[1][369] , 
        \zin[1][368] , \zin[1][367] , \zin[1][366] , \zin[1][365] , 
        \zin[1][364] , \zin[1][363] , \zin[1][362] , \zin[1][361] , 
        \zin[1][360] , \zin[1][359] , \zin[1][358] , \zin[1][357] , 
        \zin[1][356] , \zin[1][355] , \zin[1][354] , \zin[1][353] , 
        \zin[1][352] , \zin[1][351] , \zin[1][350] , \zin[1][349] , 
        \zin[1][348] , \zin[1][347] , \zin[1][346] , \zin[1][345] , 
        \zin[1][344] , \zin[1][343] , \zin[1][342] , \zin[1][341] , 
        \zin[1][340] , \zin[1][339] , \zin[1][338] , \zin[1][337] , 
        \zin[1][336] , \zin[1][335] , \zin[1][334] , \zin[1][333] , 
        \zin[1][332] , \zin[1][331] , \zin[1][330] , \zin[1][329] , 
        \zin[1][328] , \zin[1][327] , \zin[1][326] , \zin[1][325] , 
        \zin[1][324] , \zin[1][323] , \zin[1][322] , \zin[1][321] , 
        \zin[1][320] , \zin[1][319] , \zin[1][318] , \zin[1][317] , 
        \zin[1][316] , \zin[1][315] , \zin[1][314] , \zin[1][313] , 
        \zin[1][312] , \zin[1][311] , \zin[1][310] , \zin[1][309] , 
        \zin[1][308] , \zin[1][307] , \zin[1][306] , \zin[1][305] , 
        \zin[1][304] , \zin[1][303] , \zin[1][302] , \zin[1][301] , 
        \zin[1][300] , \zin[1][299] , \zin[1][298] , \zin[1][297] , 
        \zin[1][296] , \zin[1][295] , \zin[1][294] , \zin[1][293] , 
        \zin[1][292] , \zin[1][291] , \zin[1][290] , \zin[1][289] , 
        \zin[1][288] , \zin[1][287] , \zin[1][286] , \zin[1][285] , 
        \zin[1][284] , \zin[1][283] , \zin[1][282] , \zin[1][281] , 
        \zin[1][280] , \zin[1][279] , \zin[1][278] , \zin[1][277] , 
        \zin[1][276] , \zin[1][275] , \zin[1][274] , \zin[1][273] , 
        \zin[1][272] , \zin[1][271] , \zin[1][270] , \zin[1][269] , 
        \zin[1][268] , \zin[1][267] , \zin[1][266] , \zin[1][265] , 
        \zin[1][264] , \zin[1][263] , \zin[1][262] , \zin[1][261] , 
        \zin[1][260] , \zin[1][259] , \zin[1][258] , \zin[1][257] , 
        \zin[1][256] , \zin[1][255] , \zin[1][254] , \zin[1][253] , 
        \zin[1][252] , \zin[1][251] , \zin[1][250] , \zin[1][249] , 
        \zin[1][248] , \zin[1][247] , \zin[1][246] , \zin[1][245] , 
        \zin[1][244] , \zin[1][243] , \zin[1][242] , \zin[1][241] , 
        \zin[1][240] , \zin[1][239] , \zin[1][238] , \zin[1][237] , 
        \zin[1][236] , \zin[1][235] , \zin[1][234] , \zin[1][233] , 
        \zin[1][232] , \zin[1][231] , \zin[1][230] , \zin[1][229] , 
        \zin[1][228] , \zin[1][227] , \zin[1][226] , \zin[1][225] , 
        \zin[1][224] , \zin[1][223] , \zin[1][222] , \zin[1][221] , 
        \zin[1][220] , \zin[1][219] , \zin[1][218] , \zin[1][217] , 
        \zin[1][216] , \zin[1][215] , \zin[1][214] , \zin[1][213] , 
        \zin[1][212] , \zin[1][211] , \zin[1][210] , \zin[1][209] , 
        \zin[1][208] , \zin[1][207] , \zin[1][206] , \zin[1][205] , 
        \zin[1][204] , \zin[1][203] , \zin[1][202] , \zin[1][201] , 
        \zin[1][200] , \zin[1][199] , \zin[1][198] , \zin[1][197] , 
        \zin[1][196] , \zin[1][195] , \zin[1][194] , \zin[1][193] , 
        \zin[1][192] , \zin[1][191] , \zin[1][190] , \zin[1][189] , 
        \zin[1][188] , \zin[1][187] , \zin[1][186] , \zin[1][185] , 
        \zin[1][184] , \zin[1][183] , \zin[1][182] , \zin[1][181] , 
        \zin[1][180] , \zin[1][179] , \zin[1][178] , \zin[1][177] , 
        \zin[1][176] , \zin[1][175] , \zin[1][174] , \zin[1][173] , 
        \zin[1][172] , \zin[1][171] , \zin[1][170] , \zin[1][169] , 
        \zin[1][168] , \zin[1][167] , \zin[1][166] , \zin[1][165] , 
        \zin[1][164] , \zin[1][163] , \zin[1][162] , \zin[1][161] , 
        \zin[1][160] , \zin[1][159] , \zin[1][158] , \zin[1][157] , 
        \zin[1][156] , \zin[1][155] , \zin[1][154] , \zin[1][153] , 
        \zin[1][152] , \zin[1][151] , \zin[1][150] , \zin[1][149] , 
        \zin[1][148] , \zin[1][147] , \zin[1][146] , \zin[1][145] , 
        \zin[1][144] , \zin[1][143] , \zin[1][142] , \zin[1][141] , 
        \zin[1][140] , \zin[1][139] , \zin[1][138] , \zin[1][137] , 
        \zin[1][136] , \zin[1][135] , \zin[1][134] , \zin[1][133] , 
        \zin[1][132] , \zin[1][131] , \zin[1][130] , \zin[1][129] , 
        \zin[1][128] , \zin[1][127] , \zin[1][126] , \zin[1][125] , 
        \zin[1][124] , \zin[1][123] , \zin[1][122] , \zin[1][121] , 
        \zin[1][120] , \zin[1][119] , \zin[1][118] , \zin[1][117] , 
        \zin[1][116] , \zin[1][115] , \zin[1][114] , \zin[1][113] , 
        \zin[1][112] , \zin[1][111] , \zin[1][110] , \zin[1][109] , 
        \zin[1][108] , \zin[1][107] , \zin[1][106] , \zin[1][105] , 
        \zin[1][104] , \zin[1][103] , \zin[1][102] , \zin[1][101] , 
        \zin[1][100] , \zin[1][99] , \zin[1][98] , \zin[1][97] , \zin[1][96] , 
        \zin[1][95] , \zin[1][94] , \zin[1][93] , \zin[1][92] , \zin[1][91] , 
        \zin[1][90] , \zin[1][89] , \zin[1][88] , \zin[1][87] , \zin[1][86] , 
        \zin[1][85] , \zin[1][84] , \zin[1][83] , \zin[1][82] , \zin[1][81] , 
        \zin[1][80] , \zin[1][79] , \zin[1][78] , \zin[1][77] , \zin[1][76] , 
        \zin[1][75] , \zin[1][74] , \zin[1][73] , \zin[1][72] , \zin[1][71] , 
        \zin[1][70] , \zin[1][69] , \zin[1][68] , \zin[1][67] , \zin[1][66] , 
        \zin[1][65] , \zin[1][64] , \zin[1][63] , \zin[1][62] , \zin[1][61] , 
        \zin[1][60] , \zin[1][59] , \zin[1][58] , \zin[1][57] , \zin[1][56] , 
        \zin[1][55] , \zin[1][54] , \zin[1][53] , \zin[1][52] , \zin[1][51] , 
        \zin[1][50] , \zin[1][49] , \zin[1][48] , \zin[1][47] , \zin[1][46] , 
        \zin[1][45] , \zin[1][44] , \zin[1][43] , \zin[1][42] , \zin[1][41] , 
        \zin[1][40] , \zin[1][39] , \zin[1][38] , \zin[1][37] , \zin[1][36] , 
        \zin[1][35] , \zin[1][34] , \zin[1][33] , \zin[1][32] , \zin[1][31] , 
        \zin[1][30] , \zin[1][29] , \zin[1][28] , \zin[1][27] , \zin[1][26] , 
        \zin[1][25] , \zin[1][24] , \zin[1][23] , \zin[1][22] , \zin[1][21] , 
        \zin[1][20] , \zin[1][19] , \zin[1][18] , \zin[1][17] , \zin[1][16] , 
        \zin[1][15] , \zin[1][14] , \zin[1][13] , \zin[1][12] , \zin[1][11] , 
        \zin[1][10] , \zin[1][9] , \zin[1][8] , \zin[1][7] , \zin[1][6] , 
        \zin[1][5] , \zin[1][4] , \zin[1][3] , \zin[1][2] , \zin[1][1] , 
        \zin[1][0] }) );
  modmult_step_N512_1_1 \MODMULT_STEP[1].modmult_step_  ( .xregN_1(xin[510]), 
        .y(y), .n(n), .zin({1'b0, \zin[1][512] , \zin[1][511] , \zin[1][510] , 
        \zin[1][509] , \zin[1][508] , \zin[1][507] , \zin[1][506] , 
        \zin[1][505] , \zin[1][504] , \zin[1][503] , \zin[1][502] , 
        \zin[1][501] , \zin[1][500] , \zin[1][499] , \zin[1][498] , 
        \zin[1][497] , \zin[1][496] , \zin[1][495] , \zin[1][494] , 
        \zin[1][493] , \zin[1][492] , \zin[1][491] , \zin[1][490] , 
        \zin[1][489] , \zin[1][488] , \zin[1][487] , \zin[1][486] , 
        \zin[1][485] , \zin[1][484] , \zin[1][483] , \zin[1][482] , 
        \zin[1][481] , \zin[1][480] , \zin[1][479] , \zin[1][478] , 
        \zin[1][477] , \zin[1][476] , \zin[1][475] , \zin[1][474] , 
        \zin[1][473] , \zin[1][472] , \zin[1][471] , \zin[1][470] , 
        \zin[1][469] , \zin[1][468] , \zin[1][467] , \zin[1][466] , 
        \zin[1][465] , \zin[1][464] , \zin[1][463] , \zin[1][462] , 
        \zin[1][461] , \zin[1][460] , \zin[1][459] , \zin[1][458] , 
        \zin[1][457] , \zin[1][456] , \zin[1][455] , \zin[1][454] , 
        \zin[1][453] , \zin[1][452] , \zin[1][451] , \zin[1][450] , 
        \zin[1][449] , \zin[1][448] , \zin[1][447] , \zin[1][446] , 
        \zin[1][445] , \zin[1][444] , \zin[1][443] , \zin[1][442] , 
        \zin[1][441] , \zin[1][440] , \zin[1][439] , \zin[1][438] , 
        \zin[1][437] , \zin[1][436] , \zin[1][435] , \zin[1][434] , 
        \zin[1][433] , \zin[1][432] , \zin[1][431] , \zin[1][430] , 
        \zin[1][429] , \zin[1][428] , \zin[1][427] , \zin[1][426] , 
        \zin[1][425] , \zin[1][424] , \zin[1][423] , \zin[1][422] , 
        \zin[1][421] , \zin[1][420] , \zin[1][419] , \zin[1][418] , 
        \zin[1][417] , \zin[1][416] , \zin[1][415] , \zin[1][414] , 
        \zin[1][413] , \zin[1][412] , \zin[1][411] , \zin[1][410] , 
        \zin[1][409] , \zin[1][408] , \zin[1][407] , \zin[1][406] , 
        \zin[1][405] , \zin[1][404] , \zin[1][403] , \zin[1][402] , 
        \zin[1][401] , \zin[1][400] , \zin[1][399] , \zin[1][398] , 
        \zin[1][397] , \zin[1][396] , \zin[1][395] , \zin[1][394] , 
        \zin[1][393] , \zin[1][392] , \zin[1][391] , \zin[1][390] , 
        \zin[1][389] , \zin[1][388] , \zin[1][387] , \zin[1][386] , 
        \zin[1][385] , \zin[1][384] , \zin[1][383] , \zin[1][382] , 
        \zin[1][381] , \zin[1][380] , \zin[1][379] , \zin[1][378] , 
        \zin[1][377] , \zin[1][376] , \zin[1][375] , \zin[1][374] , 
        \zin[1][373] , \zin[1][372] , \zin[1][371] , \zin[1][370] , 
        \zin[1][369] , \zin[1][368] , \zin[1][367] , \zin[1][366] , 
        \zin[1][365] , \zin[1][364] , \zin[1][363] , \zin[1][362] , 
        \zin[1][361] , \zin[1][360] , \zin[1][359] , \zin[1][358] , 
        \zin[1][357] , \zin[1][356] , \zin[1][355] , \zin[1][354] , 
        \zin[1][353] , \zin[1][352] , \zin[1][351] , \zin[1][350] , 
        \zin[1][349] , \zin[1][348] , \zin[1][347] , \zin[1][346] , 
        \zin[1][345] , \zin[1][344] , \zin[1][343] , \zin[1][342] , 
        \zin[1][341] , \zin[1][340] , \zin[1][339] , \zin[1][338] , 
        \zin[1][337] , \zin[1][336] , \zin[1][335] , \zin[1][334] , 
        \zin[1][333] , \zin[1][332] , \zin[1][331] , \zin[1][330] , 
        \zin[1][329] , \zin[1][328] , \zin[1][327] , \zin[1][326] , 
        \zin[1][325] , \zin[1][324] , \zin[1][323] , \zin[1][322] , 
        \zin[1][321] , \zin[1][320] , \zin[1][319] , \zin[1][318] , 
        \zin[1][317] , \zin[1][316] , \zin[1][315] , \zin[1][314] , 
        \zin[1][313] , \zin[1][312] , \zin[1][311] , \zin[1][310] , 
        \zin[1][309] , \zin[1][308] , \zin[1][307] , \zin[1][306] , 
        \zin[1][305] , \zin[1][304] , \zin[1][303] , \zin[1][302] , 
        \zin[1][301] , \zin[1][300] , \zin[1][299] , \zin[1][298] , 
        \zin[1][297] , \zin[1][296] , \zin[1][295] , \zin[1][294] , 
        \zin[1][293] , \zin[1][292] , \zin[1][291] , \zin[1][290] , 
        \zin[1][289] , \zin[1][288] , \zin[1][287] , \zin[1][286] , 
        \zin[1][285] , \zin[1][284] , \zin[1][283] , \zin[1][282] , 
        \zin[1][281] , \zin[1][280] , \zin[1][279] , \zin[1][278] , 
        \zin[1][277] , \zin[1][276] , \zin[1][275] , \zin[1][274] , 
        \zin[1][273] , \zin[1][272] , \zin[1][271] , \zin[1][270] , 
        \zin[1][269] , \zin[1][268] , \zin[1][267] , \zin[1][266] , 
        \zin[1][265] , \zin[1][264] , \zin[1][263] , \zin[1][262] , 
        \zin[1][261] , \zin[1][260] , \zin[1][259] , \zin[1][258] , 
        \zin[1][257] , \zin[1][256] , \zin[1][255] , \zin[1][254] , 
        \zin[1][253] , \zin[1][252] , \zin[1][251] , \zin[1][250] , 
        \zin[1][249] , \zin[1][248] , \zin[1][247] , \zin[1][246] , 
        \zin[1][245] , \zin[1][244] , \zin[1][243] , \zin[1][242] , 
        \zin[1][241] , \zin[1][240] , \zin[1][239] , \zin[1][238] , 
        \zin[1][237] , \zin[1][236] , \zin[1][235] , \zin[1][234] , 
        \zin[1][233] , \zin[1][232] , \zin[1][231] , \zin[1][230] , 
        \zin[1][229] , \zin[1][228] , \zin[1][227] , \zin[1][226] , 
        \zin[1][225] , \zin[1][224] , \zin[1][223] , \zin[1][222] , 
        \zin[1][221] , \zin[1][220] , \zin[1][219] , \zin[1][218] , 
        \zin[1][217] , \zin[1][216] , \zin[1][215] , \zin[1][214] , 
        \zin[1][213] , \zin[1][212] , \zin[1][211] , \zin[1][210] , 
        \zin[1][209] , \zin[1][208] , \zin[1][207] , \zin[1][206] , 
        \zin[1][205] , \zin[1][204] , \zin[1][203] , \zin[1][202] , 
        \zin[1][201] , \zin[1][200] , \zin[1][199] , \zin[1][198] , 
        \zin[1][197] , \zin[1][196] , \zin[1][195] , \zin[1][194] , 
        \zin[1][193] , \zin[1][192] , \zin[1][191] , \zin[1][190] , 
        \zin[1][189] , \zin[1][188] , \zin[1][187] , \zin[1][186] , 
        \zin[1][185] , \zin[1][184] , \zin[1][183] , \zin[1][182] , 
        \zin[1][181] , \zin[1][180] , \zin[1][179] , \zin[1][178] , 
        \zin[1][177] , \zin[1][176] , \zin[1][175] , \zin[1][174] , 
        \zin[1][173] , \zin[1][172] , \zin[1][171] , \zin[1][170] , 
        \zin[1][169] , \zin[1][168] , \zin[1][167] , \zin[1][166] , 
        \zin[1][165] , \zin[1][164] , \zin[1][163] , \zin[1][162] , 
        \zin[1][161] , \zin[1][160] , \zin[1][159] , \zin[1][158] , 
        \zin[1][157] , \zin[1][156] , \zin[1][155] , \zin[1][154] , 
        \zin[1][153] , \zin[1][152] , \zin[1][151] , \zin[1][150] , 
        \zin[1][149] , \zin[1][148] , \zin[1][147] , \zin[1][146] , 
        \zin[1][145] , \zin[1][144] , \zin[1][143] , \zin[1][142] , 
        \zin[1][141] , \zin[1][140] , \zin[1][139] , \zin[1][138] , 
        \zin[1][137] , \zin[1][136] , \zin[1][135] , \zin[1][134] , 
        \zin[1][133] , \zin[1][132] , \zin[1][131] , \zin[1][130] , 
        \zin[1][129] , \zin[1][128] , \zin[1][127] , \zin[1][126] , 
        \zin[1][125] , \zin[1][124] , \zin[1][123] , \zin[1][122] , 
        \zin[1][121] , \zin[1][120] , \zin[1][119] , \zin[1][118] , 
        \zin[1][117] , \zin[1][116] , \zin[1][115] , \zin[1][114] , 
        \zin[1][113] , \zin[1][112] , \zin[1][111] , \zin[1][110] , 
        \zin[1][109] , \zin[1][108] , \zin[1][107] , \zin[1][106] , 
        \zin[1][105] , \zin[1][104] , \zin[1][103] , \zin[1][102] , 
        \zin[1][101] , \zin[1][100] , \zin[1][99] , \zin[1][98] , \zin[1][97] , 
        \zin[1][96] , \zin[1][95] , \zin[1][94] , \zin[1][93] , \zin[1][92] , 
        \zin[1][91] , \zin[1][90] , \zin[1][89] , \zin[1][88] , \zin[1][87] , 
        \zin[1][86] , \zin[1][85] , \zin[1][84] , \zin[1][83] , \zin[1][82] , 
        \zin[1][81] , \zin[1][80] , \zin[1][79] , \zin[1][78] , \zin[1][77] , 
        \zin[1][76] , \zin[1][75] , \zin[1][74] , \zin[1][73] , \zin[1][72] , 
        \zin[1][71] , \zin[1][70] , \zin[1][69] , \zin[1][68] , \zin[1][67] , 
        \zin[1][66] , \zin[1][65] , \zin[1][64] , \zin[1][63] , \zin[1][62] , 
        \zin[1][61] , \zin[1][60] , \zin[1][59] , \zin[1][58] , \zin[1][57] , 
        \zin[1][56] , \zin[1][55] , \zin[1][54] , \zin[1][53] , \zin[1][52] , 
        \zin[1][51] , \zin[1][50] , \zin[1][49] , \zin[1][48] , \zin[1][47] , 
        \zin[1][46] , \zin[1][45] , \zin[1][44] , \zin[1][43] , \zin[1][42] , 
        \zin[1][41] , \zin[1][40] , \zin[1][39] , \zin[1][38] , \zin[1][37] , 
        \zin[1][36] , \zin[1][35] , \zin[1][34] , \zin[1][33] , \zin[1][32] , 
        \zin[1][31] , \zin[1][30] , \zin[1][29] , \zin[1][28] , \zin[1][27] , 
        \zin[1][26] , \zin[1][25] , \zin[1][24] , \zin[1][23] , \zin[1][22] , 
        \zin[1][21] , \zin[1][20] , \zin[1][19] , \zin[1][18] , \zin[1][17] , 
        \zin[1][16] , \zin[1][15] , \zin[1][14] , \zin[1][13] , \zin[1][12] , 
        \zin[1][11] , \zin[1][10] , \zin[1][9] , \zin[1][8] , \zin[1][7] , 
        \zin[1][6] , \zin[1][5] , \zin[1][4] , \zin[1][3] , \zin[1][2] , 
        \zin[1][1] , \zin[1][0] }), .zout({SYNOPSYS_UNCONNECTED__1, 
        \zout[1][512] , o}) );
  DFF \xreg_reg[1]  ( .D(1'b0), .CLK(clk), .RST(start), .I(x[1]), .Q(xin[1])
         );
  DFF \xreg_reg[3]  ( .D(xin[1]), .CLK(clk), .RST(start), .I(x[3]), .Q(xin[3])
         );
  DFF \xreg_reg[5]  ( .D(xin[3]), .CLK(clk), .RST(start), .I(x[5]), .Q(xin[5])
         );
  DFF \xreg_reg[7]  ( .D(xin[5]), .CLK(clk), .RST(start), .I(x[7]), .Q(xin[7])
         );
  DFF \xreg_reg[9]  ( .D(xin[7]), .CLK(clk), .RST(start), .I(x[9]), .Q(xin[9])
         );
  DFF \xreg_reg[11]  ( .D(xin[9]), .CLK(clk), .RST(start), .I(x[11]), .Q(
        xin[11]) );
  DFF \xreg_reg[13]  ( .D(xin[11]), .CLK(clk), .RST(start), .I(x[13]), .Q(
        xin[13]) );
  DFF \xreg_reg[15]  ( .D(xin[13]), .CLK(clk), .RST(start), .I(x[15]), .Q(
        xin[15]) );
  DFF \xreg_reg[17]  ( .D(xin[15]), .CLK(clk), .RST(start), .I(x[17]), .Q(
        xin[17]) );
  DFF \xreg_reg[19]  ( .D(xin[17]), .CLK(clk), .RST(start), .I(x[19]), .Q(
        xin[19]) );
  DFF \xreg_reg[21]  ( .D(xin[19]), .CLK(clk), .RST(start), .I(x[21]), .Q(
        xin[21]) );
  DFF \xreg_reg[23]  ( .D(xin[21]), .CLK(clk), .RST(start), .I(x[23]), .Q(
        xin[23]) );
  DFF \xreg_reg[25]  ( .D(xin[23]), .CLK(clk), .RST(start), .I(x[25]), .Q(
        xin[25]) );
  DFF \xreg_reg[27]  ( .D(xin[25]), .CLK(clk), .RST(start), .I(x[27]), .Q(
        xin[27]) );
  DFF \xreg_reg[29]  ( .D(xin[27]), .CLK(clk), .RST(start), .I(x[29]), .Q(
        xin[29]) );
  DFF \xreg_reg[31]  ( .D(xin[29]), .CLK(clk), .RST(start), .I(x[31]), .Q(
        xin[31]) );
  DFF \xreg_reg[33]  ( .D(xin[31]), .CLK(clk), .RST(start), .I(x[33]), .Q(
        xin[33]) );
  DFF \xreg_reg[35]  ( .D(xin[33]), .CLK(clk), .RST(start), .I(x[35]), .Q(
        xin[35]) );
  DFF \xreg_reg[37]  ( .D(xin[35]), .CLK(clk), .RST(start), .I(x[37]), .Q(
        xin[37]) );
  DFF \xreg_reg[39]  ( .D(xin[37]), .CLK(clk), .RST(start), .I(x[39]), .Q(
        xin[39]) );
  DFF \xreg_reg[41]  ( .D(xin[39]), .CLK(clk), .RST(start), .I(x[41]), .Q(
        xin[41]) );
  DFF \xreg_reg[43]  ( .D(xin[41]), .CLK(clk), .RST(start), .I(x[43]), .Q(
        xin[43]) );
  DFF \xreg_reg[45]  ( .D(xin[43]), .CLK(clk), .RST(start), .I(x[45]), .Q(
        xin[45]) );
  DFF \xreg_reg[47]  ( .D(xin[45]), .CLK(clk), .RST(start), .I(x[47]), .Q(
        xin[47]) );
  DFF \xreg_reg[49]  ( .D(xin[47]), .CLK(clk), .RST(start), .I(x[49]), .Q(
        xin[49]) );
  DFF \xreg_reg[51]  ( .D(xin[49]), .CLK(clk), .RST(start), .I(x[51]), .Q(
        xin[51]) );
  DFF \xreg_reg[53]  ( .D(xin[51]), .CLK(clk), .RST(start), .I(x[53]), .Q(
        xin[53]) );
  DFF \xreg_reg[55]  ( .D(xin[53]), .CLK(clk), .RST(start), .I(x[55]), .Q(
        xin[55]) );
  DFF \xreg_reg[57]  ( .D(xin[55]), .CLK(clk), .RST(start), .I(x[57]), .Q(
        xin[57]) );
  DFF \xreg_reg[59]  ( .D(xin[57]), .CLK(clk), .RST(start), .I(x[59]), .Q(
        xin[59]) );
  DFF \xreg_reg[61]  ( .D(xin[59]), .CLK(clk), .RST(start), .I(x[61]), .Q(
        xin[61]) );
  DFF \xreg_reg[63]  ( .D(xin[61]), .CLK(clk), .RST(start), .I(x[63]), .Q(
        xin[63]) );
  DFF \xreg_reg[65]  ( .D(xin[63]), .CLK(clk), .RST(start), .I(x[65]), .Q(
        xin[65]) );
  DFF \xreg_reg[67]  ( .D(xin[65]), .CLK(clk), .RST(start), .I(x[67]), .Q(
        xin[67]) );
  DFF \xreg_reg[69]  ( .D(xin[67]), .CLK(clk), .RST(start), .I(x[69]), .Q(
        xin[69]) );
  DFF \xreg_reg[71]  ( .D(xin[69]), .CLK(clk), .RST(start), .I(x[71]), .Q(
        xin[71]) );
  DFF \xreg_reg[73]  ( .D(xin[71]), .CLK(clk), .RST(start), .I(x[73]), .Q(
        xin[73]) );
  DFF \xreg_reg[75]  ( .D(xin[73]), .CLK(clk), .RST(start), .I(x[75]), .Q(
        xin[75]) );
  DFF \xreg_reg[77]  ( .D(xin[75]), .CLK(clk), .RST(start), .I(x[77]), .Q(
        xin[77]) );
  DFF \xreg_reg[79]  ( .D(xin[77]), .CLK(clk), .RST(start), .I(x[79]), .Q(
        xin[79]) );
  DFF \xreg_reg[81]  ( .D(xin[79]), .CLK(clk), .RST(start), .I(x[81]), .Q(
        xin[81]) );
  DFF \xreg_reg[83]  ( .D(xin[81]), .CLK(clk), .RST(start), .I(x[83]), .Q(
        xin[83]) );
  DFF \xreg_reg[85]  ( .D(xin[83]), .CLK(clk), .RST(start), .I(x[85]), .Q(
        xin[85]) );
  DFF \xreg_reg[87]  ( .D(xin[85]), .CLK(clk), .RST(start), .I(x[87]), .Q(
        xin[87]) );
  DFF \xreg_reg[89]  ( .D(xin[87]), .CLK(clk), .RST(start), .I(x[89]), .Q(
        xin[89]) );
  DFF \xreg_reg[91]  ( .D(xin[89]), .CLK(clk), .RST(start), .I(x[91]), .Q(
        xin[91]) );
  DFF \xreg_reg[93]  ( .D(xin[91]), .CLK(clk), .RST(start), .I(x[93]), .Q(
        xin[93]) );
  DFF \xreg_reg[95]  ( .D(xin[93]), .CLK(clk), .RST(start), .I(x[95]), .Q(
        xin[95]) );
  DFF \xreg_reg[97]  ( .D(xin[95]), .CLK(clk), .RST(start), .I(x[97]), .Q(
        xin[97]) );
  DFF \xreg_reg[99]  ( .D(xin[97]), .CLK(clk), .RST(start), .I(x[99]), .Q(
        xin[99]) );
  DFF \xreg_reg[101]  ( .D(xin[99]), .CLK(clk), .RST(start), .I(x[101]), .Q(
        xin[101]) );
  DFF \xreg_reg[103]  ( .D(xin[101]), .CLK(clk), .RST(start), .I(x[103]), .Q(
        xin[103]) );
  DFF \xreg_reg[105]  ( .D(xin[103]), .CLK(clk), .RST(start), .I(x[105]), .Q(
        xin[105]) );
  DFF \xreg_reg[107]  ( .D(xin[105]), .CLK(clk), .RST(start), .I(x[107]), .Q(
        xin[107]) );
  DFF \xreg_reg[109]  ( .D(xin[107]), .CLK(clk), .RST(start), .I(x[109]), .Q(
        xin[109]) );
  DFF \xreg_reg[111]  ( .D(xin[109]), .CLK(clk), .RST(start), .I(x[111]), .Q(
        xin[111]) );
  DFF \xreg_reg[113]  ( .D(xin[111]), .CLK(clk), .RST(start), .I(x[113]), .Q(
        xin[113]) );
  DFF \xreg_reg[115]  ( .D(xin[113]), .CLK(clk), .RST(start), .I(x[115]), .Q(
        xin[115]) );
  DFF \xreg_reg[117]  ( .D(xin[115]), .CLK(clk), .RST(start), .I(x[117]), .Q(
        xin[117]) );
  DFF \xreg_reg[119]  ( .D(xin[117]), .CLK(clk), .RST(start), .I(x[119]), .Q(
        xin[119]) );
  DFF \xreg_reg[121]  ( .D(xin[119]), .CLK(clk), .RST(start), .I(x[121]), .Q(
        xin[121]) );
  DFF \xreg_reg[123]  ( .D(xin[121]), .CLK(clk), .RST(start), .I(x[123]), .Q(
        xin[123]) );
  DFF \xreg_reg[125]  ( .D(xin[123]), .CLK(clk), .RST(start), .I(x[125]), .Q(
        xin[125]) );
  DFF \xreg_reg[127]  ( .D(xin[125]), .CLK(clk), .RST(start), .I(x[127]), .Q(
        xin[127]) );
  DFF \xreg_reg[129]  ( .D(xin[127]), .CLK(clk), .RST(start), .I(x[129]), .Q(
        xin[129]) );
  DFF \xreg_reg[131]  ( .D(xin[129]), .CLK(clk), .RST(start), .I(x[131]), .Q(
        xin[131]) );
  DFF \xreg_reg[133]  ( .D(xin[131]), .CLK(clk), .RST(start), .I(x[133]), .Q(
        xin[133]) );
  DFF \xreg_reg[135]  ( .D(xin[133]), .CLK(clk), .RST(start), .I(x[135]), .Q(
        xin[135]) );
  DFF \xreg_reg[137]  ( .D(xin[135]), .CLK(clk), .RST(start), .I(x[137]), .Q(
        xin[137]) );
  DFF \xreg_reg[139]  ( .D(xin[137]), .CLK(clk), .RST(start), .I(x[139]), .Q(
        xin[139]) );
  DFF \xreg_reg[141]  ( .D(xin[139]), .CLK(clk), .RST(start), .I(x[141]), .Q(
        xin[141]) );
  DFF \xreg_reg[143]  ( .D(xin[141]), .CLK(clk), .RST(start), .I(x[143]), .Q(
        xin[143]) );
  DFF \xreg_reg[145]  ( .D(xin[143]), .CLK(clk), .RST(start), .I(x[145]), .Q(
        xin[145]) );
  DFF \xreg_reg[147]  ( .D(xin[145]), .CLK(clk), .RST(start), .I(x[147]), .Q(
        xin[147]) );
  DFF \xreg_reg[149]  ( .D(xin[147]), .CLK(clk), .RST(start), .I(x[149]), .Q(
        xin[149]) );
  DFF \xreg_reg[151]  ( .D(xin[149]), .CLK(clk), .RST(start), .I(x[151]), .Q(
        xin[151]) );
  DFF \xreg_reg[153]  ( .D(xin[151]), .CLK(clk), .RST(start), .I(x[153]), .Q(
        xin[153]) );
  DFF \xreg_reg[155]  ( .D(xin[153]), .CLK(clk), .RST(start), .I(x[155]), .Q(
        xin[155]) );
  DFF \xreg_reg[157]  ( .D(xin[155]), .CLK(clk), .RST(start), .I(x[157]), .Q(
        xin[157]) );
  DFF \xreg_reg[159]  ( .D(xin[157]), .CLK(clk), .RST(start), .I(x[159]), .Q(
        xin[159]) );
  DFF \xreg_reg[161]  ( .D(xin[159]), .CLK(clk), .RST(start), .I(x[161]), .Q(
        xin[161]) );
  DFF \xreg_reg[163]  ( .D(xin[161]), .CLK(clk), .RST(start), .I(x[163]), .Q(
        xin[163]) );
  DFF \xreg_reg[165]  ( .D(xin[163]), .CLK(clk), .RST(start), .I(x[165]), .Q(
        xin[165]) );
  DFF \xreg_reg[167]  ( .D(xin[165]), .CLK(clk), .RST(start), .I(x[167]), .Q(
        xin[167]) );
  DFF \xreg_reg[169]  ( .D(xin[167]), .CLK(clk), .RST(start), .I(x[169]), .Q(
        xin[169]) );
  DFF \xreg_reg[171]  ( .D(xin[169]), .CLK(clk), .RST(start), .I(x[171]), .Q(
        xin[171]) );
  DFF \xreg_reg[173]  ( .D(xin[171]), .CLK(clk), .RST(start), .I(x[173]), .Q(
        xin[173]) );
  DFF \xreg_reg[175]  ( .D(xin[173]), .CLK(clk), .RST(start), .I(x[175]), .Q(
        xin[175]) );
  DFF \xreg_reg[177]  ( .D(xin[175]), .CLK(clk), .RST(start), .I(x[177]), .Q(
        xin[177]) );
  DFF \xreg_reg[179]  ( .D(xin[177]), .CLK(clk), .RST(start), .I(x[179]), .Q(
        xin[179]) );
  DFF \xreg_reg[181]  ( .D(xin[179]), .CLK(clk), .RST(start), .I(x[181]), .Q(
        xin[181]) );
  DFF \xreg_reg[183]  ( .D(xin[181]), .CLK(clk), .RST(start), .I(x[183]), .Q(
        xin[183]) );
  DFF \xreg_reg[185]  ( .D(xin[183]), .CLK(clk), .RST(start), .I(x[185]), .Q(
        xin[185]) );
  DFF \xreg_reg[187]  ( .D(xin[185]), .CLK(clk), .RST(start), .I(x[187]), .Q(
        xin[187]) );
  DFF \xreg_reg[189]  ( .D(xin[187]), .CLK(clk), .RST(start), .I(x[189]), .Q(
        xin[189]) );
  DFF \xreg_reg[191]  ( .D(xin[189]), .CLK(clk), .RST(start), .I(x[191]), .Q(
        xin[191]) );
  DFF \xreg_reg[193]  ( .D(xin[191]), .CLK(clk), .RST(start), .I(x[193]), .Q(
        xin[193]) );
  DFF \xreg_reg[195]  ( .D(xin[193]), .CLK(clk), .RST(start), .I(x[195]), .Q(
        xin[195]) );
  DFF \xreg_reg[197]  ( .D(xin[195]), .CLK(clk), .RST(start), .I(x[197]), .Q(
        xin[197]) );
  DFF \xreg_reg[199]  ( .D(xin[197]), .CLK(clk), .RST(start), .I(x[199]), .Q(
        xin[199]) );
  DFF \xreg_reg[201]  ( .D(xin[199]), .CLK(clk), .RST(start), .I(x[201]), .Q(
        xin[201]) );
  DFF \xreg_reg[203]  ( .D(xin[201]), .CLK(clk), .RST(start), .I(x[203]), .Q(
        xin[203]) );
  DFF \xreg_reg[205]  ( .D(xin[203]), .CLK(clk), .RST(start), .I(x[205]), .Q(
        xin[205]) );
  DFF \xreg_reg[207]  ( .D(xin[205]), .CLK(clk), .RST(start), .I(x[207]), .Q(
        xin[207]) );
  DFF \xreg_reg[209]  ( .D(xin[207]), .CLK(clk), .RST(start), .I(x[209]), .Q(
        xin[209]) );
  DFF \xreg_reg[211]  ( .D(xin[209]), .CLK(clk), .RST(start), .I(x[211]), .Q(
        xin[211]) );
  DFF \xreg_reg[213]  ( .D(xin[211]), .CLK(clk), .RST(start), .I(x[213]), .Q(
        xin[213]) );
  DFF \xreg_reg[215]  ( .D(xin[213]), .CLK(clk), .RST(start), .I(x[215]), .Q(
        xin[215]) );
  DFF \xreg_reg[217]  ( .D(xin[215]), .CLK(clk), .RST(start), .I(x[217]), .Q(
        xin[217]) );
  DFF \xreg_reg[219]  ( .D(xin[217]), .CLK(clk), .RST(start), .I(x[219]), .Q(
        xin[219]) );
  DFF \xreg_reg[221]  ( .D(xin[219]), .CLK(clk), .RST(start), .I(x[221]), .Q(
        xin[221]) );
  DFF \xreg_reg[223]  ( .D(xin[221]), .CLK(clk), .RST(start), .I(x[223]), .Q(
        xin[223]) );
  DFF \xreg_reg[225]  ( .D(xin[223]), .CLK(clk), .RST(start), .I(x[225]), .Q(
        xin[225]) );
  DFF \xreg_reg[227]  ( .D(xin[225]), .CLK(clk), .RST(start), .I(x[227]), .Q(
        xin[227]) );
  DFF \xreg_reg[229]  ( .D(xin[227]), .CLK(clk), .RST(start), .I(x[229]), .Q(
        xin[229]) );
  DFF \xreg_reg[231]  ( .D(xin[229]), .CLK(clk), .RST(start), .I(x[231]), .Q(
        xin[231]) );
  DFF \xreg_reg[233]  ( .D(xin[231]), .CLK(clk), .RST(start), .I(x[233]), .Q(
        xin[233]) );
  DFF \xreg_reg[235]  ( .D(xin[233]), .CLK(clk), .RST(start), .I(x[235]), .Q(
        xin[235]) );
  DFF \xreg_reg[237]  ( .D(xin[235]), .CLK(clk), .RST(start), .I(x[237]), .Q(
        xin[237]) );
  DFF \xreg_reg[239]  ( .D(xin[237]), .CLK(clk), .RST(start), .I(x[239]), .Q(
        xin[239]) );
  DFF \xreg_reg[241]  ( .D(xin[239]), .CLK(clk), .RST(start), .I(x[241]), .Q(
        xin[241]) );
  DFF \xreg_reg[243]  ( .D(xin[241]), .CLK(clk), .RST(start), .I(x[243]), .Q(
        xin[243]) );
  DFF \xreg_reg[245]  ( .D(xin[243]), .CLK(clk), .RST(start), .I(x[245]), .Q(
        xin[245]) );
  DFF \xreg_reg[247]  ( .D(xin[245]), .CLK(clk), .RST(start), .I(x[247]), .Q(
        xin[247]) );
  DFF \xreg_reg[249]  ( .D(xin[247]), .CLK(clk), .RST(start), .I(x[249]), .Q(
        xin[249]) );
  DFF \xreg_reg[251]  ( .D(xin[249]), .CLK(clk), .RST(start), .I(x[251]), .Q(
        xin[251]) );
  DFF \xreg_reg[253]  ( .D(xin[251]), .CLK(clk), .RST(start), .I(x[253]), .Q(
        xin[253]) );
  DFF \xreg_reg[255]  ( .D(xin[253]), .CLK(clk), .RST(start), .I(x[255]), .Q(
        xin[255]) );
  DFF \xreg_reg[257]  ( .D(xin[255]), .CLK(clk), .RST(start), .I(x[257]), .Q(
        xin[257]) );
  DFF \xreg_reg[259]  ( .D(xin[257]), .CLK(clk), .RST(start), .I(x[259]), .Q(
        xin[259]) );
  DFF \xreg_reg[261]  ( .D(xin[259]), .CLK(clk), .RST(start), .I(x[261]), .Q(
        xin[261]) );
  DFF \xreg_reg[263]  ( .D(xin[261]), .CLK(clk), .RST(start), .I(x[263]), .Q(
        xin[263]) );
  DFF \xreg_reg[265]  ( .D(xin[263]), .CLK(clk), .RST(start), .I(x[265]), .Q(
        xin[265]) );
  DFF \xreg_reg[267]  ( .D(xin[265]), .CLK(clk), .RST(start), .I(x[267]), .Q(
        xin[267]) );
  DFF \xreg_reg[269]  ( .D(xin[267]), .CLK(clk), .RST(start), .I(x[269]), .Q(
        xin[269]) );
  DFF \xreg_reg[271]  ( .D(xin[269]), .CLK(clk), .RST(start), .I(x[271]), .Q(
        xin[271]) );
  DFF \xreg_reg[273]  ( .D(xin[271]), .CLK(clk), .RST(start), .I(x[273]), .Q(
        xin[273]) );
  DFF \xreg_reg[275]  ( .D(xin[273]), .CLK(clk), .RST(start), .I(x[275]), .Q(
        xin[275]) );
  DFF \xreg_reg[277]  ( .D(xin[275]), .CLK(clk), .RST(start), .I(x[277]), .Q(
        xin[277]) );
  DFF \xreg_reg[279]  ( .D(xin[277]), .CLK(clk), .RST(start), .I(x[279]), .Q(
        xin[279]) );
  DFF \xreg_reg[281]  ( .D(xin[279]), .CLK(clk), .RST(start), .I(x[281]), .Q(
        xin[281]) );
  DFF \xreg_reg[283]  ( .D(xin[281]), .CLK(clk), .RST(start), .I(x[283]), .Q(
        xin[283]) );
  DFF \xreg_reg[285]  ( .D(xin[283]), .CLK(clk), .RST(start), .I(x[285]), .Q(
        xin[285]) );
  DFF \xreg_reg[287]  ( .D(xin[285]), .CLK(clk), .RST(start), .I(x[287]), .Q(
        xin[287]) );
  DFF \xreg_reg[289]  ( .D(xin[287]), .CLK(clk), .RST(start), .I(x[289]), .Q(
        xin[289]) );
  DFF \xreg_reg[291]  ( .D(xin[289]), .CLK(clk), .RST(start), .I(x[291]), .Q(
        xin[291]) );
  DFF \xreg_reg[293]  ( .D(xin[291]), .CLK(clk), .RST(start), .I(x[293]), .Q(
        xin[293]) );
  DFF \xreg_reg[295]  ( .D(xin[293]), .CLK(clk), .RST(start), .I(x[295]), .Q(
        xin[295]) );
  DFF \xreg_reg[297]  ( .D(xin[295]), .CLK(clk), .RST(start), .I(x[297]), .Q(
        xin[297]) );
  DFF \xreg_reg[299]  ( .D(xin[297]), .CLK(clk), .RST(start), .I(x[299]), .Q(
        xin[299]) );
  DFF \xreg_reg[301]  ( .D(xin[299]), .CLK(clk), .RST(start), .I(x[301]), .Q(
        xin[301]) );
  DFF \xreg_reg[303]  ( .D(xin[301]), .CLK(clk), .RST(start), .I(x[303]), .Q(
        xin[303]) );
  DFF \xreg_reg[305]  ( .D(xin[303]), .CLK(clk), .RST(start), .I(x[305]), .Q(
        xin[305]) );
  DFF \xreg_reg[307]  ( .D(xin[305]), .CLK(clk), .RST(start), .I(x[307]), .Q(
        xin[307]) );
  DFF \xreg_reg[309]  ( .D(xin[307]), .CLK(clk), .RST(start), .I(x[309]), .Q(
        xin[309]) );
  DFF \xreg_reg[311]  ( .D(xin[309]), .CLK(clk), .RST(start), .I(x[311]), .Q(
        xin[311]) );
  DFF \xreg_reg[313]  ( .D(xin[311]), .CLK(clk), .RST(start), .I(x[313]), .Q(
        xin[313]) );
  DFF \xreg_reg[315]  ( .D(xin[313]), .CLK(clk), .RST(start), .I(x[315]), .Q(
        xin[315]) );
  DFF \xreg_reg[317]  ( .D(xin[315]), .CLK(clk), .RST(start), .I(x[317]), .Q(
        xin[317]) );
  DFF \xreg_reg[319]  ( .D(xin[317]), .CLK(clk), .RST(start), .I(x[319]), .Q(
        xin[319]) );
  DFF \xreg_reg[321]  ( .D(xin[319]), .CLK(clk), .RST(start), .I(x[321]), .Q(
        xin[321]) );
  DFF \xreg_reg[323]  ( .D(xin[321]), .CLK(clk), .RST(start), .I(x[323]), .Q(
        xin[323]) );
  DFF \xreg_reg[325]  ( .D(xin[323]), .CLK(clk), .RST(start), .I(x[325]), .Q(
        xin[325]) );
  DFF \xreg_reg[327]  ( .D(xin[325]), .CLK(clk), .RST(start), .I(x[327]), .Q(
        xin[327]) );
  DFF \xreg_reg[329]  ( .D(xin[327]), .CLK(clk), .RST(start), .I(x[329]), .Q(
        xin[329]) );
  DFF \xreg_reg[331]  ( .D(xin[329]), .CLK(clk), .RST(start), .I(x[331]), .Q(
        xin[331]) );
  DFF \xreg_reg[333]  ( .D(xin[331]), .CLK(clk), .RST(start), .I(x[333]), .Q(
        xin[333]) );
  DFF \xreg_reg[335]  ( .D(xin[333]), .CLK(clk), .RST(start), .I(x[335]), .Q(
        xin[335]) );
  DFF \xreg_reg[337]  ( .D(xin[335]), .CLK(clk), .RST(start), .I(x[337]), .Q(
        xin[337]) );
  DFF \xreg_reg[339]  ( .D(xin[337]), .CLK(clk), .RST(start), .I(x[339]), .Q(
        xin[339]) );
  DFF \xreg_reg[341]  ( .D(xin[339]), .CLK(clk), .RST(start), .I(x[341]), .Q(
        xin[341]) );
  DFF \xreg_reg[343]  ( .D(xin[341]), .CLK(clk), .RST(start), .I(x[343]), .Q(
        xin[343]) );
  DFF \xreg_reg[345]  ( .D(xin[343]), .CLK(clk), .RST(start), .I(x[345]), .Q(
        xin[345]) );
  DFF \xreg_reg[347]  ( .D(xin[345]), .CLK(clk), .RST(start), .I(x[347]), .Q(
        xin[347]) );
  DFF \xreg_reg[349]  ( .D(xin[347]), .CLK(clk), .RST(start), .I(x[349]), .Q(
        xin[349]) );
  DFF \xreg_reg[351]  ( .D(xin[349]), .CLK(clk), .RST(start), .I(x[351]), .Q(
        xin[351]) );
  DFF \xreg_reg[353]  ( .D(xin[351]), .CLK(clk), .RST(start), .I(x[353]), .Q(
        xin[353]) );
  DFF \xreg_reg[355]  ( .D(xin[353]), .CLK(clk), .RST(start), .I(x[355]), .Q(
        xin[355]) );
  DFF \xreg_reg[357]  ( .D(xin[355]), .CLK(clk), .RST(start), .I(x[357]), .Q(
        xin[357]) );
  DFF \xreg_reg[359]  ( .D(xin[357]), .CLK(clk), .RST(start), .I(x[359]), .Q(
        xin[359]) );
  DFF \xreg_reg[361]  ( .D(xin[359]), .CLK(clk), .RST(start), .I(x[361]), .Q(
        xin[361]) );
  DFF \xreg_reg[363]  ( .D(xin[361]), .CLK(clk), .RST(start), .I(x[363]), .Q(
        xin[363]) );
  DFF \xreg_reg[365]  ( .D(xin[363]), .CLK(clk), .RST(start), .I(x[365]), .Q(
        xin[365]) );
  DFF \xreg_reg[367]  ( .D(xin[365]), .CLK(clk), .RST(start), .I(x[367]), .Q(
        xin[367]) );
  DFF \xreg_reg[369]  ( .D(xin[367]), .CLK(clk), .RST(start), .I(x[369]), .Q(
        xin[369]) );
  DFF \xreg_reg[371]  ( .D(xin[369]), .CLK(clk), .RST(start), .I(x[371]), .Q(
        xin[371]) );
  DFF \xreg_reg[373]  ( .D(xin[371]), .CLK(clk), .RST(start), .I(x[373]), .Q(
        xin[373]) );
  DFF \xreg_reg[375]  ( .D(xin[373]), .CLK(clk), .RST(start), .I(x[375]), .Q(
        xin[375]) );
  DFF \xreg_reg[377]  ( .D(xin[375]), .CLK(clk), .RST(start), .I(x[377]), .Q(
        xin[377]) );
  DFF \xreg_reg[379]  ( .D(xin[377]), .CLK(clk), .RST(start), .I(x[379]), .Q(
        xin[379]) );
  DFF \xreg_reg[381]  ( .D(xin[379]), .CLK(clk), .RST(start), .I(x[381]), .Q(
        xin[381]) );
  DFF \xreg_reg[383]  ( .D(xin[381]), .CLK(clk), .RST(start), .I(x[383]), .Q(
        xin[383]) );
  DFF \xreg_reg[385]  ( .D(xin[383]), .CLK(clk), .RST(start), .I(x[385]), .Q(
        xin[385]) );
  DFF \xreg_reg[387]  ( .D(xin[385]), .CLK(clk), .RST(start), .I(x[387]), .Q(
        xin[387]) );
  DFF \xreg_reg[389]  ( .D(xin[387]), .CLK(clk), .RST(start), .I(x[389]), .Q(
        xin[389]) );
  DFF \xreg_reg[391]  ( .D(xin[389]), .CLK(clk), .RST(start), .I(x[391]), .Q(
        xin[391]) );
  DFF \xreg_reg[393]  ( .D(xin[391]), .CLK(clk), .RST(start), .I(x[393]), .Q(
        xin[393]) );
  DFF \xreg_reg[395]  ( .D(xin[393]), .CLK(clk), .RST(start), .I(x[395]), .Q(
        xin[395]) );
  DFF \xreg_reg[397]  ( .D(xin[395]), .CLK(clk), .RST(start), .I(x[397]), .Q(
        xin[397]) );
  DFF \xreg_reg[399]  ( .D(xin[397]), .CLK(clk), .RST(start), .I(x[399]), .Q(
        xin[399]) );
  DFF \xreg_reg[401]  ( .D(xin[399]), .CLK(clk), .RST(start), .I(x[401]), .Q(
        xin[401]) );
  DFF \xreg_reg[403]  ( .D(xin[401]), .CLK(clk), .RST(start), .I(x[403]), .Q(
        xin[403]) );
  DFF \xreg_reg[405]  ( .D(xin[403]), .CLK(clk), .RST(start), .I(x[405]), .Q(
        xin[405]) );
  DFF \xreg_reg[407]  ( .D(xin[405]), .CLK(clk), .RST(start), .I(x[407]), .Q(
        xin[407]) );
  DFF \xreg_reg[409]  ( .D(xin[407]), .CLK(clk), .RST(start), .I(x[409]), .Q(
        xin[409]) );
  DFF \xreg_reg[411]  ( .D(xin[409]), .CLK(clk), .RST(start), .I(x[411]), .Q(
        xin[411]) );
  DFF \xreg_reg[413]  ( .D(xin[411]), .CLK(clk), .RST(start), .I(x[413]), .Q(
        xin[413]) );
  DFF \xreg_reg[415]  ( .D(xin[413]), .CLK(clk), .RST(start), .I(x[415]), .Q(
        xin[415]) );
  DFF \xreg_reg[417]  ( .D(xin[415]), .CLK(clk), .RST(start), .I(x[417]), .Q(
        xin[417]) );
  DFF \xreg_reg[419]  ( .D(xin[417]), .CLK(clk), .RST(start), .I(x[419]), .Q(
        xin[419]) );
  DFF \xreg_reg[421]  ( .D(xin[419]), .CLK(clk), .RST(start), .I(x[421]), .Q(
        xin[421]) );
  DFF \xreg_reg[423]  ( .D(xin[421]), .CLK(clk), .RST(start), .I(x[423]), .Q(
        xin[423]) );
  DFF \xreg_reg[425]  ( .D(xin[423]), .CLK(clk), .RST(start), .I(x[425]), .Q(
        xin[425]) );
  DFF \xreg_reg[427]  ( .D(xin[425]), .CLK(clk), .RST(start), .I(x[427]), .Q(
        xin[427]) );
  DFF \xreg_reg[429]  ( .D(xin[427]), .CLK(clk), .RST(start), .I(x[429]), .Q(
        xin[429]) );
  DFF \xreg_reg[431]  ( .D(xin[429]), .CLK(clk), .RST(start), .I(x[431]), .Q(
        xin[431]) );
  DFF \xreg_reg[433]  ( .D(xin[431]), .CLK(clk), .RST(start), .I(x[433]), .Q(
        xin[433]) );
  DFF \xreg_reg[435]  ( .D(xin[433]), .CLK(clk), .RST(start), .I(x[435]), .Q(
        xin[435]) );
  DFF \xreg_reg[437]  ( .D(xin[435]), .CLK(clk), .RST(start), .I(x[437]), .Q(
        xin[437]) );
  DFF \xreg_reg[439]  ( .D(xin[437]), .CLK(clk), .RST(start), .I(x[439]), .Q(
        xin[439]) );
  DFF \xreg_reg[441]  ( .D(xin[439]), .CLK(clk), .RST(start), .I(x[441]), .Q(
        xin[441]) );
  DFF \xreg_reg[443]  ( .D(xin[441]), .CLK(clk), .RST(start), .I(x[443]), .Q(
        xin[443]) );
  DFF \xreg_reg[445]  ( .D(xin[443]), .CLK(clk), .RST(start), .I(x[445]), .Q(
        xin[445]) );
  DFF \xreg_reg[447]  ( .D(xin[445]), .CLK(clk), .RST(start), .I(x[447]), .Q(
        xin[447]) );
  DFF \xreg_reg[449]  ( .D(xin[447]), .CLK(clk), .RST(start), .I(x[449]), .Q(
        xin[449]) );
  DFF \xreg_reg[451]  ( .D(xin[449]), .CLK(clk), .RST(start), .I(x[451]), .Q(
        xin[451]) );
  DFF \xreg_reg[453]  ( .D(xin[451]), .CLK(clk), .RST(start), .I(x[453]), .Q(
        xin[453]) );
  DFF \xreg_reg[455]  ( .D(xin[453]), .CLK(clk), .RST(start), .I(x[455]), .Q(
        xin[455]) );
  DFF \xreg_reg[457]  ( .D(xin[455]), .CLK(clk), .RST(start), .I(x[457]), .Q(
        xin[457]) );
  DFF \xreg_reg[459]  ( .D(xin[457]), .CLK(clk), .RST(start), .I(x[459]), .Q(
        xin[459]) );
  DFF \xreg_reg[461]  ( .D(xin[459]), .CLK(clk), .RST(start), .I(x[461]), .Q(
        xin[461]) );
  DFF \xreg_reg[463]  ( .D(xin[461]), .CLK(clk), .RST(start), .I(x[463]), .Q(
        xin[463]) );
  DFF \xreg_reg[465]  ( .D(xin[463]), .CLK(clk), .RST(start), .I(x[465]), .Q(
        xin[465]) );
  DFF \xreg_reg[467]  ( .D(xin[465]), .CLK(clk), .RST(start), .I(x[467]), .Q(
        xin[467]) );
  DFF \xreg_reg[469]  ( .D(xin[467]), .CLK(clk), .RST(start), .I(x[469]), .Q(
        xin[469]) );
  DFF \xreg_reg[471]  ( .D(xin[469]), .CLK(clk), .RST(start), .I(x[471]), .Q(
        xin[471]) );
  DFF \xreg_reg[473]  ( .D(xin[471]), .CLK(clk), .RST(start), .I(x[473]), .Q(
        xin[473]) );
  DFF \xreg_reg[475]  ( .D(xin[473]), .CLK(clk), .RST(start), .I(x[475]), .Q(
        xin[475]) );
  DFF \xreg_reg[477]  ( .D(xin[475]), .CLK(clk), .RST(start), .I(x[477]), .Q(
        xin[477]) );
  DFF \xreg_reg[479]  ( .D(xin[477]), .CLK(clk), .RST(start), .I(x[479]), .Q(
        xin[479]) );
  DFF \xreg_reg[481]  ( .D(xin[479]), .CLK(clk), .RST(start), .I(x[481]), .Q(
        xin[481]) );
  DFF \xreg_reg[483]  ( .D(xin[481]), .CLK(clk), .RST(start), .I(x[483]), .Q(
        xin[483]) );
  DFF \xreg_reg[485]  ( .D(xin[483]), .CLK(clk), .RST(start), .I(x[485]), .Q(
        xin[485]) );
  DFF \xreg_reg[487]  ( .D(xin[485]), .CLK(clk), .RST(start), .I(x[487]), .Q(
        xin[487]) );
  DFF \xreg_reg[489]  ( .D(xin[487]), .CLK(clk), .RST(start), .I(x[489]), .Q(
        xin[489]) );
  DFF \xreg_reg[491]  ( .D(xin[489]), .CLK(clk), .RST(start), .I(x[491]), .Q(
        xin[491]) );
  DFF \xreg_reg[493]  ( .D(xin[491]), .CLK(clk), .RST(start), .I(x[493]), .Q(
        xin[493]) );
  DFF \xreg_reg[495]  ( .D(xin[493]), .CLK(clk), .RST(start), .I(x[495]), .Q(
        xin[495]) );
  DFF \xreg_reg[497]  ( .D(xin[495]), .CLK(clk), .RST(start), .I(x[497]), .Q(
        xin[497]) );
  DFF \xreg_reg[499]  ( .D(xin[497]), .CLK(clk), .RST(start), .I(x[499]), .Q(
        xin[499]) );
  DFF \xreg_reg[501]  ( .D(xin[499]), .CLK(clk), .RST(start), .I(x[501]), .Q(
        xin[501]) );
  DFF \xreg_reg[503]  ( .D(xin[501]), .CLK(clk), .RST(start), .I(x[503]), .Q(
        xin[503]) );
  DFF \xreg_reg[505]  ( .D(xin[503]), .CLK(clk), .RST(start), .I(x[505]), .Q(
        xin[505]) );
  DFF \xreg_reg[507]  ( .D(xin[505]), .CLK(clk), .RST(start), .I(x[507]), .Q(
        xin[507]) );
  DFF \xreg_reg[509]  ( .D(xin[507]), .CLK(clk), .RST(start), .I(x[509]), .Q(
        xin[509]) );
  DFF \xreg_reg[511]  ( .D(xin[509]), .CLK(clk), .RST(start), .I(x[511]), .Q(
        xin[511]) );
  DFF \xreg_reg[0]  ( .D(1'b0), .CLK(clk), .RST(start), .I(x[0]), .Q(xin[0])
         );
  DFF \xreg_reg[2]  ( .D(xin[0]), .CLK(clk), .RST(start), .I(x[2]), .Q(xin[2])
         );
  DFF \xreg_reg[4]  ( .D(xin[2]), .CLK(clk), .RST(start), .I(x[4]), .Q(xin[4])
         );
  DFF \xreg_reg[6]  ( .D(xin[4]), .CLK(clk), .RST(start), .I(x[6]), .Q(xin[6])
         );
  DFF \xreg_reg[8]  ( .D(xin[6]), .CLK(clk), .RST(start), .I(x[8]), .Q(xin[8])
         );
  DFF \xreg_reg[10]  ( .D(xin[8]), .CLK(clk), .RST(start), .I(x[10]), .Q(
        xin[10]) );
  DFF \xreg_reg[12]  ( .D(xin[10]), .CLK(clk), .RST(start), .I(x[12]), .Q(
        xin[12]) );
  DFF \xreg_reg[14]  ( .D(xin[12]), .CLK(clk), .RST(start), .I(x[14]), .Q(
        xin[14]) );
  DFF \xreg_reg[16]  ( .D(xin[14]), .CLK(clk), .RST(start), .I(x[16]), .Q(
        xin[16]) );
  DFF \xreg_reg[18]  ( .D(xin[16]), .CLK(clk), .RST(start), .I(x[18]), .Q(
        xin[18]) );
  DFF \xreg_reg[20]  ( .D(xin[18]), .CLK(clk), .RST(start), .I(x[20]), .Q(
        xin[20]) );
  DFF \xreg_reg[22]  ( .D(xin[20]), .CLK(clk), .RST(start), .I(x[22]), .Q(
        xin[22]) );
  DFF \xreg_reg[24]  ( .D(xin[22]), .CLK(clk), .RST(start), .I(x[24]), .Q(
        xin[24]) );
  DFF \xreg_reg[26]  ( .D(xin[24]), .CLK(clk), .RST(start), .I(x[26]), .Q(
        xin[26]) );
  DFF \xreg_reg[28]  ( .D(xin[26]), .CLK(clk), .RST(start), .I(x[28]), .Q(
        xin[28]) );
  DFF \xreg_reg[30]  ( .D(xin[28]), .CLK(clk), .RST(start), .I(x[30]), .Q(
        xin[30]) );
  DFF \xreg_reg[32]  ( .D(xin[30]), .CLK(clk), .RST(start), .I(x[32]), .Q(
        xin[32]) );
  DFF \xreg_reg[34]  ( .D(xin[32]), .CLK(clk), .RST(start), .I(x[34]), .Q(
        xin[34]) );
  DFF \xreg_reg[36]  ( .D(xin[34]), .CLK(clk), .RST(start), .I(x[36]), .Q(
        xin[36]) );
  DFF \xreg_reg[38]  ( .D(xin[36]), .CLK(clk), .RST(start), .I(x[38]), .Q(
        xin[38]) );
  DFF \xreg_reg[40]  ( .D(xin[38]), .CLK(clk), .RST(start), .I(x[40]), .Q(
        xin[40]) );
  DFF \xreg_reg[42]  ( .D(xin[40]), .CLK(clk), .RST(start), .I(x[42]), .Q(
        xin[42]) );
  DFF \xreg_reg[44]  ( .D(xin[42]), .CLK(clk), .RST(start), .I(x[44]), .Q(
        xin[44]) );
  DFF \xreg_reg[46]  ( .D(xin[44]), .CLK(clk), .RST(start), .I(x[46]), .Q(
        xin[46]) );
  DFF \xreg_reg[48]  ( .D(xin[46]), .CLK(clk), .RST(start), .I(x[48]), .Q(
        xin[48]) );
  DFF \xreg_reg[50]  ( .D(xin[48]), .CLK(clk), .RST(start), .I(x[50]), .Q(
        xin[50]) );
  DFF \xreg_reg[52]  ( .D(xin[50]), .CLK(clk), .RST(start), .I(x[52]), .Q(
        xin[52]) );
  DFF \xreg_reg[54]  ( .D(xin[52]), .CLK(clk), .RST(start), .I(x[54]), .Q(
        xin[54]) );
  DFF \xreg_reg[56]  ( .D(xin[54]), .CLK(clk), .RST(start), .I(x[56]), .Q(
        xin[56]) );
  DFF \xreg_reg[58]  ( .D(xin[56]), .CLK(clk), .RST(start), .I(x[58]), .Q(
        xin[58]) );
  DFF \xreg_reg[60]  ( .D(xin[58]), .CLK(clk), .RST(start), .I(x[60]), .Q(
        xin[60]) );
  DFF \xreg_reg[62]  ( .D(xin[60]), .CLK(clk), .RST(start), .I(x[62]), .Q(
        xin[62]) );
  DFF \xreg_reg[64]  ( .D(xin[62]), .CLK(clk), .RST(start), .I(x[64]), .Q(
        xin[64]) );
  DFF \xreg_reg[66]  ( .D(xin[64]), .CLK(clk), .RST(start), .I(x[66]), .Q(
        xin[66]) );
  DFF \xreg_reg[68]  ( .D(xin[66]), .CLK(clk), .RST(start), .I(x[68]), .Q(
        xin[68]) );
  DFF \xreg_reg[70]  ( .D(xin[68]), .CLK(clk), .RST(start), .I(x[70]), .Q(
        xin[70]) );
  DFF \xreg_reg[72]  ( .D(xin[70]), .CLK(clk), .RST(start), .I(x[72]), .Q(
        xin[72]) );
  DFF \xreg_reg[74]  ( .D(xin[72]), .CLK(clk), .RST(start), .I(x[74]), .Q(
        xin[74]) );
  DFF \xreg_reg[76]  ( .D(xin[74]), .CLK(clk), .RST(start), .I(x[76]), .Q(
        xin[76]) );
  DFF \xreg_reg[78]  ( .D(xin[76]), .CLK(clk), .RST(start), .I(x[78]), .Q(
        xin[78]) );
  DFF \xreg_reg[80]  ( .D(xin[78]), .CLK(clk), .RST(start), .I(x[80]), .Q(
        xin[80]) );
  DFF \xreg_reg[82]  ( .D(xin[80]), .CLK(clk), .RST(start), .I(x[82]), .Q(
        xin[82]) );
  DFF \xreg_reg[84]  ( .D(xin[82]), .CLK(clk), .RST(start), .I(x[84]), .Q(
        xin[84]) );
  DFF \xreg_reg[86]  ( .D(xin[84]), .CLK(clk), .RST(start), .I(x[86]), .Q(
        xin[86]) );
  DFF \xreg_reg[88]  ( .D(xin[86]), .CLK(clk), .RST(start), .I(x[88]), .Q(
        xin[88]) );
  DFF \xreg_reg[90]  ( .D(xin[88]), .CLK(clk), .RST(start), .I(x[90]), .Q(
        xin[90]) );
  DFF \xreg_reg[92]  ( .D(xin[90]), .CLK(clk), .RST(start), .I(x[92]), .Q(
        xin[92]) );
  DFF \xreg_reg[94]  ( .D(xin[92]), .CLK(clk), .RST(start), .I(x[94]), .Q(
        xin[94]) );
  DFF \xreg_reg[96]  ( .D(xin[94]), .CLK(clk), .RST(start), .I(x[96]), .Q(
        xin[96]) );
  DFF \xreg_reg[98]  ( .D(xin[96]), .CLK(clk), .RST(start), .I(x[98]), .Q(
        xin[98]) );
  DFF \xreg_reg[100]  ( .D(xin[98]), .CLK(clk), .RST(start), .I(x[100]), .Q(
        xin[100]) );
  DFF \xreg_reg[102]  ( .D(xin[100]), .CLK(clk), .RST(start), .I(x[102]), .Q(
        xin[102]) );
  DFF \xreg_reg[104]  ( .D(xin[102]), .CLK(clk), .RST(start), .I(x[104]), .Q(
        xin[104]) );
  DFF \xreg_reg[106]  ( .D(xin[104]), .CLK(clk), .RST(start), .I(x[106]), .Q(
        xin[106]) );
  DFF \xreg_reg[108]  ( .D(xin[106]), .CLK(clk), .RST(start), .I(x[108]), .Q(
        xin[108]) );
  DFF \xreg_reg[110]  ( .D(xin[108]), .CLK(clk), .RST(start), .I(x[110]), .Q(
        xin[110]) );
  DFF \xreg_reg[112]  ( .D(xin[110]), .CLK(clk), .RST(start), .I(x[112]), .Q(
        xin[112]) );
  DFF \xreg_reg[114]  ( .D(xin[112]), .CLK(clk), .RST(start), .I(x[114]), .Q(
        xin[114]) );
  DFF \xreg_reg[116]  ( .D(xin[114]), .CLK(clk), .RST(start), .I(x[116]), .Q(
        xin[116]) );
  DFF \xreg_reg[118]  ( .D(xin[116]), .CLK(clk), .RST(start), .I(x[118]), .Q(
        xin[118]) );
  DFF \xreg_reg[120]  ( .D(xin[118]), .CLK(clk), .RST(start), .I(x[120]), .Q(
        xin[120]) );
  DFF \xreg_reg[122]  ( .D(xin[120]), .CLK(clk), .RST(start), .I(x[122]), .Q(
        xin[122]) );
  DFF \xreg_reg[124]  ( .D(xin[122]), .CLK(clk), .RST(start), .I(x[124]), .Q(
        xin[124]) );
  DFF \xreg_reg[126]  ( .D(xin[124]), .CLK(clk), .RST(start), .I(x[126]), .Q(
        xin[126]) );
  DFF \xreg_reg[128]  ( .D(xin[126]), .CLK(clk), .RST(start), .I(x[128]), .Q(
        xin[128]) );
  DFF \xreg_reg[130]  ( .D(xin[128]), .CLK(clk), .RST(start), .I(x[130]), .Q(
        xin[130]) );
  DFF \xreg_reg[132]  ( .D(xin[130]), .CLK(clk), .RST(start), .I(x[132]), .Q(
        xin[132]) );
  DFF \xreg_reg[134]  ( .D(xin[132]), .CLK(clk), .RST(start), .I(x[134]), .Q(
        xin[134]) );
  DFF \xreg_reg[136]  ( .D(xin[134]), .CLK(clk), .RST(start), .I(x[136]), .Q(
        xin[136]) );
  DFF \xreg_reg[138]  ( .D(xin[136]), .CLK(clk), .RST(start), .I(x[138]), .Q(
        xin[138]) );
  DFF \xreg_reg[140]  ( .D(xin[138]), .CLK(clk), .RST(start), .I(x[140]), .Q(
        xin[140]) );
  DFF \xreg_reg[142]  ( .D(xin[140]), .CLK(clk), .RST(start), .I(x[142]), .Q(
        xin[142]) );
  DFF \xreg_reg[144]  ( .D(xin[142]), .CLK(clk), .RST(start), .I(x[144]), .Q(
        xin[144]) );
  DFF \xreg_reg[146]  ( .D(xin[144]), .CLK(clk), .RST(start), .I(x[146]), .Q(
        xin[146]) );
  DFF \xreg_reg[148]  ( .D(xin[146]), .CLK(clk), .RST(start), .I(x[148]), .Q(
        xin[148]) );
  DFF \xreg_reg[150]  ( .D(xin[148]), .CLK(clk), .RST(start), .I(x[150]), .Q(
        xin[150]) );
  DFF \xreg_reg[152]  ( .D(xin[150]), .CLK(clk), .RST(start), .I(x[152]), .Q(
        xin[152]) );
  DFF \xreg_reg[154]  ( .D(xin[152]), .CLK(clk), .RST(start), .I(x[154]), .Q(
        xin[154]) );
  DFF \xreg_reg[156]  ( .D(xin[154]), .CLK(clk), .RST(start), .I(x[156]), .Q(
        xin[156]) );
  DFF \xreg_reg[158]  ( .D(xin[156]), .CLK(clk), .RST(start), .I(x[158]), .Q(
        xin[158]) );
  DFF \xreg_reg[160]  ( .D(xin[158]), .CLK(clk), .RST(start), .I(x[160]), .Q(
        xin[160]) );
  DFF \xreg_reg[162]  ( .D(xin[160]), .CLK(clk), .RST(start), .I(x[162]), .Q(
        xin[162]) );
  DFF \xreg_reg[164]  ( .D(xin[162]), .CLK(clk), .RST(start), .I(x[164]), .Q(
        xin[164]) );
  DFF \xreg_reg[166]  ( .D(xin[164]), .CLK(clk), .RST(start), .I(x[166]), .Q(
        xin[166]) );
  DFF \xreg_reg[168]  ( .D(xin[166]), .CLK(clk), .RST(start), .I(x[168]), .Q(
        xin[168]) );
  DFF \xreg_reg[170]  ( .D(xin[168]), .CLK(clk), .RST(start), .I(x[170]), .Q(
        xin[170]) );
  DFF \xreg_reg[172]  ( .D(xin[170]), .CLK(clk), .RST(start), .I(x[172]), .Q(
        xin[172]) );
  DFF \xreg_reg[174]  ( .D(xin[172]), .CLK(clk), .RST(start), .I(x[174]), .Q(
        xin[174]) );
  DFF \xreg_reg[176]  ( .D(xin[174]), .CLK(clk), .RST(start), .I(x[176]), .Q(
        xin[176]) );
  DFF \xreg_reg[178]  ( .D(xin[176]), .CLK(clk), .RST(start), .I(x[178]), .Q(
        xin[178]) );
  DFF \xreg_reg[180]  ( .D(xin[178]), .CLK(clk), .RST(start), .I(x[180]), .Q(
        xin[180]) );
  DFF \xreg_reg[182]  ( .D(xin[180]), .CLK(clk), .RST(start), .I(x[182]), .Q(
        xin[182]) );
  DFF \xreg_reg[184]  ( .D(xin[182]), .CLK(clk), .RST(start), .I(x[184]), .Q(
        xin[184]) );
  DFF \xreg_reg[186]  ( .D(xin[184]), .CLK(clk), .RST(start), .I(x[186]), .Q(
        xin[186]) );
  DFF \xreg_reg[188]  ( .D(xin[186]), .CLK(clk), .RST(start), .I(x[188]), .Q(
        xin[188]) );
  DFF \xreg_reg[190]  ( .D(xin[188]), .CLK(clk), .RST(start), .I(x[190]), .Q(
        xin[190]) );
  DFF \xreg_reg[192]  ( .D(xin[190]), .CLK(clk), .RST(start), .I(x[192]), .Q(
        xin[192]) );
  DFF \xreg_reg[194]  ( .D(xin[192]), .CLK(clk), .RST(start), .I(x[194]), .Q(
        xin[194]) );
  DFF \xreg_reg[196]  ( .D(xin[194]), .CLK(clk), .RST(start), .I(x[196]), .Q(
        xin[196]) );
  DFF \xreg_reg[198]  ( .D(xin[196]), .CLK(clk), .RST(start), .I(x[198]), .Q(
        xin[198]) );
  DFF \xreg_reg[200]  ( .D(xin[198]), .CLK(clk), .RST(start), .I(x[200]), .Q(
        xin[200]) );
  DFF \xreg_reg[202]  ( .D(xin[200]), .CLK(clk), .RST(start), .I(x[202]), .Q(
        xin[202]) );
  DFF \xreg_reg[204]  ( .D(xin[202]), .CLK(clk), .RST(start), .I(x[204]), .Q(
        xin[204]) );
  DFF \xreg_reg[206]  ( .D(xin[204]), .CLK(clk), .RST(start), .I(x[206]), .Q(
        xin[206]) );
  DFF \xreg_reg[208]  ( .D(xin[206]), .CLK(clk), .RST(start), .I(x[208]), .Q(
        xin[208]) );
  DFF \xreg_reg[210]  ( .D(xin[208]), .CLK(clk), .RST(start), .I(x[210]), .Q(
        xin[210]) );
  DFF \xreg_reg[212]  ( .D(xin[210]), .CLK(clk), .RST(start), .I(x[212]), .Q(
        xin[212]) );
  DFF \xreg_reg[214]  ( .D(xin[212]), .CLK(clk), .RST(start), .I(x[214]), .Q(
        xin[214]) );
  DFF \xreg_reg[216]  ( .D(xin[214]), .CLK(clk), .RST(start), .I(x[216]), .Q(
        xin[216]) );
  DFF \xreg_reg[218]  ( .D(xin[216]), .CLK(clk), .RST(start), .I(x[218]), .Q(
        xin[218]) );
  DFF \xreg_reg[220]  ( .D(xin[218]), .CLK(clk), .RST(start), .I(x[220]), .Q(
        xin[220]) );
  DFF \xreg_reg[222]  ( .D(xin[220]), .CLK(clk), .RST(start), .I(x[222]), .Q(
        xin[222]) );
  DFF \xreg_reg[224]  ( .D(xin[222]), .CLK(clk), .RST(start), .I(x[224]), .Q(
        xin[224]) );
  DFF \xreg_reg[226]  ( .D(xin[224]), .CLK(clk), .RST(start), .I(x[226]), .Q(
        xin[226]) );
  DFF \xreg_reg[228]  ( .D(xin[226]), .CLK(clk), .RST(start), .I(x[228]), .Q(
        xin[228]) );
  DFF \xreg_reg[230]  ( .D(xin[228]), .CLK(clk), .RST(start), .I(x[230]), .Q(
        xin[230]) );
  DFF \xreg_reg[232]  ( .D(xin[230]), .CLK(clk), .RST(start), .I(x[232]), .Q(
        xin[232]) );
  DFF \xreg_reg[234]  ( .D(xin[232]), .CLK(clk), .RST(start), .I(x[234]), .Q(
        xin[234]) );
  DFF \xreg_reg[236]  ( .D(xin[234]), .CLK(clk), .RST(start), .I(x[236]), .Q(
        xin[236]) );
  DFF \xreg_reg[238]  ( .D(xin[236]), .CLK(clk), .RST(start), .I(x[238]), .Q(
        xin[238]) );
  DFF \xreg_reg[240]  ( .D(xin[238]), .CLK(clk), .RST(start), .I(x[240]), .Q(
        xin[240]) );
  DFF \xreg_reg[242]  ( .D(xin[240]), .CLK(clk), .RST(start), .I(x[242]), .Q(
        xin[242]) );
  DFF \xreg_reg[244]  ( .D(xin[242]), .CLK(clk), .RST(start), .I(x[244]), .Q(
        xin[244]) );
  DFF \xreg_reg[246]  ( .D(xin[244]), .CLK(clk), .RST(start), .I(x[246]), .Q(
        xin[246]) );
  DFF \xreg_reg[248]  ( .D(xin[246]), .CLK(clk), .RST(start), .I(x[248]), .Q(
        xin[248]) );
  DFF \xreg_reg[250]  ( .D(xin[248]), .CLK(clk), .RST(start), .I(x[250]), .Q(
        xin[250]) );
  DFF \xreg_reg[252]  ( .D(xin[250]), .CLK(clk), .RST(start), .I(x[252]), .Q(
        xin[252]) );
  DFF \xreg_reg[254]  ( .D(xin[252]), .CLK(clk), .RST(start), .I(x[254]), .Q(
        xin[254]) );
  DFF \xreg_reg[256]  ( .D(xin[254]), .CLK(clk), .RST(start), .I(x[256]), .Q(
        xin[256]) );
  DFF \xreg_reg[258]  ( .D(xin[256]), .CLK(clk), .RST(start), .I(x[258]), .Q(
        xin[258]) );
  DFF \xreg_reg[260]  ( .D(xin[258]), .CLK(clk), .RST(start), .I(x[260]), .Q(
        xin[260]) );
  DFF \xreg_reg[262]  ( .D(xin[260]), .CLK(clk), .RST(start), .I(x[262]), .Q(
        xin[262]) );
  DFF \xreg_reg[264]  ( .D(xin[262]), .CLK(clk), .RST(start), .I(x[264]), .Q(
        xin[264]) );
  DFF \xreg_reg[266]  ( .D(xin[264]), .CLK(clk), .RST(start), .I(x[266]), .Q(
        xin[266]) );
  DFF \xreg_reg[268]  ( .D(xin[266]), .CLK(clk), .RST(start), .I(x[268]), .Q(
        xin[268]) );
  DFF \xreg_reg[270]  ( .D(xin[268]), .CLK(clk), .RST(start), .I(x[270]), .Q(
        xin[270]) );
  DFF \xreg_reg[272]  ( .D(xin[270]), .CLK(clk), .RST(start), .I(x[272]), .Q(
        xin[272]) );
  DFF \xreg_reg[274]  ( .D(xin[272]), .CLK(clk), .RST(start), .I(x[274]), .Q(
        xin[274]) );
  DFF \xreg_reg[276]  ( .D(xin[274]), .CLK(clk), .RST(start), .I(x[276]), .Q(
        xin[276]) );
  DFF \xreg_reg[278]  ( .D(xin[276]), .CLK(clk), .RST(start), .I(x[278]), .Q(
        xin[278]) );
  DFF \xreg_reg[280]  ( .D(xin[278]), .CLK(clk), .RST(start), .I(x[280]), .Q(
        xin[280]) );
  DFF \xreg_reg[282]  ( .D(xin[280]), .CLK(clk), .RST(start), .I(x[282]), .Q(
        xin[282]) );
  DFF \xreg_reg[284]  ( .D(xin[282]), .CLK(clk), .RST(start), .I(x[284]), .Q(
        xin[284]) );
  DFF \xreg_reg[286]  ( .D(xin[284]), .CLK(clk), .RST(start), .I(x[286]), .Q(
        xin[286]) );
  DFF \xreg_reg[288]  ( .D(xin[286]), .CLK(clk), .RST(start), .I(x[288]), .Q(
        xin[288]) );
  DFF \xreg_reg[290]  ( .D(xin[288]), .CLK(clk), .RST(start), .I(x[290]), .Q(
        xin[290]) );
  DFF \xreg_reg[292]  ( .D(xin[290]), .CLK(clk), .RST(start), .I(x[292]), .Q(
        xin[292]) );
  DFF \xreg_reg[294]  ( .D(xin[292]), .CLK(clk), .RST(start), .I(x[294]), .Q(
        xin[294]) );
  DFF \xreg_reg[296]  ( .D(xin[294]), .CLK(clk), .RST(start), .I(x[296]), .Q(
        xin[296]) );
  DFF \xreg_reg[298]  ( .D(xin[296]), .CLK(clk), .RST(start), .I(x[298]), .Q(
        xin[298]) );
  DFF \xreg_reg[300]  ( .D(xin[298]), .CLK(clk), .RST(start), .I(x[300]), .Q(
        xin[300]) );
  DFF \xreg_reg[302]  ( .D(xin[300]), .CLK(clk), .RST(start), .I(x[302]), .Q(
        xin[302]) );
  DFF \xreg_reg[304]  ( .D(xin[302]), .CLK(clk), .RST(start), .I(x[304]), .Q(
        xin[304]) );
  DFF \xreg_reg[306]  ( .D(xin[304]), .CLK(clk), .RST(start), .I(x[306]), .Q(
        xin[306]) );
  DFF \xreg_reg[308]  ( .D(xin[306]), .CLK(clk), .RST(start), .I(x[308]), .Q(
        xin[308]) );
  DFF \xreg_reg[310]  ( .D(xin[308]), .CLK(clk), .RST(start), .I(x[310]), .Q(
        xin[310]) );
  DFF \xreg_reg[312]  ( .D(xin[310]), .CLK(clk), .RST(start), .I(x[312]), .Q(
        xin[312]) );
  DFF \xreg_reg[314]  ( .D(xin[312]), .CLK(clk), .RST(start), .I(x[314]), .Q(
        xin[314]) );
  DFF \xreg_reg[316]  ( .D(xin[314]), .CLK(clk), .RST(start), .I(x[316]), .Q(
        xin[316]) );
  DFF \xreg_reg[318]  ( .D(xin[316]), .CLK(clk), .RST(start), .I(x[318]), .Q(
        xin[318]) );
  DFF \xreg_reg[320]  ( .D(xin[318]), .CLK(clk), .RST(start), .I(x[320]), .Q(
        xin[320]) );
  DFF \xreg_reg[322]  ( .D(xin[320]), .CLK(clk), .RST(start), .I(x[322]), .Q(
        xin[322]) );
  DFF \xreg_reg[324]  ( .D(xin[322]), .CLK(clk), .RST(start), .I(x[324]), .Q(
        xin[324]) );
  DFF \xreg_reg[326]  ( .D(xin[324]), .CLK(clk), .RST(start), .I(x[326]), .Q(
        xin[326]) );
  DFF \xreg_reg[328]  ( .D(xin[326]), .CLK(clk), .RST(start), .I(x[328]), .Q(
        xin[328]) );
  DFF \xreg_reg[330]  ( .D(xin[328]), .CLK(clk), .RST(start), .I(x[330]), .Q(
        xin[330]) );
  DFF \xreg_reg[332]  ( .D(xin[330]), .CLK(clk), .RST(start), .I(x[332]), .Q(
        xin[332]) );
  DFF \xreg_reg[334]  ( .D(xin[332]), .CLK(clk), .RST(start), .I(x[334]), .Q(
        xin[334]) );
  DFF \xreg_reg[336]  ( .D(xin[334]), .CLK(clk), .RST(start), .I(x[336]), .Q(
        xin[336]) );
  DFF \xreg_reg[338]  ( .D(xin[336]), .CLK(clk), .RST(start), .I(x[338]), .Q(
        xin[338]) );
  DFF \xreg_reg[340]  ( .D(xin[338]), .CLK(clk), .RST(start), .I(x[340]), .Q(
        xin[340]) );
  DFF \xreg_reg[342]  ( .D(xin[340]), .CLK(clk), .RST(start), .I(x[342]), .Q(
        xin[342]) );
  DFF \xreg_reg[344]  ( .D(xin[342]), .CLK(clk), .RST(start), .I(x[344]), .Q(
        xin[344]) );
  DFF \xreg_reg[346]  ( .D(xin[344]), .CLK(clk), .RST(start), .I(x[346]), .Q(
        xin[346]) );
  DFF \xreg_reg[348]  ( .D(xin[346]), .CLK(clk), .RST(start), .I(x[348]), .Q(
        xin[348]) );
  DFF \xreg_reg[350]  ( .D(xin[348]), .CLK(clk), .RST(start), .I(x[350]), .Q(
        xin[350]) );
  DFF \xreg_reg[352]  ( .D(xin[350]), .CLK(clk), .RST(start), .I(x[352]), .Q(
        xin[352]) );
  DFF \xreg_reg[354]  ( .D(xin[352]), .CLK(clk), .RST(start), .I(x[354]), .Q(
        xin[354]) );
  DFF \xreg_reg[356]  ( .D(xin[354]), .CLK(clk), .RST(start), .I(x[356]), .Q(
        xin[356]) );
  DFF \xreg_reg[358]  ( .D(xin[356]), .CLK(clk), .RST(start), .I(x[358]), .Q(
        xin[358]) );
  DFF \xreg_reg[360]  ( .D(xin[358]), .CLK(clk), .RST(start), .I(x[360]), .Q(
        xin[360]) );
  DFF \xreg_reg[362]  ( .D(xin[360]), .CLK(clk), .RST(start), .I(x[362]), .Q(
        xin[362]) );
  DFF \xreg_reg[364]  ( .D(xin[362]), .CLK(clk), .RST(start), .I(x[364]), .Q(
        xin[364]) );
  DFF \xreg_reg[366]  ( .D(xin[364]), .CLK(clk), .RST(start), .I(x[366]), .Q(
        xin[366]) );
  DFF \xreg_reg[368]  ( .D(xin[366]), .CLK(clk), .RST(start), .I(x[368]), .Q(
        xin[368]) );
  DFF \xreg_reg[370]  ( .D(xin[368]), .CLK(clk), .RST(start), .I(x[370]), .Q(
        xin[370]) );
  DFF \xreg_reg[372]  ( .D(xin[370]), .CLK(clk), .RST(start), .I(x[372]), .Q(
        xin[372]) );
  DFF \xreg_reg[374]  ( .D(xin[372]), .CLK(clk), .RST(start), .I(x[374]), .Q(
        xin[374]) );
  DFF \xreg_reg[376]  ( .D(xin[374]), .CLK(clk), .RST(start), .I(x[376]), .Q(
        xin[376]) );
  DFF \xreg_reg[378]  ( .D(xin[376]), .CLK(clk), .RST(start), .I(x[378]), .Q(
        xin[378]) );
  DFF \xreg_reg[380]  ( .D(xin[378]), .CLK(clk), .RST(start), .I(x[380]), .Q(
        xin[380]) );
  DFF \xreg_reg[382]  ( .D(xin[380]), .CLK(clk), .RST(start), .I(x[382]), .Q(
        xin[382]) );
  DFF \xreg_reg[384]  ( .D(xin[382]), .CLK(clk), .RST(start), .I(x[384]), .Q(
        xin[384]) );
  DFF \xreg_reg[386]  ( .D(xin[384]), .CLK(clk), .RST(start), .I(x[386]), .Q(
        xin[386]) );
  DFF \xreg_reg[388]  ( .D(xin[386]), .CLK(clk), .RST(start), .I(x[388]), .Q(
        xin[388]) );
  DFF \xreg_reg[390]  ( .D(xin[388]), .CLK(clk), .RST(start), .I(x[390]), .Q(
        xin[390]) );
  DFF \xreg_reg[392]  ( .D(xin[390]), .CLK(clk), .RST(start), .I(x[392]), .Q(
        xin[392]) );
  DFF \xreg_reg[394]  ( .D(xin[392]), .CLK(clk), .RST(start), .I(x[394]), .Q(
        xin[394]) );
  DFF \xreg_reg[396]  ( .D(xin[394]), .CLK(clk), .RST(start), .I(x[396]), .Q(
        xin[396]) );
  DFF \xreg_reg[398]  ( .D(xin[396]), .CLK(clk), .RST(start), .I(x[398]), .Q(
        xin[398]) );
  DFF \xreg_reg[400]  ( .D(xin[398]), .CLK(clk), .RST(start), .I(x[400]), .Q(
        xin[400]) );
  DFF \xreg_reg[402]  ( .D(xin[400]), .CLK(clk), .RST(start), .I(x[402]), .Q(
        xin[402]) );
  DFF \xreg_reg[404]  ( .D(xin[402]), .CLK(clk), .RST(start), .I(x[404]), .Q(
        xin[404]) );
  DFF \xreg_reg[406]  ( .D(xin[404]), .CLK(clk), .RST(start), .I(x[406]), .Q(
        xin[406]) );
  DFF \xreg_reg[408]  ( .D(xin[406]), .CLK(clk), .RST(start), .I(x[408]), .Q(
        xin[408]) );
  DFF \xreg_reg[410]  ( .D(xin[408]), .CLK(clk), .RST(start), .I(x[410]), .Q(
        xin[410]) );
  DFF \xreg_reg[412]  ( .D(xin[410]), .CLK(clk), .RST(start), .I(x[412]), .Q(
        xin[412]) );
  DFF \xreg_reg[414]  ( .D(xin[412]), .CLK(clk), .RST(start), .I(x[414]), .Q(
        xin[414]) );
  DFF \xreg_reg[416]  ( .D(xin[414]), .CLK(clk), .RST(start), .I(x[416]), .Q(
        xin[416]) );
  DFF \xreg_reg[418]  ( .D(xin[416]), .CLK(clk), .RST(start), .I(x[418]), .Q(
        xin[418]) );
  DFF \xreg_reg[420]  ( .D(xin[418]), .CLK(clk), .RST(start), .I(x[420]), .Q(
        xin[420]) );
  DFF \xreg_reg[422]  ( .D(xin[420]), .CLK(clk), .RST(start), .I(x[422]), .Q(
        xin[422]) );
  DFF \xreg_reg[424]  ( .D(xin[422]), .CLK(clk), .RST(start), .I(x[424]), .Q(
        xin[424]) );
  DFF \xreg_reg[426]  ( .D(xin[424]), .CLK(clk), .RST(start), .I(x[426]), .Q(
        xin[426]) );
  DFF \xreg_reg[428]  ( .D(xin[426]), .CLK(clk), .RST(start), .I(x[428]), .Q(
        xin[428]) );
  DFF \xreg_reg[430]  ( .D(xin[428]), .CLK(clk), .RST(start), .I(x[430]), .Q(
        xin[430]) );
  DFF \xreg_reg[432]  ( .D(xin[430]), .CLK(clk), .RST(start), .I(x[432]), .Q(
        xin[432]) );
  DFF \xreg_reg[434]  ( .D(xin[432]), .CLK(clk), .RST(start), .I(x[434]), .Q(
        xin[434]) );
  DFF \xreg_reg[436]  ( .D(xin[434]), .CLK(clk), .RST(start), .I(x[436]), .Q(
        xin[436]) );
  DFF \xreg_reg[438]  ( .D(xin[436]), .CLK(clk), .RST(start), .I(x[438]), .Q(
        xin[438]) );
  DFF \xreg_reg[440]  ( .D(xin[438]), .CLK(clk), .RST(start), .I(x[440]), .Q(
        xin[440]) );
  DFF \xreg_reg[442]  ( .D(xin[440]), .CLK(clk), .RST(start), .I(x[442]), .Q(
        xin[442]) );
  DFF \xreg_reg[444]  ( .D(xin[442]), .CLK(clk), .RST(start), .I(x[444]), .Q(
        xin[444]) );
  DFF \xreg_reg[446]  ( .D(xin[444]), .CLK(clk), .RST(start), .I(x[446]), .Q(
        xin[446]) );
  DFF \xreg_reg[448]  ( .D(xin[446]), .CLK(clk), .RST(start), .I(x[448]), .Q(
        xin[448]) );
  DFF \xreg_reg[450]  ( .D(xin[448]), .CLK(clk), .RST(start), .I(x[450]), .Q(
        xin[450]) );
  DFF \xreg_reg[452]  ( .D(xin[450]), .CLK(clk), .RST(start), .I(x[452]), .Q(
        xin[452]) );
  DFF \xreg_reg[454]  ( .D(xin[452]), .CLK(clk), .RST(start), .I(x[454]), .Q(
        xin[454]) );
  DFF \xreg_reg[456]  ( .D(xin[454]), .CLK(clk), .RST(start), .I(x[456]), .Q(
        xin[456]) );
  DFF \xreg_reg[458]  ( .D(xin[456]), .CLK(clk), .RST(start), .I(x[458]), .Q(
        xin[458]) );
  DFF \xreg_reg[460]  ( .D(xin[458]), .CLK(clk), .RST(start), .I(x[460]), .Q(
        xin[460]) );
  DFF \xreg_reg[462]  ( .D(xin[460]), .CLK(clk), .RST(start), .I(x[462]), .Q(
        xin[462]) );
  DFF \xreg_reg[464]  ( .D(xin[462]), .CLK(clk), .RST(start), .I(x[464]), .Q(
        xin[464]) );
  DFF \xreg_reg[466]  ( .D(xin[464]), .CLK(clk), .RST(start), .I(x[466]), .Q(
        xin[466]) );
  DFF \xreg_reg[468]  ( .D(xin[466]), .CLK(clk), .RST(start), .I(x[468]), .Q(
        xin[468]) );
  DFF \xreg_reg[470]  ( .D(xin[468]), .CLK(clk), .RST(start), .I(x[470]), .Q(
        xin[470]) );
  DFF \xreg_reg[472]  ( .D(xin[470]), .CLK(clk), .RST(start), .I(x[472]), .Q(
        xin[472]) );
  DFF \xreg_reg[474]  ( .D(xin[472]), .CLK(clk), .RST(start), .I(x[474]), .Q(
        xin[474]) );
  DFF \xreg_reg[476]  ( .D(xin[474]), .CLK(clk), .RST(start), .I(x[476]), .Q(
        xin[476]) );
  DFF \xreg_reg[478]  ( .D(xin[476]), .CLK(clk), .RST(start), .I(x[478]), .Q(
        xin[478]) );
  DFF \xreg_reg[480]  ( .D(xin[478]), .CLK(clk), .RST(start), .I(x[480]), .Q(
        xin[480]) );
  DFF \xreg_reg[482]  ( .D(xin[480]), .CLK(clk), .RST(start), .I(x[482]), .Q(
        xin[482]) );
  DFF \xreg_reg[484]  ( .D(xin[482]), .CLK(clk), .RST(start), .I(x[484]), .Q(
        xin[484]) );
  DFF \xreg_reg[486]  ( .D(xin[484]), .CLK(clk), .RST(start), .I(x[486]), .Q(
        xin[486]) );
  DFF \xreg_reg[488]  ( .D(xin[486]), .CLK(clk), .RST(start), .I(x[488]), .Q(
        xin[488]) );
  DFF \xreg_reg[490]  ( .D(xin[488]), .CLK(clk), .RST(start), .I(x[490]), .Q(
        xin[490]) );
  DFF \xreg_reg[492]  ( .D(xin[490]), .CLK(clk), .RST(start), .I(x[492]), .Q(
        xin[492]) );
  DFF \xreg_reg[494]  ( .D(xin[492]), .CLK(clk), .RST(start), .I(x[494]), .Q(
        xin[494]) );
  DFF \xreg_reg[496]  ( .D(xin[494]), .CLK(clk), .RST(start), .I(x[496]), .Q(
        xin[496]) );
  DFF \xreg_reg[498]  ( .D(xin[496]), .CLK(clk), .RST(start), .I(x[498]), .Q(
        xin[498]) );
  DFF \xreg_reg[500]  ( .D(xin[498]), .CLK(clk), .RST(start), .I(x[500]), .Q(
        xin[500]) );
  DFF \xreg_reg[502]  ( .D(xin[500]), .CLK(clk), .RST(start), .I(x[502]), .Q(
        xin[502]) );
  DFF \xreg_reg[504]  ( .D(xin[502]), .CLK(clk), .RST(start), .I(x[504]), .Q(
        xin[504]) );
  DFF \xreg_reg[506]  ( .D(xin[504]), .CLK(clk), .RST(start), .I(x[506]), .Q(
        xin[506]) );
  DFF \xreg_reg[508]  ( .D(xin[506]), .CLK(clk), .RST(start), .I(x[508]), .Q(
        xin[508]) );
  DFF \xreg_reg[510]  ( .D(xin[508]), .CLK(clk), .RST(start), .I(x[510]), .Q(
        xin[510]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][0] ) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][1] ) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][2] ) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][3] ) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][4] ) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][5] ) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][6] ) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][7] ) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][8] ) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][9] ) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][10] ) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][11] ) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][12] ) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][13] ) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][14] ) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][15] ) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][16] ) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][17] ) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][18] ) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][19] ) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][20] ) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][21] ) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][22] ) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][23] ) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][24] ) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][25] ) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][26] ) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][27] ) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][28] ) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][29] ) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][30] ) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][31] ) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][32] ) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][33] ) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][34] ) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][35] ) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][36] ) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][37] ) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][38] ) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][39] ) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][40] ) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][41] ) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][42] ) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][43] ) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][44] ) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][45] ) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][46] ) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][47] ) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][48] ) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][49] ) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][50] ) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][51] ) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][52] ) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][53] ) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][54] ) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][55] ) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][56] ) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][57] ) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][58] ) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][59] ) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][60] ) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][61] ) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][62] ) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][63] ) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][64] ) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][65] ) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][66] ) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][67] ) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][68] ) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][69] ) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][70] ) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][71] ) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][72] ) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][73] ) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][74] ) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][75] ) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][76] ) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][77] ) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][78] ) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][79] ) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][80] ) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][81] ) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][82] ) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][83] ) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][84] ) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][85] ) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][86] ) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][87] ) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][88] ) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][89] ) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][90] ) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][91] ) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][92] ) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][93] ) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][94] ) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][95] ) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][96] ) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][97] ) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][98] ) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][99] ) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][100] ) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][101] ) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][102] ) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][103] ) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][104] ) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][105] ) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][106] ) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][107] ) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][108] ) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][109] ) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][110] ) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][111] ) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][112] ) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][113] ) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][114] ) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][115] ) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][116] ) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][117] ) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][118] ) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][119] ) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][120] ) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][121] ) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][122] ) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][123] ) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][124] ) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][125] ) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][126] ) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][127] ) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][128] ) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][129] ) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][130] ) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][131] ) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][132] ) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][133] ) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][134] ) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][135] ) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][136] ) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][137] ) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][138] ) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][139] ) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][140] ) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][141] ) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][142] ) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][143] ) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][144] ) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][145] ) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][146] ) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][147] ) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][148] ) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][149] ) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][150] ) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][151] ) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][152] ) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][153] ) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][154] ) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][155] ) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][156] ) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][157] ) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][158] ) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][159] ) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][160] ) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][161] ) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][162] ) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][163] ) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][164] ) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][165] ) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][166] ) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][167] ) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][168] ) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][169] ) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][170] ) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][171] ) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][172] ) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][173] ) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][174] ) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][175] ) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][176] ) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][177] ) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][178] ) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][179] ) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][180] ) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][181] ) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][182] ) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][183] ) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][184] ) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][185] ) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][186] ) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][187] ) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][188] ) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][189] ) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][190] ) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][191] ) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][192] ) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][193] ) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][194] ) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][195] ) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][196] ) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][197] ) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][198] ) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][199] ) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][200] ) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][201] ) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][202] ) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][203] ) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][204] ) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][205] ) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][206] ) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][207] ) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][208] ) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][209] ) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][210] ) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][211] ) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][212] ) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][213] ) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][214] ) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][215] ) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][216] ) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][217] ) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][218] ) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][219] ) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][220] ) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][221] ) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][222] ) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][223] ) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][224] ) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][225] ) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][226] ) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][227] ) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][228] ) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][229] ) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][230] ) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][231] ) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][232] ) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][233] ) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][234] ) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][235] ) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][236] ) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][237] ) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][238] ) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][239] ) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][240] ) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][241] ) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][242] ) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][243] ) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][244] ) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][245] ) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][246] ) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][247] ) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][248] ) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][249] ) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][250] ) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][251] ) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][252] ) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][253] ) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][254] ) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][255] ) );
  DFF \zreg_reg[256]  ( .D(o[256]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][256] ) );
  DFF \zreg_reg[257]  ( .D(o[257]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][257] ) );
  DFF \zreg_reg[258]  ( .D(o[258]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][258] ) );
  DFF \zreg_reg[259]  ( .D(o[259]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][259] ) );
  DFF \zreg_reg[260]  ( .D(o[260]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][260] ) );
  DFF \zreg_reg[261]  ( .D(o[261]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][261] ) );
  DFF \zreg_reg[262]  ( .D(o[262]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][262] ) );
  DFF \zreg_reg[263]  ( .D(o[263]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][263] ) );
  DFF \zreg_reg[264]  ( .D(o[264]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][264] ) );
  DFF \zreg_reg[265]  ( .D(o[265]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][265] ) );
  DFF \zreg_reg[266]  ( .D(o[266]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][266] ) );
  DFF \zreg_reg[267]  ( .D(o[267]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][267] ) );
  DFF \zreg_reg[268]  ( .D(o[268]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][268] ) );
  DFF \zreg_reg[269]  ( .D(o[269]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][269] ) );
  DFF \zreg_reg[270]  ( .D(o[270]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][270] ) );
  DFF \zreg_reg[271]  ( .D(o[271]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][271] ) );
  DFF \zreg_reg[272]  ( .D(o[272]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][272] ) );
  DFF \zreg_reg[273]  ( .D(o[273]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][273] ) );
  DFF \zreg_reg[274]  ( .D(o[274]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][274] ) );
  DFF \zreg_reg[275]  ( .D(o[275]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][275] ) );
  DFF \zreg_reg[276]  ( .D(o[276]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][276] ) );
  DFF \zreg_reg[277]  ( .D(o[277]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][277] ) );
  DFF \zreg_reg[278]  ( .D(o[278]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][278] ) );
  DFF \zreg_reg[279]  ( .D(o[279]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][279] ) );
  DFF \zreg_reg[280]  ( .D(o[280]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][280] ) );
  DFF \zreg_reg[281]  ( .D(o[281]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][281] ) );
  DFF \zreg_reg[282]  ( .D(o[282]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][282] ) );
  DFF \zreg_reg[283]  ( .D(o[283]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][283] ) );
  DFF \zreg_reg[284]  ( .D(o[284]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][284] ) );
  DFF \zreg_reg[285]  ( .D(o[285]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][285] ) );
  DFF \zreg_reg[286]  ( .D(o[286]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][286] ) );
  DFF \zreg_reg[287]  ( .D(o[287]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][287] ) );
  DFF \zreg_reg[288]  ( .D(o[288]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][288] ) );
  DFF \zreg_reg[289]  ( .D(o[289]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][289] ) );
  DFF \zreg_reg[290]  ( .D(o[290]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][290] ) );
  DFF \zreg_reg[291]  ( .D(o[291]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][291] ) );
  DFF \zreg_reg[292]  ( .D(o[292]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][292] ) );
  DFF \zreg_reg[293]  ( .D(o[293]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][293] ) );
  DFF \zreg_reg[294]  ( .D(o[294]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][294] ) );
  DFF \zreg_reg[295]  ( .D(o[295]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][295] ) );
  DFF \zreg_reg[296]  ( .D(o[296]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][296] ) );
  DFF \zreg_reg[297]  ( .D(o[297]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][297] ) );
  DFF \zreg_reg[298]  ( .D(o[298]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][298] ) );
  DFF \zreg_reg[299]  ( .D(o[299]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][299] ) );
  DFF \zreg_reg[300]  ( .D(o[300]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][300] ) );
  DFF \zreg_reg[301]  ( .D(o[301]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][301] ) );
  DFF \zreg_reg[302]  ( .D(o[302]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][302] ) );
  DFF \zreg_reg[303]  ( .D(o[303]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][303] ) );
  DFF \zreg_reg[304]  ( .D(o[304]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][304] ) );
  DFF \zreg_reg[305]  ( .D(o[305]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][305] ) );
  DFF \zreg_reg[306]  ( .D(o[306]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][306] ) );
  DFF \zreg_reg[307]  ( .D(o[307]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][307] ) );
  DFF \zreg_reg[308]  ( .D(o[308]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][308] ) );
  DFF \zreg_reg[309]  ( .D(o[309]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][309] ) );
  DFF \zreg_reg[310]  ( .D(o[310]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][310] ) );
  DFF \zreg_reg[311]  ( .D(o[311]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][311] ) );
  DFF \zreg_reg[312]  ( .D(o[312]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][312] ) );
  DFF \zreg_reg[313]  ( .D(o[313]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][313] ) );
  DFF \zreg_reg[314]  ( .D(o[314]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][314] ) );
  DFF \zreg_reg[315]  ( .D(o[315]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][315] ) );
  DFF \zreg_reg[316]  ( .D(o[316]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][316] ) );
  DFF \zreg_reg[317]  ( .D(o[317]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][317] ) );
  DFF \zreg_reg[318]  ( .D(o[318]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][318] ) );
  DFF \zreg_reg[319]  ( .D(o[319]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][319] ) );
  DFF \zreg_reg[320]  ( .D(o[320]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][320] ) );
  DFF \zreg_reg[321]  ( .D(o[321]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][321] ) );
  DFF \zreg_reg[322]  ( .D(o[322]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][322] ) );
  DFF \zreg_reg[323]  ( .D(o[323]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][323] ) );
  DFF \zreg_reg[324]  ( .D(o[324]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][324] ) );
  DFF \zreg_reg[325]  ( .D(o[325]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][325] ) );
  DFF \zreg_reg[326]  ( .D(o[326]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][326] ) );
  DFF \zreg_reg[327]  ( .D(o[327]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][327] ) );
  DFF \zreg_reg[328]  ( .D(o[328]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][328] ) );
  DFF \zreg_reg[329]  ( .D(o[329]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][329] ) );
  DFF \zreg_reg[330]  ( .D(o[330]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][330] ) );
  DFF \zreg_reg[331]  ( .D(o[331]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][331] ) );
  DFF \zreg_reg[332]  ( .D(o[332]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][332] ) );
  DFF \zreg_reg[333]  ( .D(o[333]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][333] ) );
  DFF \zreg_reg[334]  ( .D(o[334]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][334] ) );
  DFF \zreg_reg[335]  ( .D(o[335]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][335] ) );
  DFF \zreg_reg[336]  ( .D(o[336]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][336] ) );
  DFF \zreg_reg[337]  ( .D(o[337]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][337] ) );
  DFF \zreg_reg[338]  ( .D(o[338]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][338] ) );
  DFF \zreg_reg[339]  ( .D(o[339]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][339] ) );
  DFF \zreg_reg[340]  ( .D(o[340]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][340] ) );
  DFF \zreg_reg[341]  ( .D(o[341]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][341] ) );
  DFF \zreg_reg[342]  ( .D(o[342]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][342] ) );
  DFF \zreg_reg[343]  ( .D(o[343]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][343] ) );
  DFF \zreg_reg[344]  ( .D(o[344]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][344] ) );
  DFF \zreg_reg[345]  ( .D(o[345]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][345] ) );
  DFF \zreg_reg[346]  ( .D(o[346]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][346] ) );
  DFF \zreg_reg[347]  ( .D(o[347]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][347] ) );
  DFF \zreg_reg[348]  ( .D(o[348]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][348] ) );
  DFF \zreg_reg[349]  ( .D(o[349]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][349] ) );
  DFF \zreg_reg[350]  ( .D(o[350]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][350] ) );
  DFF \zreg_reg[351]  ( .D(o[351]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][351] ) );
  DFF \zreg_reg[352]  ( .D(o[352]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][352] ) );
  DFF \zreg_reg[353]  ( .D(o[353]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][353] ) );
  DFF \zreg_reg[354]  ( .D(o[354]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][354] ) );
  DFF \zreg_reg[355]  ( .D(o[355]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][355] ) );
  DFF \zreg_reg[356]  ( .D(o[356]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][356] ) );
  DFF \zreg_reg[357]  ( .D(o[357]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][357] ) );
  DFF \zreg_reg[358]  ( .D(o[358]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][358] ) );
  DFF \zreg_reg[359]  ( .D(o[359]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][359] ) );
  DFF \zreg_reg[360]  ( .D(o[360]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][360] ) );
  DFF \zreg_reg[361]  ( .D(o[361]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][361] ) );
  DFF \zreg_reg[362]  ( .D(o[362]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][362] ) );
  DFF \zreg_reg[363]  ( .D(o[363]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][363] ) );
  DFF \zreg_reg[364]  ( .D(o[364]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][364] ) );
  DFF \zreg_reg[365]  ( .D(o[365]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][365] ) );
  DFF \zreg_reg[366]  ( .D(o[366]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][366] ) );
  DFF \zreg_reg[367]  ( .D(o[367]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][367] ) );
  DFF \zreg_reg[368]  ( .D(o[368]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][368] ) );
  DFF \zreg_reg[369]  ( .D(o[369]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][369] ) );
  DFF \zreg_reg[370]  ( .D(o[370]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][370] ) );
  DFF \zreg_reg[371]  ( .D(o[371]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][371] ) );
  DFF \zreg_reg[372]  ( .D(o[372]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][372] ) );
  DFF \zreg_reg[373]  ( .D(o[373]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][373] ) );
  DFF \zreg_reg[374]  ( .D(o[374]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][374] ) );
  DFF \zreg_reg[375]  ( .D(o[375]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][375] ) );
  DFF \zreg_reg[376]  ( .D(o[376]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][376] ) );
  DFF \zreg_reg[377]  ( .D(o[377]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][377] ) );
  DFF \zreg_reg[378]  ( .D(o[378]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][378] ) );
  DFF \zreg_reg[379]  ( .D(o[379]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][379] ) );
  DFF \zreg_reg[380]  ( .D(o[380]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][380] ) );
  DFF \zreg_reg[381]  ( .D(o[381]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][381] ) );
  DFF \zreg_reg[382]  ( .D(o[382]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][382] ) );
  DFF \zreg_reg[383]  ( .D(o[383]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][383] ) );
  DFF \zreg_reg[384]  ( .D(o[384]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][384] ) );
  DFF \zreg_reg[385]  ( .D(o[385]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][385] ) );
  DFF \zreg_reg[386]  ( .D(o[386]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][386] ) );
  DFF \zreg_reg[387]  ( .D(o[387]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][387] ) );
  DFF \zreg_reg[388]  ( .D(o[388]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][388] ) );
  DFF \zreg_reg[389]  ( .D(o[389]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][389] ) );
  DFF \zreg_reg[390]  ( .D(o[390]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][390] ) );
  DFF \zreg_reg[391]  ( .D(o[391]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][391] ) );
  DFF \zreg_reg[392]  ( .D(o[392]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][392] ) );
  DFF \zreg_reg[393]  ( .D(o[393]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][393] ) );
  DFF \zreg_reg[394]  ( .D(o[394]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][394] ) );
  DFF \zreg_reg[395]  ( .D(o[395]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][395] ) );
  DFF \zreg_reg[396]  ( .D(o[396]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][396] ) );
  DFF \zreg_reg[397]  ( .D(o[397]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][397] ) );
  DFF \zreg_reg[398]  ( .D(o[398]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][398] ) );
  DFF \zreg_reg[399]  ( .D(o[399]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][399] ) );
  DFF \zreg_reg[400]  ( .D(o[400]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][400] ) );
  DFF \zreg_reg[401]  ( .D(o[401]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][401] ) );
  DFF \zreg_reg[402]  ( .D(o[402]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][402] ) );
  DFF \zreg_reg[403]  ( .D(o[403]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][403] ) );
  DFF \zreg_reg[404]  ( .D(o[404]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][404] ) );
  DFF \zreg_reg[405]  ( .D(o[405]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][405] ) );
  DFF \zreg_reg[406]  ( .D(o[406]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][406] ) );
  DFF \zreg_reg[407]  ( .D(o[407]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][407] ) );
  DFF \zreg_reg[408]  ( .D(o[408]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][408] ) );
  DFF \zreg_reg[409]  ( .D(o[409]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][409] ) );
  DFF \zreg_reg[410]  ( .D(o[410]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][410] ) );
  DFF \zreg_reg[411]  ( .D(o[411]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][411] ) );
  DFF \zreg_reg[412]  ( .D(o[412]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][412] ) );
  DFF \zreg_reg[413]  ( .D(o[413]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][413] ) );
  DFF \zreg_reg[414]  ( .D(o[414]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][414] ) );
  DFF \zreg_reg[415]  ( .D(o[415]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][415] ) );
  DFF \zreg_reg[416]  ( .D(o[416]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][416] ) );
  DFF \zreg_reg[417]  ( .D(o[417]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][417] ) );
  DFF \zreg_reg[418]  ( .D(o[418]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][418] ) );
  DFF \zreg_reg[419]  ( .D(o[419]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][419] ) );
  DFF \zreg_reg[420]  ( .D(o[420]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][420] ) );
  DFF \zreg_reg[421]  ( .D(o[421]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][421] ) );
  DFF \zreg_reg[422]  ( .D(o[422]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][422] ) );
  DFF \zreg_reg[423]  ( .D(o[423]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][423] ) );
  DFF \zreg_reg[424]  ( .D(o[424]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][424] ) );
  DFF \zreg_reg[425]  ( .D(o[425]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][425] ) );
  DFF \zreg_reg[426]  ( .D(o[426]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][426] ) );
  DFF \zreg_reg[427]  ( .D(o[427]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][427] ) );
  DFF \zreg_reg[428]  ( .D(o[428]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][428] ) );
  DFF \zreg_reg[429]  ( .D(o[429]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][429] ) );
  DFF \zreg_reg[430]  ( .D(o[430]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][430] ) );
  DFF \zreg_reg[431]  ( .D(o[431]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][431] ) );
  DFF \zreg_reg[432]  ( .D(o[432]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][432] ) );
  DFF \zreg_reg[433]  ( .D(o[433]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][433] ) );
  DFF \zreg_reg[434]  ( .D(o[434]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][434] ) );
  DFF \zreg_reg[435]  ( .D(o[435]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][435] ) );
  DFF \zreg_reg[436]  ( .D(o[436]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][436] ) );
  DFF \zreg_reg[437]  ( .D(o[437]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][437] ) );
  DFF \zreg_reg[438]  ( .D(o[438]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][438] ) );
  DFF \zreg_reg[439]  ( .D(o[439]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][439] ) );
  DFF \zreg_reg[440]  ( .D(o[440]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][440] ) );
  DFF \zreg_reg[441]  ( .D(o[441]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][441] ) );
  DFF \zreg_reg[442]  ( .D(o[442]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][442] ) );
  DFF \zreg_reg[443]  ( .D(o[443]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][443] ) );
  DFF \zreg_reg[444]  ( .D(o[444]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][444] ) );
  DFF \zreg_reg[445]  ( .D(o[445]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][445] ) );
  DFF \zreg_reg[446]  ( .D(o[446]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][446] ) );
  DFF \zreg_reg[447]  ( .D(o[447]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][447] ) );
  DFF \zreg_reg[448]  ( .D(o[448]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][448] ) );
  DFF \zreg_reg[449]  ( .D(o[449]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][449] ) );
  DFF \zreg_reg[450]  ( .D(o[450]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][450] ) );
  DFF \zreg_reg[451]  ( .D(o[451]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][451] ) );
  DFF \zreg_reg[452]  ( .D(o[452]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][452] ) );
  DFF \zreg_reg[453]  ( .D(o[453]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][453] ) );
  DFF \zreg_reg[454]  ( .D(o[454]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][454] ) );
  DFF \zreg_reg[455]  ( .D(o[455]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][455] ) );
  DFF \zreg_reg[456]  ( .D(o[456]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][456] ) );
  DFF \zreg_reg[457]  ( .D(o[457]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][457] ) );
  DFF \zreg_reg[458]  ( .D(o[458]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][458] ) );
  DFF \zreg_reg[459]  ( .D(o[459]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][459] ) );
  DFF \zreg_reg[460]  ( .D(o[460]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][460] ) );
  DFF \zreg_reg[461]  ( .D(o[461]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][461] ) );
  DFF \zreg_reg[462]  ( .D(o[462]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][462] ) );
  DFF \zreg_reg[463]  ( .D(o[463]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][463] ) );
  DFF \zreg_reg[464]  ( .D(o[464]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][464] ) );
  DFF \zreg_reg[465]  ( .D(o[465]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][465] ) );
  DFF \zreg_reg[466]  ( .D(o[466]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][466] ) );
  DFF \zreg_reg[467]  ( .D(o[467]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][467] ) );
  DFF \zreg_reg[468]  ( .D(o[468]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][468] ) );
  DFF \zreg_reg[469]  ( .D(o[469]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][469] ) );
  DFF \zreg_reg[470]  ( .D(o[470]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][470] ) );
  DFF \zreg_reg[471]  ( .D(o[471]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][471] ) );
  DFF \zreg_reg[472]  ( .D(o[472]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][472] ) );
  DFF \zreg_reg[473]  ( .D(o[473]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][473] ) );
  DFF \zreg_reg[474]  ( .D(o[474]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][474] ) );
  DFF \zreg_reg[475]  ( .D(o[475]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][475] ) );
  DFF \zreg_reg[476]  ( .D(o[476]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][476] ) );
  DFF \zreg_reg[477]  ( .D(o[477]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][477] ) );
  DFF \zreg_reg[478]  ( .D(o[478]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][478] ) );
  DFF \zreg_reg[479]  ( .D(o[479]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][479] ) );
  DFF \zreg_reg[480]  ( .D(o[480]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][480] ) );
  DFF \zreg_reg[481]  ( .D(o[481]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][481] ) );
  DFF \zreg_reg[482]  ( .D(o[482]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][482] ) );
  DFF \zreg_reg[483]  ( .D(o[483]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][483] ) );
  DFF \zreg_reg[484]  ( .D(o[484]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][484] ) );
  DFF \zreg_reg[485]  ( .D(o[485]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][485] ) );
  DFF \zreg_reg[486]  ( .D(o[486]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][486] ) );
  DFF \zreg_reg[487]  ( .D(o[487]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][487] ) );
  DFF \zreg_reg[488]  ( .D(o[488]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][488] ) );
  DFF \zreg_reg[489]  ( .D(o[489]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][489] ) );
  DFF \zreg_reg[490]  ( .D(o[490]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][490] ) );
  DFF \zreg_reg[491]  ( .D(o[491]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][491] ) );
  DFF \zreg_reg[492]  ( .D(o[492]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][492] ) );
  DFF \zreg_reg[493]  ( .D(o[493]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][493] ) );
  DFF \zreg_reg[494]  ( .D(o[494]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][494] ) );
  DFF \zreg_reg[495]  ( .D(o[495]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][495] ) );
  DFF \zreg_reg[496]  ( .D(o[496]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][496] ) );
  DFF \zreg_reg[497]  ( .D(o[497]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][497] ) );
  DFF \zreg_reg[498]  ( .D(o[498]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][498] ) );
  DFF \zreg_reg[499]  ( .D(o[499]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][499] ) );
  DFF \zreg_reg[500]  ( .D(o[500]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][500] ) );
  DFF \zreg_reg[501]  ( .D(o[501]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][501] ) );
  DFF \zreg_reg[502]  ( .D(o[502]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][502] ) );
  DFF \zreg_reg[503]  ( .D(o[503]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][503] ) );
  DFF \zreg_reg[504]  ( .D(o[504]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][504] ) );
  DFF \zreg_reg[505]  ( .D(o[505]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][505] ) );
  DFF \zreg_reg[506]  ( .D(o[506]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][506] ) );
  DFF \zreg_reg[507]  ( .D(o[507]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][507] ) );
  DFF \zreg_reg[508]  ( .D(o[508]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][508] ) );
  DFF \zreg_reg[509]  ( .D(o[509]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][509] ) );
  DFF \zreg_reg[510]  ( .D(o[510]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][510] ) );
  DFF \zreg_reg[511]  ( .D(o[511]), .CLK(clk), .RST(start), .I(1'b0), .Q(
        \zin[0][511] ) );
  DFF \zreg_reg[512]  ( .D(\zout[1][512] ), .CLK(clk), .RST(start), .I(1'b0), 
        .Q(\zin[0][512] ) );
endmodule


module MUX_N512_4 ( A, B, S, O );
  input [511:0] A;
  input [511:0] B;
  output [511:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024;

  XOR U1 ( .A(A[9]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XOR U4 ( .A(A[99]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U7 ( .A(A[98]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U10 ( .A(A[97]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U13 ( .A(A[96]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U16 ( .A(A[95]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U19 ( .A(A[94]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U22 ( .A(A[93]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U25 ( .A(A[92]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U28 ( .A(A[91]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U31 ( .A(A[90]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U34 ( .A(A[8]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U37 ( .A(A[89]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U40 ( .A(A[88]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U43 ( .A(A[87]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U46 ( .A(A[86]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U49 ( .A(A[85]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U52 ( .A(A[84]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U55 ( .A(A[83]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U58 ( .A(A[82]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U61 ( .A(A[81]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U64 ( .A(A[80]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U67 ( .A(A[7]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U70 ( .A(A[79]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U73 ( .A(A[78]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U76 ( .A(A[77]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U79 ( .A(A[76]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U82 ( .A(A[75]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U85 ( .A(A[74]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U88 ( .A(A[73]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U91 ( .A(A[72]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U94 ( .A(A[71]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U97 ( .A(A[70]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U100 ( .A(A[6]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U103 ( .A(A[69]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U106 ( .A(A[68]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U109 ( .A(A[67]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U112 ( .A(A[66]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U115 ( .A(A[65]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U118 ( .A(A[64]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U121 ( .A(A[63]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U124 ( .A(A[62]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U127 ( .A(A[61]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U130 ( .A(A[60]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U133 ( .A(A[5]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U136 ( .A(A[59]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U139 ( .A(A[58]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U142 ( .A(A[57]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U145 ( .A(A[56]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U148 ( .A(A[55]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U151 ( .A(A[54]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U154 ( .A(A[53]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U157 ( .A(A[52]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U160 ( .A(A[51]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U163 ( .A(A[511]), .B(n109), .Z(O[511]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[511]), .B(A[511]), .Z(n110) );
  XOR U166 ( .A(A[510]), .B(n111), .Z(O[510]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[510]), .B(A[510]), .Z(n112) );
  XOR U169 ( .A(A[50]), .B(n113), .Z(O[50]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[50]), .B(A[50]), .Z(n114) );
  XOR U172 ( .A(A[509]), .B(n115), .Z(O[509]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[509]), .B(A[509]), .Z(n116) );
  XOR U175 ( .A(A[508]), .B(n117), .Z(O[508]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[508]), .B(A[508]), .Z(n118) );
  XOR U178 ( .A(A[507]), .B(n119), .Z(O[507]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[507]), .B(A[507]), .Z(n120) );
  XOR U181 ( .A(A[506]), .B(n121), .Z(O[506]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[506]), .B(A[506]), .Z(n122) );
  XOR U184 ( .A(A[505]), .B(n123), .Z(O[505]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[505]), .B(A[505]), .Z(n124) );
  XOR U187 ( .A(A[504]), .B(n125), .Z(O[504]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[504]), .B(A[504]), .Z(n126) );
  XOR U190 ( .A(A[503]), .B(n127), .Z(O[503]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[503]), .B(A[503]), .Z(n128) );
  XOR U193 ( .A(A[502]), .B(n129), .Z(O[502]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[502]), .B(A[502]), .Z(n130) );
  XOR U196 ( .A(A[501]), .B(n131), .Z(O[501]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[501]), .B(A[501]), .Z(n132) );
  XOR U199 ( .A(A[500]), .B(n133), .Z(O[500]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[500]), .B(A[500]), .Z(n134) );
  XOR U202 ( .A(A[4]), .B(n135), .Z(O[4]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[4]), .B(A[4]), .Z(n136) );
  XOR U205 ( .A(A[49]), .B(n137), .Z(O[49]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[49]), .B(A[49]), .Z(n138) );
  XOR U208 ( .A(A[499]), .B(n139), .Z(O[499]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[499]), .B(A[499]), .Z(n140) );
  XOR U211 ( .A(A[498]), .B(n141), .Z(O[498]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[498]), .B(A[498]), .Z(n142) );
  XOR U214 ( .A(A[497]), .B(n143), .Z(O[497]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[497]), .B(A[497]), .Z(n144) );
  XOR U217 ( .A(A[496]), .B(n145), .Z(O[496]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[496]), .B(A[496]), .Z(n146) );
  XOR U220 ( .A(A[495]), .B(n147), .Z(O[495]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[495]), .B(A[495]), .Z(n148) );
  XOR U223 ( .A(A[494]), .B(n149), .Z(O[494]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[494]), .B(A[494]), .Z(n150) );
  XOR U226 ( .A(A[493]), .B(n151), .Z(O[493]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[493]), .B(A[493]), .Z(n152) );
  XOR U229 ( .A(A[492]), .B(n153), .Z(O[492]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[492]), .B(A[492]), .Z(n154) );
  XOR U232 ( .A(A[491]), .B(n155), .Z(O[491]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[491]), .B(A[491]), .Z(n156) );
  XOR U235 ( .A(A[490]), .B(n157), .Z(O[490]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[490]), .B(A[490]), .Z(n158) );
  XOR U238 ( .A(A[48]), .B(n159), .Z(O[48]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[48]), .B(A[48]), .Z(n160) );
  XOR U241 ( .A(A[489]), .B(n161), .Z(O[489]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[489]), .B(A[489]), .Z(n162) );
  XOR U244 ( .A(A[488]), .B(n163), .Z(O[488]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[488]), .B(A[488]), .Z(n164) );
  XOR U247 ( .A(A[487]), .B(n165), .Z(O[487]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[487]), .B(A[487]), .Z(n166) );
  XOR U250 ( .A(A[486]), .B(n167), .Z(O[486]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[486]), .B(A[486]), .Z(n168) );
  XOR U253 ( .A(A[485]), .B(n169), .Z(O[485]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[485]), .B(A[485]), .Z(n170) );
  XOR U256 ( .A(A[484]), .B(n171), .Z(O[484]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[484]), .B(A[484]), .Z(n172) );
  XOR U259 ( .A(A[483]), .B(n173), .Z(O[483]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[483]), .B(A[483]), .Z(n174) );
  XOR U262 ( .A(A[482]), .B(n175), .Z(O[482]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[482]), .B(A[482]), .Z(n176) );
  XOR U265 ( .A(A[481]), .B(n177), .Z(O[481]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[481]), .B(A[481]), .Z(n178) );
  XOR U268 ( .A(A[480]), .B(n179), .Z(O[480]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[480]), .B(A[480]), .Z(n180) );
  XOR U271 ( .A(A[47]), .B(n181), .Z(O[47]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[47]), .B(A[47]), .Z(n182) );
  XOR U274 ( .A(A[479]), .B(n183), .Z(O[479]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[479]), .B(A[479]), .Z(n184) );
  XOR U277 ( .A(A[478]), .B(n185), .Z(O[478]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[478]), .B(A[478]), .Z(n186) );
  XOR U280 ( .A(A[477]), .B(n187), .Z(O[477]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[477]), .B(A[477]), .Z(n188) );
  XOR U283 ( .A(A[476]), .B(n189), .Z(O[476]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[476]), .B(A[476]), .Z(n190) );
  XOR U286 ( .A(A[475]), .B(n191), .Z(O[475]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[475]), .B(A[475]), .Z(n192) );
  XOR U289 ( .A(A[474]), .B(n193), .Z(O[474]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[474]), .B(A[474]), .Z(n194) );
  XOR U292 ( .A(A[473]), .B(n195), .Z(O[473]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[473]), .B(A[473]), .Z(n196) );
  XOR U295 ( .A(A[472]), .B(n197), .Z(O[472]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[472]), .B(A[472]), .Z(n198) );
  XOR U298 ( .A(A[471]), .B(n199), .Z(O[471]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[471]), .B(A[471]), .Z(n200) );
  XOR U301 ( .A(A[470]), .B(n201), .Z(O[470]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[470]), .B(A[470]), .Z(n202) );
  XOR U304 ( .A(A[46]), .B(n203), .Z(O[46]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[46]), .B(A[46]), .Z(n204) );
  XOR U307 ( .A(A[469]), .B(n205), .Z(O[469]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[469]), .B(A[469]), .Z(n206) );
  XOR U310 ( .A(A[468]), .B(n207), .Z(O[468]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[468]), .B(A[468]), .Z(n208) );
  XOR U313 ( .A(A[467]), .B(n209), .Z(O[467]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[467]), .B(A[467]), .Z(n210) );
  XOR U316 ( .A(A[466]), .B(n211), .Z(O[466]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[466]), .B(A[466]), .Z(n212) );
  XOR U319 ( .A(A[465]), .B(n213), .Z(O[465]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[465]), .B(A[465]), .Z(n214) );
  XOR U322 ( .A(A[464]), .B(n215), .Z(O[464]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[464]), .B(A[464]), .Z(n216) );
  XOR U325 ( .A(A[463]), .B(n217), .Z(O[463]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[463]), .B(A[463]), .Z(n218) );
  XOR U328 ( .A(A[462]), .B(n219), .Z(O[462]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[462]), .B(A[462]), .Z(n220) );
  XOR U331 ( .A(A[461]), .B(n221), .Z(O[461]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[461]), .B(A[461]), .Z(n222) );
  XOR U334 ( .A(A[460]), .B(n223), .Z(O[460]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[460]), .B(A[460]), .Z(n224) );
  XOR U337 ( .A(A[45]), .B(n225), .Z(O[45]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[45]), .B(A[45]), .Z(n226) );
  XOR U340 ( .A(A[459]), .B(n227), .Z(O[459]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[459]), .B(A[459]), .Z(n228) );
  XOR U343 ( .A(A[458]), .B(n229), .Z(O[458]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[458]), .B(A[458]), .Z(n230) );
  XOR U346 ( .A(A[457]), .B(n231), .Z(O[457]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[457]), .B(A[457]), .Z(n232) );
  XOR U349 ( .A(A[456]), .B(n233), .Z(O[456]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[456]), .B(A[456]), .Z(n234) );
  XOR U352 ( .A(A[455]), .B(n235), .Z(O[455]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[455]), .B(A[455]), .Z(n236) );
  XOR U355 ( .A(A[454]), .B(n237), .Z(O[454]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[454]), .B(A[454]), .Z(n238) );
  XOR U358 ( .A(A[453]), .B(n239), .Z(O[453]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[453]), .B(A[453]), .Z(n240) );
  XOR U361 ( .A(A[452]), .B(n241), .Z(O[452]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[452]), .B(A[452]), .Z(n242) );
  XOR U364 ( .A(A[451]), .B(n243), .Z(O[451]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[451]), .B(A[451]), .Z(n244) );
  XOR U367 ( .A(A[450]), .B(n245), .Z(O[450]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[450]), .B(A[450]), .Z(n246) );
  XOR U370 ( .A(A[44]), .B(n247), .Z(O[44]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[44]), .B(A[44]), .Z(n248) );
  XOR U373 ( .A(A[449]), .B(n249), .Z(O[449]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[449]), .B(A[449]), .Z(n250) );
  XOR U376 ( .A(A[448]), .B(n251), .Z(O[448]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[448]), .B(A[448]), .Z(n252) );
  XOR U379 ( .A(A[447]), .B(n253), .Z(O[447]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[447]), .B(A[447]), .Z(n254) );
  XOR U382 ( .A(A[446]), .B(n255), .Z(O[446]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[446]), .B(A[446]), .Z(n256) );
  XOR U385 ( .A(A[445]), .B(n257), .Z(O[445]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[445]), .B(A[445]), .Z(n258) );
  XOR U388 ( .A(A[444]), .B(n259), .Z(O[444]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[444]), .B(A[444]), .Z(n260) );
  XOR U391 ( .A(A[443]), .B(n261), .Z(O[443]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[443]), .B(A[443]), .Z(n262) );
  XOR U394 ( .A(A[442]), .B(n263), .Z(O[442]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[442]), .B(A[442]), .Z(n264) );
  XOR U397 ( .A(A[441]), .B(n265), .Z(O[441]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[441]), .B(A[441]), .Z(n266) );
  XOR U400 ( .A(A[440]), .B(n267), .Z(O[440]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[440]), .B(A[440]), .Z(n268) );
  XOR U403 ( .A(A[43]), .B(n269), .Z(O[43]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[43]), .B(A[43]), .Z(n270) );
  XOR U406 ( .A(A[439]), .B(n271), .Z(O[439]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[439]), .B(A[439]), .Z(n272) );
  XOR U409 ( .A(A[438]), .B(n273), .Z(O[438]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[438]), .B(A[438]), .Z(n274) );
  XOR U412 ( .A(A[437]), .B(n275), .Z(O[437]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[437]), .B(A[437]), .Z(n276) );
  XOR U415 ( .A(A[436]), .B(n277), .Z(O[436]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[436]), .B(A[436]), .Z(n278) );
  XOR U418 ( .A(A[435]), .B(n279), .Z(O[435]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[435]), .B(A[435]), .Z(n280) );
  XOR U421 ( .A(A[434]), .B(n281), .Z(O[434]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[434]), .B(A[434]), .Z(n282) );
  XOR U424 ( .A(A[433]), .B(n283), .Z(O[433]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[433]), .B(A[433]), .Z(n284) );
  XOR U427 ( .A(A[432]), .B(n285), .Z(O[432]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[432]), .B(A[432]), .Z(n286) );
  XOR U430 ( .A(A[431]), .B(n287), .Z(O[431]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[431]), .B(A[431]), .Z(n288) );
  XOR U433 ( .A(A[430]), .B(n289), .Z(O[430]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[430]), .B(A[430]), .Z(n290) );
  XOR U436 ( .A(A[42]), .B(n291), .Z(O[42]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[42]), .B(A[42]), .Z(n292) );
  XOR U439 ( .A(A[429]), .B(n293), .Z(O[429]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[429]), .B(A[429]), .Z(n294) );
  XOR U442 ( .A(A[428]), .B(n295), .Z(O[428]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[428]), .B(A[428]), .Z(n296) );
  XOR U445 ( .A(A[427]), .B(n297), .Z(O[427]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[427]), .B(A[427]), .Z(n298) );
  XOR U448 ( .A(A[426]), .B(n299), .Z(O[426]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[426]), .B(A[426]), .Z(n300) );
  XOR U451 ( .A(A[425]), .B(n301), .Z(O[425]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[425]), .B(A[425]), .Z(n302) );
  XOR U454 ( .A(A[424]), .B(n303), .Z(O[424]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[424]), .B(A[424]), .Z(n304) );
  XOR U457 ( .A(A[423]), .B(n305), .Z(O[423]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[423]), .B(A[423]), .Z(n306) );
  XOR U460 ( .A(A[422]), .B(n307), .Z(O[422]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[422]), .B(A[422]), .Z(n308) );
  XOR U463 ( .A(A[421]), .B(n309), .Z(O[421]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[421]), .B(A[421]), .Z(n310) );
  XOR U466 ( .A(A[420]), .B(n311), .Z(O[420]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[420]), .B(A[420]), .Z(n312) );
  XOR U469 ( .A(A[41]), .B(n313), .Z(O[41]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[41]), .B(A[41]), .Z(n314) );
  XOR U472 ( .A(A[419]), .B(n315), .Z(O[419]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[419]), .B(A[419]), .Z(n316) );
  XOR U475 ( .A(A[418]), .B(n317), .Z(O[418]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[418]), .B(A[418]), .Z(n318) );
  XOR U478 ( .A(A[417]), .B(n319), .Z(O[417]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[417]), .B(A[417]), .Z(n320) );
  XOR U481 ( .A(A[416]), .B(n321), .Z(O[416]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[416]), .B(A[416]), .Z(n322) );
  XOR U484 ( .A(A[415]), .B(n323), .Z(O[415]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[415]), .B(A[415]), .Z(n324) );
  XOR U487 ( .A(A[414]), .B(n325), .Z(O[414]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[414]), .B(A[414]), .Z(n326) );
  XOR U490 ( .A(A[413]), .B(n327), .Z(O[413]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[413]), .B(A[413]), .Z(n328) );
  XOR U493 ( .A(A[412]), .B(n329), .Z(O[412]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[412]), .B(A[412]), .Z(n330) );
  XOR U496 ( .A(A[411]), .B(n331), .Z(O[411]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[411]), .B(A[411]), .Z(n332) );
  XOR U499 ( .A(A[410]), .B(n333), .Z(O[410]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[410]), .B(A[410]), .Z(n334) );
  XOR U502 ( .A(A[40]), .B(n335), .Z(O[40]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[40]), .B(A[40]), .Z(n336) );
  XOR U505 ( .A(A[409]), .B(n337), .Z(O[409]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[409]), .B(A[409]), .Z(n338) );
  XOR U508 ( .A(A[408]), .B(n339), .Z(O[408]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[408]), .B(A[408]), .Z(n340) );
  XOR U511 ( .A(A[407]), .B(n341), .Z(O[407]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[407]), .B(A[407]), .Z(n342) );
  XOR U514 ( .A(A[406]), .B(n343), .Z(O[406]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[406]), .B(A[406]), .Z(n344) );
  XOR U517 ( .A(A[405]), .B(n345), .Z(O[405]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[405]), .B(A[405]), .Z(n346) );
  XOR U520 ( .A(A[404]), .B(n347), .Z(O[404]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[404]), .B(A[404]), .Z(n348) );
  XOR U523 ( .A(A[403]), .B(n349), .Z(O[403]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[403]), .B(A[403]), .Z(n350) );
  XOR U526 ( .A(A[402]), .B(n351), .Z(O[402]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[402]), .B(A[402]), .Z(n352) );
  XOR U529 ( .A(A[401]), .B(n353), .Z(O[401]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[401]), .B(A[401]), .Z(n354) );
  XOR U532 ( .A(A[400]), .B(n355), .Z(O[400]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[400]), .B(A[400]), .Z(n356) );
  XOR U535 ( .A(A[3]), .B(n357), .Z(O[3]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[3]), .B(A[3]), .Z(n358) );
  XOR U538 ( .A(A[39]), .B(n359), .Z(O[39]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[39]), .B(A[39]), .Z(n360) );
  XOR U541 ( .A(A[399]), .B(n361), .Z(O[399]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[399]), .B(A[399]), .Z(n362) );
  XOR U544 ( .A(A[398]), .B(n363), .Z(O[398]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[398]), .B(A[398]), .Z(n364) );
  XOR U547 ( .A(A[397]), .B(n365), .Z(O[397]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[397]), .B(A[397]), .Z(n366) );
  XOR U550 ( .A(A[396]), .B(n367), .Z(O[396]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[396]), .B(A[396]), .Z(n368) );
  XOR U553 ( .A(A[395]), .B(n369), .Z(O[395]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[395]), .B(A[395]), .Z(n370) );
  XOR U556 ( .A(A[394]), .B(n371), .Z(O[394]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[394]), .B(A[394]), .Z(n372) );
  XOR U559 ( .A(A[393]), .B(n373), .Z(O[393]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[393]), .B(A[393]), .Z(n374) );
  XOR U562 ( .A(A[392]), .B(n375), .Z(O[392]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[392]), .B(A[392]), .Z(n376) );
  XOR U565 ( .A(A[391]), .B(n377), .Z(O[391]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[391]), .B(A[391]), .Z(n378) );
  XOR U568 ( .A(A[390]), .B(n379), .Z(O[390]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[390]), .B(A[390]), .Z(n380) );
  XOR U571 ( .A(A[38]), .B(n381), .Z(O[38]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[38]), .B(A[38]), .Z(n382) );
  XOR U574 ( .A(A[389]), .B(n383), .Z(O[389]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[389]), .B(A[389]), .Z(n384) );
  XOR U577 ( .A(A[388]), .B(n385), .Z(O[388]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[388]), .B(A[388]), .Z(n386) );
  XOR U580 ( .A(A[387]), .B(n387), .Z(O[387]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[387]), .B(A[387]), .Z(n388) );
  XOR U583 ( .A(A[386]), .B(n389), .Z(O[386]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[386]), .B(A[386]), .Z(n390) );
  XOR U586 ( .A(A[385]), .B(n391), .Z(O[385]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[385]), .B(A[385]), .Z(n392) );
  XOR U589 ( .A(A[384]), .B(n393), .Z(O[384]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[384]), .B(A[384]), .Z(n394) );
  XOR U592 ( .A(A[383]), .B(n395), .Z(O[383]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[383]), .B(A[383]), .Z(n396) );
  XOR U595 ( .A(A[382]), .B(n397), .Z(O[382]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[382]), .B(A[382]), .Z(n398) );
  XOR U598 ( .A(A[381]), .B(n399), .Z(O[381]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[381]), .B(A[381]), .Z(n400) );
  XOR U601 ( .A(A[380]), .B(n401), .Z(O[380]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[380]), .B(A[380]), .Z(n402) );
  XOR U604 ( .A(A[37]), .B(n403), .Z(O[37]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[37]), .B(A[37]), .Z(n404) );
  XOR U607 ( .A(A[379]), .B(n405), .Z(O[379]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[379]), .B(A[379]), .Z(n406) );
  XOR U610 ( .A(A[378]), .B(n407), .Z(O[378]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[378]), .B(A[378]), .Z(n408) );
  XOR U613 ( .A(A[377]), .B(n409), .Z(O[377]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[377]), .B(A[377]), .Z(n410) );
  XOR U616 ( .A(A[376]), .B(n411), .Z(O[376]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[376]), .B(A[376]), .Z(n412) );
  XOR U619 ( .A(A[375]), .B(n413), .Z(O[375]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[375]), .B(A[375]), .Z(n414) );
  XOR U622 ( .A(A[374]), .B(n415), .Z(O[374]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[374]), .B(A[374]), .Z(n416) );
  XOR U625 ( .A(A[373]), .B(n417), .Z(O[373]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[373]), .B(A[373]), .Z(n418) );
  XOR U628 ( .A(A[372]), .B(n419), .Z(O[372]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[372]), .B(A[372]), .Z(n420) );
  XOR U631 ( .A(A[371]), .B(n421), .Z(O[371]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[371]), .B(A[371]), .Z(n422) );
  XOR U634 ( .A(A[370]), .B(n423), .Z(O[370]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[370]), .B(A[370]), .Z(n424) );
  XOR U637 ( .A(A[36]), .B(n425), .Z(O[36]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[36]), .B(A[36]), .Z(n426) );
  XOR U640 ( .A(A[369]), .B(n427), .Z(O[369]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[369]), .B(A[369]), .Z(n428) );
  XOR U643 ( .A(A[368]), .B(n429), .Z(O[368]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[368]), .B(A[368]), .Z(n430) );
  XOR U646 ( .A(A[367]), .B(n431), .Z(O[367]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[367]), .B(A[367]), .Z(n432) );
  XOR U649 ( .A(A[366]), .B(n433), .Z(O[366]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[366]), .B(A[366]), .Z(n434) );
  XOR U652 ( .A(A[365]), .B(n435), .Z(O[365]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[365]), .B(A[365]), .Z(n436) );
  XOR U655 ( .A(A[364]), .B(n437), .Z(O[364]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[364]), .B(A[364]), .Z(n438) );
  XOR U658 ( .A(A[363]), .B(n439), .Z(O[363]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[363]), .B(A[363]), .Z(n440) );
  XOR U661 ( .A(A[362]), .B(n441), .Z(O[362]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[362]), .B(A[362]), .Z(n442) );
  XOR U664 ( .A(A[361]), .B(n443), .Z(O[361]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[361]), .B(A[361]), .Z(n444) );
  XOR U667 ( .A(A[360]), .B(n445), .Z(O[360]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[360]), .B(A[360]), .Z(n446) );
  XOR U670 ( .A(A[35]), .B(n447), .Z(O[35]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[35]), .B(A[35]), .Z(n448) );
  XOR U673 ( .A(A[359]), .B(n449), .Z(O[359]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[359]), .B(A[359]), .Z(n450) );
  XOR U676 ( .A(A[358]), .B(n451), .Z(O[358]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[358]), .B(A[358]), .Z(n452) );
  XOR U679 ( .A(A[357]), .B(n453), .Z(O[357]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[357]), .B(A[357]), .Z(n454) );
  XOR U682 ( .A(A[356]), .B(n455), .Z(O[356]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[356]), .B(A[356]), .Z(n456) );
  XOR U685 ( .A(A[355]), .B(n457), .Z(O[355]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[355]), .B(A[355]), .Z(n458) );
  XOR U688 ( .A(A[354]), .B(n459), .Z(O[354]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[354]), .B(A[354]), .Z(n460) );
  XOR U691 ( .A(A[353]), .B(n461), .Z(O[353]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[353]), .B(A[353]), .Z(n462) );
  XOR U694 ( .A(A[352]), .B(n463), .Z(O[352]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[352]), .B(A[352]), .Z(n464) );
  XOR U697 ( .A(A[351]), .B(n465), .Z(O[351]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[351]), .B(A[351]), .Z(n466) );
  XOR U700 ( .A(A[350]), .B(n467), .Z(O[350]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[350]), .B(A[350]), .Z(n468) );
  XOR U703 ( .A(A[34]), .B(n469), .Z(O[34]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[34]), .B(A[34]), .Z(n470) );
  XOR U706 ( .A(A[349]), .B(n471), .Z(O[349]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[349]), .B(A[349]), .Z(n472) );
  XOR U709 ( .A(A[348]), .B(n473), .Z(O[348]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[348]), .B(A[348]), .Z(n474) );
  XOR U712 ( .A(A[347]), .B(n475), .Z(O[347]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[347]), .B(A[347]), .Z(n476) );
  XOR U715 ( .A(A[346]), .B(n477), .Z(O[346]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[346]), .B(A[346]), .Z(n478) );
  XOR U718 ( .A(A[345]), .B(n479), .Z(O[345]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[345]), .B(A[345]), .Z(n480) );
  XOR U721 ( .A(A[344]), .B(n481), .Z(O[344]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[344]), .B(A[344]), .Z(n482) );
  XOR U724 ( .A(A[343]), .B(n483), .Z(O[343]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[343]), .B(A[343]), .Z(n484) );
  XOR U727 ( .A(A[342]), .B(n485), .Z(O[342]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[342]), .B(A[342]), .Z(n486) );
  XOR U730 ( .A(A[341]), .B(n487), .Z(O[341]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[341]), .B(A[341]), .Z(n488) );
  XOR U733 ( .A(A[340]), .B(n489), .Z(O[340]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[340]), .B(A[340]), .Z(n490) );
  XOR U736 ( .A(A[33]), .B(n491), .Z(O[33]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[33]), .B(A[33]), .Z(n492) );
  XOR U739 ( .A(A[339]), .B(n493), .Z(O[339]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[339]), .B(A[339]), .Z(n494) );
  XOR U742 ( .A(A[338]), .B(n495), .Z(O[338]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[338]), .B(A[338]), .Z(n496) );
  XOR U745 ( .A(A[337]), .B(n497), .Z(O[337]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[337]), .B(A[337]), .Z(n498) );
  XOR U748 ( .A(A[336]), .B(n499), .Z(O[336]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[336]), .B(A[336]), .Z(n500) );
  XOR U751 ( .A(A[335]), .B(n501), .Z(O[335]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[335]), .B(A[335]), .Z(n502) );
  XOR U754 ( .A(A[334]), .B(n503), .Z(O[334]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[334]), .B(A[334]), .Z(n504) );
  XOR U757 ( .A(A[333]), .B(n505), .Z(O[333]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[333]), .B(A[333]), .Z(n506) );
  XOR U760 ( .A(A[332]), .B(n507), .Z(O[332]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[332]), .B(A[332]), .Z(n508) );
  XOR U763 ( .A(A[331]), .B(n509), .Z(O[331]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[331]), .B(A[331]), .Z(n510) );
  XOR U766 ( .A(A[330]), .B(n511), .Z(O[330]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[330]), .B(A[330]), .Z(n512) );
  XOR U769 ( .A(A[32]), .B(n513), .Z(O[32]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[32]), .B(A[32]), .Z(n514) );
  XOR U772 ( .A(A[329]), .B(n515), .Z(O[329]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[329]), .B(A[329]), .Z(n516) );
  XOR U775 ( .A(A[328]), .B(n517), .Z(O[328]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[328]), .B(A[328]), .Z(n518) );
  XOR U778 ( .A(A[327]), .B(n519), .Z(O[327]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[327]), .B(A[327]), .Z(n520) );
  XOR U781 ( .A(A[326]), .B(n521), .Z(O[326]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[326]), .B(A[326]), .Z(n522) );
  XOR U784 ( .A(A[325]), .B(n523), .Z(O[325]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[325]), .B(A[325]), .Z(n524) );
  XOR U787 ( .A(A[324]), .B(n525), .Z(O[324]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[324]), .B(A[324]), .Z(n526) );
  XOR U790 ( .A(A[323]), .B(n527), .Z(O[323]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[323]), .B(A[323]), .Z(n528) );
  XOR U793 ( .A(A[322]), .B(n529), .Z(O[322]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[322]), .B(A[322]), .Z(n530) );
  XOR U796 ( .A(A[321]), .B(n531), .Z(O[321]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[321]), .B(A[321]), .Z(n532) );
  XOR U799 ( .A(A[320]), .B(n533), .Z(O[320]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[320]), .B(A[320]), .Z(n534) );
  XOR U802 ( .A(A[31]), .B(n535), .Z(O[31]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[31]), .B(A[31]), .Z(n536) );
  XOR U805 ( .A(A[319]), .B(n537), .Z(O[319]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[319]), .B(A[319]), .Z(n538) );
  XOR U808 ( .A(A[318]), .B(n539), .Z(O[318]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[318]), .B(A[318]), .Z(n540) );
  XOR U811 ( .A(A[317]), .B(n541), .Z(O[317]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[317]), .B(A[317]), .Z(n542) );
  XOR U814 ( .A(A[316]), .B(n543), .Z(O[316]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[316]), .B(A[316]), .Z(n544) );
  XOR U817 ( .A(A[315]), .B(n545), .Z(O[315]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[315]), .B(A[315]), .Z(n546) );
  XOR U820 ( .A(A[314]), .B(n547), .Z(O[314]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[314]), .B(A[314]), .Z(n548) );
  XOR U823 ( .A(A[313]), .B(n549), .Z(O[313]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[313]), .B(A[313]), .Z(n550) );
  XOR U826 ( .A(A[312]), .B(n551), .Z(O[312]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[312]), .B(A[312]), .Z(n552) );
  XOR U829 ( .A(A[311]), .B(n553), .Z(O[311]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[311]), .B(A[311]), .Z(n554) );
  XOR U832 ( .A(A[310]), .B(n555), .Z(O[310]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[310]), .B(A[310]), .Z(n556) );
  XOR U835 ( .A(A[30]), .B(n557), .Z(O[30]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[30]), .B(A[30]), .Z(n558) );
  XOR U838 ( .A(A[309]), .B(n559), .Z(O[309]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[309]), .B(A[309]), .Z(n560) );
  XOR U841 ( .A(A[308]), .B(n561), .Z(O[308]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[308]), .B(A[308]), .Z(n562) );
  XOR U844 ( .A(A[307]), .B(n563), .Z(O[307]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[307]), .B(A[307]), .Z(n564) );
  XOR U847 ( .A(A[306]), .B(n565), .Z(O[306]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[306]), .B(A[306]), .Z(n566) );
  XOR U850 ( .A(A[305]), .B(n567), .Z(O[305]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[305]), .B(A[305]), .Z(n568) );
  XOR U853 ( .A(A[304]), .B(n569), .Z(O[304]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[304]), .B(A[304]), .Z(n570) );
  XOR U856 ( .A(A[303]), .B(n571), .Z(O[303]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[303]), .B(A[303]), .Z(n572) );
  XOR U859 ( .A(A[302]), .B(n573), .Z(O[302]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[302]), .B(A[302]), .Z(n574) );
  XOR U862 ( .A(A[301]), .B(n575), .Z(O[301]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[301]), .B(A[301]), .Z(n576) );
  XOR U865 ( .A(A[300]), .B(n577), .Z(O[300]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[300]), .B(A[300]), .Z(n578) );
  XOR U868 ( .A(A[2]), .B(n579), .Z(O[2]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[2]), .B(A[2]), .Z(n580) );
  XOR U871 ( .A(A[29]), .B(n581), .Z(O[29]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[29]), .B(A[29]), .Z(n582) );
  XOR U874 ( .A(A[299]), .B(n583), .Z(O[299]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[299]), .B(A[299]), .Z(n584) );
  XOR U877 ( .A(A[298]), .B(n585), .Z(O[298]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[298]), .B(A[298]), .Z(n586) );
  XOR U880 ( .A(A[297]), .B(n587), .Z(O[297]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[297]), .B(A[297]), .Z(n588) );
  XOR U883 ( .A(A[296]), .B(n589), .Z(O[296]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[296]), .B(A[296]), .Z(n590) );
  XOR U886 ( .A(A[295]), .B(n591), .Z(O[295]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[295]), .B(A[295]), .Z(n592) );
  XOR U889 ( .A(A[294]), .B(n593), .Z(O[294]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[294]), .B(A[294]), .Z(n594) );
  XOR U892 ( .A(A[293]), .B(n595), .Z(O[293]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[293]), .B(A[293]), .Z(n596) );
  XOR U895 ( .A(A[292]), .B(n597), .Z(O[292]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[292]), .B(A[292]), .Z(n598) );
  XOR U898 ( .A(A[291]), .B(n599), .Z(O[291]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[291]), .B(A[291]), .Z(n600) );
  XOR U901 ( .A(A[290]), .B(n601), .Z(O[290]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[290]), .B(A[290]), .Z(n602) );
  XOR U904 ( .A(A[28]), .B(n603), .Z(O[28]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[28]), .B(A[28]), .Z(n604) );
  XOR U907 ( .A(A[289]), .B(n605), .Z(O[289]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[289]), .B(A[289]), .Z(n606) );
  XOR U910 ( .A(A[288]), .B(n607), .Z(O[288]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[288]), .B(A[288]), .Z(n608) );
  XOR U913 ( .A(A[287]), .B(n609), .Z(O[287]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[287]), .B(A[287]), .Z(n610) );
  XOR U916 ( .A(A[286]), .B(n611), .Z(O[286]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[286]), .B(A[286]), .Z(n612) );
  XOR U919 ( .A(A[285]), .B(n613), .Z(O[285]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[285]), .B(A[285]), .Z(n614) );
  XOR U922 ( .A(A[284]), .B(n615), .Z(O[284]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[284]), .B(A[284]), .Z(n616) );
  XOR U925 ( .A(A[283]), .B(n617), .Z(O[283]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[283]), .B(A[283]), .Z(n618) );
  XOR U928 ( .A(A[282]), .B(n619), .Z(O[282]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[282]), .B(A[282]), .Z(n620) );
  XOR U931 ( .A(A[281]), .B(n621), .Z(O[281]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[281]), .B(A[281]), .Z(n622) );
  XOR U934 ( .A(A[280]), .B(n623), .Z(O[280]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[280]), .B(A[280]), .Z(n624) );
  XOR U937 ( .A(A[27]), .B(n625), .Z(O[27]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[27]), .B(A[27]), .Z(n626) );
  XOR U940 ( .A(A[279]), .B(n627), .Z(O[279]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[279]), .B(A[279]), .Z(n628) );
  XOR U943 ( .A(A[278]), .B(n629), .Z(O[278]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[278]), .B(A[278]), .Z(n630) );
  XOR U946 ( .A(A[277]), .B(n631), .Z(O[277]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[277]), .B(A[277]), .Z(n632) );
  XOR U949 ( .A(A[276]), .B(n633), .Z(O[276]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[276]), .B(A[276]), .Z(n634) );
  XOR U952 ( .A(A[275]), .B(n635), .Z(O[275]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[275]), .B(A[275]), .Z(n636) );
  XOR U955 ( .A(A[274]), .B(n637), .Z(O[274]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[274]), .B(A[274]), .Z(n638) );
  XOR U958 ( .A(A[273]), .B(n639), .Z(O[273]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[273]), .B(A[273]), .Z(n640) );
  XOR U961 ( .A(A[272]), .B(n641), .Z(O[272]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[272]), .B(A[272]), .Z(n642) );
  XOR U964 ( .A(A[271]), .B(n643), .Z(O[271]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[271]), .B(A[271]), .Z(n644) );
  XOR U967 ( .A(A[270]), .B(n645), .Z(O[270]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[270]), .B(A[270]), .Z(n646) );
  XOR U970 ( .A(A[26]), .B(n647), .Z(O[26]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[26]), .B(A[26]), .Z(n648) );
  XOR U973 ( .A(A[269]), .B(n649), .Z(O[269]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[269]), .B(A[269]), .Z(n650) );
  XOR U976 ( .A(A[268]), .B(n651), .Z(O[268]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[268]), .B(A[268]), .Z(n652) );
  XOR U979 ( .A(A[267]), .B(n653), .Z(O[267]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[267]), .B(A[267]), .Z(n654) );
  XOR U982 ( .A(A[266]), .B(n655), .Z(O[266]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[266]), .B(A[266]), .Z(n656) );
  XOR U985 ( .A(A[265]), .B(n657), .Z(O[265]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[265]), .B(A[265]), .Z(n658) );
  XOR U988 ( .A(A[264]), .B(n659), .Z(O[264]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[264]), .B(A[264]), .Z(n660) );
  XOR U991 ( .A(A[263]), .B(n661), .Z(O[263]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[263]), .B(A[263]), .Z(n662) );
  XOR U994 ( .A(A[262]), .B(n663), .Z(O[262]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[262]), .B(A[262]), .Z(n664) );
  XOR U997 ( .A(A[261]), .B(n665), .Z(O[261]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[261]), .B(A[261]), .Z(n666) );
  XOR U1000 ( .A(A[260]), .B(n667), .Z(O[260]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[260]), .B(A[260]), .Z(n668) );
  XOR U1003 ( .A(A[25]), .B(n669), .Z(O[25]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[25]), .B(A[25]), .Z(n670) );
  XOR U1006 ( .A(A[259]), .B(n671), .Z(O[259]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[259]), .B(A[259]), .Z(n672) );
  XOR U1009 ( .A(A[258]), .B(n673), .Z(O[258]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[258]), .B(A[258]), .Z(n674) );
  XOR U1012 ( .A(A[257]), .B(n675), .Z(O[257]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[257]), .B(A[257]), .Z(n676) );
  XOR U1015 ( .A(A[256]), .B(n677), .Z(O[256]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[256]), .B(A[256]), .Z(n678) );
  XOR U1018 ( .A(A[255]), .B(n679), .Z(O[255]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[255]), .B(A[255]), .Z(n680) );
  XOR U1021 ( .A(A[254]), .B(n681), .Z(O[254]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[254]), .B(A[254]), .Z(n682) );
  XOR U1024 ( .A(A[253]), .B(n683), .Z(O[253]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[253]), .B(A[253]), .Z(n684) );
  XOR U1027 ( .A(A[252]), .B(n685), .Z(O[252]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[252]), .B(A[252]), .Z(n686) );
  XOR U1030 ( .A(A[251]), .B(n687), .Z(O[251]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[251]), .B(A[251]), .Z(n688) );
  XOR U1033 ( .A(A[250]), .B(n689), .Z(O[250]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[250]), .B(A[250]), .Z(n690) );
  XOR U1036 ( .A(A[24]), .B(n691), .Z(O[24]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[24]), .B(A[24]), .Z(n692) );
  XOR U1039 ( .A(A[249]), .B(n693), .Z(O[249]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[249]), .B(A[249]), .Z(n694) );
  XOR U1042 ( .A(A[248]), .B(n695), .Z(O[248]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[248]), .B(A[248]), .Z(n696) );
  XOR U1045 ( .A(A[247]), .B(n697), .Z(O[247]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[247]), .B(A[247]), .Z(n698) );
  XOR U1048 ( .A(A[246]), .B(n699), .Z(O[246]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[246]), .B(A[246]), .Z(n700) );
  XOR U1051 ( .A(A[245]), .B(n701), .Z(O[245]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[245]), .B(A[245]), .Z(n702) );
  XOR U1054 ( .A(A[244]), .B(n703), .Z(O[244]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[244]), .B(A[244]), .Z(n704) );
  XOR U1057 ( .A(A[243]), .B(n705), .Z(O[243]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[243]), .B(A[243]), .Z(n706) );
  XOR U1060 ( .A(A[242]), .B(n707), .Z(O[242]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[242]), .B(A[242]), .Z(n708) );
  XOR U1063 ( .A(A[241]), .B(n709), .Z(O[241]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[241]), .B(A[241]), .Z(n710) );
  XOR U1066 ( .A(A[240]), .B(n711), .Z(O[240]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[240]), .B(A[240]), .Z(n712) );
  XOR U1069 ( .A(A[23]), .B(n713), .Z(O[23]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[23]), .B(A[23]), .Z(n714) );
  XOR U1072 ( .A(A[239]), .B(n715), .Z(O[239]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[239]), .B(A[239]), .Z(n716) );
  XOR U1075 ( .A(A[238]), .B(n717), .Z(O[238]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[238]), .B(A[238]), .Z(n718) );
  XOR U1078 ( .A(A[237]), .B(n719), .Z(O[237]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[237]), .B(A[237]), .Z(n720) );
  XOR U1081 ( .A(A[236]), .B(n721), .Z(O[236]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[236]), .B(A[236]), .Z(n722) );
  XOR U1084 ( .A(A[235]), .B(n723), .Z(O[235]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[235]), .B(A[235]), .Z(n724) );
  XOR U1087 ( .A(A[234]), .B(n725), .Z(O[234]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[234]), .B(A[234]), .Z(n726) );
  XOR U1090 ( .A(A[233]), .B(n727), .Z(O[233]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[233]), .B(A[233]), .Z(n728) );
  XOR U1093 ( .A(A[232]), .B(n729), .Z(O[232]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[232]), .B(A[232]), .Z(n730) );
  XOR U1096 ( .A(A[231]), .B(n731), .Z(O[231]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[231]), .B(A[231]), .Z(n732) );
  XOR U1099 ( .A(A[230]), .B(n733), .Z(O[230]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[230]), .B(A[230]), .Z(n734) );
  XOR U1102 ( .A(A[22]), .B(n735), .Z(O[22]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[22]), .B(A[22]), .Z(n736) );
  XOR U1105 ( .A(A[229]), .B(n737), .Z(O[229]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[229]), .B(A[229]), .Z(n738) );
  XOR U1108 ( .A(A[228]), .B(n739), .Z(O[228]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[228]), .B(A[228]), .Z(n740) );
  XOR U1111 ( .A(A[227]), .B(n741), .Z(O[227]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[227]), .B(A[227]), .Z(n742) );
  XOR U1114 ( .A(A[226]), .B(n743), .Z(O[226]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[226]), .B(A[226]), .Z(n744) );
  XOR U1117 ( .A(A[225]), .B(n745), .Z(O[225]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[225]), .B(A[225]), .Z(n746) );
  XOR U1120 ( .A(A[224]), .B(n747), .Z(O[224]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[224]), .B(A[224]), .Z(n748) );
  XOR U1123 ( .A(A[223]), .B(n749), .Z(O[223]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[223]), .B(A[223]), .Z(n750) );
  XOR U1126 ( .A(A[222]), .B(n751), .Z(O[222]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[222]), .B(A[222]), .Z(n752) );
  XOR U1129 ( .A(A[221]), .B(n753), .Z(O[221]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[221]), .B(A[221]), .Z(n754) );
  XOR U1132 ( .A(A[220]), .B(n755), .Z(O[220]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[220]), .B(A[220]), .Z(n756) );
  XOR U1135 ( .A(A[21]), .B(n757), .Z(O[21]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[21]), .B(A[21]), .Z(n758) );
  XOR U1138 ( .A(A[219]), .B(n759), .Z(O[219]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[219]), .B(A[219]), .Z(n760) );
  XOR U1141 ( .A(A[218]), .B(n761), .Z(O[218]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[218]), .B(A[218]), .Z(n762) );
  XOR U1144 ( .A(A[217]), .B(n763), .Z(O[217]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[217]), .B(A[217]), .Z(n764) );
  XOR U1147 ( .A(A[216]), .B(n765), .Z(O[216]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[216]), .B(A[216]), .Z(n766) );
  XOR U1150 ( .A(A[215]), .B(n767), .Z(O[215]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[215]), .B(A[215]), .Z(n768) );
  XOR U1153 ( .A(A[214]), .B(n769), .Z(O[214]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[214]), .B(A[214]), .Z(n770) );
  XOR U1156 ( .A(A[213]), .B(n771), .Z(O[213]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[213]), .B(A[213]), .Z(n772) );
  XOR U1159 ( .A(A[212]), .B(n773), .Z(O[212]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[212]), .B(A[212]), .Z(n774) );
  XOR U1162 ( .A(A[211]), .B(n775), .Z(O[211]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[211]), .B(A[211]), .Z(n776) );
  XOR U1165 ( .A(A[210]), .B(n777), .Z(O[210]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[210]), .B(A[210]), .Z(n778) );
  XOR U1168 ( .A(A[20]), .B(n779), .Z(O[20]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[20]), .B(A[20]), .Z(n780) );
  XOR U1171 ( .A(A[209]), .B(n781), .Z(O[209]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[209]), .B(A[209]), .Z(n782) );
  XOR U1174 ( .A(A[208]), .B(n783), .Z(O[208]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[208]), .B(A[208]), .Z(n784) );
  XOR U1177 ( .A(A[207]), .B(n785), .Z(O[207]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[207]), .B(A[207]), .Z(n786) );
  XOR U1180 ( .A(A[206]), .B(n787), .Z(O[206]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[206]), .B(A[206]), .Z(n788) );
  XOR U1183 ( .A(A[205]), .B(n789), .Z(O[205]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[205]), .B(A[205]), .Z(n790) );
  XOR U1186 ( .A(A[204]), .B(n791), .Z(O[204]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[204]), .B(A[204]), .Z(n792) );
  XOR U1189 ( .A(A[203]), .B(n793), .Z(O[203]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[203]), .B(A[203]), .Z(n794) );
  XOR U1192 ( .A(A[202]), .B(n795), .Z(O[202]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[202]), .B(A[202]), .Z(n796) );
  XOR U1195 ( .A(A[201]), .B(n797), .Z(O[201]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[201]), .B(A[201]), .Z(n798) );
  XOR U1198 ( .A(A[200]), .B(n799), .Z(O[200]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[200]), .B(A[200]), .Z(n800) );
  XOR U1201 ( .A(A[1]), .B(n801), .Z(O[1]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[1]), .B(A[1]), .Z(n802) );
  XOR U1204 ( .A(A[19]), .B(n803), .Z(O[19]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[19]), .B(A[19]), .Z(n804) );
  XOR U1207 ( .A(A[199]), .B(n805), .Z(O[199]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[199]), .B(A[199]), .Z(n806) );
  XOR U1210 ( .A(A[198]), .B(n807), .Z(O[198]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[198]), .B(A[198]), .Z(n808) );
  XOR U1213 ( .A(A[197]), .B(n809), .Z(O[197]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[197]), .B(A[197]), .Z(n810) );
  XOR U1216 ( .A(A[196]), .B(n811), .Z(O[196]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[196]), .B(A[196]), .Z(n812) );
  XOR U1219 ( .A(A[195]), .B(n813), .Z(O[195]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[195]), .B(A[195]), .Z(n814) );
  XOR U1222 ( .A(A[194]), .B(n815), .Z(O[194]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[194]), .B(A[194]), .Z(n816) );
  XOR U1225 ( .A(A[193]), .B(n817), .Z(O[193]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[193]), .B(A[193]), .Z(n818) );
  XOR U1228 ( .A(A[192]), .B(n819), .Z(O[192]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[192]), .B(A[192]), .Z(n820) );
  XOR U1231 ( .A(A[191]), .B(n821), .Z(O[191]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[191]), .B(A[191]), .Z(n822) );
  XOR U1234 ( .A(A[190]), .B(n823), .Z(O[190]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[190]), .B(A[190]), .Z(n824) );
  XOR U1237 ( .A(A[18]), .B(n825), .Z(O[18]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[18]), .B(A[18]), .Z(n826) );
  XOR U1240 ( .A(A[189]), .B(n827), .Z(O[189]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[189]), .B(A[189]), .Z(n828) );
  XOR U1243 ( .A(A[188]), .B(n829), .Z(O[188]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[188]), .B(A[188]), .Z(n830) );
  XOR U1246 ( .A(A[187]), .B(n831), .Z(O[187]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[187]), .B(A[187]), .Z(n832) );
  XOR U1249 ( .A(A[186]), .B(n833), .Z(O[186]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[186]), .B(A[186]), .Z(n834) );
  XOR U1252 ( .A(A[185]), .B(n835), .Z(O[185]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[185]), .B(A[185]), .Z(n836) );
  XOR U1255 ( .A(A[184]), .B(n837), .Z(O[184]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[184]), .B(A[184]), .Z(n838) );
  XOR U1258 ( .A(A[183]), .B(n839), .Z(O[183]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[183]), .B(A[183]), .Z(n840) );
  XOR U1261 ( .A(A[182]), .B(n841), .Z(O[182]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[182]), .B(A[182]), .Z(n842) );
  XOR U1264 ( .A(A[181]), .B(n843), .Z(O[181]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[181]), .B(A[181]), .Z(n844) );
  XOR U1267 ( .A(A[180]), .B(n845), .Z(O[180]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[180]), .B(A[180]), .Z(n846) );
  XOR U1270 ( .A(A[17]), .B(n847), .Z(O[17]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[17]), .B(A[17]), .Z(n848) );
  XOR U1273 ( .A(A[179]), .B(n849), .Z(O[179]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[179]), .B(A[179]), .Z(n850) );
  XOR U1276 ( .A(A[178]), .B(n851), .Z(O[178]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[178]), .B(A[178]), .Z(n852) );
  XOR U1279 ( .A(A[177]), .B(n853), .Z(O[177]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[177]), .B(A[177]), .Z(n854) );
  XOR U1282 ( .A(A[176]), .B(n855), .Z(O[176]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[176]), .B(A[176]), .Z(n856) );
  XOR U1285 ( .A(A[175]), .B(n857), .Z(O[175]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[175]), .B(A[175]), .Z(n858) );
  XOR U1288 ( .A(A[174]), .B(n859), .Z(O[174]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[174]), .B(A[174]), .Z(n860) );
  XOR U1291 ( .A(A[173]), .B(n861), .Z(O[173]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[173]), .B(A[173]), .Z(n862) );
  XOR U1294 ( .A(A[172]), .B(n863), .Z(O[172]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[172]), .B(A[172]), .Z(n864) );
  XOR U1297 ( .A(A[171]), .B(n865), .Z(O[171]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[171]), .B(A[171]), .Z(n866) );
  XOR U1300 ( .A(A[170]), .B(n867), .Z(O[170]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[170]), .B(A[170]), .Z(n868) );
  XOR U1303 ( .A(A[16]), .B(n869), .Z(O[16]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[16]), .B(A[16]), .Z(n870) );
  XOR U1306 ( .A(A[169]), .B(n871), .Z(O[169]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[169]), .B(A[169]), .Z(n872) );
  XOR U1309 ( .A(A[168]), .B(n873), .Z(O[168]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[168]), .B(A[168]), .Z(n874) );
  XOR U1312 ( .A(A[167]), .B(n875), .Z(O[167]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[167]), .B(A[167]), .Z(n876) );
  XOR U1315 ( .A(A[166]), .B(n877), .Z(O[166]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[166]), .B(A[166]), .Z(n878) );
  XOR U1318 ( .A(A[165]), .B(n879), .Z(O[165]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[165]), .B(A[165]), .Z(n880) );
  XOR U1321 ( .A(A[164]), .B(n881), .Z(O[164]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[164]), .B(A[164]), .Z(n882) );
  XOR U1324 ( .A(A[163]), .B(n883), .Z(O[163]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[163]), .B(A[163]), .Z(n884) );
  XOR U1327 ( .A(A[162]), .B(n885), .Z(O[162]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[162]), .B(A[162]), .Z(n886) );
  XOR U1330 ( .A(A[161]), .B(n887), .Z(O[161]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[161]), .B(A[161]), .Z(n888) );
  XOR U1333 ( .A(A[160]), .B(n889), .Z(O[160]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[160]), .B(A[160]), .Z(n890) );
  XOR U1336 ( .A(A[15]), .B(n891), .Z(O[15]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[15]), .B(A[15]), .Z(n892) );
  XOR U1339 ( .A(A[159]), .B(n893), .Z(O[159]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[159]), .B(A[159]), .Z(n894) );
  XOR U1342 ( .A(A[158]), .B(n895), .Z(O[158]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[158]), .B(A[158]), .Z(n896) );
  XOR U1345 ( .A(A[157]), .B(n897), .Z(O[157]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[157]), .B(A[157]), .Z(n898) );
  XOR U1348 ( .A(A[156]), .B(n899), .Z(O[156]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[156]), .B(A[156]), .Z(n900) );
  XOR U1351 ( .A(A[155]), .B(n901), .Z(O[155]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[155]), .B(A[155]), .Z(n902) );
  XOR U1354 ( .A(A[154]), .B(n903), .Z(O[154]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[154]), .B(A[154]), .Z(n904) );
  XOR U1357 ( .A(A[153]), .B(n905), .Z(O[153]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[153]), .B(A[153]), .Z(n906) );
  XOR U1360 ( .A(A[152]), .B(n907), .Z(O[152]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[152]), .B(A[152]), .Z(n908) );
  XOR U1363 ( .A(A[151]), .B(n909), .Z(O[151]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[151]), .B(A[151]), .Z(n910) );
  XOR U1366 ( .A(A[150]), .B(n911), .Z(O[150]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[150]), .B(A[150]), .Z(n912) );
  XOR U1369 ( .A(A[14]), .B(n913), .Z(O[14]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[14]), .B(A[14]), .Z(n914) );
  XOR U1372 ( .A(A[149]), .B(n915), .Z(O[149]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[149]), .B(A[149]), .Z(n916) );
  XOR U1375 ( .A(A[148]), .B(n917), .Z(O[148]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[148]), .B(A[148]), .Z(n918) );
  XOR U1378 ( .A(A[147]), .B(n919), .Z(O[147]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[147]), .B(A[147]), .Z(n920) );
  XOR U1381 ( .A(A[146]), .B(n921), .Z(O[146]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[146]), .B(A[146]), .Z(n922) );
  XOR U1384 ( .A(A[145]), .B(n923), .Z(O[145]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[145]), .B(A[145]), .Z(n924) );
  XOR U1387 ( .A(A[144]), .B(n925), .Z(O[144]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[144]), .B(A[144]), .Z(n926) );
  XOR U1390 ( .A(A[143]), .B(n927), .Z(O[143]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[143]), .B(A[143]), .Z(n928) );
  XOR U1393 ( .A(A[142]), .B(n929), .Z(O[142]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[142]), .B(A[142]), .Z(n930) );
  XOR U1396 ( .A(A[141]), .B(n931), .Z(O[141]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[141]), .B(A[141]), .Z(n932) );
  XOR U1399 ( .A(A[140]), .B(n933), .Z(O[140]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[140]), .B(A[140]), .Z(n934) );
  XOR U1402 ( .A(A[13]), .B(n935), .Z(O[13]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[13]), .B(A[13]), .Z(n936) );
  XOR U1405 ( .A(A[139]), .B(n937), .Z(O[139]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[139]), .B(A[139]), .Z(n938) );
  XOR U1408 ( .A(A[138]), .B(n939), .Z(O[138]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[138]), .B(A[138]), .Z(n940) );
  XOR U1411 ( .A(A[137]), .B(n941), .Z(O[137]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[137]), .B(A[137]), .Z(n942) );
  XOR U1414 ( .A(A[136]), .B(n943), .Z(O[136]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[136]), .B(A[136]), .Z(n944) );
  XOR U1417 ( .A(A[135]), .B(n945), .Z(O[135]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[135]), .B(A[135]), .Z(n946) );
  XOR U1420 ( .A(A[134]), .B(n947), .Z(O[134]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[134]), .B(A[134]), .Z(n948) );
  XOR U1423 ( .A(A[133]), .B(n949), .Z(O[133]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[133]), .B(A[133]), .Z(n950) );
  XOR U1426 ( .A(A[132]), .B(n951), .Z(O[132]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[132]), .B(A[132]), .Z(n952) );
  XOR U1429 ( .A(A[131]), .B(n953), .Z(O[131]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[131]), .B(A[131]), .Z(n954) );
  XOR U1432 ( .A(A[130]), .B(n955), .Z(O[130]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[130]), .B(A[130]), .Z(n956) );
  XOR U1435 ( .A(A[12]), .B(n957), .Z(O[12]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[12]), .B(A[12]), .Z(n958) );
  XOR U1438 ( .A(A[129]), .B(n959), .Z(O[129]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[129]), .B(A[129]), .Z(n960) );
  XOR U1441 ( .A(A[128]), .B(n961), .Z(O[128]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[128]), .B(A[128]), .Z(n962) );
  XOR U1444 ( .A(A[127]), .B(n963), .Z(O[127]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[127]), .B(A[127]), .Z(n964) );
  XOR U1447 ( .A(A[126]), .B(n965), .Z(O[126]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[126]), .B(A[126]), .Z(n966) );
  XOR U1450 ( .A(A[125]), .B(n967), .Z(O[125]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[125]), .B(A[125]), .Z(n968) );
  XOR U1453 ( .A(A[124]), .B(n969), .Z(O[124]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[124]), .B(A[124]), .Z(n970) );
  XOR U1456 ( .A(A[123]), .B(n971), .Z(O[123]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[123]), .B(A[123]), .Z(n972) );
  XOR U1459 ( .A(A[122]), .B(n973), .Z(O[122]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[122]), .B(A[122]), .Z(n974) );
  XOR U1462 ( .A(A[121]), .B(n975), .Z(O[121]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[121]), .B(A[121]), .Z(n976) );
  XOR U1465 ( .A(A[120]), .B(n977), .Z(O[120]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[120]), .B(A[120]), .Z(n978) );
  XOR U1468 ( .A(A[11]), .B(n979), .Z(O[11]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[11]), .B(A[11]), .Z(n980) );
  XOR U1471 ( .A(A[119]), .B(n981), .Z(O[119]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[119]), .B(A[119]), .Z(n982) );
  XOR U1474 ( .A(A[118]), .B(n983), .Z(O[118]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[118]), .B(A[118]), .Z(n984) );
  XOR U1477 ( .A(A[117]), .B(n985), .Z(O[117]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[117]), .B(A[117]), .Z(n986) );
  XOR U1480 ( .A(A[116]), .B(n987), .Z(O[116]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[116]), .B(A[116]), .Z(n988) );
  XOR U1483 ( .A(A[115]), .B(n989), .Z(O[115]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[115]), .B(A[115]), .Z(n990) );
  XOR U1486 ( .A(A[114]), .B(n991), .Z(O[114]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[114]), .B(A[114]), .Z(n992) );
  XOR U1489 ( .A(A[113]), .B(n993), .Z(O[113]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[113]), .B(A[113]), .Z(n994) );
  XOR U1492 ( .A(A[112]), .B(n995), .Z(O[112]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[112]), .B(A[112]), .Z(n996) );
  XOR U1495 ( .A(A[111]), .B(n997), .Z(O[111]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[111]), .B(A[111]), .Z(n998) );
  XOR U1498 ( .A(A[110]), .B(n999), .Z(O[110]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[110]), .B(A[110]), .Z(n1000) );
  XOR U1501 ( .A(A[10]), .B(n1001), .Z(O[10]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[10]), .B(A[10]), .Z(n1002) );
  XOR U1504 ( .A(A[109]), .B(n1003), .Z(O[109]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[109]), .B(A[109]), .Z(n1004) );
  XOR U1507 ( .A(A[108]), .B(n1005), .Z(O[108]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[108]), .B(A[108]), .Z(n1006) );
  XOR U1510 ( .A(A[107]), .B(n1007), .Z(O[107]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[107]), .B(A[107]), .Z(n1008) );
  XOR U1513 ( .A(A[106]), .B(n1009), .Z(O[106]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[106]), .B(A[106]), .Z(n1010) );
  XOR U1516 ( .A(A[105]), .B(n1011), .Z(O[105]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[105]), .B(A[105]), .Z(n1012) );
  XOR U1519 ( .A(A[104]), .B(n1013), .Z(O[104]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[104]), .B(A[104]), .Z(n1014) );
  XOR U1522 ( .A(A[103]), .B(n1015), .Z(O[103]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[103]), .B(A[103]), .Z(n1016) );
  XOR U1525 ( .A(A[102]), .B(n1017), .Z(O[102]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[102]), .B(A[102]), .Z(n1018) );
  XOR U1528 ( .A(A[101]), .B(n1019), .Z(O[101]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[101]), .B(A[101]), .Z(n1020) );
  XOR U1531 ( .A(A[100]), .B(n1021), .Z(O[100]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[100]), .B(A[100]), .Z(n1022) );
  XOR U1534 ( .A(A[0]), .B(n1023), .Z(O[0]) );
  AND U1535 ( .A(S), .B(n1024), .Z(n1023) );
  XOR U1536 ( .A(B[0]), .B(A[0]), .Z(n1024) );
endmodule


module MUX_N512_5 ( A, B, S, O );
  input [511:0] A;
  input [511:0] B;
  output [511:0] O;
  input S;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  XOR U1 ( .A(B[8]), .B(n1), .Z(O[9]) );
  AND U2 ( .A(S), .B(n2), .Z(n1) );
  XOR U3 ( .A(B[9]), .B(B[8]), .Z(n2) );
  XOR U4 ( .A(B[98]), .B(n3), .Z(O[99]) );
  AND U5 ( .A(S), .B(n4), .Z(n3) );
  XOR U6 ( .A(B[99]), .B(B[98]), .Z(n4) );
  XOR U7 ( .A(B[97]), .B(n5), .Z(O[98]) );
  AND U8 ( .A(S), .B(n6), .Z(n5) );
  XOR U9 ( .A(B[98]), .B(B[97]), .Z(n6) );
  XOR U10 ( .A(B[96]), .B(n7), .Z(O[97]) );
  AND U11 ( .A(S), .B(n8), .Z(n7) );
  XOR U12 ( .A(B[97]), .B(B[96]), .Z(n8) );
  XOR U13 ( .A(B[95]), .B(n9), .Z(O[96]) );
  AND U14 ( .A(S), .B(n10), .Z(n9) );
  XOR U15 ( .A(B[96]), .B(B[95]), .Z(n10) );
  XOR U16 ( .A(B[94]), .B(n11), .Z(O[95]) );
  AND U17 ( .A(S), .B(n12), .Z(n11) );
  XOR U18 ( .A(B[95]), .B(B[94]), .Z(n12) );
  XOR U19 ( .A(B[93]), .B(n13), .Z(O[94]) );
  AND U20 ( .A(S), .B(n14), .Z(n13) );
  XOR U21 ( .A(B[94]), .B(B[93]), .Z(n14) );
  XOR U22 ( .A(B[92]), .B(n15), .Z(O[93]) );
  AND U23 ( .A(S), .B(n16), .Z(n15) );
  XOR U24 ( .A(B[93]), .B(B[92]), .Z(n16) );
  XOR U25 ( .A(B[91]), .B(n17), .Z(O[92]) );
  AND U26 ( .A(S), .B(n18), .Z(n17) );
  XOR U27 ( .A(B[92]), .B(B[91]), .Z(n18) );
  XOR U28 ( .A(B[90]), .B(n19), .Z(O[91]) );
  AND U29 ( .A(S), .B(n20), .Z(n19) );
  XOR U30 ( .A(B[91]), .B(B[90]), .Z(n20) );
  XOR U31 ( .A(B[89]), .B(n21), .Z(O[90]) );
  AND U32 ( .A(S), .B(n22), .Z(n21) );
  XOR U33 ( .A(B[90]), .B(B[89]), .Z(n22) );
  XOR U34 ( .A(B[7]), .B(n23), .Z(O[8]) );
  AND U35 ( .A(S), .B(n24), .Z(n23) );
  XOR U36 ( .A(B[8]), .B(B[7]), .Z(n24) );
  XOR U37 ( .A(B[88]), .B(n25), .Z(O[89]) );
  AND U38 ( .A(S), .B(n26), .Z(n25) );
  XOR U39 ( .A(B[89]), .B(B[88]), .Z(n26) );
  XOR U40 ( .A(B[87]), .B(n27), .Z(O[88]) );
  AND U41 ( .A(S), .B(n28), .Z(n27) );
  XOR U42 ( .A(B[88]), .B(B[87]), .Z(n28) );
  XOR U43 ( .A(B[86]), .B(n29), .Z(O[87]) );
  AND U44 ( .A(S), .B(n30), .Z(n29) );
  XOR U45 ( .A(B[87]), .B(B[86]), .Z(n30) );
  XOR U46 ( .A(B[85]), .B(n31), .Z(O[86]) );
  AND U47 ( .A(S), .B(n32), .Z(n31) );
  XOR U48 ( .A(B[86]), .B(B[85]), .Z(n32) );
  XOR U49 ( .A(B[84]), .B(n33), .Z(O[85]) );
  AND U50 ( .A(S), .B(n34), .Z(n33) );
  XOR U51 ( .A(B[85]), .B(B[84]), .Z(n34) );
  XOR U52 ( .A(B[83]), .B(n35), .Z(O[84]) );
  AND U53 ( .A(S), .B(n36), .Z(n35) );
  XOR U54 ( .A(B[84]), .B(B[83]), .Z(n36) );
  XOR U55 ( .A(B[82]), .B(n37), .Z(O[83]) );
  AND U56 ( .A(S), .B(n38), .Z(n37) );
  XOR U57 ( .A(B[83]), .B(B[82]), .Z(n38) );
  XOR U58 ( .A(B[81]), .B(n39), .Z(O[82]) );
  AND U59 ( .A(S), .B(n40), .Z(n39) );
  XOR U60 ( .A(B[82]), .B(B[81]), .Z(n40) );
  XOR U61 ( .A(B[80]), .B(n41), .Z(O[81]) );
  AND U62 ( .A(S), .B(n42), .Z(n41) );
  XOR U63 ( .A(B[81]), .B(B[80]), .Z(n42) );
  XOR U64 ( .A(B[79]), .B(n43), .Z(O[80]) );
  AND U65 ( .A(S), .B(n44), .Z(n43) );
  XOR U66 ( .A(B[80]), .B(B[79]), .Z(n44) );
  XOR U67 ( .A(B[6]), .B(n45), .Z(O[7]) );
  AND U68 ( .A(S), .B(n46), .Z(n45) );
  XOR U69 ( .A(B[7]), .B(B[6]), .Z(n46) );
  XOR U70 ( .A(B[78]), .B(n47), .Z(O[79]) );
  AND U71 ( .A(S), .B(n48), .Z(n47) );
  XOR U72 ( .A(B[79]), .B(B[78]), .Z(n48) );
  XOR U73 ( .A(B[77]), .B(n49), .Z(O[78]) );
  AND U74 ( .A(S), .B(n50), .Z(n49) );
  XOR U75 ( .A(B[78]), .B(B[77]), .Z(n50) );
  XOR U76 ( .A(B[76]), .B(n51), .Z(O[77]) );
  AND U77 ( .A(S), .B(n52), .Z(n51) );
  XOR U78 ( .A(B[77]), .B(B[76]), .Z(n52) );
  XOR U79 ( .A(B[75]), .B(n53), .Z(O[76]) );
  AND U80 ( .A(S), .B(n54), .Z(n53) );
  XOR U81 ( .A(B[76]), .B(B[75]), .Z(n54) );
  XOR U82 ( .A(B[74]), .B(n55), .Z(O[75]) );
  AND U83 ( .A(S), .B(n56), .Z(n55) );
  XOR U84 ( .A(B[75]), .B(B[74]), .Z(n56) );
  XOR U85 ( .A(B[73]), .B(n57), .Z(O[74]) );
  AND U86 ( .A(S), .B(n58), .Z(n57) );
  XOR U87 ( .A(B[74]), .B(B[73]), .Z(n58) );
  XOR U88 ( .A(B[72]), .B(n59), .Z(O[73]) );
  AND U89 ( .A(S), .B(n60), .Z(n59) );
  XOR U90 ( .A(B[73]), .B(B[72]), .Z(n60) );
  XOR U91 ( .A(B[71]), .B(n61), .Z(O[72]) );
  AND U92 ( .A(S), .B(n62), .Z(n61) );
  XOR U93 ( .A(B[72]), .B(B[71]), .Z(n62) );
  XOR U94 ( .A(B[70]), .B(n63), .Z(O[71]) );
  AND U95 ( .A(S), .B(n64), .Z(n63) );
  XOR U96 ( .A(B[71]), .B(B[70]), .Z(n64) );
  XOR U97 ( .A(B[69]), .B(n65), .Z(O[70]) );
  AND U98 ( .A(S), .B(n66), .Z(n65) );
  XOR U99 ( .A(B[70]), .B(B[69]), .Z(n66) );
  XOR U100 ( .A(B[5]), .B(n67), .Z(O[6]) );
  AND U101 ( .A(S), .B(n68), .Z(n67) );
  XOR U102 ( .A(B[6]), .B(B[5]), .Z(n68) );
  XOR U103 ( .A(B[68]), .B(n69), .Z(O[69]) );
  AND U104 ( .A(S), .B(n70), .Z(n69) );
  XOR U105 ( .A(B[69]), .B(B[68]), .Z(n70) );
  XOR U106 ( .A(B[67]), .B(n71), .Z(O[68]) );
  AND U107 ( .A(S), .B(n72), .Z(n71) );
  XOR U108 ( .A(B[68]), .B(B[67]), .Z(n72) );
  XOR U109 ( .A(B[66]), .B(n73), .Z(O[67]) );
  AND U110 ( .A(S), .B(n74), .Z(n73) );
  XOR U111 ( .A(B[67]), .B(B[66]), .Z(n74) );
  XOR U112 ( .A(B[65]), .B(n75), .Z(O[66]) );
  AND U113 ( .A(S), .B(n76), .Z(n75) );
  XOR U114 ( .A(B[66]), .B(B[65]), .Z(n76) );
  XOR U115 ( .A(B[64]), .B(n77), .Z(O[65]) );
  AND U116 ( .A(S), .B(n78), .Z(n77) );
  XOR U117 ( .A(B[65]), .B(B[64]), .Z(n78) );
  XOR U118 ( .A(B[63]), .B(n79), .Z(O[64]) );
  AND U119 ( .A(S), .B(n80), .Z(n79) );
  XOR U120 ( .A(B[64]), .B(B[63]), .Z(n80) );
  XOR U121 ( .A(B[62]), .B(n81), .Z(O[63]) );
  AND U122 ( .A(S), .B(n82), .Z(n81) );
  XOR U123 ( .A(B[63]), .B(B[62]), .Z(n82) );
  XOR U124 ( .A(B[61]), .B(n83), .Z(O[62]) );
  AND U125 ( .A(S), .B(n84), .Z(n83) );
  XOR U126 ( .A(B[62]), .B(B[61]), .Z(n84) );
  XOR U127 ( .A(B[60]), .B(n85), .Z(O[61]) );
  AND U128 ( .A(S), .B(n86), .Z(n85) );
  XOR U129 ( .A(B[61]), .B(B[60]), .Z(n86) );
  XOR U130 ( .A(B[59]), .B(n87), .Z(O[60]) );
  AND U131 ( .A(S), .B(n88), .Z(n87) );
  XOR U132 ( .A(B[60]), .B(B[59]), .Z(n88) );
  XOR U133 ( .A(B[4]), .B(n89), .Z(O[5]) );
  AND U134 ( .A(S), .B(n90), .Z(n89) );
  XOR U135 ( .A(B[5]), .B(B[4]), .Z(n90) );
  XOR U136 ( .A(B[58]), .B(n91), .Z(O[59]) );
  AND U137 ( .A(S), .B(n92), .Z(n91) );
  XOR U138 ( .A(B[59]), .B(B[58]), .Z(n92) );
  XOR U139 ( .A(B[57]), .B(n93), .Z(O[58]) );
  AND U140 ( .A(S), .B(n94), .Z(n93) );
  XOR U141 ( .A(B[58]), .B(B[57]), .Z(n94) );
  XOR U142 ( .A(B[56]), .B(n95), .Z(O[57]) );
  AND U143 ( .A(S), .B(n96), .Z(n95) );
  XOR U144 ( .A(B[57]), .B(B[56]), .Z(n96) );
  XOR U145 ( .A(B[55]), .B(n97), .Z(O[56]) );
  AND U146 ( .A(S), .B(n98), .Z(n97) );
  XOR U147 ( .A(B[56]), .B(B[55]), .Z(n98) );
  XOR U148 ( .A(B[54]), .B(n99), .Z(O[55]) );
  AND U149 ( .A(S), .B(n100), .Z(n99) );
  XOR U150 ( .A(B[55]), .B(B[54]), .Z(n100) );
  XOR U151 ( .A(B[53]), .B(n101), .Z(O[54]) );
  AND U152 ( .A(S), .B(n102), .Z(n101) );
  XOR U153 ( .A(B[54]), .B(B[53]), .Z(n102) );
  XOR U154 ( .A(B[52]), .B(n103), .Z(O[53]) );
  AND U155 ( .A(S), .B(n104), .Z(n103) );
  XOR U156 ( .A(B[53]), .B(B[52]), .Z(n104) );
  XOR U157 ( .A(B[51]), .B(n105), .Z(O[52]) );
  AND U158 ( .A(S), .B(n106), .Z(n105) );
  XOR U159 ( .A(B[52]), .B(B[51]), .Z(n106) );
  XOR U160 ( .A(B[50]), .B(n107), .Z(O[51]) );
  AND U161 ( .A(S), .B(n108), .Z(n107) );
  XOR U162 ( .A(B[51]), .B(B[50]), .Z(n108) );
  XOR U163 ( .A(B[510]), .B(n109), .Z(O[511]) );
  AND U164 ( .A(S), .B(n110), .Z(n109) );
  XOR U165 ( .A(B[511]), .B(B[510]), .Z(n110) );
  XOR U166 ( .A(B[509]), .B(n111), .Z(O[510]) );
  AND U167 ( .A(S), .B(n112), .Z(n111) );
  XOR U168 ( .A(B[510]), .B(B[509]), .Z(n112) );
  XOR U169 ( .A(B[49]), .B(n113), .Z(O[50]) );
  AND U170 ( .A(S), .B(n114), .Z(n113) );
  XOR U171 ( .A(B[50]), .B(B[49]), .Z(n114) );
  XOR U172 ( .A(B[508]), .B(n115), .Z(O[509]) );
  AND U173 ( .A(S), .B(n116), .Z(n115) );
  XOR U174 ( .A(B[509]), .B(B[508]), .Z(n116) );
  XOR U175 ( .A(B[507]), .B(n117), .Z(O[508]) );
  AND U176 ( .A(S), .B(n118), .Z(n117) );
  XOR U177 ( .A(B[508]), .B(B[507]), .Z(n118) );
  XOR U178 ( .A(B[506]), .B(n119), .Z(O[507]) );
  AND U179 ( .A(S), .B(n120), .Z(n119) );
  XOR U180 ( .A(B[507]), .B(B[506]), .Z(n120) );
  XOR U181 ( .A(B[505]), .B(n121), .Z(O[506]) );
  AND U182 ( .A(S), .B(n122), .Z(n121) );
  XOR U183 ( .A(B[506]), .B(B[505]), .Z(n122) );
  XOR U184 ( .A(B[504]), .B(n123), .Z(O[505]) );
  AND U185 ( .A(S), .B(n124), .Z(n123) );
  XOR U186 ( .A(B[505]), .B(B[504]), .Z(n124) );
  XOR U187 ( .A(B[503]), .B(n125), .Z(O[504]) );
  AND U188 ( .A(S), .B(n126), .Z(n125) );
  XOR U189 ( .A(B[504]), .B(B[503]), .Z(n126) );
  XOR U190 ( .A(B[502]), .B(n127), .Z(O[503]) );
  AND U191 ( .A(S), .B(n128), .Z(n127) );
  XOR U192 ( .A(B[503]), .B(B[502]), .Z(n128) );
  XOR U193 ( .A(B[501]), .B(n129), .Z(O[502]) );
  AND U194 ( .A(S), .B(n130), .Z(n129) );
  XOR U195 ( .A(B[502]), .B(B[501]), .Z(n130) );
  XOR U196 ( .A(B[500]), .B(n131), .Z(O[501]) );
  AND U197 ( .A(S), .B(n132), .Z(n131) );
  XOR U198 ( .A(B[501]), .B(B[500]), .Z(n132) );
  XOR U199 ( .A(B[499]), .B(n133), .Z(O[500]) );
  AND U200 ( .A(S), .B(n134), .Z(n133) );
  XOR U201 ( .A(B[500]), .B(B[499]), .Z(n134) );
  XOR U202 ( .A(B[3]), .B(n135), .Z(O[4]) );
  AND U203 ( .A(S), .B(n136), .Z(n135) );
  XOR U204 ( .A(B[4]), .B(B[3]), .Z(n136) );
  XOR U205 ( .A(B[48]), .B(n137), .Z(O[49]) );
  AND U206 ( .A(S), .B(n138), .Z(n137) );
  XOR U207 ( .A(B[49]), .B(B[48]), .Z(n138) );
  XOR U208 ( .A(B[498]), .B(n139), .Z(O[499]) );
  AND U209 ( .A(S), .B(n140), .Z(n139) );
  XOR U210 ( .A(B[499]), .B(B[498]), .Z(n140) );
  XOR U211 ( .A(B[497]), .B(n141), .Z(O[498]) );
  AND U212 ( .A(S), .B(n142), .Z(n141) );
  XOR U213 ( .A(B[498]), .B(B[497]), .Z(n142) );
  XOR U214 ( .A(B[496]), .B(n143), .Z(O[497]) );
  AND U215 ( .A(S), .B(n144), .Z(n143) );
  XOR U216 ( .A(B[497]), .B(B[496]), .Z(n144) );
  XOR U217 ( .A(B[495]), .B(n145), .Z(O[496]) );
  AND U218 ( .A(S), .B(n146), .Z(n145) );
  XOR U219 ( .A(B[496]), .B(B[495]), .Z(n146) );
  XOR U220 ( .A(B[494]), .B(n147), .Z(O[495]) );
  AND U221 ( .A(S), .B(n148), .Z(n147) );
  XOR U222 ( .A(B[495]), .B(B[494]), .Z(n148) );
  XOR U223 ( .A(B[493]), .B(n149), .Z(O[494]) );
  AND U224 ( .A(S), .B(n150), .Z(n149) );
  XOR U225 ( .A(B[494]), .B(B[493]), .Z(n150) );
  XOR U226 ( .A(B[492]), .B(n151), .Z(O[493]) );
  AND U227 ( .A(S), .B(n152), .Z(n151) );
  XOR U228 ( .A(B[493]), .B(B[492]), .Z(n152) );
  XOR U229 ( .A(B[491]), .B(n153), .Z(O[492]) );
  AND U230 ( .A(S), .B(n154), .Z(n153) );
  XOR U231 ( .A(B[492]), .B(B[491]), .Z(n154) );
  XOR U232 ( .A(B[490]), .B(n155), .Z(O[491]) );
  AND U233 ( .A(S), .B(n156), .Z(n155) );
  XOR U234 ( .A(B[491]), .B(B[490]), .Z(n156) );
  XOR U235 ( .A(B[489]), .B(n157), .Z(O[490]) );
  AND U236 ( .A(S), .B(n158), .Z(n157) );
  XOR U237 ( .A(B[490]), .B(B[489]), .Z(n158) );
  XOR U238 ( .A(B[47]), .B(n159), .Z(O[48]) );
  AND U239 ( .A(S), .B(n160), .Z(n159) );
  XOR U240 ( .A(B[48]), .B(B[47]), .Z(n160) );
  XOR U241 ( .A(B[488]), .B(n161), .Z(O[489]) );
  AND U242 ( .A(S), .B(n162), .Z(n161) );
  XOR U243 ( .A(B[489]), .B(B[488]), .Z(n162) );
  XOR U244 ( .A(B[487]), .B(n163), .Z(O[488]) );
  AND U245 ( .A(S), .B(n164), .Z(n163) );
  XOR U246 ( .A(B[488]), .B(B[487]), .Z(n164) );
  XOR U247 ( .A(B[486]), .B(n165), .Z(O[487]) );
  AND U248 ( .A(S), .B(n166), .Z(n165) );
  XOR U249 ( .A(B[487]), .B(B[486]), .Z(n166) );
  XOR U250 ( .A(B[485]), .B(n167), .Z(O[486]) );
  AND U251 ( .A(S), .B(n168), .Z(n167) );
  XOR U252 ( .A(B[486]), .B(B[485]), .Z(n168) );
  XOR U253 ( .A(B[484]), .B(n169), .Z(O[485]) );
  AND U254 ( .A(S), .B(n170), .Z(n169) );
  XOR U255 ( .A(B[485]), .B(B[484]), .Z(n170) );
  XOR U256 ( .A(B[483]), .B(n171), .Z(O[484]) );
  AND U257 ( .A(S), .B(n172), .Z(n171) );
  XOR U258 ( .A(B[484]), .B(B[483]), .Z(n172) );
  XOR U259 ( .A(B[482]), .B(n173), .Z(O[483]) );
  AND U260 ( .A(S), .B(n174), .Z(n173) );
  XOR U261 ( .A(B[483]), .B(B[482]), .Z(n174) );
  XOR U262 ( .A(B[481]), .B(n175), .Z(O[482]) );
  AND U263 ( .A(S), .B(n176), .Z(n175) );
  XOR U264 ( .A(B[482]), .B(B[481]), .Z(n176) );
  XOR U265 ( .A(B[480]), .B(n177), .Z(O[481]) );
  AND U266 ( .A(S), .B(n178), .Z(n177) );
  XOR U267 ( .A(B[481]), .B(B[480]), .Z(n178) );
  XOR U268 ( .A(B[479]), .B(n179), .Z(O[480]) );
  AND U269 ( .A(S), .B(n180), .Z(n179) );
  XOR U270 ( .A(B[480]), .B(B[479]), .Z(n180) );
  XOR U271 ( .A(B[46]), .B(n181), .Z(O[47]) );
  AND U272 ( .A(S), .B(n182), .Z(n181) );
  XOR U273 ( .A(B[47]), .B(B[46]), .Z(n182) );
  XOR U274 ( .A(B[478]), .B(n183), .Z(O[479]) );
  AND U275 ( .A(S), .B(n184), .Z(n183) );
  XOR U276 ( .A(B[479]), .B(B[478]), .Z(n184) );
  XOR U277 ( .A(B[477]), .B(n185), .Z(O[478]) );
  AND U278 ( .A(S), .B(n186), .Z(n185) );
  XOR U279 ( .A(B[478]), .B(B[477]), .Z(n186) );
  XOR U280 ( .A(B[476]), .B(n187), .Z(O[477]) );
  AND U281 ( .A(S), .B(n188), .Z(n187) );
  XOR U282 ( .A(B[477]), .B(B[476]), .Z(n188) );
  XOR U283 ( .A(B[475]), .B(n189), .Z(O[476]) );
  AND U284 ( .A(S), .B(n190), .Z(n189) );
  XOR U285 ( .A(B[476]), .B(B[475]), .Z(n190) );
  XOR U286 ( .A(B[474]), .B(n191), .Z(O[475]) );
  AND U287 ( .A(S), .B(n192), .Z(n191) );
  XOR U288 ( .A(B[475]), .B(B[474]), .Z(n192) );
  XOR U289 ( .A(B[473]), .B(n193), .Z(O[474]) );
  AND U290 ( .A(S), .B(n194), .Z(n193) );
  XOR U291 ( .A(B[474]), .B(B[473]), .Z(n194) );
  XOR U292 ( .A(B[472]), .B(n195), .Z(O[473]) );
  AND U293 ( .A(S), .B(n196), .Z(n195) );
  XOR U294 ( .A(B[473]), .B(B[472]), .Z(n196) );
  XOR U295 ( .A(B[471]), .B(n197), .Z(O[472]) );
  AND U296 ( .A(S), .B(n198), .Z(n197) );
  XOR U297 ( .A(B[472]), .B(B[471]), .Z(n198) );
  XOR U298 ( .A(B[470]), .B(n199), .Z(O[471]) );
  AND U299 ( .A(S), .B(n200), .Z(n199) );
  XOR U300 ( .A(B[471]), .B(B[470]), .Z(n200) );
  XOR U301 ( .A(B[469]), .B(n201), .Z(O[470]) );
  AND U302 ( .A(S), .B(n202), .Z(n201) );
  XOR U303 ( .A(B[470]), .B(B[469]), .Z(n202) );
  XOR U304 ( .A(B[45]), .B(n203), .Z(O[46]) );
  AND U305 ( .A(S), .B(n204), .Z(n203) );
  XOR U306 ( .A(B[46]), .B(B[45]), .Z(n204) );
  XOR U307 ( .A(B[468]), .B(n205), .Z(O[469]) );
  AND U308 ( .A(S), .B(n206), .Z(n205) );
  XOR U309 ( .A(B[469]), .B(B[468]), .Z(n206) );
  XOR U310 ( .A(B[467]), .B(n207), .Z(O[468]) );
  AND U311 ( .A(S), .B(n208), .Z(n207) );
  XOR U312 ( .A(B[468]), .B(B[467]), .Z(n208) );
  XOR U313 ( .A(B[466]), .B(n209), .Z(O[467]) );
  AND U314 ( .A(S), .B(n210), .Z(n209) );
  XOR U315 ( .A(B[467]), .B(B[466]), .Z(n210) );
  XOR U316 ( .A(B[465]), .B(n211), .Z(O[466]) );
  AND U317 ( .A(S), .B(n212), .Z(n211) );
  XOR U318 ( .A(B[466]), .B(B[465]), .Z(n212) );
  XOR U319 ( .A(B[464]), .B(n213), .Z(O[465]) );
  AND U320 ( .A(S), .B(n214), .Z(n213) );
  XOR U321 ( .A(B[465]), .B(B[464]), .Z(n214) );
  XOR U322 ( .A(B[463]), .B(n215), .Z(O[464]) );
  AND U323 ( .A(S), .B(n216), .Z(n215) );
  XOR U324 ( .A(B[464]), .B(B[463]), .Z(n216) );
  XOR U325 ( .A(B[462]), .B(n217), .Z(O[463]) );
  AND U326 ( .A(S), .B(n218), .Z(n217) );
  XOR U327 ( .A(B[463]), .B(B[462]), .Z(n218) );
  XOR U328 ( .A(B[461]), .B(n219), .Z(O[462]) );
  AND U329 ( .A(S), .B(n220), .Z(n219) );
  XOR U330 ( .A(B[462]), .B(B[461]), .Z(n220) );
  XOR U331 ( .A(B[460]), .B(n221), .Z(O[461]) );
  AND U332 ( .A(S), .B(n222), .Z(n221) );
  XOR U333 ( .A(B[461]), .B(B[460]), .Z(n222) );
  XOR U334 ( .A(B[459]), .B(n223), .Z(O[460]) );
  AND U335 ( .A(S), .B(n224), .Z(n223) );
  XOR U336 ( .A(B[460]), .B(B[459]), .Z(n224) );
  XOR U337 ( .A(B[44]), .B(n225), .Z(O[45]) );
  AND U338 ( .A(S), .B(n226), .Z(n225) );
  XOR U339 ( .A(B[45]), .B(B[44]), .Z(n226) );
  XOR U340 ( .A(B[458]), .B(n227), .Z(O[459]) );
  AND U341 ( .A(S), .B(n228), .Z(n227) );
  XOR U342 ( .A(B[459]), .B(B[458]), .Z(n228) );
  XOR U343 ( .A(B[457]), .B(n229), .Z(O[458]) );
  AND U344 ( .A(S), .B(n230), .Z(n229) );
  XOR U345 ( .A(B[458]), .B(B[457]), .Z(n230) );
  XOR U346 ( .A(B[456]), .B(n231), .Z(O[457]) );
  AND U347 ( .A(S), .B(n232), .Z(n231) );
  XOR U348 ( .A(B[457]), .B(B[456]), .Z(n232) );
  XOR U349 ( .A(B[455]), .B(n233), .Z(O[456]) );
  AND U350 ( .A(S), .B(n234), .Z(n233) );
  XOR U351 ( .A(B[456]), .B(B[455]), .Z(n234) );
  XOR U352 ( .A(B[454]), .B(n235), .Z(O[455]) );
  AND U353 ( .A(S), .B(n236), .Z(n235) );
  XOR U354 ( .A(B[455]), .B(B[454]), .Z(n236) );
  XOR U355 ( .A(B[453]), .B(n237), .Z(O[454]) );
  AND U356 ( .A(S), .B(n238), .Z(n237) );
  XOR U357 ( .A(B[454]), .B(B[453]), .Z(n238) );
  XOR U358 ( .A(B[452]), .B(n239), .Z(O[453]) );
  AND U359 ( .A(S), .B(n240), .Z(n239) );
  XOR U360 ( .A(B[453]), .B(B[452]), .Z(n240) );
  XOR U361 ( .A(B[451]), .B(n241), .Z(O[452]) );
  AND U362 ( .A(S), .B(n242), .Z(n241) );
  XOR U363 ( .A(B[452]), .B(B[451]), .Z(n242) );
  XOR U364 ( .A(B[450]), .B(n243), .Z(O[451]) );
  AND U365 ( .A(S), .B(n244), .Z(n243) );
  XOR U366 ( .A(B[451]), .B(B[450]), .Z(n244) );
  XOR U367 ( .A(B[449]), .B(n245), .Z(O[450]) );
  AND U368 ( .A(S), .B(n246), .Z(n245) );
  XOR U369 ( .A(B[450]), .B(B[449]), .Z(n246) );
  XOR U370 ( .A(B[43]), .B(n247), .Z(O[44]) );
  AND U371 ( .A(S), .B(n248), .Z(n247) );
  XOR U372 ( .A(B[44]), .B(B[43]), .Z(n248) );
  XOR U373 ( .A(B[448]), .B(n249), .Z(O[449]) );
  AND U374 ( .A(S), .B(n250), .Z(n249) );
  XOR U375 ( .A(B[449]), .B(B[448]), .Z(n250) );
  XOR U376 ( .A(B[447]), .B(n251), .Z(O[448]) );
  AND U377 ( .A(S), .B(n252), .Z(n251) );
  XOR U378 ( .A(B[448]), .B(B[447]), .Z(n252) );
  XOR U379 ( .A(B[446]), .B(n253), .Z(O[447]) );
  AND U380 ( .A(S), .B(n254), .Z(n253) );
  XOR U381 ( .A(B[447]), .B(B[446]), .Z(n254) );
  XOR U382 ( .A(B[445]), .B(n255), .Z(O[446]) );
  AND U383 ( .A(S), .B(n256), .Z(n255) );
  XOR U384 ( .A(B[446]), .B(B[445]), .Z(n256) );
  XOR U385 ( .A(B[444]), .B(n257), .Z(O[445]) );
  AND U386 ( .A(S), .B(n258), .Z(n257) );
  XOR U387 ( .A(B[445]), .B(B[444]), .Z(n258) );
  XOR U388 ( .A(B[443]), .B(n259), .Z(O[444]) );
  AND U389 ( .A(S), .B(n260), .Z(n259) );
  XOR U390 ( .A(B[444]), .B(B[443]), .Z(n260) );
  XOR U391 ( .A(B[442]), .B(n261), .Z(O[443]) );
  AND U392 ( .A(S), .B(n262), .Z(n261) );
  XOR U393 ( .A(B[443]), .B(B[442]), .Z(n262) );
  XOR U394 ( .A(B[441]), .B(n263), .Z(O[442]) );
  AND U395 ( .A(S), .B(n264), .Z(n263) );
  XOR U396 ( .A(B[442]), .B(B[441]), .Z(n264) );
  XOR U397 ( .A(B[440]), .B(n265), .Z(O[441]) );
  AND U398 ( .A(S), .B(n266), .Z(n265) );
  XOR U399 ( .A(B[441]), .B(B[440]), .Z(n266) );
  XOR U400 ( .A(B[439]), .B(n267), .Z(O[440]) );
  AND U401 ( .A(S), .B(n268), .Z(n267) );
  XOR U402 ( .A(B[440]), .B(B[439]), .Z(n268) );
  XOR U403 ( .A(B[42]), .B(n269), .Z(O[43]) );
  AND U404 ( .A(S), .B(n270), .Z(n269) );
  XOR U405 ( .A(B[43]), .B(B[42]), .Z(n270) );
  XOR U406 ( .A(B[438]), .B(n271), .Z(O[439]) );
  AND U407 ( .A(S), .B(n272), .Z(n271) );
  XOR U408 ( .A(B[439]), .B(B[438]), .Z(n272) );
  XOR U409 ( .A(B[437]), .B(n273), .Z(O[438]) );
  AND U410 ( .A(S), .B(n274), .Z(n273) );
  XOR U411 ( .A(B[438]), .B(B[437]), .Z(n274) );
  XOR U412 ( .A(B[436]), .B(n275), .Z(O[437]) );
  AND U413 ( .A(S), .B(n276), .Z(n275) );
  XOR U414 ( .A(B[437]), .B(B[436]), .Z(n276) );
  XOR U415 ( .A(B[435]), .B(n277), .Z(O[436]) );
  AND U416 ( .A(S), .B(n278), .Z(n277) );
  XOR U417 ( .A(B[436]), .B(B[435]), .Z(n278) );
  XOR U418 ( .A(B[434]), .B(n279), .Z(O[435]) );
  AND U419 ( .A(S), .B(n280), .Z(n279) );
  XOR U420 ( .A(B[435]), .B(B[434]), .Z(n280) );
  XOR U421 ( .A(B[433]), .B(n281), .Z(O[434]) );
  AND U422 ( .A(S), .B(n282), .Z(n281) );
  XOR U423 ( .A(B[434]), .B(B[433]), .Z(n282) );
  XOR U424 ( .A(B[432]), .B(n283), .Z(O[433]) );
  AND U425 ( .A(S), .B(n284), .Z(n283) );
  XOR U426 ( .A(B[433]), .B(B[432]), .Z(n284) );
  XOR U427 ( .A(B[431]), .B(n285), .Z(O[432]) );
  AND U428 ( .A(S), .B(n286), .Z(n285) );
  XOR U429 ( .A(B[432]), .B(B[431]), .Z(n286) );
  XOR U430 ( .A(B[430]), .B(n287), .Z(O[431]) );
  AND U431 ( .A(S), .B(n288), .Z(n287) );
  XOR U432 ( .A(B[431]), .B(B[430]), .Z(n288) );
  XOR U433 ( .A(B[429]), .B(n289), .Z(O[430]) );
  AND U434 ( .A(S), .B(n290), .Z(n289) );
  XOR U435 ( .A(B[430]), .B(B[429]), .Z(n290) );
  XOR U436 ( .A(B[41]), .B(n291), .Z(O[42]) );
  AND U437 ( .A(S), .B(n292), .Z(n291) );
  XOR U438 ( .A(B[42]), .B(B[41]), .Z(n292) );
  XOR U439 ( .A(B[428]), .B(n293), .Z(O[429]) );
  AND U440 ( .A(S), .B(n294), .Z(n293) );
  XOR U441 ( .A(B[429]), .B(B[428]), .Z(n294) );
  XOR U442 ( .A(B[427]), .B(n295), .Z(O[428]) );
  AND U443 ( .A(S), .B(n296), .Z(n295) );
  XOR U444 ( .A(B[428]), .B(B[427]), .Z(n296) );
  XOR U445 ( .A(B[426]), .B(n297), .Z(O[427]) );
  AND U446 ( .A(S), .B(n298), .Z(n297) );
  XOR U447 ( .A(B[427]), .B(B[426]), .Z(n298) );
  XOR U448 ( .A(B[425]), .B(n299), .Z(O[426]) );
  AND U449 ( .A(S), .B(n300), .Z(n299) );
  XOR U450 ( .A(B[426]), .B(B[425]), .Z(n300) );
  XOR U451 ( .A(B[424]), .B(n301), .Z(O[425]) );
  AND U452 ( .A(S), .B(n302), .Z(n301) );
  XOR U453 ( .A(B[425]), .B(B[424]), .Z(n302) );
  XOR U454 ( .A(B[423]), .B(n303), .Z(O[424]) );
  AND U455 ( .A(S), .B(n304), .Z(n303) );
  XOR U456 ( .A(B[424]), .B(B[423]), .Z(n304) );
  XOR U457 ( .A(B[422]), .B(n305), .Z(O[423]) );
  AND U458 ( .A(S), .B(n306), .Z(n305) );
  XOR U459 ( .A(B[423]), .B(B[422]), .Z(n306) );
  XOR U460 ( .A(B[421]), .B(n307), .Z(O[422]) );
  AND U461 ( .A(S), .B(n308), .Z(n307) );
  XOR U462 ( .A(B[422]), .B(B[421]), .Z(n308) );
  XOR U463 ( .A(B[420]), .B(n309), .Z(O[421]) );
  AND U464 ( .A(S), .B(n310), .Z(n309) );
  XOR U465 ( .A(B[421]), .B(B[420]), .Z(n310) );
  XOR U466 ( .A(B[419]), .B(n311), .Z(O[420]) );
  AND U467 ( .A(S), .B(n312), .Z(n311) );
  XOR U468 ( .A(B[420]), .B(B[419]), .Z(n312) );
  XOR U469 ( .A(B[40]), .B(n313), .Z(O[41]) );
  AND U470 ( .A(S), .B(n314), .Z(n313) );
  XOR U471 ( .A(B[41]), .B(B[40]), .Z(n314) );
  XOR U472 ( .A(B[418]), .B(n315), .Z(O[419]) );
  AND U473 ( .A(S), .B(n316), .Z(n315) );
  XOR U474 ( .A(B[419]), .B(B[418]), .Z(n316) );
  XOR U475 ( .A(B[417]), .B(n317), .Z(O[418]) );
  AND U476 ( .A(S), .B(n318), .Z(n317) );
  XOR U477 ( .A(B[418]), .B(B[417]), .Z(n318) );
  XOR U478 ( .A(B[416]), .B(n319), .Z(O[417]) );
  AND U479 ( .A(S), .B(n320), .Z(n319) );
  XOR U480 ( .A(B[417]), .B(B[416]), .Z(n320) );
  XOR U481 ( .A(B[415]), .B(n321), .Z(O[416]) );
  AND U482 ( .A(S), .B(n322), .Z(n321) );
  XOR U483 ( .A(B[416]), .B(B[415]), .Z(n322) );
  XOR U484 ( .A(B[414]), .B(n323), .Z(O[415]) );
  AND U485 ( .A(S), .B(n324), .Z(n323) );
  XOR U486 ( .A(B[415]), .B(B[414]), .Z(n324) );
  XOR U487 ( .A(B[413]), .B(n325), .Z(O[414]) );
  AND U488 ( .A(S), .B(n326), .Z(n325) );
  XOR U489 ( .A(B[414]), .B(B[413]), .Z(n326) );
  XOR U490 ( .A(B[412]), .B(n327), .Z(O[413]) );
  AND U491 ( .A(S), .B(n328), .Z(n327) );
  XOR U492 ( .A(B[413]), .B(B[412]), .Z(n328) );
  XOR U493 ( .A(B[411]), .B(n329), .Z(O[412]) );
  AND U494 ( .A(S), .B(n330), .Z(n329) );
  XOR U495 ( .A(B[412]), .B(B[411]), .Z(n330) );
  XOR U496 ( .A(B[410]), .B(n331), .Z(O[411]) );
  AND U497 ( .A(S), .B(n332), .Z(n331) );
  XOR U498 ( .A(B[411]), .B(B[410]), .Z(n332) );
  XOR U499 ( .A(B[409]), .B(n333), .Z(O[410]) );
  AND U500 ( .A(S), .B(n334), .Z(n333) );
  XOR U501 ( .A(B[410]), .B(B[409]), .Z(n334) );
  XOR U502 ( .A(B[39]), .B(n335), .Z(O[40]) );
  AND U503 ( .A(S), .B(n336), .Z(n335) );
  XOR U504 ( .A(B[40]), .B(B[39]), .Z(n336) );
  XOR U505 ( .A(B[408]), .B(n337), .Z(O[409]) );
  AND U506 ( .A(S), .B(n338), .Z(n337) );
  XOR U507 ( .A(B[409]), .B(B[408]), .Z(n338) );
  XOR U508 ( .A(B[407]), .B(n339), .Z(O[408]) );
  AND U509 ( .A(S), .B(n340), .Z(n339) );
  XOR U510 ( .A(B[408]), .B(B[407]), .Z(n340) );
  XOR U511 ( .A(B[406]), .B(n341), .Z(O[407]) );
  AND U512 ( .A(S), .B(n342), .Z(n341) );
  XOR U513 ( .A(B[407]), .B(B[406]), .Z(n342) );
  XOR U514 ( .A(B[405]), .B(n343), .Z(O[406]) );
  AND U515 ( .A(S), .B(n344), .Z(n343) );
  XOR U516 ( .A(B[406]), .B(B[405]), .Z(n344) );
  XOR U517 ( .A(B[404]), .B(n345), .Z(O[405]) );
  AND U518 ( .A(S), .B(n346), .Z(n345) );
  XOR U519 ( .A(B[405]), .B(B[404]), .Z(n346) );
  XOR U520 ( .A(B[403]), .B(n347), .Z(O[404]) );
  AND U521 ( .A(S), .B(n348), .Z(n347) );
  XOR U522 ( .A(B[404]), .B(B[403]), .Z(n348) );
  XOR U523 ( .A(B[402]), .B(n349), .Z(O[403]) );
  AND U524 ( .A(S), .B(n350), .Z(n349) );
  XOR U525 ( .A(B[403]), .B(B[402]), .Z(n350) );
  XOR U526 ( .A(B[401]), .B(n351), .Z(O[402]) );
  AND U527 ( .A(S), .B(n352), .Z(n351) );
  XOR U528 ( .A(B[402]), .B(B[401]), .Z(n352) );
  XOR U529 ( .A(B[400]), .B(n353), .Z(O[401]) );
  AND U530 ( .A(S), .B(n354), .Z(n353) );
  XOR U531 ( .A(B[401]), .B(B[400]), .Z(n354) );
  XOR U532 ( .A(B[399]), .B(n355), .Z(O[400]) );
  AND U533 ( .A(S), .B(n356), .Z(n355) );
  XOR U534 ( .A(B[400]), .B(B[399]), .Z(n356) );
  XOR U535 ( .A(B[2]), .B(n357), .Z(O[3]) );
  AND U536 ( .A(S), .B(n358), .Z(n357) );
  XOR U537 ( .A(B[3]), .B(B[2]), .Z(n358) );
  XOR U538 ( .A(B[38]), .B(n359), .Z(O[39]) );
  AND U539 ( .A(S), .B(n360), .Z(n359) );
  XOR U540 ( .A(B[39]), .B(B[38]), .Z(n360) );
  XOR U541 ( .A(B[398]), .B(n361), .Z(O[399]) );
  AND U542 ( .A(S), .B(n362), .Z(n361) );
  XOR U543 ( .A(B[399]), .B(B[398]), .Z(n362) );
  XOR U544 ( .A(B[397]), .B(n363), .Z(O[398]) );
  AND U545 ( .A(S), .B(n364), .Z(n363) );
  XOR U546 ( .A(B[398]), .B(B[397]), .Z(n364) );
  XOR U547 ( .A(B[396]), .B(n365), .Z(O[397]) );
  AND U548 ( .A(S), .B(n366), .Z(n365) );
  XOR U549 ( .A(B[397]), .B(B[396]), .Z(n366) );
  XOR U550 ( .A(B[395]), .B(n367), .Z(O[396]) );
  AND U551 ( .A(S), .B(n368), .Z(n367) );
  XOR U552 ( .A(B[396]), .B(B[395]), .Z(n368) );
  XOR U553 ( .A(B[394]), .B(n369), .Z(O[395]) );
  AND U554 ( .A(S), .B(n370), .Z(n369) );
  XOR U555 ( .A(B[395]), .B(B[394]), .Z(n370) );
  XOR U556 ( .A(B[393]), .B(n371), .Z(O[394]) );
  AND U557 ( .A(S), .B(n372), .Z(n371) );
  XOR U558 ( .A(B[394]), .B(B[393]), .Z(n372) );
  XOR U559 ( .A(B[392]), .B(n373), .Z(O[393]) );
  AND U560 ( .A(S), .B(n374), .Z(n373) );
  XOR U561 ( .A(B[393]), .B(B[392]), .Z(n374) );
  XOR U562 ( .A(B[391]), .B(n375), .Z(O[392]) );
  AND U563 ( .A(S), .B(n376), .Z(n375) );
  XOR U564 ( .A(B[392]), .B(B[391]), .Z(n376) );
  XOR U565 ( .A(B[390]), .B(n377), .Z(O[391]) );
  AND U566 ( .A(S), .B(n378), .Z(n377) );
  XOR U567 ( .A(B[391]), .B(B[390]), .Z(n378) );
  XOR U568 ( .A(B[389]), .B(n379), .Z(O[390]) );
  AND U569 ( .A(S), .B(n380), .Z(n379) );
  XOR U570 ( .A(B[390]), .B(B[389]), .Z(n380) );
  XOR U571 ( .A(B[37]), .B(n381), .Z(O[38]) );
  AND U572 ( .A(S), .B(n382), .Z(n381) );
  XOR U573 ( .A(B[38]), .B(B[37]), .Z(n382) );
  XOR U574 ( .A(B[388]), .B(n383), .Z(O[389]) );
  AND U575 ( .A(S), .B(n384), .Z(n383) );
  XOR U576 ( .A(B[389]), .B(B[388]), .Z(n384) );
  XOR U577 ( .A(B[387]), .B(n385), .Z(O[388]) );
  AND U578 ( .A(S), .B(n386), .Z(n385) );
  XOR U579 ( .A(B[388]), .B(B[387]), .Z(n386) );
  XOR U580 ( .A(B[386]), .B(n387), .Z(O[387]) );
  AND U581 ( .A(S), .B(n388), .Z(n387) );
  XOR U582 ( .A(B[387]), .B(B[386]), .Z(n388) );
  XOR U583 ( .A(B[385]), .B(n389), .Z(O[386]) );
  AND U584 ( .A(S), .B(n390), .Z(n389) );
  XOR U585 ( .A(B[386]), .B(B[385]), .Z(n390) );
  XOR U586 ( .A(B[384]), .B(n391), .Z(O[385]) );
  AND U587 ( .A(S), .B(n392), .Z(n391) );
  XOR U588 ( .A(B[385]), .B(B[384]), .Z(n392) );
  XOR U589 ( .A(B[383]), .B(n393), .Z(O[384]) );
  AND U590 ( .A(S), .B(n394), .Z(n393) );
  XOR U591 ( .A(B[384]), .B(B[383]), .Z(n394) );
  XOR U592 ( .A(B[382]), .B(n395), .Z(O[383]) );
  AND U593 ( .A(S), .B(n396), .Z(n395) );
  XOR U594 ( .A(B[383]), .B(B[382]), .Z(n396) );
  XOR U595 ( .A(B[381]), .B(n397), .Z(O[382]) );
  AND U596 ( .A(S), .B(n398), .Z(n397) );
  XOR U597 ( .A(B[382]), .B(B[381]), .Z(n398) );
  XOR U598 ( .A(B[380]), .B(n399), .Z(O[381]) );
  AND U599 ( .A(S), .B(n400), .Z(n399) );
  XOR U600 ( .A(B[381]), .B(B[380]), .Z(n400) );
  XOR U601 ( .A(B[379]), .B(n401), .Z(O[380]) );
  AND U602 ( .A(S), .B(n402), .Z(n401) );
  XOR U603 ( .A(B[380]), .B(B[379]), .Z(n402) );
  XOR U604 ( .A(B[36]), .B(n403), .Z(O[37]) );
  AND U605 ( .A(S), .B(n404), .Z(n403) );
  XOR U606 ( .A(B[37]), .B(B[36]), .Z(n404) );
  XOR U607 ( .A(B[378]), .B(n405), .Z(O[379]) );
  AND U608 ( .A(S), .B(n406), .Z(n405) );
  XOR U609 ( .A(B[379]), .B(B[378]), .Z(n406) );
  XOR U610 ( .A(B[377]), .B(n407), .Z(O[378]) );
  AND U611 ( .A(S), .B(n408), .Z(n407) );
  XOR U612 ( .A(B[378]), .B(B[377]), .Z(n408) );
  XOR U613 ( .A(B[376]), .B(n409), .Z(O[377]) );
  AND U614 ( .A(S), .B(n410), .Z(n409) );
  XOR U615 ( .A(B[377]), .B(B[376]), .Z(n410) );
  XOR U616 ( .A(B[375]), .B(n411), .Z(O[376]) );
  AND U617 ( .A(S), .B(n412), .Z(n411) );
  XOR U618 ( .A(B[376]), .B(B[375]), .Z(n412) );
  XOR U619 ( .A(B[374]), .B(n413), .Z(O[375]) );
  AND U620 ( .A(S), .B(n414), .Z(n413) );
  XOR U621 ( .A(B[375]), .B(B[374]), .Z(n414) );
  XOR U622 ( .A(B[373]), .B(n415), .Z(O[374]) );
  AND U623 ( .A(S), .B(n416), .Z(n415) );
  XOR U624 ( .A(B[374]), .B(B[373]), .Z(n416) );
  XOR U625 ( .A(B[372]), .B(n417), .Z(O[373]) );
  AND U626 ( .A(S), .B(n418), .Z(n417) );
  XOR U627 ( .A(B[373]), .B(B[372]), .Z(n418) );
  XOR U628 ( .A(B[371]), .B(n419), .Z(O[372]) );
  AND U629 ( .A(S), .B(n420), .Z(n419) );
  XOR U630 ( .A(B[372]), .B(B[371]), .Z(n420) );
  XOR U631 ( .A(B[370]), .B(n421), .Z(O[371]) );
  AND U632 ( .A(S), .B(n422), .Z(n421) );
  XOR U633 ( .A(B[371]), .B(B[370]), .Z(n422) );
  XOR U634 ( .A(B[369]), .B(n423), .Z(O[370]) );
  AND U635 ( .A(S), .B(n424), .Z(n423) );
  XOR U636 ( .A(B[370]), .B(B[369]), .Z(n424) );
  XOR U637 ( .A(B[35]), .B(n425), .Z(O[36]) );
  AND U638 ( .A(S), .B(n426), .Z(n425) );
  XOR U639 ( .A(B[36]), .B(B[35]), .Z(n426) );
  XOR U640 ( .A(B[368]), .B(n427), .Z(O[369]) );
  AND U641 ( .A(S), .B(n428), .Z(n427) );
  XOR U642 ( .A(B[369]), .B(B[368]), .Z(n428) );
  XOR U643 ( .A(B[367]), .B(n429), .Z(O[368]) );
  AND U644 ( .A(S), .B(n430), .Z(n429) );
  XOR U645 ( .A(B[368]), .B(B[367]), .Z(n430) );
  XOR U646 ( .A(B[366]), .B(n431), .Z(O[367]) );
  AND U647 ( .A(S), .B(n432), .Z(n431) );
  XOR U648 ( .A(B[367]), .B(B[366]), .Z(n432) );
  XOR U649 ( .A(B[365]), .B(n433), .Z(O[366]) );
  AND U650 ( .A(S), .B(n434), .Z(n433) );
  XOR U651 ( .A(B[366]), .B(B[365]), .Z(n434) );
  XOR U652 ( .A(B[364]), .B(n435), .Z(O[365]) );
  AND U653 ( .A(S), .B(n436), .Z(n435) );
  XOR U654 ( .A(B[365]), .B(B[364]), .Z(n436) );
  XOR U655 ( .A(B[363]), .B(n437), .Z(O[364]) );
  AND U656 ( .A(S), .B(n438), .Z(n437) );
  XOR U657 ( .A(B[364]), .B(B[363]), .Z(n438) );
  XOR U658 ( .A(B[362]), .B(n439), .Z(O[363]) );
  AND U659 ( .A(S), .B(n440), .Z(n439) );
  XOR U660 ( .A(B[363]), .B(B[362]), .Z(n440) );
  XOR U661 ( .A(B[361]), .B(n441), .Z(O[362]) );
  AND U662 ( .A(S), .B(n442), .Z(n441) );
  XOR U663 ( .A(B[362]), .B(B[361]), .Z(n442) );
  XOR U664 ( .A(B[360]), .B(n443), .Z(O[361]) );
  AND U665 ( .A(S), .B(n444), .Z(n443) );
  XOR U666 ( .A(B[361]), .B(B[360]), .Z(n444) );
  XOR U667 ( .A(B[359]), .B(n445), .Z(O[360]) );
  AND U668 ( .A(S), .B(n446), .Z(n445) );
  XOR U669 ( .A(B[360]), .B(B[359]), .Z(n446) );
  XOR U670 ( .A(B[34]), .B(n447), .Z(O[35]) );
  AND U671 ( .A(S), .B(n448), .Z(n447) );
  XOR U672 ( .A(B[35]), .B(B[34]), .Z(n448) );
  XOR U673 ( .A(B[358]), .B(n449), .Z(O[359]) );
  AND U674 ( .A(S), .B(n450), .Z(n449) );
  XOR U675 ( .A(B[359]), .B(B[358]), .Z(n450) );
  XOR U676 ( .A(B[357]), .B(n451), .Z(O[358]) );
  AND U677 ( .A(S), .B(n452), .Z(n451) );
  XOR U678 ( .A(B[358]), .B(B[357]), .Z(n452) );
  XOR U679 ( .A(B[356]), .B(n453), .Z(O[357]) );
  AND U680 ( .A(S), .B(n454), .Z(n453) );
  XOR U681 ( .A(B[357]), .B(B[356]), .Z(n454) );
  XOR U682 ( .A(B[355]), .B(n455), .Z(O[356]) );
  AND U683 ( .A(S), .B(n456), .Z(n455) );
  XOR U684 ( .A(B[356]), .B(B[355]), .Z(n456) );
  XOR U685 ( .A(B[354]), .B(n457), .Z(O[355]) );
  AND U686 ( .A(S), .B(n458), .Z(n457) );
  XOR U687 ( .A(B[355]), .B(B[354]), .Z(n458) );
  XOR U688 ( .A(B[353]), .B(n459), .Z(O[354]) );
  AND U689 ( .A(S), .B(n460), .Z(n459) );
  XOR U690 ( .A(B[354]), .B(B[353]), .Z(n460) );
  XOR U691 ( .A(B[352]), .B(n461), .Z(O[353]) );
  AND U692 ( .A(S), .B(n462), .Z(n461) );
  XOR U693 ( .A(B[353]), .B(B[352]), .Z(n462) );
  XOR U694 ( .A(B[351]), .B(n463), .Z(O[352]) );
  AND U695 ( .A(S), .B(n464), .Z(n463) );
  XOR U696 ( .A(B[352]), .B(B[351]), .Z(n464) );
  XOR U697 ( .A(B[350]), .B(n465), .Z(O[351]) );
  AND U698 ( .A(S), .B(n466), .Z(n465) );
  XOR U699 ( .A(B[351]), .B(B[350]), .Z(n466) );
  XOR U700 ( .A(B[349]), .B(n467), .Z(O[350]) );
  AND U701 ( .A(S), .B(n468), .Z(n467) );
  XOR U702 ( .A(B[350]), .B(B[349]), .Z(n468) );
  XOR U703 ( .A(B[33]), .B(n469), .Z(O[34]) );
  AND U704 ( .A(S), .B(n470), .Z(n469) );
  XOR U705 ( .A(B[34]), .B(B[33]), .Z(n470) );
  XOR U706 ( .A(B[348]), .B(n471), .Z(O[349]) );
  AND U707 ( .A(S), .B(n472), .Z(n471) );
  XOR U708 ( .A(B[349]), .B(B[348]), .Z(n472) );
  XOR U709 ( .A(B[347]), .B(n473), .Z(O[348]) );
  AND U710 ( .A(S), .B(n474), .Z(n473) );
  XOR U711 ( .A(B[348]), .B(B[347]), .Z(n474) );
  XOR U712 ( .A(B[346]), .B(n475), .Z(O[347]) );
  AND U713 ( .A(S), .B(n476), .Z(n475) );
  XOR U714 ( .A(B[347]), .B(B[346]), .Z(n476) );
  XOR U715 ( .A(B[345]), .B(n477), .Z(O[346]) );
  AND U716 ( .A(S), .B(n478), .Z(n477) );
  XOR U717 ( .A(B[346]), .B(B[345]), .Z(n478) );
  XOR U718 ( .A(B[344]), .B(n479), .Z(O[345]) );
  AND U719 ( .A(S), .B(n480), .Z(n479) );
  XOR U720 ( .A(B[345]), .B(B[344]), .Z(n480) );
  XOR U721 ( .A(B[343]), .B(n481), .Z(O[344]) );
  AND U722 ( .A(S), .B(n482), .Z(n481) );
  XOR U723 ( .A(B[344]), .B(B[343]), .Z(n482) );
  XOR U724 ( .A(B[342]), .B(n483), .Z(O[343]) );
  AND U725 ( .A(S), .B(n484), .Z(n483) );
  XOR U726 ( .A(B[343]), .B(B[342]), .Z(n484) );
  XOR U727 ( .A(B[341]), .B(n485), .Z(O[342]) );
  AND U728 ( .A(S), .B(n486), .Z(n485) );
  XOR U729 ( .A(B[342]), .B(B[341]), .Z(n486) );
  XOR U730 ( .A(B[340]), .B(n487), .Z(O[341]) );
  AND U731 ( .A(S), .B(n488), .Z(n487) );
  XOR U732 ( .A(B[341]), .B(B[340]), .Z(n488) );
  XOR U733 ( .A(B[339]), .B(n489), .Z(O[340]) );
  AND U734 ( .A(S), .B(n490), .Z(n489) );
  XOR U735 ( .A(B[340]), .B(B[339]), .Z(n490) );
  XOR U736 ( .A(B[32]), .B(n491), .Z(O[33]) );
  AND U737 ( .A(S), .B(n492), .Z(n491) );
  XOR U738 ( .A(B[33]), .B(B[32]), .Z(n492) );
  XOR U739 ( .A(B[338]), .B(n493), .Z(O[339]) );
  AND U740 ( .A(S), .B(n494), .Z(n493) );
  XOR U741 ( .A(B[339]), .B(B[338]), .Z(n494) );
  XOR U742 ( .A(B[337]), .B(n495), .Z(O[338]) );
  AND U743 ( .A(S), .B(n496), .Z(n495) );
  XOR U744 ( .A(B[338]), .B(B[337]), .Z(n496) );
  XOR U745 ( .A(B[336]), .B(n497), .Z(O[337]) );
  AND U746 ( .A(S), .B(n498), .Z(n497) );
  XOR U747 ( .A(B[337]), .B(B[336]), .Z(n498) );
  XOR U748 ( .A(B[335]), .B(n499), .Z(O[336]) );
  AND U749 ( .A(S), .B(n500), .Z(n499) );
  XOR U750 ( .A(B[336]), .B(B[335]), .Z(n500) );
  XOR U751 ( .A(B[334]), .B(n501), .Z(O[335]) );
  AND U752 ( .A(S), .B(n502), .Z(n501) );
  XOR U753 ( .A(B[335]), .B(B[334]), .Z(n502) );
  XOR U754 ( .A(B[333]), .B(n503), .Z(O[334]) );
  AND U755 ( .A(S), .B(n504), .Z(n503) );
  XOR U756 ( .A(B[334]), .B(B[333]), .Z(n504) );
  XOR U757 ( .A(B[332]), .B(n505), .Z(O[333]) );
  AND U758 ( .A(S), .B(n506), .Z(n505) );
  XOR U759 ( .A(B[333]), .B(B[332]), .Z(n506) );
  XOR U760 ( .A(B[331]), .B(n507), .Z(O[332]) );
  AND U761 ( .A(S), .B(n508), .Z(n507) );
  XOR U762 ( .A(B[332]), .B(B[331]), .Z(n508) );
  XOR U763 ( .A(B[330]), .B(n509), .Z(O[331]) );
  AND U764 ( .A(S), .B(n510), .Z(n509) );
  XOR U765 ( .A(B[331]), .B(B[330]), .Z(n510) );
  XOR U766 ( .A(B[329]), .B(n511), .Z(O[330]) );
  AND U767 ( .A(S), .B(n512), .Z(n511) );
  XOR U768 ( .A(B[330]), .B(B[329]), .Z(n512) );
  XOR U769 ( .A(B[31]), .B(n513), .Z(O[32]) );
  AND U770 ( .A(S), .B(n514), .Z(n513) );
  XOR U771 ( .A(B[32]), .B(B[31]), .Z(n514) );
  XOR U772 ( .A(B[328]), .B(n515), .Z(O[329]) );
  AND U773 ( .A(S), .B(n516), .Z(n515) );
  XOR U774 ( .A(B[329]), .B(B[328]), .Z(n516) );
  XOR U775 ( .A(B[327]), .B(n517), .Z(O[328]) );
  AND U776 ( .A(S), .B(n518), .Z(n517) );
  XOR U777 ( .A(B[328]), .B(B[327]), .Z(n518) );
  XOR U778 ( .A(B[326]), .B(n519), .Z(O[327]) );
  AND U779 ( .A(S), .B(n520), .Z(n519) );
  XOR U780 ( .A(B[327]), .B(B[326]), .Z(n520) );
  XOR U781 ( .A(B[325]), .B(n521), .Z(O[326]) );
  AND U782 ( .A(S), .B(n522), .Z(n521) );
  XOR U783 ( .A(B[326]), .B(B[325]), .Z(n522) );
  XOR U784 ( .A(B[324]), .B(n523), .Z(O[325]) );
  AND U785 ( .A(S), .B(n524), .Z(n523) );
  XOR U786 ( .A(B[325]), .B(B[324]), .Z(n524) );
  XOR U787 ( .A(B[323]), .B(n525), .Z(O[324]) );
  AND U788 ( .A(S), .B(n526), .Z(n525) );
  XOR U789 ( .A(B[324]), .B(B[323]), .Z(n526) );
  XOR U790 ( .A(B[322]), .B(n527), .Z(O[323]) );
  AND U791 ( .A(S), .B(n528), .Z(n527) );
  XOR U792 ( .A(B[323]), .B(B[322]), .Z(n528) );
  XOR U793 ( .A(B[321]), .B(n529), .Z(O[322]) );
  AND U794 ( .A(S), .B(n530), .Z(n529) );
  XOR U795 ( .A(B[322]), .B(B[321]), .Z(n530) );
  XOR U796 ( .A(B[320]), .B(n531), .Z(O[321]) );
  AND U797 ( .A(S), .B(n532), .Z(n531) );
  XOR U798 ( .A(B[321]), .B(B[320]), .Z(n532) );
  XOR U799 ( .A(B[319]), .B(n533), .Z(O[320]) );
  AND U800 ( .A(S), .B(n534), .Z(n533) );
  XOR U801 ( .A(B[320]), .B(B[319]), .Z(n534) );
  XOR U802 ( .A(B[30]), .B(n535), .Z(O[31]) );
  AND U803 ( .A(S), .B(n536), .Z(n535) );
  XOR U804 ( .A(B[31]), .B(B[30]), .Z(n536) );
  XOR U805 ( .A(B[318]), .B(n537), .Z(O[319]) );
  AND U806 ( .A(S), .B(n538), .Z(n537) );
  XOR U807 ( .A(B[319]), .B(B[318]), .Z(n538) );
  XOR U808 ( .A(B[317]), .B(n539), .Z(O[318]) );
  AND U809 ( .A(S), .B(n540), .Z(n539) );
  XOR U810 ( .A(B[318]), .B(B[317]), .Z(n540) );
  XOR U811 ( .A(B[316]), .B(n541), .Z(O[317]) );
  AND U812 ( .A(S), .B(n542), .Z(n541) );
  XOR U813 ( .A(B[317]), .B(B[316]), .Z(n542) );
  XOR U814 ( .A(B[315]), .B(n543), .Z(O[316]) );
  AND U815 ( .A(S), .B(n544), .Z(n543) );
  XOR U816 ( .A(B[316]), .B(B[315]), .Z(n544) );
  XOR U817 ( .A(B[314]), .B(n545), .Z(O[315]) );
  AND U818 ( .A(S), .B(n546), .Z(n545) );
  XOR U819 ( .A(B[315]), .B(B[314]), .Z(n546) );
  XOR U820 ( .A(B[313]), .B(n547), .Z(O[314]) );
  AND U821 ( .A(S), .B(n548), .Z(n547) );
  XOR U822 ( .A(B[314]), .B(B[313]), .Z(n548) );
  XOR U823 ( .A(B[312]), .B(n549), .Z(O[313]) );
  AND U824 ( .A(S), .B(n550), .Z(n549) );
  XOR U825 ( .A(B[313]), .B(B[312]), .Z(n550) );
  XOR U826 ( .A(B[311]), .B(n551), .Z(O[312]) );
  AND U827 ( .A(S), .B(n552), .Z(n551) );
  XOR U828 ( .A(B[312]), .B(B[311]), .Z(n552) );
  XOR U829 ( .A(B[310]), .B(n553), .Z(O[311]) );
  AND U830 ( .A(S), .B(n554), .Z(n553) );
  XOR U831 ( .A(B[311]), .B(B[310]), .Z(n554) );
  XOR U832 ( .A(B[309]), .B(n555), .Z(O[310]) );
  AND U833 ( .A(S), .B(n556), .Z(n555) );
  XOR U834 ( .A(B[310]), .B(B[309]), .Z(n556) );
  XOR U835 ( .A(B[29]), .B(n557), .Z(O[30]) );
  AND U836 ( .A(S), .B(n558), .Z(n557) );
  XOR U837 ( .A(B[30]), .B(B[29]), .Z(n558) );
  XOR U838 ( .A(B[308]), .B(n559), .Z(O[309]) );
  AND U839 ( .A(S), .B(n560), .Z(n559) );
  XOR U840 ( .A(B[309]), .B(B[308]), .Z(n560) );
  XOR U841 ( .A(B[307]), .B(n561), .Z(O[308]) );
  AND U842 ( .A(S), .B(n562), .Z(n561) );
  XOR U843 ( .A(B[308]), .B(B[307]), .Z(n562) );
  XOR U844 ( .A(B[306]), .B(n563), .Z(O[307]) );
  AND U845 ( .A(S), .B(n564), .Z(n563) );
  XOR U846 ( .A(B[307]), .B(B[306]), .Z(n564) );
  XOR U847 ( .A(B[305]), .B(n565), .Z(O[306]) );
  AND U848 ( .A(S), .B(n566), .Z(n565) );
  XOR U849 ( .A(B[306]), .B(B[305]), .Z(n566) );
  XOR U850 ( .A(B[304]), .B(n567), .Z(O[305]) );
  AND U851 ( .A(S), .B(n568), .Z(n567) );
  XOR U852 ( .A(B[305]), .B(B[304]), .Z(n568) );
  XOR U853 ( .A(B[303]), .B(n569), .Z(O[304]) );
  AND U854 ( .A(S), .B(n570), .Z(n569) );
  XOR U855 ( .A(B[304]), .B(B[303]), .Z(n570) );
  XOR U856 ( .A(B[302]), .B(n571), .Z(O[303]) );
  AND U857 ( .A(S), .B(n572), .Z(n571) );
  XOR U858 ( .A(B[303]), .B(B[302]), .Z(n572) );
  XOR U859 ( .A(B[301]), .B(n573), .Z(O[302]) );
  AND U860 ( .A(S), .B(n574), .Z(n573) );
  XOR U861 ( .A(B[302]), .B(B[301]), .Z(n574) );
  XOR U862 ( .A(B[300]), .B(n575), .Z(O[301]) );
  AND U863 ( .A(S), .B(n576), .Z(n575) );
  XOR U864 ( .A(B[301]), .B(B[300]), .Z(n576) );
  XOR U865 ( .A(B[299]), .B(n577), .Z(O[300]) );
  AND U866 ( .A(S), .B(n578), .Z(n577) );
  XOR U867 ( .A(B[300]), .B(B[299]), .Z(n578) );
  XOR U868 ( .A(B[1]), .B(n579), .Z(O[2]) );
  AND U869 ( .A(S), .B(n580), .Z(n579) );
  XOR U870 ( .A(B[2]), .B(B[1]), .Z(n580) );
  XOR U871 ( .A(B[28]), .B(n581), .Z(O[29]) );
  AND U872 ( .A(S), .B(n582), .Z(n581) );
  XOR U873 ( .A(B[29]), .B(B[28]), .Z(n582) );
  XOR U874 ( .A(B[298]), .B(n583), .Z(O[299]) );
  AND U875 ( .A(S), .B(n584), .Z(n583) );
  XOR U876 ( .A(B[299]), .B(B[298]), .Z(n584) );
  XOR U877 ( .A(B[297]), .B(n585), .Z(O[298]) );
  AND U878 ( .A(S), .B(n586), .Z(n585) );
  XOR U879 ( .A(B[298]), .B(B[297]), .Z(n586) );
  XOR U880 ( .A(B[296]), .B(n587), .Z(O[297]) );
  AND U881 ( .A(S), .B(n588), .Z(n587) );
  XOR U882 ( .A(B[297]), .B(B[296]), .Z(n588) );
  XOR U883 ( .A(B[295]), .B(n589), .Z(O[296]) );
  AND U884 ( .A(S), .B(n590), .Z(n589) );
  XOR U885 ( .A(B[296]), .B(B[295]), .Z(n590) );
  XOR U886 ( .A(B[294]), .B(n591), .Z(O[295]) );
  AND U887 ( .A(S), .B(n592), .Z(n591) );
  XOR U888 ( .A(B[295]), .B(B[294]), .Z(n592) );
  XOR U889 ( .A(B[293]), .B(n593), .Z(O[294]) );
  AND U890 ( .A(S), .B(n594), .Z(n593) );
  XOR U891 ( .A(B[294]), .B(B[293]), .Z(n594) );
  XOR U892 ( .A(B[292]), .B(n595), .Z(O[293]) );
  AND U893 ( .A(S), .B(n596), .Z(n595) );
  XOR U894 ( .A(B[293]), .B(B[292]), .Z(n596) );
  XOR U895 ( .A(B[291]), .B(n597), .Z(O[292]) );
  AND U896 ( .A(S), .B(n598), .Z(n597) );
  XOR U897 ( .A(B[292]), .B(B[291]), .Z(n598) );
  XOR U898 ( .A(B[290]), .B(n599), .Z(O[291]) );
  AND U899 ( .A(S), .B(n600), .Z(n599) );
  XOR U900 ( .A(B[291]), .B(B[290]), .Z(n600) );
  XOR U901 ( .A(B[289]), .B(n601), .Z(O[290]) );
  AND U902 ( .A(S), .B(n602), .Z(n601) );
  XOR U903 ( .A(B[290]), .B(B[289]), .Z(n602) );
  XOR U904 ( .A(B[27]), .B(n603), .Z(O[28]) );
  AND U905 ( .A(S), .B(n604), .Z(n603) );
  XOR U906 ( .A(B[28]), .B(B[27]), .Z(n604) );
  XOR U907 ( .A(B[288]), .B(n605), .Z(O[289]) );
  AND U908 ( .A(S), .B(n606), .Z(n605) );
  XOR U909 ( .A(B[289]), .B(B[288]), .Z(n606) );
  XOR U910 ( .A(B[287]), .B(n607), .Z(O[288]) );
  AND U911 ( .A(S), .B(n608), .Z(n607) );
  XOR U912 ( .A(B[288]), .B(B[287]), .Z(n608) );
  XOR U913 ( .A(B[286]), .B(n609), .Z(O[287]) );
  AND U914 ( .A(S), .B(n610), .Z(n609) );
  XOR U915 ( .A(B[287]), .B(B[286]), .Z(n610) );
  XOR U916 ( .A(B[285]), .B(n611), .Z(O[286]) );
  AND U917 ( .A(S), .B(n612), .Z(n611) );
  XOR U918 ( .A(B[286]), .B(B[285]), .Z(n612) );
  XOR U919 ( .A(B[284]), .B(n613), .Z(O[285]) );
  AND U920 ( .A(S), .B(n614), .Z(n613) );
  XOR U921 ( .A(B[285]), .B(B[284]), .Z(n614) );
  XOR U922 ( .A(B[283]), .B(n615), .Z(O[284]) );
  AND U923 ( .A(S), .B(n616), .Z(n615) );
  XOR U924 ( .A(B[284]), .B(B[283]), .Z(n616) );
  XOR U925 ( .A(B[282]), .B(n617), .Z(O[283]) );
  AND U926 ( .A(S), .B(n618), .Z(n617) );
  XOR U927 ( .A(B[283]), .B(B[282]), .Z(n618) );
  XOR U928 ( .A(B[281]), .B(n619), .Z(O[282]) );
  AND U929 ( .A(S), .B(n620), .Z(n619) );
  XOR U930 ( .A(B[282]), .B(B[281]), .Z(n620) );
  XOR U931 ( .A(B[280]), .B(n621), .Z(O[281]) );
  AND U932 ( .A(S), .B(n622), .Z(n621) );
  XOR U933 ( .A(B[281]), .B(B[280]), .Z(n622) );
  XOR U934 ( .A(B[279]), .B(n623), .Z(O[280]) );
  AND U935 ( .A(S), .B(n624), .Z(n623) );
  XOR U936 ( .A(B[280]), .B(B[279]), .Z(n624) );
  XOR U937 ( .A(B[26]), .B(n625), .Z(O[27]) );
  AND U938 ( .A(S), .B(n626), .Z(n625) );
  XOR U939 ( .A(B[27]), .B(B[26]), .Z(n626) );
  XOR U940 ( .A(B[278]), .B(n627), .Z(O[279]) );
  AND U941 ( .A(S), .B(n628), .Z(n627) );
  XOR U942 ( .A(B[279]), .B(B[278]), .Z(n628) );
  XOR U943 ( .A(B[277]), .B(n629), .Z(O[278]) );
  AND U944 ( .A(S), .B(n630), .Z(n629) );
  XOR U945 ( .A(B[278]), .B(B[277]), .Z(n630) );
  XOR U946 ( .A(B[276]), .B(n631), .Z(O[277]) );
  AND U947 ( .A(S), .B(n632), .Z(n631) );
  XOR U948 ( .A(B[277]), .B(B[276]), .Z(n632) );
  XOR U949 ( .A(B[275]), .B(n633), .Z(O[276]) );
  AND U950 ( .A(S), .B(n634), .Z(n633) );
  XOR U951 ( .A(B[276]), .B(B[275]), .Z(n634) );
  XOR U952 ( .A(B[274]), .B(n635), .Z(O[275]) );
  AND U953 ( .A(S), .B(n636), .Z(n635) );
  XOR U954 ( .A(B[275]), .B(B[274]), .Z(n636) );
  XOR U955 ( .A(B[273]), .B(n637), .Z(O[274]) );
  AND U956 ( .A(S), .B(n638), .Z(n637) );
  XOR U957 ( .A(B[274]), .B(B[273]), .Z(n638) );
  XOR U958 ( .A(B[272]), .B(n639), .Z(O[273]) );
  AND U959 ( .A(S), .B(n640), .Z(n639) );
  XOR U960 ( .A(B[273]), .B(B[272]), .Z(n640) );
  XOR U961 ( .A(B[271]), .B(n641), .Z(O[272]) );
  AND U962 ( .A(S), .B(n642), .Z(n641) );
  XOR U963 ( .A(B[272]), .B(B[271]), .Z(n642) );
  XOR U964 ( .A(B[270]), .B(n643), .Z(O[271]) );
  AND U965 ( .A(S), .B(n644), .Z(n643) );
  XOR U966 ( .A(B[271]), .B(B[270]), .Z(n644) );
  XOR U967 ( .A(B[269]), .B(n645), .Z(O[270]) );
  AND U968 ( .A(S), .B(n646), .Z(n645) );
  XOR U969 ( .A(B[270]), .B(B[269]), .Z(n646) );
  XOR U970 ( .A(B[25]), .B(n647), .Z(O[26]) );
  AND U971 ( .A(S), .B(n648), .Z(n647) );
  XOR U972 ( .A(B[26]), .B(B[25]), .Z(n648) );
  XOR U973 ( .A(B[268]), .B(n649), .Z(O[269]) );
  AND U974 ( .A(S), .B(n650), .Z(n649) );
  XOR U975 ( .A(B[269]), .B(B[268]), .Z(n650) );
  XOR U976 ( .A(B[267]), .B(n651), .Z(O[268]) );
  AND U977 ( .A(S), .B(n652), .Z(n651) );
  XOR U978 ( .A(B[268]), .B(B[267]), .Z(n652) );
  XOR U979 ( .A(B[266]), .B(n653), .Z(O[267]) );
  AND U980 ( .A(S), .B(n654), .Z(n653) );
  XOR U981 ( .A(B[267]), .B(B[266]), .Z(n654) );
  XOR U982 ( .A(B[265]), .B(n655), .Z(O[266]) );
  AND U983 ( .A(S), .B(n656), .Z(n655) );
  XOR U984 ( .A(B[266]), .B(B[265]), .Z(n656) );
  XOR U985 ( .A(B[264]), .B(n657), .Z(O[265]) );
  AND U986 ( .A(S), .B(n658), .Z(n657) );
  XOR U987 ( .A(B[265]), .B(B[264]), .Z(n658) );
  XOR U988 ( .A(B[263]), .B(n659), .Z(O[264]) );
  AND U989 ( .A(S), .B(n660), .Z(n659) );
  XOR U990 ( .A(B[264]), .B(B[263]), .Z(n660) );
  XOR U991 ( .A(B[262]), .B(n661), .Z(O[263]) );
  AND U992 ( .A(S), .B(n662), .Z(n661) );
  XOR U993 ( .A(B[263]), .B(B[262]), .Z(n662) );
  XOR U994 ( .A(B[261]), .B(n663), .Z(O[262]) );
  AND U995 ( .A(S), .B(n664), .Z(n663) );
  XOR U996 ( .A(B[262]), .B(B[261]), .Z(n664) );
  XOR U997 ( .A(B[260]), .B(n665), .Z(O[261]) );
  AND U998 ( .A(S), .B(n666), .Z(n665) );
  XOR U999 ( .A(B[261]), .B(B[260]), .Z(n666) );
  XOR U1000 ( .A(B[259]), .B(n667), .Z(O[260]) );
  AND U1001 ( .A(S), .B(n668), .Z(n667) );
  XOR U1002 ( .A(B[260]), .B(B[259]), .Z(n668) );
  XOR U1003 ( .A(B[24]), .B(n669), .Z(O[25]) );
  AND U1004 ( .A(S), .B(n670), .Z(n669) );
  XOR U1005 ( .A(B[25]), .B(B[24]), .Z(n670) );
  XOR U1006 ( .A(B[258]), .B(n671), .Z(O[259]) );
  AND U1007 ( .A(S), .B(n672), .Z(n671) );
  XOR U1008 ( .A(B[259]), .B(B[258]), .Z(n672) );
  XOR U1009 ( .A(B[257]), .B(n673), .Z(O[258]) );
  AND U1010 ( .A(S), .B(n674), .Z(n673) );
  XOR U1011 ( .A(B[258]), .B(B[257]), .Z(n674) );
  XOR U1012 ( .A(B[256]), .B(n675), .Z(O[257]) );
  AND U1013 ( .A(S), .B(n676), .Z(n675) );
  XOR U1014 ( .A(B[257]), .B(B[256]), .Z(n676) );
  XOR U1015 ( .A(B[255]), .B(n677), .Z(O[256]) );
  AND U1016 ( .A(S), .B(n678), .Z(n677) );
  XOR U1017 ( .A(B[256]), .B(B[255]), .Z(n678) );
  XOR U1018 ( .A(B[254]), .B(n679), .Z(O[255]) );
  AND U1019 ( .A(S), .B(n680), .Z(n679) );
  XOR U1020 ( .A(B[255]), .B(B[254]), .Z(n680) );
  XOR U1021 ( .A(B[253]), .B(n681), .Z(O[254]) );
  AND U1022 ( .A(S), .B(n682), .Z(n681) );
  XOR U1023 ( .A(B[254]), .B(B[253]), .Z(n682) );
  XOR U1024 ( .A(B[252]), .B(n683), .Z(O[253]) );
  AND U1025 ( .A(S), .B(n684), .Z(n683) );
  XOR U1026 ( .A(B[253]), .B(B[252]), .Z(n684) );
  XOR U1027 ( .A(B[251]), .B(n685), .Z(O[252]) );
  AND U1028 ( .A(S), .B(n686), .Z(n685) );
  XOR U1029 ( .A(B[252]), .B(B[251]), .Z(n686) );
  XOR U1030 ( .A(B[250]), .B(n687), .Z(O[251]) );
  AND U1031 ( .A(S), .B(n688), .Z(n687) );
  XOR U1032 ( .A(B[251]), .B(B[250]), .Z(n688) );
  XOR U1033 ( .A(B[249]), .B(n689), .Z(O[250]) );
  AND U1034 ( .A(S), .B(n690), .Z(n689) );
  XOR U1035 ( .A(B[250]), .B(B[249]), .Z(n690) );
  XOR U1036 ( .A(B[23]), .B(n691), .Z(O[24]) );
  AND U1037 ( .A(S), .B(n692), .Z(n691) );
  XOR U1038 ( .A(B[24]), .B(B[23]), .Z(n692) );
  XOR U1039 ( .A(B[248]), .B(n693), .Z(O[249]) );
  AND U1040 ( .A(S), .B(n694), .Z(n693) );
  XOR U1041 ( .A(B[249]), .B(B[248]), .Z(n694) );
  XOR U1042 ( .A(B[247]), .B(n695), .Z(O[248]) );
  AND U1043 ( .A(S), .B(n696), .Z(n695) );
  XOR U1044 ( .A(B[248]), .B(B[247]), .Z(n696) );
  XOR U1045 ( .A(B[246]), .B(n697), .Z(O[247]) );
  AND U1046 ( .A(S), .B(n698), .Z(n697) );
  XOR U1047 ( .A(B[247]), .B(B[246]), .Z(n698) );
  XOR U1048 ( .A(B[245]), .B(n699), .Z(O[246]) );
  AND U1049 ( .A(S), .B(n700), .Z(n699) );
  XOR U1050 ( .A(B[246]), .B(B[245]), .Z(n700) );
  XOR U1051 ( .A(B[244]), .B(n701), .Z(O[245]) );
  AND U1052 ( .A(S), .B(n702), .Z(n701) );
  XOR U1053 ( .A(B[245]), .B(B[244]), .Z(n702) );
  XOR U1054 ( .A(B[243]), .B(n703), .Z(O[244]) );
  AND U1055 ( .A(S), .B(n704), .Z(n703) );
  XOR U1056 ( .A(B[244]), .B(B[243]), .Z(n704) );
  XOR U1057 ( .A(B[242]), .B(n705), .Z(O[243]) );
  AND U1058 ( .A(S), .B(n706), .Z(n705) );
  XOR U1059 ( .A(B[243]), .B(B[242]), .Z(n706) );
  XOR U1060 ( .A(B[241]), .B(n707), .Z(O[242]) );
  AND U1061 ( .A(S), .B(n708), .Z(n707) );
  XOR U1062 ( .A(B[242]), .B(B[241]), .Z(n708) );
  XOR U1063 ( .A(B[240]), .B(n709), .Z(O[241]) );
  AND U1064 ( .A(S), .B(n710), .Z(n709) );
  XOR U1065 ( .A(B[241]), .B(B[240]), .Z(n710) );
  XOR U1066 ( .A(B[239]), .B(n711), .Z(O[240]) );
  AND U1067 ( .A(S), .B(n712), .Z(n711) );
  XOR U1068 ( .A(B[240]), .B(B[239]), .Z(n712) );
  XOR U1069 ( .A(B[22]), .B(n713), .Z(O[23]) );
  AND U1070 ( .A(S), .B(n714), .Z(n713) );
  XOR U1071 ( .A(B[23]), .B(B[22]), .Z(n714) );
  XOR U1072 ( .A(B[238]), .B(n715), .Z(O[239]) );
  AND U1073 ( .A(S), .B(n716), .Z(n715) );
  XOR U1074 ( .A(B[239]), .B(B[238]), .Z(n716) );
  XOR U1075 ( .A(B[237]), .B(n717), .Z(O[238]) );
  AND U1076 ( .A(S), .B(n718), .Z(n717) );
  XOR U1077 ( .A(B[238]), .B(B[237]), .Z(n718) );
  XOR U1078 ( .A(B[236]), .B(n719), .Z(O[237]) );
  AND U1079 ( .A(S), .B(n720), .Z(n719) );
  XOR U1080 ( .A(B[237]), .B(B[236]), .Z(n720) );
  XOR U1081 ( .A(B[235]), .B(n721), .Z(O[236]) );
  AND U1082 ( .A(S), .B(n722), .Z(n721) );
  XOR U1083 ( .A(B[236]), .B(B[235]), .Z(n722) );
  XOR U1084 ( .A(B[234]), .B(n723), .Z(O[235]) );
  AND U1085 ( .A(S), .B(n724), .Z(n723) );
  XOR U1086 ( .A(B[235]), .B(B[234]), .Z(n724) );
  XOR U1087 ( .A(B[233]), .B(n725), .Z(O[234]) );
  AND U1088 ( .A(S), .B(n726), .Z(n725) );
  XOR U1089 ( .A(B[234]), .B(B[233]), .Z(n726) );
  XOR U1090 ( .A(B[232]), .B(n727), .Z(O[233]) );
  AND U1091 ( .A(S), .B(n728), .Z(n727) );
  XOR U1092 ( .A(B[233]), .B(B[232]), .Z(n728) );
  XOR U1093 ( .A(B[231]), .B(n729), .Z(O[232]) );
  AND U1094 ( .A(S), .B(n730), .Z(n729) );
  XOR U1095 ( .A(B[232]), .B(B[231]), .Z(n730) );
  XOR U1096 ( .A(B[230]), .B(n731), .Z(O[231]) );
  AND U1097 ( .A(S), .B(n732), .Z(n731) );
  XOR U1098 ( .A(B[231]), .B(B[230]), .Z(n732) );
  XOR U1099 ( .A(B[229]), .B(n733), .Z(O[230]) );
  AND U1100 ( .A(S), .B(n734), .Z(n733) );
  XOR U1101 ( .A(B[230]), .B(B[229]), .Z(n734) );
  XOR U1102 ( .A(B[21]), .B(n735), .Z(O[22]) );
  AND U1103 ( .A(S), .B(n736), .Z(n735) );
  XOR U1104 ( .A(B[22]), .B(B[21]), .Z(n736) );
  XOR U1105 ( .A(B[228]), .B(n737), .Z(O[229]) );
  AND U1106 ( .A(S), .B(n738), .Z(n737) );
  XOR U1107 ( .A(B[229]), .B(B[228]), .Z(n738) );
  XOR U1108 ( .A(B[227]), .B(n739), .Z(O[228]) );
  AND U1109 ( .A(S), .B(n740), .Z(n739) );
  XOR U1110 ( .A(B[228]), .B(B[227]), .Z(n740) );
  XOR U1111 ( .A(B[226]), .B(n741), .Z(O[227]) );
  AND U1112 ( .A(S), .B(n742), .Z(n741) );
  XOR U1113 ( .A(B[227]), .B(B[226]), .Z(n742) );
  XOR U1114 ( .A(B[225]), .B(n743), .Z(O[226]) );
  AND U1115 ( .A(S), .B(n744), .Z(n743) );
  XOR U1116 ( .A(B[226]), .B(B[225]), .Z(n744) );
  XOR U1117 ( .A(B[224]), .B(n745), .Z(O[225]) );
  AND U1118 ( .A(S), .B(n746), .Z(n745) );
  XOR U1119 ( .A(B[225]), .B(B[224]), .Z(n746) );
  XOR U1120 ( .A(B[223]), .B(n747), .Z(O[224]) );
  AND U1121 ( .A(S), .B(n748), .Z(n747) );
  XOR U1122 ( .A(B[224]), .B(B[223]), .Z(n748) );
  XOR U1123 ( .A(B[222]), .B(n749), .Z(O[223]) );
  AND U1124 ( .A(S), .B(n750), .Z(n749) );
  XOR U1125 ( .A(B[223]), .B(B[222]), .Z(n750) );
  XOR U1126 ( .A(B[221]), .B(n751), .Z(O[222]) );
  AND U1127 ( .A(S), .B(n752), .Z(n751) );
  XOR U1128 ( .A(B[222]), .B(B[221]), .Z(n752) );
  XOR U1129 ( .A(B[220]), .B(n753), .Z(O[221]) );
  AND U1130 ( .A(S), .B(n754), .Z(n753) );
  XOR U1131 ( .A(B[221]), .B(B[220]), .Z(n754) );
  XOR U1132 ( .A(B[219]), .B(n755), .Z(O[220]) );
  AND U1133 ( .A(S), .B(n756), .Z(n755) );
  XOR U1134 ( .A(B[220]), .B(B[219]), .Z(n756) );
  XOR U1135 ( .A(B[20]), .B(n757), .Z(O[21]) );
  AND U1136 ( .A(S), .B(n758), .Z(n757) );
  XOR U1137 ( .A(B[21]), .B(B[20]), .Z(n758) );
  XOR U1138 ( .A(B[218]), .B(n759), .Z(O[219]) );
  AND U1139 ( .A(S), .B(n760), .Z(n759) );
  XOR U1140 ( .A(B[219]), .B(B[218]), .Z(n760) );
  XOR U1141 ( .A(B[217]), .B(n761), .Z(O[218]) );
  AND U1142 ( .A(S), .B(n762), .Z(n761) );
  XOR U1143 ( .A(B[218]), .B(B[217]), .Z(n762) );
  XOR U1144 ( .A(B[216]), .B(n763), .Z(O[217]) );
  AND U1145 ( .A(S), .B(n764), .Z(n763) );
  XOR U1146 ( .A(B[217]), .B(B[216]), .Z(n764) );
  XOR U1147 ( .A(B[215]), .B(n765), .Z(O[216]) );
  AND U1148 ( .A(S), .B(n766), .Z(n765) );
  XOR U1149 ( .A(B[216]), .B(B[215]), .Z(n766) );
  XOR U1150 ( .A(B[214]), .B(n767), .Z(O[215]) );
  AND U1151 ( .A(S), .B(n768), .Z(n767) );
  XOR U1152 ( .A(B[215]), .B(B[214]), .Z(n768) );
  XOR U1153 ( .A(B[213]), .B(n769), .Z(O[214]) );
  AND U1154 ( .A(S), .B(n770), .Z(n769) );
  XOR U1155 ( .A(B[214]), .B(B[213]), .Z(n770) );
  XOR U1156 ( .A(B[212]), .B(n771), .Z(O[213]) );
  AND U1157 ( .A(S), .B(n772), .Z(n771) );
  XOR U1158 ( .A(B[213]), .B(B[212]), .Z(n772) );
  XOR U1159 ( .A(B[211]), .B(n773), .Z(O[212]) );
  AND U1160 ( .A(S), .B(n774), .Z(n773) );
  XOR U1161 ( .A(B[212]), .B(B[211]), .Z(n774) );
  XOR U1162 ( .A(B[210]), .B(n775), .Z(O[211]) );
  AND U1163 ( .A(S), .B(n776), .Z(n775) );
  XOR U1164 ( .A(B[211]), .B(B[210]), .Z(n776) );
  XOR U1165 ( .A(B[209]), .B(n777), .Z(O[210]) );
  AND U1166 ( .A(S), .B(n778), .Z(n777) );
  XOR U1167 ( .A(B[210]), .B(B[209]), .Z(n778) );
  XOR U1168 ( .A(B[19]), .B(n779), .Z(O[20]) );
  AND U1169 ( .A(S), .B(n780), .Z(n779) );
  XOR U1170 ( .A(B[20]), .B(B[19]), .Z(n780) );
  XOR U1171 ( .A(B[208]), .B(n781), .Z(O[209]) );
  AND U1172 ( .A(S), .B(n782), .Z(n781) );
  XOR U1173 ( .A(B[209]), .B(B[208]), .Z(n782) );
  XOR U1174 ( .A(B[207]), .B(n783), .Z(O[208]) );
  AND U1175 ( .A(S), .B(n784), .Z(n783) );
  XOR U1176 ( .A(B[208]), .B(B[207]), .Z(n784) );
  XOR U1177 ( .A(B[206]), .B(n785), .Z(O[207]) );
  AND U1178 ( .A(S), .B(n786), .Z(n785) );
  XOR U1179 ( .A(B[207]), .B(B[206]), .Z(n786) );
  XOR U1180 ( .A(B[205]), .B(n787), .Z(O[206]) );
  AND U1181 ( .A(S), .B(n788), .Z(n787) );
  XOR U1182 ( .A(B[206]), .B(B[205]), .Z(n788) );
  XOR U1183 ( .A(B[204]), .B(n789), .Z(O[205]) );
  AND U1184 ( .A(S), .B(n790), .Z(n789) );
  XOR U1185 ( .A(B[205]), .B(B[204]), .Z(n790) );
  XOR U1186 ( .A(B[203]), .B(n791), .Z(O[204]) );
  AND U1187 ( .A(S), .B(n792), .Z(n791) );
  XOR U1188 ( .A(B[204]), .B(B[203]), .Z(n792) );
  XOR U1189 ( .A(B[202]), .B(n793), .Z(O[203]) );
  AND U1190 ( .A(S), .B(n794), .Z(n793) );
  XOR U1191 ( .A(B[203]), .B(B[202]), .Z(n794) );
  XOR U1192 ( .A(B[201]), .B(n795), .Z(O[202]) );
  AND U1193 ( .A(S), .B(n796), .Z(n795) );
  XOR U1194 ( .A(B[202]), .B(B[201]), .Z(n796) );
  XOR U1195 ( .A(B[200]), .B(n797), .Z(O[201]) );
  AND U1196 ( .A(S), .B(n798), .Z(n797) );
  XOR U1197 ( .A(B[201]), .B(B[200]), .Z(n798) );
  XOR U1198 ( .A(B[199]), .B(n799), .Z(O[200]) );
  AND U1199 ( .A(S), .B(n800), .Z(n799) );
  XOR U1200 ( .A(B[200]), .B(B[199]), .Z(n800) );
  XOR U1201 ( .A(B[0]), .B(n801), .Z(O[1]) );
  AND U1202 ( .A(S), .B(n802), .Z(n801) );
  XOR U1203 ( .A(B[1]), .B(B[0]), .Z(n802) );
  XOR U1204 ( .A(B[18]), .B(n803), .Z(O[19]) );
  AND U1205 ( .A(S), .B(n804), .Z(n803) );
  XOR U1206 ( .A(B[19]), .B(B[18]), .Z(n804) );
  XOR U1207 ( .A(B[198]), .B(n805), .Z(O[199]) );
  AND U1208 ( .A(S), .B(n806), .Z(n805) );
  XOR U1209 ( .A(B[199]), .B(B[198]), .Z(n806) );
  XOR U1210 ( .A(B[197]), .B(n807), .Z(O[198]) );
  AND U1211 ( .A(S), .B(n808), .Z(n807) );
  XOR U1212 ( .A(B[198]), .B(B[197]), .Z(n808) );
  XOR U1213 ( .A(B[196]), .B(n809), .Z(O[197]) );
  AND U1214 ( .A(S), .B(n810), .Z(n809) );
  XOR U1215 ( .A(B[197]), .B(B[196]), .Z(n810) );
  XOR U1216 ( .A(B[195]), .B(n811), .Z(O[196]) );
  AND U1217 ( .A(S), .B(n812), .Z(n811) );
  XOR U1218 ( .A(B[196]), .B(B[195]), .Z(n812) );
  XOR U1219 ( .A(B[194]), .B(n813), .Z(O[195]) );
  AND U1220 ( .A(S), .B(n814), .Z(n813) );
  XOR U1221 ( .A(B[195]), .B(B[194]), .Z(n814) );
  XOR U1222 ( .A(B[193]), .B(n815), .Z(O[194]) );
  AND U1223 ( .A(S), .B(n816), .Z(n815) );
  XOR U1224 ( .A(B[194]), .B(B[193]), .Z(n816) );
  XOR U1225 ( .A(B[192]), .B(n817), .Z(O[193]) );
  AND U1226 ( .A(S), .B(n818), .Z(n817) );
  XOR U1227 ( .A(B[193]), .B(B[192]), .Z(n818) );
  XOR U1228 ( .A(B[191]), .B(n819), .Z(O[192]) );
  AND U1229 ( .A(S), .B(n820), .Z(n819) );
  XOR U1230 ( .A(B[192]), .B(B[191]), .Z(n820) );
  XOR U1231 ( .A(B[190]), .B(n821), .Z(O[191]) );
  AND U1232 ( .A(S), .B(n822), .Z(n821) );
  XOR U1233 ( .A(B[191]), .B(B[190]), .Z(n822) );
  XOR U1234 ( .A(B[189]), .B(n823), .Z(O[190]) );
  AND U1235 ( .A(S), .B(n824), .Z(n823) );
  XOR U1236 ( .A(B[190]), .B(B[189]), .Z(n824) );
  XOR U1237 ( .A(B[17]), .B(n825), .Z(O[18]) );
  AND U1238 ( .A(S), .B(n826), .Z(n825) );
  XOR U1239 ( .A(B[18]), .B(B[17]), .Z(n826) );
  XOR U1240 ( .A(B[188]), .B(n827), .Z(O[189]) );
  AND U1241 ( .A(S), .B(n828), .Z(n827) );
  XOR U1242 ( .A(B[189]), .B(B[188]), .Z(n828) );
  XOR U1243 ( .A(B[187]), .B(n829), .Z(O[188]) );
  AND U1244 ( .A(S), .B(n830), .Z(n829) );
  XOR U1245 ( .A(B[188]), .B(B[187]), .Z(n830) );
  XOR U1246 ( .A(B[186]), .B(n831), .Z(O[187]) );
  AND U1247 ( .A(S), .B(n832), .Z(n831) );
  XOR U1248 ( .A(B[187]), .B(B[186]), .Z(n832) );
  XOR U1249 ( .A(B[185]), .B(n833), .Z(O[186]) );
  AND U1250 ( .A(S), .B(n834), .Z(n833) );
  XOR U1251 ( .A(B[186]), .B(B[185]), .Z(n834) );
  XOR U1252 ( .A(B[184]), .B(n835), .Z(O[185]) );
  AND U1253 ( .A(S), .B(n836), .Z(n835) );
  XOR U1254 ( .A(B[185]), .B(B[184]), .Z(n836) );
  XOR U1255 ( .A(B[183]), .B(n837), .Z(O[184]) );
  AND U1256 ( .A(S), .B(n838), .Z(n837) );
  XOR U1257 ( .A(B[184]), .B(B[183]), .Z(n838) );
  XOR U1258 ( .A(B[182]), .B(n839), .Z(O[183]) );
  AND U1259 ( .A(S), .B(n840), .Z(n839) );
  XOR U1260 ( .A(B[183]), .B(B[182]), .Z(n840) );
  XOR U1261 ( .A(B[181]), .B(n841), .Z(O[182]) );
  AND U1262 ( .A(S), .B(n842), .Z(n841) );
  XOR U1263 ( .A(B[182]), .B(B[181]), .Z(n842) );
  XOR U1264 ( .A(B[180]), .B(n843), .Z(O[181]) );
  AND U1265 ( .A(S), .B(n844), .Z(n843) );
  XOR U1266 ( .A(B[181]), .B(B[180]), .Z(n844) );
  XOR U1267 ( .A(B[179]), .B(n845), .Z(O[180]) );
  AND U1268 ( .A(S), .B(n846), .Z(n845) );
  XOR U1269 ( .A(B[180]), .B(B[179]), .Z(n846) );
  XOR U1270 ( .A(B[16]), .B(n847), .Z(O[17]) );
  AND U1271 ( .A(S), .B(n848), .Z(n847) );
  XOR U1272 ( .A(B[17]), .B(B[16]), .Z(n848) );
  XOR U1273 ( .A(B[178]), .B(n849), .Z(O[179]) );
  AND U1274 ( .A(S), .B(n850), .Z(n849) );
  XOR U1275 ( .A(B[179]), .B(B[178]), .Z(n850) );
  XOR U1276 ( .A(B[177]), .B(n851), .Z(O[178]) );
  AND U1277 ( .A(S), .B(n852), .Z(n851) );
  XOR U1278 ( .A(B[178]), .B(B[177]), .Z(n852) );
  XOR U1279 ( .A(B[176]), .B(n853), .Z(O[177]) );
  AND U1280 ( .A(S), .B(n854), .Z(n853) );
  XOR U1281 ( .A(B[177]), .B(B[176]), .Z(n854) );
  XOR U1282 ( .A(B[175]), .B(n855), .Z(O[176]) );
  AND U1283 ( .A(S), .B(n856), .Z(n855) );
  XOR U1284 ( .A(B[176]), .B(B[175]), .Z(n856) );
  XOR U1285 ( .A(B[174]), .B(n857), .Z(O[175]) );
  AND U1286 ( .A(S), .B(n858), .Z(n857) );
  XOR U1287 ( .A(B[175]), .B(B[174]), .Z(n858) );
  XOR U1288 ( .A(B[173]), .B(n859), .Z(O[174]) );
  AND U1289 ( .A(S), .B(n860), .Z(n859) );
  XOR U1290 ( .A(B[174]), .B(B[173]), .Z(n860) );
  XOR U1291 ( .A(B[172]), .B(n861), .Z(O[173]) );
  AND U1292 ( .A(S), .B(n862), .Z(n861) );
  XOR U1293 ( .A(B[173]), .B(B[172]), .Z(n862) );
  XOR U1294 ( .A(B[171]), .B(n863), .Z(O[172]) );
  AND U1295 ( .A(S), .B(n864), .Z(n863) );
  XOR U1296 ( .A(B[172]), .B(B[171]), .Z(n864) );
  XOR U1297 ( .A(B[170]), .B(n865), .Z(O[171]) );
  AND U1298 ( .A(S), .B(n866), .Z(n865) );
  XOR U1299 ( .A(B[171]), .B(B[170]), .Z(n866) );
  XOR U1300 ( .A(B[169]), .B(n867), .Z(O[170]) );
  AND U1301 ( .A(S), .B(n868), .Z(n867) );
  XOR U1302 ( .A(B[170]), .B(B[169]), .Z(n868) );
  XOR U1303 ( .A(B[15]), .B(n869), .Z(O[16]) );
  AND U1304 ( .A(S), .B(n870), .Z(n869) );
  XOR U1305 ( .A(B[16]), .B(B[15]), .Z(n870) );
  XOR U1306 ( .A(B[168]), .B(n871), .Z(O[169]) );
  AND U1307 ( .A(S), .B(n872), .Z(n871) );
  XOR U1308 ( .A(B[169]), .B(B[168]), .Z(n872) );
  XOR U1309 ( .A(B[167]), .B(n873), .Z(O[168]) );
  AND U1310 ( .A(S), .B(n874), .Z(n873) );
  XOR U1311 ( .A(B[168]), .B(B[167]), .Z(n874) );
  XOR U1312 ( .A(B[166]), .B(n875), .Z(O[167]) );
  AND U1313 ( .A(S), .B(n876), .Z(n875) );
  XOR U1314 ( .A(B[167]), .B(B[166]), .Z(n876) );
  XOR U1315 ( .A(B[165]), .B(n877), .Z(O[166]) );
  AND U1316 ( .A(S), .B(n878), .Z(n877) );
  XOR U1317 ( .A(B[166]), .B(B[165]), .Z(n878) );
  XOR U1318 ( .A(B[164]), .B(n879), .Z(O[165]) );
  AND U1319 ( .A(S), .B(n880), .Z(n879) );
  XOR U1320 ( .A(B[165]), .B(B[164]), .Z(n880) );
  XOR U1321 ( .A(B[163]), .B(n881), .Z(O[164]) );
  AND U1322 ( .A(S), .B(n882), .Z(n881) );
  XOR U1323 ( .A(B[164]), .B(B[163]), .Z(n882) );
  XOR U1324 ( .A(B[162]), .B(n883), .Z(O[163]) );
  AND U1325 ( .A(S), .B(n884), .Z(n883) );
  XOR U1326 ( .A(B[163]), .B(B[162]), .Z(n884) );
  XOR U1327 ( .A(B[161]), .B(n885), .Z(O[162]) );
  AND U1328 ( .A(S), .B(n886), .Z(n885) );
  XOR U1329 ( .A(B[162]), .B(B[161]), .Z(n886) );
  XOR U1330 ( .A(B[160]), .B(n887), .Z(O[161]) );
  AND U1331 ( .A(S), .B(n888), .Z(n887) );
  XOR U1332 ( .A(B[161]), .B(B[160]), .Z(n888) );
  XOR U1333 ( .A(B[159]), .B(n889), .Z(O[160]) );
  AND U1334 ( .A(S), .B(n890), .Z(n889) );
  XOR U1335 ( .A(B[160]), .B(B[159]), .Z(n890) );
  XOR U1336 ( .A(B[14]), .B(n891), .Z(O[15]) );
  AND U1337 ( .A(S), .B(n892), .Z(n891) );
  XOR U1338 ( .A(B[15]), .B(B[14]), .Z(n892) );
  XOR U1339 ( .A(B[158]), .B(n893), .Z(O[159]) );
  AND U1340 ( .A(S), .B(n894), .Z(n893) );
  XOR U1341 ( .A(B[159]), .B(B[158]), .Z(n894) );
  XOR U1342 ( .A(B[157]), .B(n895), .Z(O[158]) );
  AND U1343 ( .A(S), .B(n896), .Z(n895) );
  XOR U1344 ( .A(B[158]), .B(B[157]), .Z(n896) );
  XOR U1345 ( .A(B[156]), .B(n897), .Z(O[157]) );
  AND U1346 ( .A(S), .B(n898), .Z(n897) );
  XOR U1347 ( .A(B[157]), .B(B[156]), .Z(n898) );
  XOR U1348 ( .A(B[155]), .B(n899), .Z(O[156]) );
  AND U1349 ( .A(S), .B(n900), .Z(n899) );
  XOR U1350 ( .A(B[156]), .B(B[155]), .Z(n900) );
  XOR U1351 ( .A(B[154]), .B(n901), .Z(O[155]) );
  AND U1352 ( .A(S), .B(n902), .Z(n901) );
  XOR U1353 ( .A(B[155]), .B(B[154]), .Z(n902) );
  XOR U1354 ( .A(B[153]), .B(n903), .Z(O[154]) );
  AND U1355 ( .A(S), .B(n904), .Z(n903) );
  XOR U1356 ( .A(B[154]), .B(B[153]), .Z(n904) );
  XOR U1357 ( .A(B[152]), .B(n905), .Z(O[153]) );
  AND U1358 ( .A(S), .B(n906), .Z(n905) );
  XOR U1359 ( .A(B[153]), .B(B[152]), .Z(n906) );
  XOR U1360 ( .A(B[151]), .B(n907), .Z(O[152]) );
  AND U1361 ( .A(S), .B(n908), .Z(n907) );
  XOR U1362 ( .A(B[152]), .B(B[151]), .Z(n908) );
  XOR U1363 ( .A(B[150]), .B(n909), .Z(O[151]) );
  AND U1364 ( .A(S), .B(n910), .Z(n909) );
  XOR U1365 ( .A(B[151]), .B(B[150]), .Z(n910) );
  XOR U1366 ( .A(B[149]), .B(n911), .Z(O[150]) );
  AND U1367 ( .A(S), .B(n912), .Z(n911) );
  XOR U1368 ( .A(B[150]), .B(B[149]), .Z(n912) );
  XOR U1369 ( .A(B[13]), .B(n913), .Z(O[14]) );
  AND U1370 ( .A(S), .B(n914), .Z(n913) );
  XOR U1371 ( .A(B[14]), .B(B[13]), .Z(n914) );
  XOR U1372 ( .A(B[148]), .B(n915), .Z(O[149]) );
  AND U1373 ( .A(S), .B(n916), .Z(n915) );
  XOR U1374 ( .A(B[149]), .B(B[148]), .Z(n916) );
  XOR U1375 ( .A(B[147]), .B(n917), .Z(O[148]) );
  AND U1376 ( .A(S), .B(n918), .Z(n917) );
  XOR U1377 ( .A(B[148]), .B(B[147]), .Z(n918) );
  XOR U1378 ( .A(B[146]), .B(n919), .Z(O[147]) );
  AND U1379 ( .A(S), .B(n920), .Z(n919) );
  XOR U1380 ( .A(B[147]), .B(B[146]), .Z(n920) );
  XOR U1381 ( .A(B[145]), .B(n921), .Z(O[146]) );
  AND U1382 ( .A(S), .B(n922), .Z(n921) );
  XOR U1383 ( .A(B[146]), .B(B[145]), .Z(n922) );
  XOR U1384 ( .A(B[144]), .B(n923), .Z(O[145]) );
  AND U1385 ( .A(S), .B(n924), .Z(n923) );
  XOR U1386 ( .A(B[145]), .B(B[144]), .Z(n924) );
  XOR U1387 ( .A(B[143]), .B(n925), .Z(O[144]) );
  AND U1388 ( .A(S), .B(n926), .Z(n925) );
  XOR U1389 ( .A(B[144]), .B(B[143]), .Z(n926) );
  XOR U1390 ( .A(B[142]), .B(n927), .Z(O[143]) );
  AND U1391 ( .A(S), .B(n928), .Z(n927) );
  XOR U1392 ( .A(B[143]), .B(B[142]), .Z(n928) );
  XOR U1393 ( .A(B[141]), .B(n929), .Z(O[142]) );
  AND U1394 ( .A(S), .B(n930), .Z(n929) );
  XOR U1395 ( .A(B[142]), .B(B[141]), .Z(n930) );
  XOR U1396 ( .A(B[140]), .B(n931), .Z(O[141]) );
  AND U1397 ( .A(S), .B(n932), .Z(n931) );
  XOR U1398 ( .A(B[141]), .B(B[140]), .Z(n932) );
  XOR U1399 ( .A(B[139]), .B(n933), .Z(O[140]) );
  AND U1400 ( .A(S), .B(n934), .Z(n933) );
  XOR U1401 ( .A(B[140]), .B(B[139]), .Z(n934) );
  XOR U1402 ( .A(B[12]), .B(n935), .Z(O[13]) );
  AND U1403 ( .A(S), .B(n936), .Z(n935) );
  XOR U1404 ( .A(B[13]), .B(B[12]), .Z(n936) );
  XOR U1405 ( .A(B[138]), .B(n937), .Z(O[139]) );
  AND U1406 ( .A(S), .B(n938), .Z(n937) );
  XOR U1407 ( .A(B[139]), .B(B[138]), .Z(n938) );
  XOR U1408 ( .A(B[137]), .B(n939), .Z(O[138]) );
  AND U1409 ( .A(S), .B(n940), .Z(n939) );
  XOR U1410 ( .A(B[138]), .B(B[137]), .Z(n940) );
  XOR U1411 ( .A(B[136]), .B(n941), .Z(O[137]) );
  AND U1412 ( .A(S), .B(n942), .Z(n941) );
  XOR U1413 ( .A(B[137]), .B(B[136]), .Z(n942) );
  XOR U1414 ( .A(B[135]), .B(n943), .Z(O[136]) );
  AND U1415 ( .A(S), .B(n944), .Z(n943) );
  XOR U1416 ( .A(B[136]), .B(B[135]), .Z(n944) );
  XOR U1417 ( .A(B[134]), .B(n945), .Z(O[135]) );
  AND U1418 ( .A(S), .B(n946), .Z(n945) );
  XOR U1419 ( .A(B[135]), .B(B[134]), .Z(n946) );
  XOR U1420 ( .A(B[133]), .B(n947), .Z(O[134]) );
  AND U1421 ( .A(S), .B(n948), .Z(n947) );
  XOR U1422 ( .A(B[134]), .B(B[133]), .Z(n948) );
  XOR U1423 ( .A(B[132]), .B(n949), .Z(O[133]) );
  AND U1424 ( .A(S), .B(n950), .Z(n949) );
  XOR U1425 ( .A(B[133]), .B(B[132]), .Z(n950) );
  XOR U1426 ( .A(B[131]), .B(n951), .Z(O[132]) );
  AND U1427 ( .A(S), .B(n952), .Z(n951) );
  XOR U1428 ( .A(B[132]), .B(B[131]), .Z(n952) );
  XOR U1429 ( .A(B[130]), .B(n953), .Z(O[131]) );
  AND U1430 ( .A(S), .B(n954), .Z(n953) );
  XOR U1431 ( .A(B[131]), .B(B[130]), .Z(n954) );
  XOR U1432 ( .A(B[129]), .B(n955), .Z(O[130]) );
  AND U1433 ( .A(S), .B(n956), .Z(n955) );
  XOR U1434 ( .A(B[130]), .B(B[129]), .Z(n956) );
  XOR U1435 ( .A(B[11]), .B(n957), .Z(O[12]) );
  AND U1436 ( .A(S), .B(n958), .Z(n957) );
  XOR U1437 ( .A(B[12]), .B(B[11]), .Z(n958) );
  XOR U1438 ( .A(B[128]), .B(n959), .Z(O[129]) );
  AND U1439 ( .A(S), .B(n960), .Z(n959) );
  XOR U1440 ( .A(B[129]), .B(B[128]), .Z(n960) );
  XOR U1441 ( .A(B[127]), .B(n961), .Z(O[128]) );
  AND U1442 ( .A(S), .B(n962), .Z(n961) );
  XOR U1443 ( .A(B[128]), .B(B[127]), .Z(n962) );
  XOR U1444 ( .A(B[126]), .B(n963), .Z(O[127]) );
  AND U1445 ( .A(S), .B(n964), .Z(n963) );
  XOR U1446 ( .A(B[127]), .B(B[126]), .Z(n964) );
  XOR U1447 ( .A(B[125]), .B(n965), .Z(O[126]) );
  AND U1448 ( .A(S), .B(n966), .Z(n965) );
  XOR U1449 ( .A(B[126]), .B(B[125]), .Z(n966) );
  XOR U1450 ( .A(B[124]), .B(n967), .Z(O[125]) );
  AND U1451 ( .A(S), .B(n968), .Z(n967) );
  XOR U1452 ( .A(B[125]), .B(B[124]), .Z(n968) );
  XOR U1453 ( .A(B[123]), .B(n969), .Z(O[124]) );
  AND U1454 ( .A(S), .B(n970), .Z(n969) );
  XOR U1455 ( .A(B[124]), .B(B[123]), .Z(n970) );
  XOR U1456 ( .A(B[122]), .B(n971), .Z(O[123]) );
  AND U1457 ( .A(S), .B(n972), .Z(n971) );
  XOR U1458 ( .A(B[123]), .B(B[122]), .Z(n972) );
  XOR U1459 ( .A(B[121]), .B(n973), .Z(O[122]) );
  AND U1460 ( .A(S), .B(n974), .Z(n973) );
  XOR U1461 ( .A(B[122]), .B(B[121]), .Z(n974) );
  XOR U1462 ( .A(B[120]), .B(n975), .Z(O[121]) );
  AND U1463 ( .A(S), .B(n976), .Z(n975) );
  XOR U1464 ( .A(B[121]), .B(B[120]), .Z(n976) );
  XOR U1465 ( .A(B[119]), .B(n977), .Z(O[120]) );
  AND U1466 ( .A(S), .B(n978), .Z(n977) );
  XOR U1467 ( .A(B[120]), .B(B[119]), .Z(n978) );
  XOR U1468 ( .A(B[10]), .B(n979), .Z(O[11]) );
  AND U1469 ( .A(S), .B(n980), .Z(n979) );
  XOR U1470 ( .A(B[11]), .B(B[10]), .Z(n980) );
  XOR U1471 ( .A(B[118]), .B(n981), .Z(O[119]) );
  AND U1472 ( .A(S), .B(n982), .Z(n981) );
  XOR U1473 ( .A(B[119]), .B(B[118]), .Z(n982) );
  XOR U1474 ( .A(B[117]), .B(n983), .Z(O[118]) );
  AND U1475 ( .A(S), .B(n984), .Z(n983) );
  XOR U1476 ( .A(B[118]), .B(B[117]), .Z(n984) );
  XOR U1477 ( .A(B[116]), .B(n985), .Z(O[117]) );
  AND U1478 ( .A(S), .B(n986), .Z(n985) );
  XOR U1479 ( .A(B[117]), .B(B[116]), .Z(n986) );
  XOR U1480 ( .A(B[115]), .B(n987), .Z(O[116]) );
  AND U1481 ( .A(S), .B(n988), .Z(n987) );
  XOR U1482 ( .A(B[116]), .B(B[115]), .Z(n988) );
  XOR U1483 ( .A(B[114]), .B(n989), .Z(O[115]) );
  AND U1484 ( .A(S), .B(n990), .Z(n989) );
  XOR U1485 ( .A(B[115]), .B(B[114]), .Z(n990) );
  XOR U1486 ( .A(B[113]), .B(n991), .Z(O[114]) );
  AND U1487 ( .A(S), .B(n992), .Z(n991) );
  XOR U1488 ( .A(B[114]), .B(B[113]), .Z(n992) );
  XOR U1489 ( .A(B[112]), .B(n993), .Z(O[113]) );
  AND U1490 ( .A(S), .B(n994), .Z(n993) );
  XOR U1491 ( .A(B[113]), .B(B[112]), .Z(n994) );
  XOR U1492 ( .A(B[111]), .B(n995), .Z(O[112]) );
  AND U1493 ( .A(S), .B(n996), .Z(n995) );
  XOR U1494 ( .A(B[112]), .B(B[111]), .Z(n996) );
  XOR U1495 ( .A(B[110]), .B(n997), .Z(O[111]) );
  AND U1496 ( .A(S), .B(n998), .Z(n997) );
  XOR U1497 ( .A(B[111]), .B(B[110]), .Z(n998) );
  XOR U1498 ( .A(B[109]), .B(n999), .Z(O[110]) );
  AND U1499 ( .A(S), .B(n1000), .Z(n999) );
  XOR U1500 ( .A(B[110]), .B(B[109]), .Z(n1000) );
  XOR U1501 ( .A(B[9]), .B(n1001), .Z(O[10]) );
  AND U1502 ( .A(S), .B(n1002), .Z(n1001) );
  XOR U1503 ( .A(B[9]), .B(B[10]), .Z(n1002) );
  XOR U1504 ( .A(B[108]), .B(n1003), .Z(O[109]) );
  AND U1505 ( .A(S), .B(n1004), .Z(n1003) );
  XOR U1506 ( .A(B[109]), .B(B[108]), .Z(n1004) );
  XOR U1507 ( .A(B[107]), .B(n1005), .Z(O[108]) );
  AND U1508 ( .A(S), .B(n1006), .Z(n1005) );
  XOR U1509 ( .A(B[108]), .B(B[107]), .Z(n1006) );
  XOR U1510 ( .A(B[106]), .B(n1007), .Z(O[107]) );
  AND U1511 ( .A(S), .B(n1008), .Z(n1007) );
  XOR U1512 ( .A(B[107]), .B(B[106]), .Z(n1008) );
  XOR U1513 ( .A(B[105]), .B(n1009), .Z(O[106]) );
  AND U1514 ( .A(S), .B(n1010), .Z(n1009) );
  XOR U1515 ( .A(B[106]), .B(B[105]), .Z(n1010) );
  XOR U1516 ( .A(B[104]), .B(n1011), .Z(O[105]) );
  AND U1517 ( .A(S), .B(n1012), .Z(n1011) );
  XOR U1518 ( .A(B[105]), .B(B[104]), .Z(n1012) );
  XOR U1519 ( .A(B[103]), .B(n1013), .Z(O[104]) );
  AND U1520 ( .A(S), .B(n1014), .Z(n1013) );
  XOR U1521 ( .A(B[104]), .B(B[103]), .Z(n1014) );
  XOR U1522 ( .A(B[102]), .B(n1015), .Z(O[103]) );
  AND U1523 ( .A(S), .B(n1016), .Z(n1015) );
  XOR U1524 ( .A(B[103]), .B(B[102]), .Z(n1016) );
  XOR U1525 ( .A(B[101]), .B(n1017), .Z(O[102]) );
  AND U1526 ( .A(S), .B(n1018), .Z(n1017) );
  XOR U1527 ( .A(B[102]), .B(B[101]), .Z(n1018) );
  XOR U1528 ( .A(B[100]), .B(n1019), .Z(O[101]) );
  AND U1529 ( .A(S), .B(n1020), .Z(n1019) );
  XOR U1530 ( .A(B[101]), .B(B[100]), .Z(n1020) );
  XOR U1531 ( .A(B[99]), .B(n1021), .Z(O[100]) );
  AND U1532 ( .A(S), .B(n1022), .Z(n1021) );
  XOR U1533 ( .A(B[99]), .B(B[100]), .Z(n1022) );
  AND U1534 ( .A(B[0]), .B(S), .Z(O[0]) );
endmodule


module modexp_2N_NN_N512_CC262144 ( clk, rst, m, e, n, c );
  input [511:0] m;
  input [511:0] e;
  input [511:0] n;
  output [511:0] c;
  input clk, rst;
  wire   _0_net_, first_one, mul_pow, n6, n8, n265, n266, n267, n268;
  wire   [255:0] start_in;
  wire   [511:0] ein;
  wire   [511:0] creg_next;
  wire   [511:0] o;
  wire   [511:0] ereg_next;
  wire   [511:0] y;

  MUX_N512_3 MUX_4 ( .A(o), .B(c), .S(_0_net_), .O(creg_next) );
  MUX_N512_5 MUX_6 ( .A({ein[510:0], 1'b0}), .B(ein), .S(mul_pow), .O(
        ereg_next) );
  MUX_N512_4 MUX_9 ( .A(m), .B(c), .S(mul_pow), .O(y) );
  modmult_N512_CC256 modmult_1 ( .clk(clk), .rst(1'b0), .start(start_in[0]), 
        .x(c), .y(y), .n(n), .o(o) );
  DFF \start_reg_reg[0]  ( .D(start_in[255]), .CLK(clk), .RST(rst), .I(1'b1), 
        .Q(start_in[0]) );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[63]) );
  DFF \start_reg_reg[64]  ( .D(start_in[63]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[64]) );
  DFF \start_reg_reg[65]  ( .D(start_in[64]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[65]) );
  DFF \start_reg_reg[66]  ( .D(start_in[65]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[66]) );
  DFF \start_reg_reg[67]  ( .D(start_in[66]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[67]) );
  DFF \start_reg_reg[68]  ( .D(start_in[67]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[68]) );
  DFF \start_reg_reg[69]  ( .D(start_in[68]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[69]) );
  DFF \start_reg_reg[70]  ( .D(start_in[69]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[70]) );
  DFF \start_reg_reg[71]  ( .D(start_in[70]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[71]) );
  DFF \start_reg_reg[72]  ( .D(start_in[71]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[72]) );
  DFF \start_reg_reg[73]  ( .D(start_in[72]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[73]) );
  DFF \start_reg_reg[74]  ( .D(start_in[73]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[74]) );
  DFF \start_reg_reg[75]  ( .D(start_in[74]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[75]) );
  DFF \start_reg_reg[76]  ( .D(start_in[75]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[76]) );
  DFF \start_reg_reg[77]  ( .D(start_in[76]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[77]) );
  DFF \start_reg_reg[78]  ( .D(start_in[77]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[78]) );
  DFF \start_reg_reg[79]  ( .D(start_in[78]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[79]) );
  DFF \start_reg_reg[80]  ( .D(start_in[79]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[80]) );
  DFF \start_reg_reg[81]  ( .D(start_in[80]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[81]) );
  DFF \start_reg_reg[82]  ( .D(start_in[81]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[82]) );
  DFF \start_reg_reg[83]  ( .D(start_in[82]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[83]) );
  DFF \start_reg_reg[84]  ( .D(start_in[83]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[84]) );
  DFF \start_reg_reg[85]  ( .D(start_in[84]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[85]) );
  DFF \start_reg_reg[86]  ( .D(start_in[85]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[86]) );
  DFF \start_reg_reg[87]  ( .D(start_in[86]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[87]) );
  DFF \start_reg_reg[88]  ( .D(start_in[87]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[88]) );
  DFF \start_reg_reg[89]  ( .D(start_in[88]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[89]) );
  DFF \start_reg_reg[90]  ( .D(start_in[89]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[90]) );
  DFF \start_reg_reg[91]  ( .D(start_in[90]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[91]) );
  DFF \start_reg_reg[92]  ( .D(start_in[91]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[92]) );
  DFF \start_reg_reg[93]  ( .D(start_in[92]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[93]) );
  DFF \start_reg_reg[94]  ( .D(start_in[93]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[94]) );
  DFF \start_reg_reg[95]  ( .D(start_in[94]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[95]) );
  DFF \start_reg_reg[96]  ( .D(start_in[95]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[96]) );
  DFF \start_reg_reg[97]  ( .D(start_in[96]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[97]) );
  DFF \start_reg_reg[98]  ( .D(start_in[97]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[98]) );
  DFF \start_reg_reg[99]  ( .D(start_in[98]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[99]) );
  DFF \start_reg_reg[100]  ( .D(start_in[99]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[100]) );
  DFF \start_reg_reg[101]  ( .D(start_in[100]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[101]) );
  DFF \start_reg_reg[102]  ( .D(start_in[101]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[102]) );
  DFF \start_reg_reg[103]  ( .D(start_in[102]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[103]) );
  DFF \start_reg_reg[104]  ( .D(start_in[103]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[104]) );
  DFF \start_reg_reg[105]  ( .D(start_in[104]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[105]) );
  DFF \start_reg_reg[106]  ( .D(start_in[105]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[106]) );
  DFF \start_reg_reg[107]  ( .D(start_in[106]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[107]) );
  DFF \start_reg_reg[108]  ( .D(start_in[107]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[108]) );
  DFF \start_reg_reg[109]  ( .D(start_in[108]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[109]) );
  DFF \start_reg_reg[110]  ( .D(start_in[109]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[110]) );
  DFF \start_reg_reg[111]  ( .D(start_in[110]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[111]) );
  DFF \start_reg_reg[112]  ( .D(start_in[111]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[112]) );
  DFF \start_reg_reg[113]  ( .D(start_in[112]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[113]) );
  DFF \start_reg_reg[114]  ( .D(start_in[113]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[114]) );
  DFF \start_reg_reg[115]  ( .D(start_in[114]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[115]) );
  DFF \start_reg_reg[116]  ( .D(start_in[115]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[116]) );
  DFF \start_reg_reg[117]  ( .D(start_in[116]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[117]) );
  DFF \start_reg_reg[118]  ( .D(start_in[117]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[118]) );
  DFF \start_reg_reg[119]  ( .D(start_in[118]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[119]) );
  DFF \start_reg_reg[120]  ( .D(start_in[119]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[120]) );
  DFF \start_reg_reg[121]  ( .D(start_in[120]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[121]) );
  DFF \start_reg_reg[122]  ( .D(start_in[121]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[122]) );
  DFF \start_reg_reg[123]  ( .D(start_in[122]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[123]) );
  DFF \start_reg_reg[124]  ( .D(start_in[123]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[124]) );
  DFF \start_reg_reg[125]  ( .D(start_in[124]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[125]) );
  DFF \start_reg_reg[126]  ( .D(start_in[125]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[126]) );
  DFF \start_reg_reg[127]  ( .D(start_in[126]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[127]) );
  DFF \start_reg_reg[128]  ( .D(start_in[127]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[128]) );
  DFF \start_reg_reg[129]  ( .D(start_in[128]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[129]) );
  DFF \start_reg_reg[130]  ( .D(start_in[129]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[130]) );
  DFF \start_reg_reg[131]  ( .D(start_in[130]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[131]) );
  DFF \start_reg_reg[132]  ( .D(start_in[131]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[132]) );
  DFF \start_reg_reg[133]  ( .D(start_in[132]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[133]) );
  DFF \start_reg_reg[134]  ( .D(start_in[133]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[134]) );
  DFF \start_reg_reg[135]  ( .D(start_in[134]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[135]) );
  DFF \start_reg_reg[136]  ( .D(start_in[135]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[136]) );
  DFF \start_reg_reg[137]  ( .D(start_in[136]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[137]) );
  DFF \start_reg_reg[138]  ( .D(start_in[137]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[138]) );
  DFF \start_reg_reg[139]  ( .D(start_in[138]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[139]) );
  DFF \start_reg_reg[140]  ( .D(start_in[139]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[140]) );
  DFF \start_reg_reg[141]  ( .D(start_in[140]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[141]) );
  DFF \start_reg_reg[142]  ( .D(start_in[141]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[142]) );
  DFF \start_reg_reg[143]  ( .D(start_in[142]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[143]) );
  DFF \start_reg_reg[144]  ( .D(start_in[143]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[144]) );
  DFF \start_reg_reg[145]  ( .D(start_in[144]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[145]) );
  DFF \start_reg_reg[146]  ( .D(start_in[145]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[146]) );
  DFF \start_reg_reg[147]  ( .D(start_in[146]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[147]) );
  DFF \start_reg_reg[148]  ( .D(start_in[147]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[148]) );
  DFF \start_reg_reg[149]  ( .D(start_in[148]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[149]) );
  DFF \start_reg_reg[150]  ( .D(start_in[149]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[150]) );
  DFF \start_reg_reg[151]  ( .D(start_in[150]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[151]) );
  DFF \start_reg_reg[152]  ( .D(start_in[151]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[152]) );
  DFF \start_reg_reg[153]  ( .D(start_in[152]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[153]) );
  DFF \start_reg_reg[154]  ( .D(start_in[153]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[154]) );
  DFF \start_reg_reg[155]  ( .D(start_in[154]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[155]) );
  DFF \start_reg_reg[156]  ( .D(start_in[155]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[156]) );
  DFF \start_reg_reg[157]  ( .D(start_in[156]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[157]) );
  DFF \start_reg_reg[158]  ( .D(start_in[157]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[158]) );
  DFF \start_reg_reg[159]  ( .D(start_in[158]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[159]) );
  DFF \start_reg_reg[160]  ( .D(start_in[159]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[160]) );
  DFF \start_reg_reg[161]  ( .D(start_in[160]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[161]) );
  DFF \start_reg_reg[162]  ( .D(start_in[161]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[162]) );
  DFF \start_reg_reg[163]  ( .D(start_in[162]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[163]) );
  DFF \start_reg_reg[164]  ( .D(start_in[163]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[164]) );
  DFF \start_reg_reg[165]  ( .D(start_in[164]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[165]) );
  DFF \start_reg_reg[166]  ( .D(start_in[165]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[166]) );
  DFF \start_reg_reg[167]  ( .D(start_in[166]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[167]) );
  DFF \start_reg_reg[168]  ( .D(start_in[167]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[168]) );
  DFF \start_reg_reg[169]  ( .D(start_in[168]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[169]) );
  DFF \start_reg_reg[170]  ( .D(start_in[169]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[170]) );
  DFF \start_reg_reg[171]  ( .D(start_in[170]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[171]) );
  DFF \start_reg_reg[172]  ( .D(start_in[171]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[172]) );
  DFF \start_reg_reg[173]  ( .D(start_in[172]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[173]) );
  DFF \start_reg_reg[174]  ( .D(start_in[173]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[174]) );
  DFF \start_reg_reg[175]  ( .D(start_in[174]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[175]) );
  DFF \start_reg_reg[176]  ( .D(start_in[175]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[176]) );
  DFF \start_reg_reg[177]  ( .D(start_in[176]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[177]) );
  DFF \start_reg_reg[178]  ( .D(start_in[177]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[178]) );
  DFF \start_reg_reg[179]  ( .D(start_in[178]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[179]) );
  DFF \start_reg_reg[180]  ( .D(start_in[179]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[180]) );
  DFF \start_reg_reg[181]  ( .D(start_in[180]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[181]) );
  DFF \start_reg_reg[182]  ( .D(start_in[181]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[182]) );
  DFF \start_reg_reg[183]  ( .D(start_in[182]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[183]) );
  DFF \start_reg_reg[184]  ( .D(start_in[183]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[184]) );
  DFF \start_reg_reg[185]  ( .D(start_in[184]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[185]) );
  DFF \start_reg_reg[186]  ( .D(start_in[185]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[186]) );
  DFF \start_reg_reg[187]  ( .D(start_in[186]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[187]) );
  DFF \start_reg_reg[188]  ( .D(start_in[187]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[188]) );
  DFF \start_reg_reg[189]  ( .D(start_in[188]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[189]) );
  DFF \start_reg_reg[190]  ( .D(start_in[189]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[190]) );
  DFF \start_reg_reg[191]  ( .D(start_in[190]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[191]) );
  DFF \start_reg_reg[192]  ( .D(start_in[191]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[192]) );
  DFF \start_reg_reg[193]  ( .D(start_in[192]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[193]) );
  DFF \start_reg_reg[194]  ( .D(start_in[193]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[194]) );
  DFF \start_reg_reg[195]  ( .D(start_in[194]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[195]) );
  DFF \start_reg_reg[196]  ( .D(start_in[195]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[196]) );
  DFF \start_reg_reg[197]  ( .D(start_in[196]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[197]) );
  DFF \start_reg_reg[198]  ( .D(start_in[197]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[198]) );
  DFF \start_reg_reg[199]  ( .D(start_in[198]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[199]) );
  DFF \start_reg_reg[200]  ( .D(start_in[199]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[200]) );
  DFF \start_reg_reg[201]  ( .D(start_in[200]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[201]) );
  DFF \start_reg_reg[202]  ( .D(start_in[201]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[202]) );
  DFF \start_reg_reg[203]  ( .D(start_in[202]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[203]) );
  DFF \start_reg_reg[204]  ( .D(start_in[203]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[204]) );
  DFF \start_reg_reg[205]  ( .D(start_in[204]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[205]) );
  DFF \start_reg_reg[206]  ( .D(start_in[205]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[206]) );
  DFF \start_reg_reg[207]  ( .D(start_in[206]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[207]) );
  DFF \start_reg_reg[208]  ( .D(start_in[207]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[208]) );
  DFF \start_reg_reg[209]  ( .D(start_in[208]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[209]) );
  DFF \start_reg_reg[210]  ( .D(start_in[209]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[210]) );
  DFF \start_reg_reg[211]  ( .D(start_in[210]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[211]) );
  DFF \start_reg_reg[212]  ( .D(start_in[211]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[212]) );
  DFF \start_reg_reg[213]  ( .D(start_in[212]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[213]) );
  DFF \start_reg_reg[214]  ( .D(start_in[213]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[214]) );
  DFF \start_reg_reg[215]  ( .D(start_in[214]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[215]) );
  DFF \start_reg_reg[216]  ( .D(start_in[215]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[216]) );
  DFF \start_reg_reg[217]  ( .D(start_in[216]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[217]) );
  DFF \start_reg_reg[218]  ( .D(start_in[217]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[218]) );
  DFF \start_reg_reg[219]  ( .D(start_in[218]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[219]) );
  DFF \start_reg_reg[220]  ( .D(start_in[219]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[220]) );
  DFF \start_reg_reg[221]  ( .D(start_in[220]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[221]) );
  DFF \start_reg_reg[222]  ( .D(start_in[221]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[222]) );
  DFF \start_reg_reg[223]  ( .D(start_in[222]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[223]) );
  DFF \start_reg_reg[224]  ( .D(start_in[223]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[224]) );
  DFF \start_reg_reg[225]  ( .D(start_in[224]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[225]) );
  DFF \start_reg_reg[226]  ( .D(start_in[225]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[226]) );
  DFF \start_reg_reg[227]  ( .D(start_in[226]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[227]) );
  DFF \start_reg_reg[228]  ( .D(start_in[227]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[228]) );
  DFF \start_reg_reg[229]  ( .D(start_in[228]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[229]) );
  DFF \start_reg_reg[230]  ( .D(start_in[229]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[230]) );
  DFF \start_reg_reg[231]  ( .D(start_in[230]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[231]) );
  DFF \start_reg_reg[232]  ( .D(start_in[231]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[232]) );
  DFF \start_reg_reg[233]  ( .D(start_in[232]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[233]) );
  DFF \start_reg_reg[234]  ( .D(start_in[233]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[234]) );
  DFF \start_reg_reg[235]  ( .D(start_in[234]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[235]) );
  DFF \start_reg_reg[236]  ( .D(start_in[235]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[236]) );
  DFF \start_reg_reg[237]  ( .D(start_in[236]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[237]) );
  DFF \start_reg_reg[238]  ( .D(start_in[237]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[238]) );
  DFF \start_reg_reg[239]  ( .D(start_in[238]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[239]) );
  DFF \start_reg_reg[240]  ( .D(start_in[239]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[240]) );
  DFF \start_reg_reg[241]  ( .D(start_in[240]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[241]) );
  DFF \start_reg_reg[242]  ( .D(start_in[241]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[242]) );
  DFF \start_reg_reg[243]  ( .D(start_in[242]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[243]) );
  DFF \start_reg_reg[244]  ( .D(start_in[243]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[244]) );
  DFF \start_reg_reg[245]  ( .D(start_in[244]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[245]) );
  DFF \start_reg_reg[246]  ( .D(start_in[245]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[246]) );
  DFF \start_reg_reg[247]  ( .D(start_in[246]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[247]) );
  DFF \start_reg_reg[248]  ( .D(start_in[247]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[248]) );
  DFF \start_reg_reg[249]  ( .D(start_in[248]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[249]) );
  DFF \start_reg_reg[250]  ( .D(start_in[249]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[250]) );
  DFF \start_reg_reg[251]  ( .D(start_in[250]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[251]) );
  DFF \start_reg_reg[252]  ( .D(start_in[251]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[252]) );
  DFF \start_reg_reg[253]  ( .D(start_in[252]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[253]) );
  DFF \start_reg_reg[254]  ( .D(start_in[253]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[254]) );
  DFF \start_reg_reg[255]  ( .D(start_in[254]), .CLK(clk), .RST(rst), .I(1'b0), 
        .Q(start_in[255]) );
  DFF mul_pow_reg ( .D(n8), .CLK(clk), .RST(rst), .I(1'b0), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(ereg_next[0]), .CLK(clk), .RST(rst), .I(e[0]), .Q(
        ein[0]) );
  DFF \ereg_reg[1]  ( .D(ereg_next[1]), .CLK(clk), .RST(rst), .I(e[1]), .Q(
        ein[1]) );
  DFF \ereg_reg[2]  ( .D(ereg_next[2]), .CLK(clk), .RST(rst), .I(e[2]), .Q(
        ein[2]) );
  DFF \ereg_reg[3]  ( .D(ereg_next[3]), .CLK(clk), .RST(rst), .I(e[3]), .Q(
        ein[3]) );
  DFF \ereg_reg[4]  ( .D(ereg_next[4]), .CLK(clk), .RST(rst), .I(e[4]), .Q(
        ein[4]) );
  DFF \ereg_reg[5]  ( .D(ereg_next[5]), .CLK(clk), .RST(rst), .I(e[5]), .Q(
        ein[5]) );
  DFF \ereg_reg[6]  ( .D(ereg_next[6]), .CLK(clk), .RST(rst), .I(e[6]), .Q(
        ein[6]) );
  DFF \ereg_reg[7]  ( .D(ereg_next[7]), .CLK(clk), .RST(rst), .I(e[7]), .Q(
        ein[7]) );
  DFF \ereg_reg[8]  ( .D(ereg_next[8]), .CLK(clk), .RST(rst), .I(e[8]), .Q(
        ein[8]) );
  DFF \ereg_reg[9]  ( .D(ereg_next[9]), .CLK(clk), .RST(rst), .I(e[9]), .Q(
        ein[9]) );
  DFF \ereg_reg[10]  ( .D(ereg_next[10]), .CLK(clk), .RST(rst), .I(e[10]), .Q(
        ein[10]) );
  DFF \ereg_reg[11]  ( .D(ereg_next[11]), .CLK(clk), .RST(rst), .I(e[11]), .Q(
        ein[11]) );
  DFF \ereg_reg[12]  ( .D(ereg_next[12]), .CLK(clk), .RST(rst), .I(e[12]), .Q(
        ein[12]) );
  DFF \ereg_reg[13]  ( .D(ereg_next[13]), .CLK(clk), .RST(rst), .I(e[13]), .Q(
        ein[13]) );
  DFF \ereg_reg[14]  ( .D(ereg_next[14]), .CLK(clk), .RST(rst), .I(e[14]), .Q(
        ein[14]) );
  DFF \ereg_reg[15]  ( .D(ereg_next[15]), .CLK(clk), .RST(rst), .I(e[15]), .Q(
        ein[15]) );
  DFF \ereg_reg[16]  ( .D(ereg_next[16]), .CLK(clk), .RST(rst), .I(e[16]), .Q(
        ein[16]) );
  DFF \ereg_reg[17]  ( .D(ereg_next[17]), .CLK(clk), .RST(rst), .I(e[17]), .Q(
        ein[17]) );
  DFF \ereg_reg[18]  ( .D(ereg_next[18]), .CLK(clk), .RST(rst), .I(e[18]), .Q(
        ein[18]) );
  DFF \ereg_reg[19]  ( .D(ereg_next[19]), .CLK(clk), .RST(rst), .I(e[19]), .Q(
        ein[19]) );
  DFF \ereg_reg[20]  ( .D(ereg_next[20]), .CLK(clk), .RST(rst), .I(e[20]), .Q(
        ein[20]) );
  DFF \ereg_reg[21]  ( .D(ereg_next[21]), .CLK(clk), .RST(rst), .I(e[21]), .Q(
        ein[21]) );
  DFF \ereg_reg[22]  ( .D(ereg_next[22]), .CLK(clk), .RST(rst), .I(e[22]), .Q(
        ein[22]) );
  DFF \ereg_reg[23]  ( .D(ereg_next[23]), .CLK(clk), .RST(rst), .I(e[23]), .Q(
        ein[23]) );
  DFF \ereg_reg[24]  ( .D(ereg_next[24]), .CLK(clk), .RST(rst), .I(e[24]), .Q(
        ein[24]) );
  DFF \ereg_reg[25]  ( .D(ereg_next[25]), .CLK(clk), .RST(rst), .I(e[25]), .Q(
        ein[25]) );
  DFF \ereg_reg[26]  ( .D(ereg_next[26]), .CLK(clk), .RST(rst), .I(e[26]), .Q(
        ein[26]) );
  DFF \ereg_reg[27]  ( .D(ereg_next[27]), .CLK(clk), .RST(rst), .I(e[27]), .Q(
        ein[27]) );
  DFF \ereg_reg[28]  ( .D(ereg_next[28]), .CLK(clk), .RST(rst), .I(e[28]), .Q(
        ein[28]) );
  DFF \ereg_reg[29]  ( .D(ereg_next[29]), .CLK(clk), .RST(rst), .I(e[29]), .Q(
        ein[29]) );
  DFF \ereg_reg[30]  ( .D(ereg_next[30]), .CLK(clk), .RST(rst), .I(e[30]), .Q(
        ein[30]) );
  DFF \ereg_reg[31]  ( .D(ereg_next[31]), .CLK(clk), .RST(rst), .I(e[31]), .Q(
        ein[31]) );
  DFF \ereg_reg[32]  ( .D(ereg_next[32]), .CLK(clk), .RST(rst), .I(e[32]), .Q(
        ein[32]) );
  DFF \ereg_reg[33]  ( .D(ereg_next[33]), .CLK(clk), .RST(rst), .I(e[33]), .Q(
        ein[33]) );
  DFF \ereg_reg[34]  ( .D(ereg_next[34]), .CLK(clk), .RST(rst), .I(e[34]), .Q(
        ein[34]) );
  DFF \ereg_reg[35]  ( .D(ereg_next[35]), .CLK(clk), .RST(rst), .I(e[35]), .Q(
        ein[35]) );
  DFF \ereg_reg[36]  ( .D(ereg_next[36]), .CLK(clk), .RST(rst), .I(e[36]), .Q(
        ein[36]) );
  DFF \ereg_reg[37]  ( .D(ereg_next[37]), .CLK(clk), .RST(rst), .I(e[37]), .Q(
        ein[37]) );
  DFF \ereg_reg[38]  ( .D(ereg_next[38]), .CLK(clk), .RST(rst), .I(e[38]), .Q(
        ein[38]) );
  DFF \ereg_reg[39]  ( .D(ereg_next[39]), .CLK(clk), .RST(rst), .I(e[39]), .Q(
        ein[39]) );
  DFF \ereg_reg[40]  ( .D(ereg_next[40]), .CLK(clk), .RST(rst), .I(e[40]), .Q(
        ein[40]) );
  DFF \ereg_reg[41]  ( .D(ereg_next[41]), .CLK(clk), .RST(rst), .I(e[41]), .Q(
        ein[41]) );
  DFF \ereg_reg[42]  ( .D(ereg_next[42]), .CLK(clk), .RST(rst), .I(e[42]), .Q(
        ein[42]) );
  DFF \ereg_reg[43]  ( .D(ereg_next[43]), .CLK(clk), .RST(rst), .I(e[43]), .Q(
        ein[43]) );
  DFF \ereg_reg[44]  ( .D(ereg_next[44]), .CLK(clk), .RST(rst), .I(e[44]), .Q(
        ein[44]) );
  DFF \ereg_reg[45]  ( .D(ereg_next[45]), .CLK(clk), .RST(rst), .I(e[45]), .Q(
        ein[45]) );
  DFF \ereg_reg[46]  ( .D(ereg_next[46]), .CLK(clk), .RST(rst), .I(e[46]), .Q(
        ein[46]) );
  DFF \ereg_reg[47]  ( .D(ereg_next[47]), .CLK(clk), .RST(rst), .I(e[47]), .Q(
        ein[47]) );
  DFF \ereg_reg[48]  ( .D(ereg_next[48]), .CLK(clk), .RST(rst), .I(e[48]), .Q(
        ein[48]) );
  DFF \ereg_reg[49]  ( .D(ereg_next[49]), .CLK(clk), .RST(rst), .I(e[49]), .Q(
        ein[49]) );
  DFF \ereg_reg[50]  ( .D(ereg_next[50]), .CLK(clk), .RST(rst), .I(e[50]), .Q(
        ein[50]) );
  DFF \ereg_reg[51]  ( .D(ereg_next[51]), .CLK(clk), .RST(rst), .I(e[51]), .Q(
        ein[51]) );
  DFF \ereg_reg[52]  ( .D(ereg_next[52]), .CLK(clk), .RST(rst), .I(e[52]), .Q(
        ein[52]) );
  DFF \ereg_reg[53]  ( .D(ereg_next[53]), .CLK(clk), .RST(rst), .I(e[53]), .Q(
        ein[53]) );
  DFF \ereg_reg[54]  ( .D(ereg_next[54]), .CLK(clk), .RST(rst), .I(e[54]), .Q(
        ein[54]) );
  DFF \ereg_reg[55]  ( .D(ereg_next[55]), .CLK(clk), .RST(rst), .I(e[55]), .Q(
        ein[55]) );
  DFF \ereg_reg[56]  ( .D(ereg_next[56]), .CLK(clk), .RST(rst), .I(e[56]), .Q(
        ein[56]) );
  DFF \ereg_reg[57]  ( .D(ereg_next[57]), .CLK(clk), .RST(rst), .I(e[57]), .Q(
        ein[57]) );
  DFF \ereg_reg[58]  ( .D(ereg_next[58]), .CLK(clk), .RST(rst), .I(e[58]), .Q(
        ein[58]) );
  DFF \ereg_reg[59]  ( .D(ereg_next[59]), .CLK(clk), .RST(rst), .I(e[59]), .Q(
        ein[59]) );
  DFF \ereg_reg[60]  ( .D(ereg_next[60]), .CLK(clk), .RST(rst), .I(e[60]), .Q(
        ein[60]) );
  DFF \ereg_reg[61]  ( .D(ereg_next[61]), .CLK(clk), .RST(rst), .I(e[61]), .Q(
        ein[61]) );
  DFF \ereg_reg[62]  ( .D(ereg_next[62]), .CLK(clk), .RST(rst), .I(e[62]), .Q(
        ein[62]) );
  DFF \ereg_reg[63]  ( .D(ereg_next[63]), .CLK(clk), .RST(rst), .I(e[63]), .Q(
        ein[63]) );
  DFF \ereg_reg[64]  ( .D(ereg_next[64]), .CLK(clk), .RST(rst), .I(e[64]), .Q(
        ein[64]) );
  DFF \ereg_reg[65]  ( .D(ereg_next[65]), .CLK(clk), .RST(rst), .I(e[65]), .Q(
        ein[65]) );
  DFF \ereg_reg[66]  ( .D(ereg_next[66]), .CLK(clk), .RST(rst), .I(e[66]), .Q(
        ein[66]) );
  DFF \ereg_reg[67]  ( .D(ereg_next[67]), .CLK(clk), .RST(rst), .I(e[67]), .Q(
        ein[67]) );
  DFF \ereg_reg[68]  ( .D(ereg_next[68]), .CLK(clk), .RST(rst), .I(e[68]), .Q(
        ein[68]) );
  DFF \ereg_reg[69]  ( .D(ereg_next[69]), .CLK(clk), .RST(rst), .I(e[69]), .Q(
        ein[69]) );
  DFF \ereg_reg[70]  ( .D(ereg_next[70]), .CLK(clk), .RST(rst), .I(e[70]), .Q(
        ein[70]) );
  DFF \ereg_reg[71]  ( .D(ereg_next[71]), .CLK(clk), .RST(rst), .I(e[71]), .Q(
        ein[71]) );
  DFF \ereg_reg[72]  ( .D(ereg_next[72]), .CLK(clk), .RST(rst), .I(e[72]), .Q(
        ein[72]) );
  DFF \ereg_reg[73]  ( .D(ereg_next[73]), .CLK(clk), .RST(rst), .I(e[73]), .Q(
        ein[73]) );
  DFF \ereg_reg[74]  ( .D(ereg_next[74]), .CLK(clk), .RST(rst), .I(e[74]), .Q(
        ein[74]) );
  DFF \ereg_reg[75]  ( .D(ereg_next[75]), .CLK(clk), .RST(rst), .I(e[75]), .Q(
        ein[75]) );
  DFF \ereg_reg[76]  ( .D(ereg_next[76]), .CLK(clk), .RST(rst), .I(e[76]), .Q(
        ein[76]) );
  DFF \ereg_reg[77]  ( .D(ereg_next[77]), .CLK(clk), .RST(rst), .I(e[77]), .Q(
        ein[77]) );
  DFF \ereg_reg[78]  ( .D(ereg_next[78]), .CLK(clk), .RST(rst), .I(e[78]), .Q(
        ein[78]) );
  DFF \ereg_reg[79]  ( .D(ereg_next[79]), .CLK(clk), .RST(rst), .I(e[79]), .Q(
        ein[79]) );
  DFF \ereg_reg[80]  ( .D(ereg_next[80]), .CLK(clk), .RST(rst), .I(e[80]), .Q(
        ein[80]) );
  DFF \ereg_reg[81]  ( .D(ereg_next[81]), .CLK(clk), .RST(rst), .I(e[81]), .Q(
        ein[81]) );
  DFF \ereg_reg[82]  ( .D(ereg_next[82]), .CLK(clk), .RST(rst), .I(e[82]), .Q(
        ein[82]) );
  DFF \ereg_reg[83]  ( .D(ereg_next[83]), .CLK(clk), .RST(rst), .I(e[83]), .Q(
        ein[83]) );
  DFF \ereg_reg[84]  ( .D(ereg_next[84]), .CLK(clk), .RST(rst), .I(e[84]), .Q(
        ein[84]) );
  DFF \ereg_reg[85]  ( .D(ereg_next[85]), .CLK(clk), .RST(rst), .I(e[85]), .Q(
        ein[85]) );
  DFF \ereg_reg[86]  ( .D(ereg_next[86]), .CLK(clk), .RST(rst), .I(e[86]), .Q(
        ein[86]) );
  DFF \ereg_reg[87]  ( .D(ereg_next[87]), .CLK(clk), .RST(rst), .I(e[87]), .Q(
        ein[87]) );
  DFF \ereg_reg[88]  ( .D(ereg_next[88]), .CLK(clk), .RST(rst), .I(e[88]), .Q(
        ein[88]) );
  DFF \ereg_reg[89]  ( .D(ereg_next[89]), .CLK(clk), .RST(rst), .I(e[89]), .Q(
        ein[89]) );
  DFF \ereg_reg[90]  ( .D(ereg_next[90]), .CLK(clk), .RST(rst), .I(e[90]), .Q(
        ein[90]) );
  DFF \ereg_reg[91]  ( .D(ereg_next[91]), .CLK(clk), .RST(rst), .I(e[91]), .Q(
        ein[91]) );
  DFF \ereg_reg[92]  ( .D(ereg_next[92]), .CLK(clk), .RST(rst), .I(e[92]), .Q(
        ein[92]) );
  DFF \ereg_reg[93]  ( .D(ereg_next[93]), .CLK(clk), .RST(rst), .I(e[93]), .Q(
        ein[93]) );
  DFF \ereg_reg[94]  ( .D(ereg_next[94]), .CLK(clk), .RST(rst), .I(e[94]), .Q(
        ein[94]) );
  DFF \ereg_reg[95]  ( .D(ereg_next[95]), .CLK(clk), .RST(rst), .I(e[95]), .Q(
        ein[95]) );
  DFF \ereg_reg[96]  ( .D(ereg_next[96]), .CLK(clk), .RST(rst), .I(e[96]), .Q(
        ein[96]) );
  DFF \ereg_reg[97]  ( .D(ereg_next[97]), .CLK(clk), .RST(rst), .I(e[97]), .Q(
        ein[97]) );
  DFF \ereg_reg[98]  ( .D(ereg_next[98]), .CLK(clk), .RST(rst), .I(e[98]), .Q(
        ein[98]) );
  DFF \ereg_reg[99]  ( .D(ereg_next[99]), .CLK(clk), .RST(rst), .I(e[99]), .Q(
        ein[99]) );
  DFF \ereg_reg[100]  ( .D(ereg_next[100]), .CLK(clk), .RST(rst), .I(e[100]), 
        .Q(ein[100]) );
  DFF \ereg_reg[101]  ( .D(ereg_next[101]), .CLK(clk), .RST(rst), .I(e[101]), 
        .Q(ein[101]) );
  DFF \ereg_reg[102]  ( .D(ereg_next[102]), .CLK(clk), .RST(rst), .I(e[102]), 
        .Q(ein[102]) );
  DFF \ereg_reg[103]  ( .D(ereg_next[103]), .CLK(clk), .RST(rst), .I(e[103]), 
        .Q(ein[103]) );
  DFF \ereg_reg[104]  ( .D(ereg_next[104]), .CLK(clk), .RST(rst), .I(e[104]), 
        .Q(ein[104]) );
  DFF \ereg_reg[105]  ( .D(ereg_next[105]), .CLK(clk), .RST(rst), .I(e[105]), 
        .Q(ein[105]) );
  DFF \ereg_reg[106]  ( .D(ereg_next[106]), .CLK(clk), .RST(rst), .I(e[106]), 
        .Q(ein[106]) );
  DFF \ereg_reg[107]  ( .D(ereg_next[107]), .CLK(clk), .RST(rst), .I(e[107]), 
        .Q(ein[107]) );
  DFF \ereg_reg[108]  ( .D(ereg_next[108]), .CLK(clk), .RST(rst), .I(e[108]), 
        .Q(ein[108]) );
  DFF \ereg_reg[109]  ( .D(ereg_next[109]), .CLK(clk), .RST(rst), .I(e[109]), 
        .Q(ein[109]) );
  DFF \ereg_reg[110]  ( .D(ereg_next[110]), .CLK(clk), .RST(rst), .I(e[110]), 
        .Q(ein[110]) );
  DFF \ereg_reg[111]  ( .D(ereg_next[111]), .CLK(clk), .RST(rst), .I(e[111]), 
        .Q(ein[111]) );
  DFF \ereg_reg[112]  ( .D(ereg_next[112]), .CLK(clk), .RST(rst), .I(e[112]), 
        .Q(ein[112]) );
  DFF \ereg_reg[113]  ( .D(ereg_next[113]), .CLK(clk), .RST(rst), .I(e[113]), 
        .Q(ein[113]) );
  DFF \ereg_reg[114]  ( .D(ereg_next[114]), .CLK(clk), .RST(rst), .I(e[114]), 
        .Q(ein[114]) );
  DFF \ereg_reg[115]  ( .D(ereg_next[115]), .CLK(clk), .RST(rst), .I(e[115]), 
        .Q(ein[115]) );
  DFF \ereg_reg[116]  ( .D(ereg_next[116]), .CLK(clk), .RST(rst), .I(e[116]), 
        .Q(ein[116]) );
  DFF \ereg_reg[117]  ( .D(ereg_next[117]), .CLK(clk), .RST(rst), .I(e[117]), 
        .Q(ein[117]) );
  DFF \ereg_reg[118]  ( .D(ereg_next[118]), .CLK(clk), .RST(rst), .I(e[118]), 
        .Q(ein[118]) );
  DFF \ereg_reg[119]  ( .D(ereg_next[119]), .CLK(clk), .RST(rst), .I(e[119]), 
        .Q(ein[119]) );
  DFF \ereg_reg[120]  ( .D(ereg_next[120]), .CLK(clk), .RST(rst), .I(e[120]), 
        .Q(ein[120]) );
  DFF \ereg_reg[121]  ( .D(ereg_next[121]), .CLK(clk), .RST(rst), .I(e[121]), 
        .Q(ein[121]) );
  DFF \ereg_reg[122]  ( .D(ereg_next[122]), .CLK(clk), .RST(rst), .I(e[122]), 
        .Q(ein[122]) );
  DFF \ereg_reg[123]  ( .D(ereg_next[123]), .CLK(clk), .RST(rst), .I(e[123]), 
        .Q(ein[123]) );
  DFF \ereg_reg[124]  ( .D(ereg_next[124]), .CLK(clk), .RST(rst), .I(e[124]), 
        .Q(ein[124]) );
  DFF \ereg_reg[125]  ( .D(ereg_next[125]), .CLK(clk), .RST(rst), .I(e[125]), 
        .Q(ein[125]) );
  DFF \ereg_reg[126]  ( .D(ereg_next[126]), .CLK(clk), .RST(rst), .I(e[126]), 
        .Q(ein[126]) );
  DFF \ereg_reg[127]  ( .D(ereg_next[127]), .CLK(clk), .RST(rst), .I(e[127]), 
        .Q(ein[127]) );
  DFF \ereg_reg[128]  ( .D(ereg_next[128]), .CLK(clk), .RST(rst), .I(e[128]), 
        .Q(ein[128]) );
  DFF \ereg_reg[129]  ( .D(ereg_next[129]), .CLK(clk), .RST(rst), .I(e[129]), 
        .Q(ein[129]) );
  DFF \ereg_reg[130]  ( .D(ereg_next[130]), .CLK(clk), .RST(rst), .I(e[130]), 
        .Q(ein[130]) );
  DFF \ereg_reg[131]  ( .D(ereg_next[131]), .CLK(clk), .RST(rst), .I(e[131]), 
        .Q(ein[131]) );
  DFF \ereg_reg[132]  ( .D(ereg_next[132]), .CLK(clk), .RST(rst), .I(e[132]), 
        .Q(ein[132]) );
  DFF \ereg_reg[133]  ( .D(ereg_next[133]), .CLK(clk), .RST(rst), .I(e[133]), 
        .Q(ein[133]) );
  DFF \ereg_reg[134]  ( .D(ereg_next[134]), .CLK(clk), .RST(rst), .I(e[134]), 
        .Q(ein[134]) );
  DFF \ereg_reg[135]  ( .D(ereg_next[135]), .CLK(clk), .RST(rst), .I(e[135]), 
        .Q(ein[135]) );
  DFF \ereg_reg[136]  ( .D(ereg_next[136]), .CLK(clk), .RST(rst), .I(e[136]), 
        .Q(ein[136]) );
  DFF \ereg_reg[137]  ( .D(ereg_next[137]), .CLK(clk), .RST(rst), .I(e[137]), 
        .Q(ein[137]) );
  DFF \ereg_reg[138]  ( .D(ereg_next[138]), .CLK(clk), .RST(rst), .I(e[138]), 
        .Q(ein[138]) );
  DFF \ereg_reg[139]  ( .D(ereg_next[139]), .CLK(clk), .RST(rst), .I(e[139]), 
        .Q(ein[139]) );
  DFF \ereg_reg[140]  ( .D(ereg_next[140]), .CLK(clk), .RST(rst), .I(e[140]), 
        .Q(ein[140]) );
  DFF \ereg_reg[141]  ( .D(ereg_next[141]), .CLK(clk), .RST(rst), .I(e[141]), 
        .Q(ein[141]) );
  DFF \ereg_reg[142]  ( .D(ereg_next[142]), .CLK(clk), .RST(rst), .I(e[142]), 
        .Q(ein[142]) );
  DFF \ereg_reg[143]  ( .D(ereg_next[143]), .CLK(clk), .RST(rst), .I(e[143]), 
        .Q(ein[143]) );
  DFF \ereg_reg[144]  ( .D(ereg_next[144]), .CLK(clk), .RST(rst), .I(e[144]), 
        .Q(ein[144]) );
  DFF \ereg_reg[145]  ( .D(ereg_next[145]), .CLK(clk), .RST(rst), .I(e[145]), 
        .Q(ein[145]) );
  DFF \ereg_reg[146]  ( .D(ereg_next[146]), .CLK(clk), .RST(rst), .I(e[146]), 
        .Q(ein[146]) );
  DFF \ereg_reg[147]  ( .D(ereg_next[147]), .CLK(clk), .RST(rst), .I(e[147]), 
        .Q(ein[147]) );
  DFF \ereg_reg[148]  ( .D(ereg_next[148]), .CLK(clk), .RST(rst), .I(e[148]), 
        .Q(ein[148]) );
  DFF \ereg_reg[149]  ( .D(ereg_next[149]), .CLK(clk), .RST(rst), .I(e[149]), 
        .Q(ein[149]) );
  DFF \ereg_reg[150]  ( .D(ereg_next[150]), .CLK(clk), .RST(rst), .I(e[150]), 
        .Q(ein[150]) );
  DFF \ereg_reg[151]  ( .D(ereg_next[151]), .CLK(clk), .RST(rst), .I(e[151]), 
        .Q(ein[151]) );
  DFF \ereg_reg[152]  ( .D(ereg_next[152]), .CLK(clk), .RST(rst), .I(e[152]), 
        .Q(ein[152]) );
  DFF \ereg_reg[153]  ( .D(ereg_next[153]), .CLK(clk), .RST(rst), .I(e[153]), 
        .Q(ein[153]) );
  DFF \ereg_reg[154]  ( .D(ereg_next[154]), .CLK(clk), .RST(rst), .I(e[154]), 
        .Q(ein[154]) );
  DFF \ereg_reg[155]  ( .D(ereg_next[155]), .CLK(clk), .RST(rst), .I(e[155]), 
        .Q(ein[155]) );
  DFF \ereg_reg[156]  ( .D(ereg_next[156]), .CLK(clk), .RST(rst), .I(e[156]), 
        .Q(ein[156]) );
  DFF \ereg_reg[157]  ( .D(ereg_next[157]), .CLK(clk), .RST(rst), .I(e[157]), 
        .Q(ein[157]) );
  DFF \ereg_reg[158]  ( .D(ereg_next[158]), .CLK(clk), .RST(rst), .I(e[158]), 
        .Q(ein[158]) );
  DFF \ereg_reg[159]  ( .D(ereg_next[159]), .CLK(clk), .RST(rst), .I(e[159]), 
        .Q(ein[159]) );
  DFF \ereg_reg[160]  ( .D(ereg_next[160]), .CLK(clk), .RST(rst), .I(e[160]), 
        .Q(ein[160]) );
  DFF \ereg_reg[161]  ( .D(ereg_next[161]), .CLK(clk), .RST(rst), .I(e[161]), 
        .Q(ein[161]) );
  DFF \ereg_reg[162]  ( .D(ereg_next[162]), .CLK(clk), .RST(rst), .I(e[162]), 
        .Q(ein[162]) );
  DFF \ereg_reg[163]  ( .D(ereg_next[163]), .CLK(clk), .RST(rst), .I(e[163]), 
        .Q(ein[163]) );
  DFF \ereg_reg[164]  ( .D(ereg_next[164]), .CLK(clk), .RST(rst), .I(e[164]), 
        .Q(ein[164]) );
  DFF \ereg_reg[165]  ( .D(ereg_next[165]), .CLK(clk), .RST(rst), .I(e[165]), 
        .Q(ein[165]) );
  DFF \ereg_reg[166]  ( .D(ereg_next[166]), .CLK(clk), .RST(rst), .I(e[166]), 
        .Q(ein[166]) );
  DFF \ereg_reg[167]  ( .D(ereg_next[167]), .CLK(clk), .RST(rst), .I(e[167]), 
        .Q(ein[167]) );
  DFF \ereg_reg[168]  ( .D(ereg_next[168]), .CLK(clk), .RST(rst), .I(e[168]), 
        .Q(ein[168]) );
  DFF \ereg_reg[169]  ( .D(ereg_next[169]), .CLK(clk), .RST(rst), .I(e[169]), 
        .Q(ein[169]) );
  DFF \ereg_reg[170]  ( .D(ereg_next[170]), .CLK(clk), .RST(rst), .I(e[170]), 
        .Q(ein[170]) );
  DFF \ereg_reg[171]  ( .D(ereg_next[171]), .CLK(clk), .RST(rst), .I(e[171]), 
        .Q(ein[171]) );
  DFF \ereg_reg[172]  ( .D(ereg_next[172]), .CLK(clk), .RST(rst), .I(e[172]), 
        .Q(ein[172]) );
  DFF \ereg_reg[173]  ( .D(ereg_next[173]), .CLK(clk), .RST(rst), .I(e[173]), 
        .Q(ein[173]) );
  DFF \ereg_reg[174]  ( .D(ereg_next[174]), .CLK(clk), .RST(rst), .I(e[174]), 
        .Q(ein[174]) );
  DFF \ereg_reg[175]  ( .D(ereg_next[175]), .CLK(clk), .RST(rst), .I(e[175]), 
        .Q(ein[175]) );
  DFF \ereg_reg[176]  ( .D(ereg_next[176]), .CLK(clk), .RST(rst), .I(e[176]), 
        .Q(ein[176]) );
  DFF \ereg_reg[177]  ( .D(ereg_next[177]), .CLK(clk), .RST(rst), .I(e[177]), 
        .Q(ein[177]) );
  DFF \ereg_reg[178]  ( .D(ereg_next[178]), .CLK(clk), .RST(rst), .I(e[178]), 
        .Q(ein[178]) );
  DFF \ereg_reg[179]  ( .D(ereg_next[179]), .CLK(clk), .RST(rst), .I(e[179]), 
        .Q(ein[179]) );
  DFF \ereg_reg[180]  ( .D(ereg_next[180]), .CLK(clk), .RST(rst), .I(e[180]), 
        .Q(ein[180]) );
  DFF \ereg_reg[181]  ( .D(ereg_next[181]), .CLK(clk), .RST(rst), .I(e[181]), 
        .Q(ein[181]) );
  DFF \ereg_reg[182]  ( .D(ereg_next[182]), .CLK(clk), .RST(rst), .I(e[182]), 
        .Q(ein[182]) );
  DFF \ereg_reg[183]  ( .D(ereg_next[183]), .CLK(clk), .RST(rst), .I(e[183]), 
        .Q(ein[183]) );
  DFF \ereg_reg[184]  ( .D(ereg_next[184]), .CLK(clk), .RST(rst), .I(e[184]), 
        .Q(ein[184]) );
  DFF \ereg_reg[185]  ( .D(ereg_next[185]), .CLK(clk), .RST(rst), .I(e[185]), 
        .Q(ein[185]) );
  DFF \ereg_reg[186]  ( .D(ereg_next[186]), .CLK(clk), .RST(rst), .I(e[186]), 
        .Q(ein[186]) );
  DFF \ereg_reg[187]  ( .D(ereg_next[187]), .CLK(clk), .RST(rst), .I(e[187]), 
        .Q(ein[187]) );
  DFF \ereg_reg[188]  ( .D(ereg_next[188]), .CLK(clk), .RST(rst), .I(e[188]), 
        .Q(ein[188]) );
  DFF \ereg_reg[189]  ( .D(ereg_next[189]), .CLK(clk), .RST(rst), .I(e[189]), 
        .Q(ein[189]) );
  DFF \ereg_reg[190]  ( .D(ereg_next[190]), .CLK(clk), .RST(rst), .I(e[190]), 
        .Q(ein[190]) );
  DFF \ereg_reg[191]  ( .D(ereg_next[191]), .CLK(clk), .RST(rst), .I(e[191]), 
        .Q(ein[191]) );
  DFF \ereg_reg[192]  ( .D(ereg_next[192]), .CLK(clk), .RST(rst), .I(e[192]), 
        .Q(ein[192]) );
  DFF \ereg_reg[193]  ( .D(ereg_next[193]), .CLK(clk), .RST(rst), .I(e[193]), 
        .Q(ein[193]) );
  DFF \ereg_reg[194]  ( .D(ereg_next[194]), .CLK(clk), .RST(rst), .I(e[194]), 
        .Q(ein[194]) );
  DFF \ereg_reg[195]  ( .D(ereg_next[195]), .CLK(clk), .RST(rst), .I(e[195]), 
        .Q(ein[195]) );
  DFF \ereg_reg[196]  ( .D(ereg_next[196]), .CLK(clk), .RST(rst), .I(e[196]), 
        .Q(ein[196]) );
  DFF \ereg_reg[197]  ( .D(ereg_next[197]), .CLK(clk), .RST(rst), .I(e[197]), 
        .Q(ein[197]) );
  DFF \ereg_reg[198]  ( .D(ereg_next[198]), .CLK(clk), .RST(rst), .I(e[198]), 
        .Q(ein[198]) );
  DFF \ereg_reg[199]  ( .D(ereg_next[199]), .CLK(clk), .RST(rst), .I(e[199]), 
        .Q(ein[199]) );
  DFF \ereg_reg[200]  ( .D(ereg_next[200]), .CLK(clk), .RST(rst), .I(e[200]), 
        .Q(ein[200]) );
  DFF \ereg_reg[201]  ( .D(ereg_next[201]), .CLK(clk), .RST(rst), .I(e[201]), 
        .Q(ein[201]) );
  DFF \ereg_reg[202]  ( .D(ereg_next[202]), .CLK(clk), .RST(rst), .I(e[202]), 
        .Q(ein[202]) );
  DFF \ereg_reg[203]  ( .D(ereg_next[203]), .CLK(clk), .RST(rst), .I(e[203]), 
        .Q(ein[203]) );
  DFF \ereg_reg[204]  ( .D(ereg_next[204]), .CLK(clk), .RST(rst), .I(e[204]), 
        .Q(ein[204]) );
  DFF \ereg_reg[205]  ( .D(ereg_next[205]), .CLK(clk), .RST(rst), .I(e[205]), 
        .Q(ein[205]) );
  DFF \ereg_reg[206]  ( .D(ereg_next[206]), .CLK(clk), .RST(rst), .I(e[206]), 
        .Q(ein[206]) );
  DFF \ereg_reg[207]  ( .D(ereg_next[207]), .CLK(clk), .RST(rst), .I(e[207]), 
        .Q(ein[207]) );
  DFF \ereg_reg[208]  ( .D(ereg_next[208]), .CLK(clk), .RST(rst), .I(e[208]), 
        .Q(ein[208]) );
  DFF \ereg_reg[209]  ( .D(ereg_next[209]), .CLK(clk), .RST(rst), .I(e[209]), 
        .Q(ein[209]) );
  DFF \ereg_reg[210]  ( .D(ereg_next[210]), .CLK(clk), .RST(rst), .I(e[210]), 
        .Q(ein[210]) );
  DFF \ereg_reg[211]  ( .D(ereg_next[211]), .CLK(clk), .RST(rst), .I(e[211]), 
        .Q(ein[211]) );
  DFF \ereg_reg[212]  ( .D(ereg_next[212]), .CLK(clk), .RST(rst), .I(e[212]), 
        .Q(ein[212]) );
  DFF \ereg_reg[213]  ( .D(ereg_next[213]), .CLK(clk), .RST(rst), .I(e[213]), 
        .Q(ein[213]) );
  DFF \ereg_reg[214]  ( .D(ereg_next[214]), .CLK(clk), .RST(rst), .I(e[214]), 
        .Q(ein[214]) );
  DFF \ereg_reg[215]  ( .D(ereg_next[215]), .CLK(clk), .RST(rst), .I(e[215]), 
        .Q(ein[215]) );
  DFF \ereg_reg[216]  ( .D(ereg_next[216]), .CLK(clk), .RST(rst), .I(e[216]), 
        .Q(ein[216]) );
  DFF \ereg_reg[217]  ( .D(ereg_next[217]), .CLK(clk), .RST(rst), .I(e[217]), 
        .Q(ein[217]) );
  DFF \ereg_reg[218]  ( .D(ereg_next[218]), .CLK(clk), .RST(rst), .I(e[218]), 
        .Q(ein[218]) );
  DFF \ereg_reg[219]  ( .D(ereg_next[219]), .CLK(clk), .RST(rst), .I(e[219]), 
        .Q(ein[219]) );
  DFF \ereg_reg[220]  ( .D(ereg_next[220]), .CLK(clk), .RST(rst), .I(e[220]), 
        .Q(ein[220]) );
  DFF \ereg_reg[221]  ( .D(ereg_next[221]), .CLK(clk), .RST(rst), .I(e[221]), 
        .Q(ein[221]) );
  DFF \ereg_reg[222]  ( .D(ereg_next[222]), .CLK(clk), .RST(rst), .I(e[222]), 
        .Q(ein[222]) );
  DFF \ereg_reg[223]  ( .D(ereg_next[223]), .CLK(clk), .RST(rst), .I(e[223]), 
        .Q(ein[223]) );
  DFF \ereg_reg[224]  ( .D(ereg_next[224]), .CLK(clk), .RST(rst), .I(e[224]), 
        .Q(ein[224]) );
  DFF \ereg_reg[225]  ( .D(ereg_next[225]), .CLK(clk), .RST(rst), .I(e[225]), 
        .Q(ein[225]) );
  DFF \ereg_reg[226]  ( .D(ereg_next[226]), .CLK(clk), .RST(rst), .I(e[226]), 
        .Q(ein[226]) );
  DFF \ereg_reg[227]  ( .D(ereg_next[227]), .CLK(clk), .RST(rst), .I(e[227]), 
        .Q(ein[227]) );
  DFF \ereg_reg[228]  ( .D(ereg_next[228]), .CLK(clk), .RST(rst), .I(e[228]), 
        .Q(ein[228]) );
  DFF \ereg_reg[229]  ( .D(ereg_next[229]), .CLK(clk), .RST(rst), .I(e[229]), 
        .Q(ein[229]) );
  DFF \ereg_reg[230]  ( .D(ereg_next[230]), .CLK(clk), .RST(rst), .I(e[230]), 
        .Q(ein[230]) );
  DFF \ereg_reg[231]  ( .D(ereg_next[231]), .CLK(clk), .RST(rst), .I(e[231]), 
        .Q(ein[231]) );
  DFF \ereg_reg[232]  ( .D(ereg_next[232]), .CLK(clk), .RST(rst), .I(e[232]), 
        .Q(ein[232]) );
  DFF \ereg_reg[233]  ( .D(ereg_next[233]), .CLK(clk), .RST(rst), .I(e[233]), 
        .Q(ein[233]) );
  DFF \ereg_reg[234]  ( .D(ereg_next[234]), .CLK(clk), .RST(rst), .I(e[234]), 
        .Q(ein[234]) );
  DFF \ereg_reg[235]  ( .D(ereg_next[235]), .CLK(clk), .RST(rst), .I(e[235]), 
        .Q(ein[235]) );
  DFF \ereg_reg[236]  ( .D(ereg_next[236]), .CLK(clk), .RST(rst), .I(e[236]), 
        .Q(ein[236]) );
  DFF \ereg_reg[237]  ( .D(ereg_next[237]), .CLK(clk), .RST(rst), .I(e[237]), 
        .Q(ein[237]) );
  DFF \ereg_reg[238]  ( .D(ereg_next[238]), .CLK(clk), .RST(rst), .I(e[238]), 
        .Q(ein[238]) );
  DFF \ereg_reg[239]  ( .D(ereg_next[239]), .CLK(clk), .RST(rst), .I(e[239]), 
        .Q(ein[239]) );
  DFF \ereg_reg[240]  ( .D(ereg_next[240]), .CLK(clk), .RST(rst), .I(e[240]), 
        .Q(ein[240]) );
  DFF \ereg_reg[241]  ( .D(ereg_next[241]), .CLK(clk), .RST(rst), .I(e[241]), 
        .Q(ein[241]) );
  DFF \ereg_reg[242]  ( .D(ereg_next[242]), .CLK(clk), .RST(rst), .I(e[242]), 
        .Q(ein[242]) );
  DFF \ereg_reg[243]  ( .D(ereg_next[243]), .CLK(clk), .RST(rst), .I(e[243]), 
        .Q(ein[243]) );
  DFF \ereg_reg[244]  ( .D(ereg_next[244]), .CLK(clk), .RST(rst), .I(e[244]), 
        .Q(ein[244]) );
  DFF \ereg_reg[245]  ( .D(ereg_next[245]), .CLK(clk), .RST(rst), .I(e[245]), 
        .Q(ein[245]) );
  DFF \ereg_reg[246]  ( .D(ereg_next[246]), .CLK(clk), .RST(rst), .I(e[246]), 
        .Q(ein[246]) );
  DFF \ereg_reg[247]  ( .D(ereg_next[247]), .CLK(clk), .RST(rst), .I(e[247]), 
        .Q(ein[247]) );
  DFF \ereg_reg[248]  ( .D(ereg_next[248]), .CLK(clk), .RST(rst), .I(e[248]), 
        .Q(ein[248]) );
  DFF \ereg_reg[249]  ( .D(ereg_next[249]), .CLK(clk), .RST(rst), .I(e[249]), 
        .Q(ein[249]) );
  DFF \ereg_reg[250]  ( .D(ereg_next[250]), .CLK(clk), .RST(rst), .I(e[250]), 
        .Q(ein[250]) );
  DFF \ereg_reg[251]  ( .D(ereg_next[251]), .CLK(clk), .RST(rst), .I(e[251]), 
        .Q(ein[251]) );
  DFF \ereg_reg[252]  ( .D(ereg_next[252]), .CLK(clk), .RST(rst), .I(e[252]), 
        .Q(ein[252]) );
  DFF \ereg_reg[253]  ( .D(ereg_next[253]), .CLK(clk), .RST(rst), .I(e[253]), 
        .Q(ein[253]) );
  DFF \ereg_reg[254]  ( .D(ereg_next[254]), .CLK(clk), .RST(rst), .I(e[254]), 
        .Q(ein[254]) );
  DFF \ereg_reg[255]  ( .D(ereg_next[255]), .CLK(clk), .RST(rst), .I(e[255]), 
        .Q(ein[255]) );
  DFF \ereg_reg[256]  ( .D(ereg_next[256]), .CLK(clk), .RST(rst), .I(e[256]), 
        .Q(ein[256]) );
  DFF \ereg_reg[257]  ( .D(ereg_next[257]), .CLK(clk), .RST(rst), .I(e[257]), 
        .Q(ein[257]) );
  DFF \ereg_reg[258]  ( .D(ereg_next[258]), .CLK(clk), .RST(rst), .I(e[258]), 
        .Q(ein[258]) );
  DFF \ereg_reg[259]  ( .D(ereg_next[259]), .CLK(clk), .RST(rst), .I(e[259]), 
        .Q(ein[259]) );
  DFF \ereg_reg[260]  ( .D(ereg_next[260]), .CLK(clk), .RST(rst), .I(e[260]), 
        .Q(ein[260]) );
  DFF \ereg_reg[261]  ( .D(ereg_next[261]), .CLK(clk), .RST(rst), .I(e[261]), 
        .Q(ein[261]) );
  DFF \ereg_reg[262]  ( .D(ereg_next[262]), .CLK(clk), .RST(rst), .I(e[262]), 
        .Q(ein[262]) );
  DFF \ereg_reg[263]  ( .D(ereg_next[263]), .CLK(clk), .RST(rst), .I(e[263]), 
        .Q(ein[263]) );
  DFF \ereg_reg[264]  ( .D(ereg_next[264]), .CLK(clk), .RST(rst), .I(e[264]), 
        .Q(ein[264]) );
  DFF \ereg_reg[265]  ( .D(ereg_next[265]), .CLK(clk), .RST(rst), .I(e[265]), 
        .Q(ein[265]) );
  DFF \ereg_reg[266]  ( .D(ereg_next[266]), .CLK(clk), .RST(rst), .I(e[266]), 
        .Q(ein[266]) );
  DFF \ereg_reg[267]  ( .D(ereg_next[267]), .CLK(clk), .RST(rst), .I(e[267]), 
        .Q(ein[267]) );
  DFF \ereg_reg[268]  ( .D(ereg_next[268]), .CLK(clk), .RST(rst), .I(e[268]), 
        .Q(ein[268]) );
  DFF \ereg_reg[269]  ( .D(ereg_next[269]), .CLK(clk), .RST(rst), .I(e[269]), 
        .Q(ein[269]) );
  DFF \ereg_reg[270]  ( .D(ereg_next[270]), .CLK(clk), .RST(rst), .I(e[270]), 
        .Q(ein[270]) );
  DFF \ereg_reg[271]  ( .D(ereg_next[271]), .CLK(clk), .RST(rst), .I(e[271]), 
        .Q(ein[271]) );
  DFF \ereg_reg[272]  ( .D(ereg_next[272]), .CLK(clk), .RST(rst), .I(e[272]), 
        .Q(ein[272]) );
  DFF \ereg_reg[273]  ( .D(ereg_next[273]), .CLK(clk), .RST(rst), .I(e[273]), 
        .Q(ein[273]) );
  DFF \ereg_reg[274]  ( .D(ereg_next[274]), .CLK(clk), .RST(rst), .I(e[274]), 
        .Q(ein[274]) );
  DFF \ereg_reg[275]  ( .D(ereg_next[275]), .CLK(clk), .RST(rst), .I(e[275]), 
        .Q(ein[275]) );
  DFF \ereg_reg[276]  ( .D(ereg_next[276]), .CLK(clk), .RST(rst), .I(e[276]), 
        .Q(ein[276]) );
  DFF \ereg_reg[277]  ( .D(ereg_next[277]), .CLK(clk), .RST(rst), .I(e[277]), 
        .Q(ein[277]) );
  DFF \ereg_reg[278]  ( .D(ereg_next[278]), .CLK(clk), .RST(rst), .I(e[278]), 
        .Q(ein[278]) );
  DFF \ereg_reg[279]  ( .D(ereg_next[279]), .CLK(clk), .RST(rst), .I(e[279]), 
        .Q(ein[279]) );
  DFF \ereg_reg[280]  ( .D(ereg_next[280]), .CLK(clk), .RST(rst), .I(e[280]), 
        .Q(ein[280]) );
  DFF \ereg_reg[281]  ( .D(ereg_next[281]), .CLK(clk), .RST(rst), .I(e[281]), 
        .Q(ein[281]) );
  DFF \ereg_reg[282]  ( .D(ereg_next[282]), .CLK(clk), .RST(rst), .I(e[282]), 
        .Q(ein[282]) );
  DFF \ereg_reg[283]  ( .D(ereg_next[283]), .CLK(clk), .RST(rst), .I(e[283]), 
        .Q(ein[283]) );
  DFF \ereg_reg[284]  ( .D(ereg_next[284]), .CLK(clk), .RST(rst), .I(e[284]), 
        .Q(ein[284]) );
  DFF \ereg_reg[285]  ( .D(ereg_next[285]), .CLK(clk), .RST(rst), .I(e[285]), 
        .Q(ein[285]) );
  DFF \ereg_reg[286]  ( .D(ereg_next[286]), .CLK(clk), .RST(rst), .I(e[286]), 
        .Q(ein[286]) );
  DFF \ereg_reg[287]  ( .D(ereg_next[287]), .CLK(clk), .RST(rst), .I(e[287]), 
        .Q(ein[287]) );
  DFF \ereg_reg[288]  ( .D(ereg_next[288]), .CLK(clk), .RST(rst), .I(e[288]), 
        .Q(ein[288]) );
  DFF \ereg_reg[289]  ( .D(ereg_next[289]), .CLK(clk), .RST(rst), .I(e[289]), 
        .Q(ein[289]) );
  DFF \ereg_reg[290]  ( .D(ereg_next[290]), .CLK(clk), .RST(rst), .I(e[290]), 
        .Q(ein[290]) );
  DFF \ereg_reg[291]  ( .D(ereg_next[291]), .CLK(clk), .RST(rst), .I(e[291]), 
        .Q(ein[291]) );
  DFF \ereg_reg[292]  ( .D(ereg_next[292]), .CLK(clk), .RST(rst), .I(e[292]), 
        .Q(ein[292]) );
  DFF \ereg_reg[293]  ( .D(ereg_next[293]), .CLK(clk), .RST(rst), .I(e[293]), 
        .Q(ein[293]) );
  DFF \ereg_reg[294]  ( .D(ereg_next[294]), .CLK(clk), .RST(rst), .I(e[294]), 
        .Q(ein[294]) );
  DFF \ereg_reg[295]  ( .D(ereg_next[295]), .CLK(clk), .RST(rst), .I(e[295]), 
        .Q(ein[295]) );
  DFF \ereg_reg[296]  ( .D(ereg_next[296]), .CLK(clk), .RST(rst), .I(e[296]), 
        .Q(ein[296]) );
  DFF \ereg_reg[297]  ( .D(ereg_next[297]), .CLK(clk), .RST(rst), .I(e[297]), 
        .Q(ein[297]) );
  DFF \ereg_reg[298]  ( .D(ereg_next[298]), .CLK(clk), .RST(rst), .I(e[298]), 
        .Q(ein[298]) );
  DFF \ereg_reg[299]  ( .D(ereg_next[299]), .CLK(clk), .RST(rst), .I(e[299]), 
        .Q(ein[299]) );
  DFF \ereg_reg[300]  ( .D(ereg_next[300]), .CLK(clk), .RST(rst), .I(e[300]), 
        .Q(ein[300]) );
  DFF \ereg_reg[301]  ( .D(ereg_next[301]), .CLK(clk), .RST(rst), .I(e[301]), 
        .Q(ein[301]) );
  DFF \ereg_reg[302]  ( .D(ereg_next[302]), .CLK(clk), .RST(rst), .I(e[302]), 
        .Q(ein[302]) );
  DFF \ereg_reg[303]  ( .D(ereg_next[303]), .CLK(clk), .RST(rst), .I(e[303]), 
        .Q(ein[303]) );
  DFF \ereg_reg[304]  ( .D(ereg_next[304]), .CLK(clk), .RST(rst), .I(e[304]), 
        .Q(ein[304]) );
  DFF \ereg_reg[305]  ( .D(ereg_next[305]), .CLK(clk), .RST(rst), .I(e[305]), 
        .Q(ein[305]) );
  DFF \ereg_reg[306]  ( .D(ereg_next[306]), .CLK(clk), .RST(rst), .I(e[306]), 
        .Q(ein[306]) );
  DFF \ereg_reg[307]  ( .D(ereg_next[307]), .CLK(clk), .RST(rst), .I(e[307]), 
        .Q(ein[307]) );
  DFF \ereg_reg[308]  ( .D(ereg_next[308]), .CLK(clk), .RST(rst), .I(e[308]), 
        .Q(ein[308]) );
  DFF \ereg_reg[309]  ( .D(ereg_next[309]), .CLK(clk), .RST(rst), .I(e[309]), 
        .Q(ein[309]) );
  DFF \ereg_reg[310]  ( .D(ereg_next[310]), .CLK(clk), .RST(rst), .I(e[310]), 
        .Q(ein[310]) );
  DFF \ereg_reg[311]  ( .D(ereg_next[311]), .CLK(clk), .RST(rst), .I(e[311]), 
        .Q(ein[311]) );
  DFF \ereg_reg[312]  ( .D(ereg_next[312]), .CLK(clk), .RST(rst), .I(e[312]), 
        .Q(ein[312]) );
  DFF \ereg_reg[313]  ( .D(ereg_next[313]), .CLK(clk), .RST(rst), .I(e[313]), 
        .Q(ein[313]) );
  DFF \ereg_reg[314]  ( .D(ereg_next[314]), .CLK(clk), .RST(rst), .I(e[314]), 
        .Q(ein[314]) );
  DFF \ereg_reg[315]  ( .D(ereg_next[315]), .CLK(clk), .RST(rst), .I(e[315]), 
        .Q(ein[315]) );
  DFF \ereg_reg[316]  ( .D(ereg_next[316]), .CLK(clk), .RST(rst), .I(e[316]), 
        .Q(ein[316]) );
  DFF \ereg_reg[317]  ( .D(ereg_next[317]), .CLK(clk), .RST(rst), .I(e[317]), 
        .Q(ein[317]) );
  DFF \ereg_reg[318]  ( .D(ereg_next[318]), .CLK(clk), .RST(rst), .I(e[318]), 
        .Q(ein[318]) );
  DFF \ereg_reg[319]  ( .D(ereg_next[319]), .CLK(clk), .RST(rst), .I(e[319]), 
        .Q(ein[319]) );
  DFF \ereg_reg[320]  ( .D(ereg_next[320]), .CLK(clk), .RST(rst), .I(e[320]), 
        .Q(ein[320]) );
  DFF \ereg_reg[321]  ( .D(ereg_next[321]), .CLK(clk), .RST(rst), .I(e[321]), 
        .Q(ein[321]) );
  DFF \ereg_reg[322]  ( .D(ereg_next[322]), .CLK(clk), .RST(rst), .I(e[322]), 
        .Q(ein[322]) );
  DFF \ereg_reg[323]  ( .D(ereg_next[323]), .CLK(clk), .RST(rst), .I(e[323]), 
        .Q(ein[323]) );
  DFF \ereg_reg[324]  ( .D(ereg_next[324]), .CLK(clk), .RST(rst), .I(e[324]), 
        .Q(ein[324]) );
  DFF \ereg_reg[325]  ( .D(ereg_next[325]), .CLK(clk), .RST(rst), .I(e[325]), 
        .Q(ein[325]) );
  DFF \ereg_reg[326]  ( .D(ereg_next[326]), .CLK(clk), .RST(rst), .I(e[326]), 
        .Q(ein[326]) );
  DFF \ereg_reg[327]  ( .D(ereg_next[327]), .CLK(clk), .RST(rst), .I(e[327]), 
        .Q(ein[327]) );
  DFF \ereg_reg[328]  ( .D(ereg_next[328]), .CLK(clk), .RST(rst), .I(e[328]), 
        .Q(ein[328]) );
  DFF \ereg_reg[329]  ( .D(ereg_next[329]), .CLK(clk), .RST(rst), .I(e[329]), 
        .Q(ein[329]) );
  DFF \ereg_reg[330]  ( .D(ereg_next[330]), .CLK(clk), .RST(rst), .I(e[330]), 
        .Q(ein[330]) );
  DFF \ereg_reg[331]  ( .D(ereg_next[331]), .CLK(clk), .RST(rst), .I(e[331]), 
        .Q(ein[331]) );
  DFF \ereg_reg[332]  ( .D(ereg_next[332]), .CLK(clk), .RST(rst), .I(e[332]), 
        .Q(ein[332]) );
  DFF \ereg_reg[333]  ( .D(ereg_next[333]), .CLK(clk), .RST(rst), .I(e[333]), 
        .Q(ein[333]) );
  DFF \ereg_reg[334]  ( .D(ereg_next[334]), .CLK(clk), .RST(rst), .I(e[334]), 
        .Q(ein[334]) );
  DFF \ereg_reg[335]  ( .D(ereg_next[335]), .CLK(clk), .RST(rst), .I(e[335]), 
        .Q(ein[335]) );
  DFF \ereg_reg[336]  ( .D(ereg_next[336]), .CLK(clk), .RST(rst), .I(e[336]), 
        .Q(ein[336]) );
  DFF \ereg_reg[337]  ( .D(ereg_next[337]), .CLK(clk), .RST(rst), .I(e[337]), 
        .Q(ein[337]) );
  DFF \ereg_reg[338]  ( .D(ereg_next[338]), .CLK(clk), .RST(rst), .I(e[338]), 
        .Q(ein[338]) );
  DFF \ereg_reg[339]  ( .D(ereg_next[339]), .CLK(clk), .RST(rst), .I(e[339]), 
        .Q(ein[339]) );
  DFF \ereg_reg[340]  ( .D(ereg_next[340]), .CLK(clk), .RST(rst), .I(e[340]), 
        .Q(ein[340]) );
  DFF \ereg_reg[341]  ( .D(ereg_next[341]), .CLK(clk), .RST(rst), .I(e[341]), 
        .Q(ein[341]) );
  DFF \ereg_reg[342]  ( .D(ereg_next[342]), .CLK(clk), .RST(rst), .I(e[342]), 
        .Q(ein[342]) );
  DFF \ereg_reg[343]  ( .D(ereg_next[343]), .CLK(clk), .RST(rst), .I(e[343]), 
        .Q(ein[343]) );
  DFF \ereg_reg[344]  ( .D(ereg_next[344]), .CLK(clk), .RST(rst), .I(e[344]), 
        .Q(ein[344]) );
  DFF \ereg_reg[345]  ( .D(ereg_next[345]), .CLK(clk), .RST(rst), .I(e[345]), 
        .Q(ein[345]) );
  DFF \ereg_reg[346]  ( .D(ereg_next[346]), .CLK(clk), .RST(rst), .I(e[346]), 
        .Q(ein[346]) );
  DFF \ereg_reg[347]  ( .D(ereg_next[347]), .CLK(clk), .RST(rst), .I(e[347]), 
        .Q(ein[347]) );
  DFF \ereg_reg[348]  ( .D(ereg_next[348]), .CLK(clk), .RST(rst), .I(e[348]), 
        .Q(ein[348]) );
  DFF \ereg_reg[349]  ( .D(ereg_next[349]), .CLK(clk), .RST(rst), .I(e[349]), 
        .Q(ein[349]) );
  DFF \ereg_reg[350]  ( .D(ereg_next[350]), .CLK(clk), .RST(rst), .I(e[350]), 
        .Q(ein[350]) );
  DFF \ereg_reg[351]  ( .D(ereg_next[351]), .CLK(clk), .RST(rst), .I(e[351]), 
        .Q(ein[351]) );
  DFF \ereg_reg[352]  ( .D(ereg_next[352]), .CLK(clk), .RST(rst), .I(e[352]), 
        .Q(ein[352]) );
  DFF \ereg_reg[353]  ( .D(ereg_next[353]), .CLK(clk), .RST(rst), .I(e[353]), 
        .Q(ein[353]) );
  DFF \ereg_reg[354]  ( .D(ereg_next[354]), .CLK(clk), .RST(rst), .I(e[354]), 
        .Q(ein[354]) );
  DFF \ereg_reg[355]  ( .D(ereg_next[355]), .CLK(clk), .RST(rst), .I(e[355]), 
        .Q(ein[355]) );
  DFF \ereg_reg[356]  ( .D(ereg_next[356]), .CLK(clk), .RST(rst), .I(e[356]), 
        .Q(ein[356]) );
  DFF \ereg_reg[357]  ( .D(ereg_next[357]), .CLK(clk), .RST(rst), .I(e[357]), 
        .Q(ein[357]) );
  DFF \ereg_reg[358]  ( .D(ereg_next[358]), .CLK(clk), .RST(rst), .I(e[358]), 
        .Q(ein[358]) );
  DFF \ereg_reg[359]  ( .D(ereg_next[359]), .CLK(clk), .RST(rst), .I(e[359]), 
        .Q(ein[359]) );
  DFF \ereg_reg[360]  ( .D(ereg_next[360]), .CLK(clk), .RST(rst), .I(e[360]), 
        .Q(ein[360]) );
  DFF \ereg_reg[361]  ( .D(ereg_next[361]), .CLK(clk), .RST(rst), .I(e[361]), 
        .Q(ein[361]) );
  DFF \ereg_reg[362]  ( .D(ereg_next[362]), .CLK(clk), .RST(rst), .I(e[362]), 
        .Q(ein[362]) );
  DFF \ereg_reg[363]  ( .D(ereg_next[363]), .CLK(clk), .RST(rst), .I(e[363]), 
        .Q(ein[363]) );
  DFF \ereg_reg[364]  ( .D(ereg_next[364]), .CLK(clk), .RST(rst), .I(e[364]), 
        .Q(ein[364]) );
  DFF \ereg_reg[365]  ( .D(ereg_next[365]), .CLK(clk), .RST(rst), .I(e[365]), 
        .Q(ein[365]) );
  DFF \ereg_reg[366]  ( .D(ereg_next[366]), .CLK(clk), .RST(rst), .I(e[366]), 
        .Q(ein[366]) );
  DFF \ereg_reg[367]  ( .D(ereg_next[367]), .CLK(clk), .RST(rst), .I(e[367]), 
        .Q(ein[367]) );
  DFF \ereg_reg[368]  ( .D(ereg_next[368]), .CLK(clk), .RST(rst), .I(e[368]), 
        .Q(ein[368]) );
  DFF \ereg_reg[369]  ( .D(ereg_next[369]), .CLK(clk), .RST(rst), .I(e[369]), 
        .Q(ein[369]) );
  DFF \ereg_reg[370]  ( .D(ereg_next[370]), .CLK(clk), .RST(rst), .I(e[370]), 
        .Q(ein[370]) );
  DFF \ereg_reg[371]  ( .D(ereg_next[371]), .CLK(clk), .RST(rst), .I(e[371]), 
        .Q(ein[371]) );
  DFF \ereg_reg[372]  ( .D(ereg_next[372]), .CLK(clk), .RST(rst), .I(e[372]), 
        .Q(ein[372]) );
  DFF \ereg_reg[373]  ( .D(ereg_next[373]), .CLK(clk), .RST(rst), .I(e[373]), 
        .Q(ein[373]) );
  DFF \ereg_reg[374]  ( .D(ereg_next[374]), .CLK(clk), .RST(rst), .I(e[374]), 
        .Q(ein[374]) );
  DFF \ereg_reg[375]  ( .D(ereg_next[375]), .CLK(clk), .RST(rst), .I(e[375]), 
        .Q(ein[375]) );
  DFF \ereg_reg[376]  ( .D(ereg_next[376]), .CLK(clk), .RST(rst), .I(e[376]), 
        .Q(ein[376]) );
  DFF \ereg_reg[377]  ( .D(ereg_next[377]), .CLK(clk), .RST(rst), .I(e[377]), 
        .Q(ein[377]) );
  DFF \ereg_reg[378]  ( .D(ereg_next[378]), .CLK(clk), .RST(rst), .I(e[378]), 
        .Q(ein[378]) );
  DFF \ereg_reg[379]  ( .D(ereg_next[379]), .CLK(clk), .RST(rst), .I(e[379]), 
        .Q(ein[379]) );
  DFF \ereg_reg[380]  ( .D(ereg_next[380]), .CLK(clk), .RST(rst), .I(e[380]), 
        .Q(ein[380]) );
  DFF \ereg_reg[381]  ( .D(ereg_next[381]), .CLK(clk), .RST(rst), .I(e[381]), 
        .Q(ein[381]) );
  DFF \ereg_reg[382]  ( .D(ereg_next[382]), .CLK(clk), .RST(rst), .I(e[382]), 
        .Q(ein[382]) );
  DFF \ereg_reg[383]  ( .D(ereg_next[383]), .CLK(clk), .RST(rst), .I(e[383]), 
        .Q(ein[383]) );
  DFF \ereg_reg[384]  ( .D(ereg_next[384]), .CLK(clk), .RST(rst), .I(e[384]), 
        .Q(ein[384]) );
  DFF \ereg_reg[385]  ( .D(ereg_next[385]), .CLK(clk), .RST(rst), .I(e[385]), 
        .Q(ein[385]) );
  DFF \ereg_reg[386]  ( .D(ereg_next[386]), .CLK(clk), .RST(rst), .I(e[386]), 
        .Q(ein[386]) );
  DFF \ereg_reg[387]  ( .D(ereg_next[387]), .CLK(clk), .RST(rst), .I(e[387]), 
        .Q(ein[387]) );
  DFF \ereg_reg[388]  ( .D(ereg_next[388]), .CLK(clk), .RST(rst), .I(e[388]), 
        .Q(ein[388]) );
  DFF \ereg_reg[389]  ( .D(ereg_next[389]), .CLK(clk), .RST(rst), .I(e[389]), 
        .Q(ein[389]) );
  DFF \ereg_reg[390]  ( .D(ereg_next[390]), .CLK(clk), .RST(rst), .I(e[390]), 
        .Q(ein[390]) );
  DFF \ereg_reg[391]  ( .D(ereg_next[391]), .CLK(clk), .RST(rst), .I(e[391]), 
        .Q(ein[391]) );
  DFF \ereg_reg[392]  ( .D(ereg_next[392]), .CLK(clk), .RST(rst), .I(e[392]), 
        .Q(ein[392]) );
  DFF \ereg_reg[393]  ( .D(ereg_next[393]), .CLK(clk), .RST(rst), .I(e[393]), 
        .Q(ein[393]) );
  DFF \ereg_reg[394]  ( .D(ereg_next[394]), .CLK(clk), .RST(rst), .I(e[394]), 
        .Q(ein[394]) );
  DFF \ereg_reg[395]  ( .D(ereg_next[395]), .CLK(clk), .RST(rst), .I(e[395]), 
        .Q(ein[395]) );
  DFF \ereg_reg[396]  ( .D(ereg_next[396]), .CLK(clk), .RST(rst), .I(e[396]), 
        .Q(ein[396]) );
  DFF \ereg_reg[397]  ( .D(ereg_next[397]), .CLK(clk), .RST(rst), .I(e[397]), 
        .Q(ein[397]) );
  DFF \ereg_reg[398]  ( .D(ereg_next[398]), .CLK(clk), .RST(rst), .I(e[398]), 
        .Q(ein[398]) );
  DFF \ereg_reg[399]  ( .D(ereg_next[399]), .CLK(clk), .RST(rst), .I(e[399]), 
        .Q(ein[399]) );
  DFF \ereg_reg[400]  ( .D(ereg_next[400]), .CLK(clk), .RST(rst), .I(e[400]), 
        .Q(ein[400]) );
  DFF \ereg_reg[401]  ( .D(ereg_next[401]), .CLK(clk), .RST(rst), .I(e[401]), 
        .Q(ein[401]) );
  DFF \ereg_reg[402]  ( .D(ereg_next[402]), .CLK(clk), .RST(rst), .I(e[402]), 
        .Q(ein[402]) );
  DFF \ereg_reg[403]  ( .D(ereg_next[403]), .CLK(clk), .RST(rst), .I(e[403]), 
        .Q(ein[403]) );
  DFF \ereg_reg[404]  ( .D(ereg_next[404]), .CLK(clk), .RST(rst), .I(e[404]), 
        .Q(ein[404]) );
  DFF \ereg_reg[405]  ( .D(ereg_next[405]), .CLK(clk), .RST(rst), .I(e[405]), 
        .Q(ein[405]) );
  DFF \ereg_reg[406]  ( .D(ereg_next[406]), .CLK(clk), .RST(rst), .I(e[406]), 
        .Q(ein[406]) );
  DFF \ereg_reg[407]  ( .D(ereg_next[407]), .CLK(clk), .RST(rst), .I(e[407]), 
        .Q(ein[407]) );
  DFF \ereg_reg[408]  ( .D(ereg_next[408]), .CLK(clk), .RST(rst), .I(e[408]), 
        .Q(ein[408]) );
  DFF \ereg_reg[409]  ( .D(ereg_next[409]), .CLK(clk), .RST(rst), .I(e[409]), 
        .Q(ein[409]) );
  DFF \ereg_reg[410]  ( .D(ereg_next[410]), .CLK(clk), .RST(rst), .I(e[410]), 
        .Q(ein[410]) );
  DFF \ereg_reg[411]  ( .D(ereg_next[411]), .CLK(clk), .RST(rst), .I(e[411]), 
        .Q(ein[411]) );
  DFF \ereg_reg[412]  ( .D(ereg_next[412]), .CLK(clk), .RST(rst), .I(e[412]), 
        .Q(ein[412]) );
  DFF \ereg_reg[413]  ( .D(ereg_next[413]), .CLK(clk), .RST(rst), .I(e[413]), 
        .Q(ein[413]) );
  DFF \ereg_reg[414]  ( .D(ereg_next[414]), .CLK(clk), .RST(rst), .I(e[414]), 
        .Q(ein[414]) );
  DFF \ereg_reg[415]  ( .D(ereg_next[415]), .CLK(clk), .RST(rst), .I(e[415]), 
        .Q(ein[415]) );
  DFF \ereg_reg[416]  ( .D(ereg_next[416]), .CLK(clk), .RST(rst), .I(e[416]), 
        .Q(ein[416]) );
  DFF \ereg_reg[417]  ( .D(ereg_next[417]), .CLK(clk), .RST(rst), .I(e[417]), 
        .Q(ein[417]) );
  DFF \ereg_reg[418]  ( .D(ereg_next[418]), .CLK(clk), .RST(rst), .I(e[418]), 
        .Q(ein[418]) );
  DFF \ereg_reg[419]  ( .D(ereg_next[419]), .CLK(clk), .RST(rst), .I(e[419]), 
        .Q(ein[419]) );
  DFF \ereg_reg[420]  ( .D(ereg_next[420]), .CLK(clk), .RST(rst), .I(e[420]), 
        .Q(ein[420]) );
  DFF \ereg_reg[421]  ( .D(ereg_next[421]), .CLK(clk), .RST(rst), .I(e[421]), 
        .Q(ein[421]) );
  DFF \ereg_reg[422]  ( .D(ereg_next[422]), .CLK(clk), .RST(rst), .I(e[422]), 
        .Q(ein[422]) );
  DFF \ereg_reg[423]  ( .D(ereg_next[423]), .CLK(clk), .RST(rst), .I(e[423]), 
        .Q(ein[423]) );
  DFF \ereg_reg[424]  ( .D(ereg_next[424]), .CLK(clk), .RST(rst), .I(e[424]), 
        .Q(ein[424]) );
  DFF \ereg_reg[425]  ( .D(ereg_next[425]), .CLK(clk), .RST(rst), .I(e[425]), 
        .Q(ein[425]) );
  DFF \ereg_reg[426]  ( .D(ereg_next[426]), .CLK(clk), .RST(rst), .I(e[426]), 
        .Q(ein[426]) );
  DFF \ereg_reg[427]  ( .D(ereg_next[427]), .CLK(clk), .RST(rst), .I(e[427]), 
        .Q(ein[427]) );
  DFF \ereg_reg[428]  ( .D(ereg_next[428]), .CLK(clk), .RST(rst), .I(e[428]), 
        .Q(ein[428]) );
  DFF \ereg_reg[429]  ( .D(ereg_next[429]), .CLK(clk), .RST(rst), .I(e[429]), 
        .Q(ein[429]) );
  DFF \ereg_reg[430]  ( .D(ereg_next[430]), .CLK(clk), .RST(rst), .I(e[430]), 
        .Q(ein[430]) );
  DFF \ereg_reg[431]  ( .D(ereg_next[431]), .CLK(clk), .RST(rst), .I(e[431]), 
        .Q(ein[431]) );
  DFF \ereg_reg[432]  ( .D(ereg_next[432]), .CLK(clk), .RST(rst), .I(e[432]), 
        .Q(ein[432]) );
  DFF \ereg_reg[433]  ( .D(ereg_next[433]), .CLK(clk), .RST(rst), .I(e[433]), 
        .Q(ein[433]) );
  DFF \ereg_reg[434]  ( .D(ereg_next[434]), .CLK(clk), .RST(rst), .I(e[434]), 
        .Q(ein[434]) );
  DFF \ereg_reg[435]  ( .D(ereg_next[435]), .CLK(clk), .RST(rst), .I(e[435]), 
        .Q(ein[435]) );
  DFF \ereg_reg[436]  ( .D(ereg_next[436]), .CLK(clk), .RST(rst), .I(e[436]), 
        .Q(ein[436]) );
  DFF \ereg_reg[437]  ( .D(ereg_next[437]), .CLK(clk), .RST(rst), .I(e[437]), 
        .Q(ein[437]) );
  DFF \ereg_reg[438]  ( .D(ereg_next[438]), .CLK(clk), .RST(rst), .I(e[438]), 
        .Q(ein[438]) );
  DFF \ereg_reg[439]  ( .D(ereg_next[439]), .CLK(clk), .RST(rst), .I(e[439]), 
        .Q(ein[439]) );
  DFF \ereg_reg[440]  ( .D(ereg_next[440]), .CLK(clk), .RST(rst), .I(e[440]), 
        .Q(ein[440]) );
  DFF \ereg_reg[441]  ( .D(ereg_next[441]), .CLK(clk), .RST(rst), .I(e[441]), 
        .Q(ein[441]) );
  DFF \ereg_reg[442]  ( .D(ereg_next[442]), .CLK(clk), .RST(rst), .I(e[442]), 
        .Q(ein[442]) );
  DFF \ereg_reg[443]  ( .D(ereg_next[443]), .CLK(clk), .RST(rst), .I(e[443]), 
        .Q(ein[443]) );
  DFF \ereg_reg[444]  ( .D(ereg_next[444]), .CLK(clk), .RST(rst), .I(e[444]), 
        .Q(ein[444]) );
  DFF \ereg_reg[445]  ( .D(ereg_next[445]), .CLK(clk), .RST(rst), .I(e[445]), 
        .Q(ein[445]) );
  DFF \ereg_reg[446]  ( .D(ereg_next[446]), .CLK(clk), .RST(rst), .I(e[446]), 
        .Q(ein[446]) );
  DFF \ereg_reg[447]  ( .D(ereg_next[447]), .CLK(clk), .RST(rst), .I(e[447]), 
        .Q(ein[447]) );
  DFF \ereg_reg[448]  ( .D(ereg_next[448]), .CLK(clk), .RST(rst), .I(e[448]), 
        .Q(ein[448]) );
  DFF \ereg_reg[449]  ( .D(ereg_next[449]), .CLK(clk), .RST(rst), .I(e[449]), 
        .Q(ein[449]) );
  DFF \ereg_reg[450]  ( .D(ereg_next[450]), .CLK(clk), .RST(rst), .I(e[450]), 
        .Q(ein[450]) );
  DFF \ereg_reg[451]  ( .D(ereg_next[451]), .CLK(clk), .RST(rst), .I(e[451]), 
        .Q(ein[451]) );
  DFF \ereg_reg[452]  ( .D(ereg_next[452]), .CLK(clk), .RST(rst), .I(e[452]), 
        .Q(ein[452]) );
  DFF \ereg_reg[453]  ( .D(ereg_next[453]), .CLK(clk), .RST(rst), .I(e[453]), 
        .Q(ein[453]) );
  DFF \ereg_reg[454]  ( .D(ereg_next[454]), .CLK(clk), .RST(rst), .I(e[454]), 
        .Q(ein[454]) );
  DFF \ereg_reg[455]  ( .D(ereg_next[455]), .CLK(clk), .RST(rst), .I(e[455]), 
        .Q(ein[455]) );
  DFF \ereg_reg[456]  ( .D(ereg_next[456]), .CLK(clk), .RST(rst), .I(e[456]), 
        .Q(ein[456]) );
  DFF \ereg_reg[457]  ( .D(ereg_next[457]), .CLK(clk), .RST(rst), .I(e[457]), 
        .Q(ein[457]) );
  DFF \ereg_reg[458]  ( .D(ereg_next[458]), .CLK(clk), .RST(rst), .I(e[458]), 
        .Q(ein[458]) );
  DFF \ereg_reg[459]  ( .D(ereg_next[459]), .CLK(clk), .RST(rst), .I(e[459]), 
        .Q(ein[459]) );
  DFF \ereg_reg[460]  ( .D(ereg_next[460]), .CLK(clk), .RST(rst), .I(e[460]), 
        .Q(ein[460]) );
  DFF \ereg_reg[461]  ( .D(ereg_next[461]), .CLK(clk), .RST(rst), .I(e[461]), 
        .Q(ein[461]) );
  DFF \ereg_reg[462]  ( .D(ereg_next[462]), .CLK(clk), .RST(rst), .I(e[462]), 
        .Q(ein[462]) );
  DFF \ereg_reg[463]  ( .D(ereg_next[463]), .CLK(clk), .RST(rst), .I(e[463]), 
        .Q(ein[463]) );
  DFF \ereg_reg[464]  ( .D(ereg_next[464]), .CLK(clk), .RST(rst), .I(e[464]), 
        .Q(ein[464]) );
  DFF \ereg_reg[465]  ( .D(ereg_next[465]), .CLK(clk), .RST(rst), .I(e[465]), 
        .Q(ein[465]) );
  DFF \ereg_reg[466]  ( .D(ereg_next[466]), .CLK(clk), .RST(rst), .I(e[466]), 
        .Q(ein[466]) );
  DFF \ereg_reg[467]  ( .D(ereg_next[467]), .CLK(clk), .RST(rst), .I(e[467]), 
        .Q(ein[467]) );
  DFF \ereg_reg[468]  ( .D(ereg_next[468]), .CLK(clk), .RST(rst), .I(e[468]), 
        .Q(ein[468]) );
  DFF \ereg_reg[469]  ( .D(ereg_next[469]), .CLK(clk), .RST(rst), .I(e[469]), 
        .Q(ein[469]) );
  DFF \ereg_reg[470]  ( .D(ereg_next[470]), .CLK(clk), .RST(rst), .I(e[470]), 
        .Q(ein[470]) );
  DFF \ereg_reg[471]  ( .D(ereg_next[471]), .CLK(clk), .RST(rst), .I(e[471]), 
        .Q(ein[471]) );
  DFF \ereg_reg[472]  ( .D(ereg_next[472]), .CLK(clk), .RST(rst), .I(e[472]), 
        .Q(ein[472]) );
  DFF \ereg_reg[473]  ( .D(ereg_next[473]), .CLK(clk), .RST(rst), .I(e[473]), 
        .Q(ein[473]) );
  DFF \ereg_reg[474]  ( .D(ereg_next[474]), .CLK(clk), .RST(rst), .I(e[474]), 
        .Q(ein[474]) );
  DFF \ereg_reg[475]  ( .D(ereg_next[475]), .CLK(clk), .RST(rst), .I(e[475]), 
        .Q(ein[475]) );
  DFF \ereg_reg[476]  ( .D(ereg_next[476]), .CLK(clk), .RST(rst), .I(e[476]), 
        .Q(ein[476]) );
  DFF \ereg_reg[477]  ( .D(ereg_next[477]), .CLK(clk), .RST(rst), .I(e[477]), 
        .Q(ein[477]) );
  DFF \ereg_reg[478]  ( .D(ereg_next[478]), .CLK(clk), .RST(rst), .I(e[478]), 
        .Q(ein[478]) );
  DFF \ereg_reg[479]  ( .D(ereg_next[479]), .CLK(clk), .RST(rst), .I(e[479]), 
        .Q(ein[479]) );
  DFF \ereg_reg[480]  ( .D(ereg_next[480]), .CLK(clk), .RST(rst), .I(e[480]), 
        .Q(ein[480]) );
  DFF \ereg_reg[481]  ( .D(ereg_next[481]), .CLK(clk), .RST(rst), .I(e[481]), 
        .Q(ein[481]) );
  DFF \ereg_reg[482]  ( .D(ereg_next[482]), .CLK(clk), .RST(rst), .I(e[482]), 
        .Q(ein[482]) );
  DFF \ereg_reg[483]  ( .D(ereg_next[483]), .CLK(clk), .RST(rst), .I(e[483]), 
        .Q(ein[483]) );
  DFF \ereg_reg[484]  ( .D(ereg_next[484]), .CLK(clk), .RST(rst), .I(e[484]), 
        .Q(ein[484]) );
  DFF \ereg_reg[485]  ( .D(ereg_next[485]), .CLK(clk), .RST(rst), .I(e[485]), 
        .Q(ein[485]) );
  DFF \ereg_reg[486]  ( .D(ereg_next[486]), .CLK(clk), .RST(rst), .I(e[486]), 
        .Q(ein[486]) );
  DFF \ereg_reg[487]  ( .D(ereg_next[487]), .CLK(clk), .RST(rst), .I(e[487]), 
        .Q(ein[487]) );
  DFF \ereg_reg[488]  ( .D(ereg_next[488]), .CLK(clk), .RST(rst), .I(e[488]), 
        .Q(ein[488]) );
  DFF \ereg_reg[489]  ( .D(ereg_next[489]), .CLK(clk), .RST(rst), .I(e[489]), 
        .Q(ein[489]) );
  DFF \ereg_reg[490]  ( .D(ereg_next[490]), .CLK(clk), .RST(rst), .I(e[490]), 
        .Q(ein[490]) );
  DFF \ereg_reg[491]  ( .D(ereg_next[491]), .CLK(clk), .RST(rst), .I(e[491]), 
        .Q(ein[491]) );
  DFF \ereg_reg[492]  ( .D(ereg_next[492]), .CLK(clk), .RST(rst), .I(e[492]), 
        .Q(ein[492]) );
  DFF \ereg_reg[493]  ( .D(ereg_next[493]), .CLK(clk), .RST(rst), .I(e[493]), 
        .Q(ein[493]) );
  DFF \ereg_reg[494]  ( .D(ereg_next[494]), .CLK(clk), .RST(rst), .I(e[494]), 
        .Q(ein[494]) );
  DFF \ereg_reg[495]  ( .D(ereg_next[495]), .CLK(clk), .RST(rst), .I(e[495]), 
        .Q(ein[495]) );
  DFF \ereg_reg[496]  ( .D(ereg_next[496]), .CLK(clk), .RST(rst), .I(e[496]), 
        .Q(ein[496]) );
  DFF \ereg_reg[497]  ( .D(ereg_next[497]), .CLK(clk), .RST(rst), .I(e[497]), 
        .Q(ein[497]) );
  DFF \ereg_reg[498]  ( .D(ereg_next[498]), .CLK(clk), .RST(rst), .I(e[498]), 
        .Q(ein[498]) );
  DFF \ereg_reg[499]  ( .D(ereg_next[499]), .CLK(clk), .RST(rst), .I(e[499]), 
        .Q(ein[499]) );
  DFF \ereg_reg[500]  ( .D(ereg_next[500]), .CLK(clk), .RST(rst), .I(e[500]), 
        .Q(ein[500]) );
  DFF \ereg_reg[501]  ( .D(ereg_next[501]), .CLK(clk), .RST(rst), .I(e[501]), 
        .Q(ein[501]) );
  DFF \ereg_reg[502]  ( .D(ereg_next[502]), .CLK(clk), .RST(rst), .I(e[502]), 
        .Q(ein[502]) );
  DFF \ereg_reg[503]  ( .D(ereg_next[503]), .CLK(clk), .RST(rst), .I(e[503]), 
        .Q(ein[503]) );
  DFF \ereg_reg[504]  ( .D(ereg_next[504]), .CLK(clk), .RST(rst), .I(e[504]), 
        .Q(ein[504]) );
  DFF \ereg_reg[505]  ( .D(ereg_next[505]), .CLK(clk), .RST(rst), .I(e[505]), 
        .Q(ein[505]) );
  DFF \ereg_reg[506]  ( .D(ereg_next[506]), .CLK(clk), .RST(rst), .I(e[506]), 
        .Q(ein[506]) );
  DFF \ereg_reg[507]  ( .D(ereg_next[507]), .CLK(clk), .RST(rst), .I(e[507]), 
        .Q(ein[507]) );
  DFF \ereg_reg[508]  ( .D(ereg_next[508]), .CLK(clk), .RST(rst), .I(e[508]), 
        .Q(ein[508]) );
  DFF \ereg_reg[509]  ( .D(ereg_next[509]), .CLK(clk), .RST(rst), .I(e[509]), 
        .Q(ein[509]) );
  DFF \ereg_reg[510]  ( .D(ereg_next[510]), .CLK(clk), .RST(rst), .I(e[510]), 
        .Q(ein[510]) );
  DFF \ereg_reg[511]  ( .D(ereg_next[511]), .CLK(clk), .RST(rst), .I(e[511]), 
        .Q(ein[511]) );
  DFF first_one_reg ( .D(n6), .CLK(clk), .RST(rst), .I(1'b0), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(creg_next[0]), .CLK(clk), .RST(rst), .I(m[0]), .Q(
        c[0]) );
  DFF \creg_reg[1]  ( .D(creg_next[1]), .CLK(clk), .RST(rst), .I(m[1]), .Q(
        c[1]) );
  DFF \creg_reg[2]  ( .D(creg_next[2]), .CLK(clk), .RST(rst), .I(m[2]), .Q(
        c[2]) );
  DFF \creg_reg[3]  ( .D(creg_next[3]), .CLK(clk), .RST(rst), .I(m[3]), .Q(
        c[3]) );
  DFF \creg_reg[4]  ( .D(creg_next[4]), .CLK(clk), .RST(rst), .I(m[4]), .Q(
        c[4]) );
  DFF \creg_reg[5]  ( .D(creg_next[5]), .CLK(clk), .RST(rst), .I(m[5]), .Q(
        c[5]) );
  DFF \creg_reg[6]  ( .D(creg_next[6]), .CLK(clk), .RST(rst), .I(m[6]), .Q(
        c[6]) );
  DFF \creg_reg[7]  ( .D(creg_next[7]), .CLK(clk), .RST(rst), .I(m[7]), .Q(
        c[7]) );
  DFF \creg_reg[8]  ( .D(creg_next[8]), .CLK(clk), .RST(rst), .I(m[8]), .Q(
        c[8]) );
  DFF \creg_reg[9]  ( .D(creg_next[9]), .CLK(clk), .RST(rst), .I(m[9]), .Q(
        c[9]) );
  DFF \creg_reg[10]  ( .D(creg_next[10]), .CLK(clk), .RST(rst), .I(m[10]), .Q(
        c[10]) );
  DFF \creg_reg[11]  ( .D(creg_next[11]), .CLK(clk), .RST(rst), .I(m[11]), .Q(
        c[11]) );
  DFF \creg_reg[12]  ( .D(creg_next[12]), .CLK(clk), .RST(rst), .I(m[12]), .Q(
        c[12]) );
  DFF \creg_reg[13]  ( .D(creg_next[13]), .CLK(clk), .RST(rst), .I(m[13]), .Q(
        c[13]) );
  DFF \creg_reg[14]  ( .D(creg_next[14]), .CLK(clk), .RST(rst), .I(m[14]), .Q(
        c[14]) );
  DFF \creg_reg[15]  ( .D(creg_next[15]), .CLK(clk), .RST(rst), .I(m[15]), .Q(
        c[15]) );
  DFF \creg_reg[16]  ( .D(creg_next[16]), .CLK(clk), .RST(rst), .I(m[16]), .Q(
        c[16]) );
  DFF \creg_reg[17]  ( .D(creg_next[17]), .CLK(clk), .RST(rst), .I(m[17]), .Q(
        c[17]) );
  DFF \creg_reg[18]  ( .D(creg_next[18]), .CLK(clk), .RST(rst), .I(m[18]), .Q(
        c[18]) );
  DFF \creg_reg[19]  ( .D(creg_next[19]), .CLK(clk), .RST(rst), .I(m[19]), .Q(
        c[19]) );
  DFF \creg_reg[20]  ( .D(creg_next[20]), .CLK(clk), .RST(rst), .I(m[20]), .Q(
        c[20]) );
  DFF \creg_reg[21]  ( .D(creg_next[21]), .CLK(clk), .RST(rst), .I(m[21]), .Q(
        c[21]) );
  DFF \creg_reg[22]  ( .D(creg_next[22]), .CLK(clk), .RST(rst), .I(m[22]), .Q(
        c[22]) );
  DFF \creg_reg[23]  ( .D(creg_next[23]), .CLK(clk), .RST(rst), .I(m[23]), .Q(
        c[23]) );
  DFF \creg_reg[24]  ( .D(creg_next[24]), .CLK(clk), .RST(rst), .I(m[24]), .Q(
        c[24]) );
  DFF \creg_reg[25]  ( .D(creg_next[25]), .CLK(clk), .RST(rst), .I(m[25]), .Q(
        c[25]) );
  DFF \creg_reg[26]  ( .D(creg_next[26]), .CLK(clk), .RST(rst), .I(m[26]), .Q(
        c[26]) );
  DFF \creg_reg[27]  ( .D(creg_next[27]), .CLK(clk), .RST(rst), .I(m[27]), .Q(
        c[27]) );
  DFF \creg_reg[28]  ( .D(creg_next[28]), .CLK(clk), .RST(rst), .I(m[28]), .Q(
        c[28]) );
  DFF \creg_reg[29]  ( .D(creg_next[29]), .CLK(clk), .RST(rst), .I(m[29]), .Q(
        c[29]) );
  DFF \creg_reg[30]  ( .D(creg_next[30]), .CLK(clk), .RST(rst), .I(m[30]), .Q(
        c[30]) );
  DFF \creg_reg[31]  ( .D(creg_next[31]), .CLK(clk), .RST(rst), .I(m[31]), .Q(
        c[31]) );
  DFF \creg_reg[32]  ( .D(creg_next[32]), .CLK(clk), .RST(rst), .I(m[32]), .Q(
        c[32]) );
  DFF \creg_reg[33]  ( .D(creg_next[33]), .CLK(clk), .RST(rst), .I(m[33]), .Q(
        c[33]) );
  DFF \creg_reg[34]  ( .D(creg_next[34]), .CLK(clk), .RST(rst), .I(m[34]), .Q(
        c[34]) );
  DFF \creg_reg[35]  ( .D(creg_next[35]), .CLK(clk), .RST(rst), .I(m[35]), .Q(
        c[35]) );
  DFF \creg_reg[36]  ( .D(creg_next[36]), .CLK(clk), .RST(rst), .I(m[36]), .Q(
        c[36]) );
  DFF \creg_reg[37]  ( .D(creg_next[37]), .CLK(clk), .RST(rst), .I(m[37]), .Q(
        c[37]) );
  DFF \creg_reg[38]  ( .D(creg_next[38]), .CLK(clk), .RST(rst), .I(m[38]), .Q(
        c[38]) );
  DFF \creg_reg[39]  ( .D(creg_next[39]), .CLK(clk), .RST(rst), .I(m[39]), .Q(
        c[39]) );
  DFF \creg_reg[40]  ( .D(creg_next[40]), .CLK(clk), .RST(rst), .I(m[40]), .Q(
        c[40]) );
  DFF \creg_reg[41]  ( .D(creg_next[41]), .CLK(clk), .RST(rst), .I(m[41]), .Q(
        c[41]) );
  DFF \creg_reg[42]  ( .D(creg_next[42]), .CLK(clk), .RST(rst), .I(m[42]), .Q(
        c[42]) );
  DFF \creg_reg[43]  ( .D(creg_next[43]), .CLK(clk), .RST(rst), .I(m[43]), .Q(
        c[43]) );
  DFF \creg_reg[44]  ( .D(creg_next[44]), .CLK(clk), .RST(rst), .I(m[44]), .Q(
        c[44]) );
  DFF \creg_reg[45]  ( .D(creg_next[45]), .CLK(clk), .RST(rst), .I(m[45]), .Q(
        c[45]) );
  DFF \creg_reg[46]  ( .D(creg_next[46]), .CLK(clk), .RST(rst), .I(m[46]), .Q(
        c[46]) );
  DFF \creg_reg[47]  ( .D(creg_next[47]), .CLK(clk), .RST(rst), .I(m[47]), .Q(
        c[47]) );
  DFF \creg_reg[48]  ( .D(creg_next[48]), .CLK(clk), .RST(rst), .I(m[48]), .Q(
        c[48]) );
  DFF \creg_reg[49]  ( .D(creg_next[49]), .CLK(clk), .RST(rst), .I(m[49]), .Q(
        c[49]) );
  DFF \creg_reg[50]  ( .D(creg_next[50]), .CLK(clk), .RST(rst), .I(m[50]), .Q(
        c[50]) );
  DFF \creg_reg[51]  ( .D(creg_next[51]), .CLK(clk), .RST(rst), .I(m[51]), .Q(
        c[51]) );
  DFF \creg_reg[52]  ( .D(creg_next[52]), .CLK(clk), .RST(rst), .I(m[52]), .Q(
        c[52]) );
  DFF \creg_reg[53]  ( .D(creg_next[53]), .CLK(clk), .RST(rst), .I(m[53]), .Q(
        c[53]) );
  DFF \creg_reg[54]  ( .D(creg_next[54]), .CLK(clk), .RST(rst), .I(m[54]), .Q(
        c[54]) );
  DFF \creg_reg[55]  ( .D(creg_next[55]), .CLK(clk), .RST(rst), .I(m[55]), .Q(
        c[55]) );
  DFF \creg_reg[56]  ( .D(creg_next[56]), .CLK(clk), .RST(rst), .I(m[56]), .Q(
        c[56]) );
  DFF \creg_reg[57]  ( .D(creg_next[57]), .CLK(clk), .RST(rst), .I(m[57]), .Q(
        c[57]) );
  DFF \creg_reg[58]  ( .D(creg_next[58]), .CLK(clk), .RST(rst), .I(m[58]), .Q(
        c[58]) );
  DFF \creg_reg[59]  ( .D(creg_next[59]), .CLK(clk), .RST(rst), .I(m[59]), .Q(
        c[59]) );
  DFF \creg_reg[60]  ( .D(creg_next[60]), .CLK(clk), .RST(rst), .I(m[60]), .Q(
        c[60]) );
  DFF \creg_reg[61]  ( .D(creg_next[61]), .CLK(clk), .RST(rst), .I(m[61]), .Q(
        c[61]) );
  DFF \creg_reg[62]  ( .D(creg_next[62]), .CLK(clk), .RST(rst), .I(m[62]), .Q(
        c[62]) );
  DFF \creg_reg[63]  ( .D(creg_next[63]), .CLK(clk), .RST(rst), .I(m[63]), .Q(
        c[63]) );
  DFF \creg_reg[64]  ( .D(creg_next[64]), .CLK(clk), .RST(rst), .I(m[64]), .Q(
        c[64]) );
  DFF \creg_reg[65]  ( .D(creg_next[65]), .CLK(clk), .RST(rst), .I(m[65]), .Q(
        c[65]) );
  DFF \creg_reg[66]  ( .D(creg_next[66]), .CLK(clk), .RST(rst), .I(m[66]), .Q(
        c[66]) );
  DFF \creg_reg[67]  ( .D(creg_next[67]), .CLK(clk), .RST(rst), .I(m[67]), .Q(
        c[67]) );
  DFF \creg_reg[68]  ( .D(creg_next[68]), .CLK(clk), .RST(rst), .I(m[68]), .Q(
        c[68]) );
  DFF \creg_reg[69]  ( .D(creg_next[69]), .CLK(clk), .RST(rst), .I(m[69]), .Q(
        c[69]) );
  DFF \creg_reg[70]  ( .D(creg_next[70]), .CLK(clk), .RST(rst), .I(m[70]), .Q(
        c[70]) );
  DFF \creg_reg[71]  ( .D(creg_next[71]), .CLK(clk), .RST(rst), .I(m[71]), .Q(
        c[71]) );
  DFF \creg_reg[72]  ( .D(creg_next[72]), .CLK(clk), .RST(rst), .I(m[72]), .Q(
        c[72]) );
  DFF \creg_reg[73]  ( .D(creg_next[73]), .CLK(clk), .RST(rst), .I(m[73]), .Q(
        c[73]) );
  DFF \creg_reg[74]  ( .D(creg_next[74]), .CLK(clk), .RST(rst), .I(m[74]), .Q(
        c[74]) );
  DFF \creg_reg[75]  ( .D(creg_next[75]), .CLK(clk), .RST(rst), .I(m[75]), .Q(
        c[75]) );
  DFF \creg_reg[76]  ( .D(creg_next[76]), .CLK(clk), .RST(rst), .I(m[76]), .Q(
        c[76]) );
  DFF \creg_reg[77]  ( .D(creg_next[77]), .CLK(clk), .RST(rst), .I(m[77]), .Q(
        c[77]) );
  DFF \creg_reg[78]  ( .D(creg_next[78]), .CLK(clk), .RST(rst), .I(m[78]), .Q(
        c[78]) );
  DFF \creg_reg[79]  ( .D(creg_next[79]), .CLK(clk), .RST(rst), .I(m[79]), .Q(
        c[79]) );
  DFF \creg_reg[80]  ( .D(creg_next[80]), .CLK(clk), .RST(rst), .I(m[80]), .Q(
        c[80]) );
  DFF \creg_reg[81]  ( .D(creg_next[81]), .CLK(clk), .RST(rst), .I(m[81]), .Q(
        c[81]) );
  DFF \creg_reg[82]  ( .D(creg_next[82]), .CLK(clk), .RST(rst), .I(m[82]), .Q(
        c[82]) );
  DFF \creg_reg[83]  ( .D(creg_next[83]), .CLK(clk), .RST(rst), .I(m[83]), .Q(
        c[83]) );
  DFF \creg_reg[84]  ( .D(creg_next[84]), .CLK(clk), .RST(rst), .I(m[84]), .Q(
        c[84]) );
  DFF \creg_reg[85]  ( .D(creg_next[85]), .CLK(clk), .RST(rst), .I(m[85]), .Q(
        c[85]) );
  DFF \creg_reg[86]  ( .D(creg_next[86]), .CLK(clk), .RST(rst), .I(m[86]), .Q(
        c[86]) );
  DFF \creg_reg[87]  ( .D(creg_next[87]), .CLK(clk), .RST(rst), .I(m[87]), .Q(
        c[87]) );
  DFF \creg_reg[88]  ( .D(creg_next[88]), .CLK(clk), .RST(rst), .I(m[88]), .Q(
        c[88]) );
  DFF \creg_reg[89]  ( .D(creg_next[89]), .CLK(clk), .RST(rst), .I(m[89]), .Q(
        c[89]) );
  DFF \creg_reg[90]  ( .D(creg_next[90]), .CLK(clk), .RST(rst), .I(m[90]), .Q(
        c[90]) );
  DFF \creg_reg[91]  ( .D(creg_next[91]), .CLK(clk), .RST(rst), .I(m[91]), .Q(
        c[91]) );
  DFF \creg_reg[92]  ( .D(creg_next[92]), .CLK(clk), .RST(rst), .I(m[92]), .Q(
        c[92]) );
  DFF \creg_reg[93]  ( .D(creg_next[93]), .CLK(clk), .RST(rst), .I(m[93]), .Q(
        c[93]) );
  DFF \creg_reg[94]  ( .D(creg_next[94]), .CLK(clk), .RST(rst), .I(m[94]), .Q(
        c[94]) );
  DFF \creg_reg[95]  ( .D(creg_next[95]), .CLK(clk), .RST(rst), .I(m[95]), .Q(
        c[95]) );
  DFF \creg_reg[96]  ( .D(creg_next[96]), .CLK(clk), .RST(rst), .I(m[96]), .Q(
        c[96]) );
  DFF \creg_reg[97]  ( .D(creg_next[97]), .CLK(clk), .RST(rst), .I(m[97]), .Q(
        c[97]) );
  DFF \creg_reg[98]  ( .D(creg_next[98]), .CLK(clk), .RST(rst), .I(m[98]), .Q(
        c[98]) );
  DFF \creg_reg[99]  ( .D(creg_next[99]), .CLK(clk), .RST(rst), .I(m[99]), .Q(
        c[99]) );
  DFF \creg_reg[100]  ( .D(creg_next[100]), .CLK(clk), .RST(rst), .I(m[100]), 
        .Q(c[100]) );
  DFF \creg_reg[101]  ( .D(creg_next[101]), .CLK(clk), .RST(rst), .I(m[101]), 
        .Q(c[101]) );
  DFF \creg_reg[102]  ( .D(creg_next[102]), .CLK(clk), .RST(rst), .I(m[102]), 
        .Q(c[102]) );
  DFF \creg_reg[103]  ( .D(creg_next[103]), .CLK(clk), .RST(rst), .I(m[103]), 
        .Q(c[103]) );
  DFF \creg_reg[104]  ( .D(creg_next[104]), .CLK(clk), .RST(rst), .I(m[104]), 
        .Q(c[104]) );
  DFF \creg_reg[105]  ( .D(creg_next[105]), .CLK(clk), .RST(rst), .I(m[105]), 
        .Q(c[105]) );
  DFF \creg_reg[106]  ( .D(creg_next[106]), .CLK(clk), .RST(rst), .I(m[106]), 
        .Q(c[106]) );
  DFF \creg_reg[107]  ( .D(creg_next[107]), .CLK(clk), .RST(rst), .I(m[107]), 
        .Q(c[107]) );
  DFF \creg_reg[108]  ( .D(creg_next[108]), .CLK(clk), .RST(rst), .I(m[108]), 
        .Q(c[108]) );
  DFF \creg_reg[109]  ( .D(creg_next[109]), .CLK(clk), .RST(rst), .I(m[109]), 
        .Q(c[109]) );
  DFF \creg_reg[110]  ( .D(creg_next[110]), .CLK(clk), .RST(rst), .I(m[110]), 
        .Q(c[110]) );
  DFF \creg_reg[111]  ( .D(creg_next[111]), .CLK(clk), .RST(rst), .I(m[111]), 
        .Q(c[111]) );
  DFF \creg_reg[112]  ( .D(creg_next[112]), .CLK(clk), .RST(rst), .I(m[112]), 
        .Q(c[112]) );
  DFF \creg_reg[113]  ( .D(creg_next[113]), .CLK(clk), .RST(rst), .I(m[113]), 
        .Q(c[113]) );
  DFF \creg_reg[114]  ( .D(creg_next[114]), .CLK(clk), .RST(rst), .I(m[114]), 
        .Q(c[114]) );
  DFF \creg_reg[115]  ( .D(creg_next[115]), .CLK(clk), .RST(rst), .I(m[115]), 
        .Q(c[115]) );
  DFF \creg_reg[116]  ( .D(creg_next[116]), .CLK(clk), .RST(rst), .I(m[116]), 
        .Q(c[116]) );
  DFF \creg_reg[117]  ( .D(creg_next[117]), .CLK(clk), .RST(rst), .I(m[117]), 
        .Q(c[117]) );
  DFF \creg_reg[118]  ( .D(creg_next[118]), .CLK(clk), .RST(rst), .I(m[118]), 
        .Q(c[118]) );
  DFF \creg_reg[119]  ( .D(creg_next[119]), .CLK(clk), .RST(rst), .I(m[119]), 
        .Q(c[119]) );
  DFF \creg_reg[120]  ( .D(creg_next[120]), .CLK(clk), .RST(rst), .I(m[120]), 
        .Q(c[120]) );
  DFF \creg_reg[121]  ( .D(creg_next[121]), .CLK(clk), .RST(rst), .I(m[121]), 
        .Q(c[121]) );
  DFF \creg_reg[122]  ( .D(creg_next[122]), .CLK(clk), .RST(rst), .I(m[122]), 
        .Q(c[122]) );
  DFF \creg_reg[123]  ( .D(creg_next[123]), .CLK(clk), .RST(rst), .I(m[123]), 
        .Q(c[123]) );
  DFF \creg_reg[124]  ( .D(creg_next[124]), .CLK(clk), .RST(rst), .I(m[124]), 
        .Q(c[124]) );
  DFF \creg_reg[125]  ( .D(creg_next[125]), .CLK(clk), .RST(rst), .I(m[125]), 
        .Q(c[125]) );
  DFF \creg_reg[126]  ( .D(creg_next[126]), .CLK(clk), .RST(rst), .I(m[126]), 
        .Q(c[126]) );
  DFF \creg_reg[127]  ( .D(creg_next[127]), .CLK(clk), .RST(rst), .I(m[127]), 
        .Q(c[127]) );
  DFF \creg_reg[128]  ( .D(creg_next[128]), .CLK(clk), .RST(rst), .I(m[128]), 
        .Q(c[128]) );
  DFF \creg_reg[129]  ( .D(creg_next[129]), .CLK(clk), .RST(rst), .I(m[129]), 
        .Q(c[129]) );
  DFF \creg_reg[130]  ( .D(creg_next[130]), .CLK(clk), .RST(rst), .I(m[130]), 
        .Q(c[130]) );
  DFF \creg_reg[131]  ( .D(creg_next[131]), .CLK(clk), .RST(rst), .I(m[131]), 
        .Q(c[131]) );
  DFF \creg_reg[132]  ( .D(creg_next[132]), .CLK(clk), .RST(rst), .I(m[132]), 
        .Q(c[132]) );
  DFF \creg_reg[133]  ( .D(creg_next[133]), .CLK(clk), .RST(rst), .I(m[133]), 
        .Q(c[133]) );
  DFF \creg_reg[134]  ( .D(creg_next[134]), .CLK(clk), .RST(rst), .I(m[134]), 
        .Q(c[134]) );
  DFF \creg_reg[135]  ( .D(creg_next[135]), .CLK(clk), .RST(rst), .I(m[135]), 
        .Q(c[135]) );
  DFF \creg_reg[136]  ( .D(creg_next[136]), .CLK(clk), .RST(rst), .I(m[136]), 
        .Q(c[136]) );
  DFF \creg_reg[137]  ( .D(creg_next[137]), .CLK(clk), .RST(rst), .I(m[137]), 
        .Q(c[137]) );
  DFF \creg_reg[138]  ( .D(creg_next[138]), .CLK(clk), .RST(rst), .I(m[138]), 
        .Q(c[138]) );
  DFF \creg_reg[139]  ( .D(creg_next[139]), .CLK(clk), .RST(rst), .I(m[139]), 
        .Q(c[139]) );
  DFF \creg_reg[140]  ( .D(creg_next[140]), .CLK(clk), .RST(rst), .I(m[140]), 
        .Q(c[140]) );
  DFF \creg_reg[141]  ( .D(creg_next[141]), .CLK(clk), .RST(rst), .I(m[141]), 
        .Q(c[141]) );
  DFF \creg_reg[142]  ( .D(creg_next[142]), .CLK(clk), .RST(rst), .I(m[142]), 
        .Q(c[142]) );
  DFF \creg_reg[143]  ( .D(creg_next[143]), .CLK(clk), .RST(rst), .I(m[143]), 
        .Q(c[143]) );
  DFF \creg_reg[144]  ( .D(creg_next[144]), .CLK(clk), .RST(rst), .I(m[144]), 
        .Q(c[144]) );
  DFF \creg_reg[145]  ( .D(creg_next[145]), .CLK(clk), .RST(rst), .I(m[145]), 
        .Q(c[145]) );
  DFF \creg_reg[146]  ( .D(creg_next[146]), .CLK(clk), .RST(rst), .I(m[146]), 
        .Q(c[146]) );
  DFF \creg_reg[147]  ( .D(creg_next[147]), .CLK(clk), .RST(rst), .I(m[147]), 
        .Q(c[147]) );
  DFF \creg_reg[148]  ( .D(creg_next[148]), .CLK(clk), .RST(rst), .I(m[148]), 
        .Q(c[148]) );
  DFF \creg_reg[149]  ( .D(creg_next[149]), .CLK(clk), .RST(rst), .I(m[149]), 
        .Q(c[149]) );
  DFF \creg_reg[150]  ( .D(creg_next[150]), .CLK(clk), .RST(rst), .I(m[150]), 
        .Q(c[150]) );
  DFF \creg_reg[151]  ( .D(creg_next[151]), .CLK(clk), .RST(rst), .I(m[151]), 
        .Q(c[151]) );
  DFF \creg_reg[152]  ( .D(creg_next[152]), .CLK(clk), .RST(rst), .I(m[152]), 
        .Q(c[152]) );
  DFF \creg_reg[153]  ( .D(creg_next[153]), .CLK(clk), .RST(rst), .I(m[153]), 
        .Q(c[153]) );
  DFF \creg_reg[154]  ( .D(creg_next[154]), .CLK(clk), .RST(rst), .I(m[154]), 
        .Q(c[154]) );
  DFF \creg_reg[155]  ( .D(creg_next[155]), .CLK(clk), .RST(rst), .I(m[155]), 
        .Q(c[155]) );
  DFF \creg_reg[156]  ( .D(creg_next[156]), .CLK(clk), .RST(rst), .I(m[156]), 
        .Q(c[156]) );
  DFF \creg_reg[157]  ( .D(creg_next[157]), .CLK(clk), .RST(rst), .I(m[157]), 
        .Q(c[157]) );
  DFF \creg_reg[158]  ( .D(creg_next[158]), .CLK(clk), .RST(rst), .I(m[158]), 
        .Q(c[158]) );
  DFF \creg_reg[159]  ( .D(creg_next[159]), .CLK(clk), .RST(rst), .I(m[159]), 
        .Q(c[159]) );
  DFF \creg_reg[160]  ( .D(creg_next[160]), .CLK(clk), .RST(rst), .I(m[160]), 
        .Q(c[160]) );
  DFF \creg_reg[161]  ( .D(creg_next[161]), .CLK(clk), .RST(rst), .I(m[161]), 
        .Q(c[161]) );
  DFF \creg_reg[162]  ( .D(creg_next[162]), .CLK(clk), .RST(rst), .I(m[162]), 
        .Q(c[162]) );
  DFF \creg_reg[163]  ( .D(creg_next[163]), .CLK(clk), .RST(rst), .I(m[163]), 
        .Q(c[163]) );
  DFF \creg_reg[164]  ( .D(creg_next[164]), .CLK(clk), .RST(rst), .I(m[164]), 
        .Q(c[164]) );
  DFF \creg_reg[165]  ( .D(creg_next[165]), .CLK(clk), .RST(rst), .I(m[165]), 
        .Q(c[165]) );
  DFF \creg_reg[166]  ( .D(creg_next[166]), .CLK(clk), .RST(rst), .I(m[166]), 
        .Q(c[166]) );
  DFF \creg_reg[167]  ( .D(creg_next[167]), .CLK(clk), .RST(rst), .I(m[167]), 
        .Q(c[167]) );
  DFF \creg_reg[168]  ( .D(creg_next[168]), .CLK(clk), .RST(rst), .I(m[168]), 
        .Q(c[168]) );
  DFF \creg_reg[169]  ( .D(creg_next[169]), .CLK(clk), .RST(rst), .I(m[169]), 
        .Q(c[169]) );
  DFF \creg_reg[170]  ( .D(creg_next[170]), .CLK(clk), .RST(rst), .I(m[170]), 
        .Q(c[170]) );
  DFF \creg_reg[171]  ( .D(creg_next[171]), .CLK(clk), .RST(rst), .I(m[171]), 
        .Q(c[171]) );
  DFF \creg_reg[172]  ( .D(creg_next[172]), .CLK(clk), .RST(rst), .I(m[172]), 
        .Q(c[172]) );
  DFF \creg_reg[173]  ( .D(creg_next[173]), .CLK(clk), .RST(rst), .I(m[173]), 
        .Q(c[173]) );
  DFF \creg_reg[174]  ( .D(creg_next[174]), .CLK(clk), .RST(rst), .I(m[174]), 
        .Q(c[174]) );
  DFF \creg_reg[175]  ( .D(creg_next[175]), .CLK(clk), .RST(rst), .I(m[175]), 
        .Q(c[175]) );
  DFF \creg_reg[176]  ( .D(creg_next[176]), .CLK(clk), .RST(rst), .I(m[176]), 
        .Q(c[176]) );
  DFF \creg_reg[177]  ( .D(creg_next[177]), .CLK(clk), .RST(rst), .I(m[177]), 
        .Q(c[177]) );
  DFF \creg_reg[178]  ( .D(creg_next[178]), .CLK(clk), .RST(rst), .I(m[178]), 
        .Q(c[178]) );
  DFF \creg_reg[179]  ( .D(creg_next[179]), .CLK(clk), .RST(rst), .I(m[179]), 
        .Q(c[179]) );
  DFF \creg_reg[180]  ( .D(creg_next[180]), .CLK(clk), .RST(rst), .I(m[180]), 
        .Q(c[180]) );
  DFF \creg_reg[181]  ( .D(creg_next[181]), .CLK(clk), .RST(rst), .I(m[181]), 
        .Q(c[181]) );
  DFF \creg_reg[182]  ( .D(creg_next[182]), .CLK(clk), .RST(rst), .I(m[182]), 
        .Q(c[182]) );
  DFF \creg_reg[183]  ( .D(creg_next[183]), .CLK(clk), .RST(rst), .I(m[183]), 
        .Q(c[183]) );
  DFF \creg_reg[184]  ( .D(creg_next[184]), .CLK(clk), .RST(rst), .I(m[184]), 
        .Q(c[184]) );
  DFF \creg_reg[185]  ( .D(creg_next[185]), .CLK(clk), .RST(rst), .I(m[185]), 
        .Q(c[185]) );
  DFF \creg_reg[186]  ( .D(creg_next[186]), .CLK(clk), .RST(rst), .I(m[186]), 
        .Q(c[186]) );
  DFF \creg_reg[187]  ( .D(creg_next[187]), .CLK(clk), .RST(rst), .I(m[187]), 
        .Q(c[187]) );
  DFF \creg_reg[188]  ( .D(creg_next[188]), .CLK(clk), .RST(rst), .I(m[188]), 
        .Q(c[188]) );
  DFF \creg_reg[189]  ( .D(creg_next[189]), .CLK(clk), .RST(rst), .I(m[189]), 
        .Q(c[189]) );
  DFF \creg_reg[190]  ( .D(creg_next[190]), .CLK(clk), .RST(rst), .I(m[190]), 
        .Q(c[190]) );
  DFF \creg_reg[191]  ( .D(creg_next[191]), .CLK(clk), .RST(rst), .I(m[191]), 
        .Q(c[191]) );
  DFF \creg_reg[192]  ( .D(creg_next[192]), .CLK(clk), .RST(rst), .I(m[192]), 
        .Q(c[192]) );
  DFF \creg_reg[193]  ( .D(creg_next[193]), .CLK(clk), .RST(rst), .I(m[193]), 
        .Q(c[193]) );
  DFF \creg_reg[194]  ( .D(creg_next[194]), .CLK(clk), .RST(rst), .I(m[194]), 
        .Q(c[194]) );
  DFF \creg_reg[195]  ( .D(creg_next[195]), .CLK(clk), .RST(rst), .I(m[195]), 
        .Q(c[195]) );
  DFF \creg_reg[196]  ( .D(creg_next[196]), .CLK(clk), .RST(rst), .I(m[196]), 
        .Q(c[196]) );
  DFF \creg_reg[197]  ( .D(creg_next[197]), .CLK(clk), .RST(rst), .I(m[197]), 
        .Q(c[197]) );
  DFF \creg_reg[198]  ( .D(creg_next[198]), .CLK(clk), .RST(rst), .I(m[198]), 
        .Q(c[198]) );
  DFF \creg_reg[199]  ( .D(creg_next[199]), .CLK(clk), .RST(rst), .I(m[199]), 
        .Q(c[199]) );
  DFF \creg_reg[200]  ( .D(creg_next[200]), .CLK(clk), .RST(rst), .I(m[200]), 
        .Q(c[200]) );
  DFF \creg_reg[201]  ( .D(creg_next[201]), .CLK(clk), .RST(rst), .I(m[201]), 
        .Q(c[201]) );
  DFF \creg_reg[202]  ( .D(creg_next[202]), .CLK(clk), .RST(rst), .I(m[202]), 
        .Q(c[202]) );
  DFF \creg_reg[203]  ( .D(creg_next[203]), .CLK(clk), .RST(rst), .I(m[203]), 
        .Q(c[203]) );
  DFF \creg_reg[204]  ( .D(creg_next[204]), .CLK(clk), .RST(rst), .I(m[204]), 
        .Q(c[204]) );
  DFF \creg_reg[205]  ( .D(creg_next[205]), .CLK(clk), .RST(rst), .I(m[205]), 
        .Q(c[205]) );
  DFF \creg_reg[206]  ( .D(creg_next[206]), .CLK(clk), .RST(rst), .I(m[206]), 
        .Q(c[206]) );
  DFF \creg_reg[207]  ( .D(creg_next[207]), .CLK(clk), .RST(rst), .I(m[207]), 
        .Q(c[207]) );
  DFF \creg_reg[208]  ( .D(creg_next[208]), .CLK(clk), .RST(rst), .I(m[208]), 
        .Q(c[208]) );
  DFF \creg_reg[209]  ( .D(creg_next[209]), .CLK(clk), .RST(rst), .I(m[209]), 
        .Q(c[209]) );
  DFF \creg_reg[210]  ( .D(creg_next[210]), .CLK(clk), .RST(rst), .I(m[210]), 
        .Q(c[210]) );
  DFF \creg_reg[211]  ( .D(creg_next[211]), .CLK(clk), .RST(rst), .I(m[211]), 
        .Q(c[211]) );
  DFF \creg_reg[212]  ( .D(creg_next[212]), .CLK(clk), .RST(rst), .I(m[212]), 
        .Q(c[212]) );
  DFF \creg_reg[213]  ( .D(creg_next[213]), .CLK(clk), .RST(rst), .I(m[213]), 
        .Q(c[213]) );
  DFF \creg_reg[214]  ( .D(creg_next[214]), .CLK(clk), .RST(rst), .I(m[214]), 
        .Q(c[214]) );
  DFF \creg_reg[215]  ( .D(creg_next[215]), .CLK(clk), .RST(rst), .I(m[215]), 
        .Q(c[215]) );
  DFF \creg_reg[216]  ( .D(creg_next[216]), .CLK(clk), .RST(rst), .I(m[216]), 
        .Q(c[216]) );
  DFF \creg_reg[217]  ( .D(creg_next[217]), .CLK(clk), .RST(rst), .I(m[217]), 
        .Q(c[217]) );
  DFF \creg_reg[218]  ( .D(creg_next[218]), .CLK(clk), .RST(rst), .I(m[218]), 
        .Q(c[218]) );
  DFF \creg_reg[219]  ( .D(creg_next[219]), .CLK(clk), .RST(rst), .I(m[219]), 
        .Q(c[219]) );
  DFF \creg_reg[220]  ( .D(creg_next[220]), .CLK(clk), .RST(rst), .I(m[220]), 
        .Q(c[220]) );
  DFF \creg_reg[221]  ( .D(creg_next[221]), .CLK(clk), .RST(rst), .I(m[221]), 
        .Q(c[221]) );
  DFF \creg_reg[222]  ( .D(creg_next[222]), .CLK(clk), .RST(rst), .I(m[222]), 
        .Q(c[222]) );
  DFF \creg_reg[223]  ( .D(creg_next[223]), .CLK(clk), .RST(rst), .I(m[223]), 
        .Q(c[223]) );
  DFF \creg_reg[224]  ( .D(creg_next[224]), .CLK(clk), .RST(rst), .I(m[224]), 
        .Q(c[224]) );
  DFF \creg_reg[225]  ( .D(creg_next[225]), .CLK(clk), .RST(rst), .I(m[225]), 
        .Q(c[225]) );
  DFF \creg_reg[226]  ( .D(creg_next[226]), .CLK(clk), .RST(rst), .I(m[226]), 
        .Q(c[226]) );
  DFF \creg_reg[227]  ( .D(creg_next[227]), .CLK(clk), .RST(rst), .I(m[227]), 
        .Q(c[227]) );
  DFF \creg_reg[228]  ( .D(creg_next[228]), .CLK(clk), .RST(rst), .I(m[228]), 
        .Q(c[228]) );
  DFF \creg_reg[229]  ( .D(creg_next[229]), .CLK(clk), .RST(rst), .I(m[229]), 
        .Q(c[229]) );
  DFF \creg_reg[230]  ( .D(creg_next[230]), .CLK(clk), .RST(rst), .I(m[230]), 
        .Q(c[230]) );
  DFF \creg_reg[231]  ( .D(creg_next[231]), .CLK(clk), .RST(rst), .I(m[231]), 
        .Q(c[231]) );
  DFF \creg_reg[232]  ( .D(creg_next[232]), .CLK(clk), .RST(rst), .I(m[232]), 
        .Q(c[232]) );
  DFF \creg_reg[233]  ( .D(creg_next[233]), .CLK(clk), .RST(rst), .I(m[233]), 
        .Q(c[233]) );
  DFF \creg_reg[234]  ( .D(creg_next[234]), .CLK(clk), .RST(rst), .I(m[234]), 
        .Q(c[234]) );
  DFF \creg_reg[235]  ( .D(creg_next[235]), .CLK(clk), .RST(rst), .I(m[235]), 
        .Q(c[235]) );
  DFF \creg_reg[236]  ( .D(creg_next[236]), .CLK(clk), .RST(rst), .I(m[236]), 
        .Q(c[236]) );
  DFF \creg_reg[237]  ( .D(creg_next[237]), .CLK(clk), .RST(rst), .I(m[237]), 
        .Q(c[237]) );
  DFF \creg_reg[238]  ( .D(creg_next[238]), .CLK(clk), .RST(rst), .I(m[238]), 
        .Q(c[238]) );
  DFF \creg_reg[239]  ( .D(creg_next[239]), .CLK(clk), .RST(rst), .I(m[239]), 
        .Q(c[239]) );
  DFF \creg_reg[240]  ( .D(creg_next[240]), .CLK(clk), .RST(rst), .I(m[240]), 
        .Q(c[240]) );
  DFF \creg_reg[241]  ( .D(creg_next[241]), .CLK(clk), .RST(rst), .I(m[241]), 
        .Q(c[241]) );
  DFF \creg_reg[242]  ( .D(creg_next[242]), .CLK(clk), .RST(rst), .I(m[242]), 
        .Q(c[242]) );
  DFF \creg_reg[243]  ( .D(creg_next[243]), .CLK(clk), .RST(rst), .I(m[243]), 
        .Q(c[243]) );
  DFF \creg_reg[244]  ( .D(creg_next[244]), .CLK(clk), .RST(rst), .I(m[244]), 
        .Q(c[244]) );
  DFF \creg_reg[245]  ( .D(creg_next[245]), .CLK(clk), .RST(rst), .I(m[245]), 
        .Q(c[245]) );
  DFF \creg_reg[246]  ( .D(creg_next[246]), .CLK(clk), .RST(rst), .I(m[246]), 
        .Q(c[246]) );
  DFF \creg_reg[247]  ( .D(creg_next[247]), .CLK(clk), .RST(rst), .I(m[247]), 
        .Q(c[247]) );
  DFF \creg_reg[248]  ( .D(creg_next[248]), .CLK(clk), .RST(rst), .I(m[248]), 
        .Q(c[248]) );
  DFF \creg_reg[249]  ( .D(creg_next[249]), .CLK(clk), .RST(rst), .I(m[249]), 
        .Q(c[249]) );
  DFF \creg_reg[250]  ( .D(creg_next[250]), .CLK(clk), .RST(rst), .I(m[250]), 
        .Q(c[250]) );
  DFF \creg_reg[251]  ( .D(creg_next[251]), .CLK(clk), .RST(rst), .I(m[251]), 
        .Q(c[251]) );
  DFF \creg_reg[252]  ( .D(creg_next[252]), .CLK(clk), .RST(rst), .I(m[252]), 
        .Q(c[252]) );
  DFF \creg_reg[253]  ( .D(creg_next[253]), .CLK(clk), .RST(rst), .I(m[253]), 
        .Q(c[253]) );
  DFF \creg_reg[254]  ( .D(creg_next[254]), .CLK(clk), .RST(rst), .I(m[254]), 
        .Q(c[254]) );
  DFF \creg_reg[255]  ( .D(creg_next[255]), .CLK(clk), .RST(rst), .I(m[255]), 
        .Q(c[255]) );
  DFF \creg_reg[256]  ( .D(creg_next[256]), .CLK(clk), .RST(rst), .I(m[256]), 
        .Q(c[256]) );
  DFF \creg_reg[257]  ( .D(creg_next[257]), .CLK(clk), .RST(rst), .I(m[257]), 
        .Q(c[257]) );
  DFF \creg_reg[258]  ( .D(creg_next[258]), .CLK(clk), .RST(rst), .I(m[258]), 
        .Q(c[258]) );
  DFF \creg_reg[259]  ( .D(creg_next[259]), .CLK(clk), .RST(rst), .I(m[259]), 
        .Q(c[259]) );
  DFF \creg_reg[260]  ( .D(creg_next[260]), .CLK(clk), .RST(rst), .I(m[260]), 
        .Q(c[260]) );
  DFF \creg_reg[261]  ( .D(creg_next[261]), .CLK(clk), .RST(rst), .I(m[261]), 
        .Q(c[261]) );
  DFF \creg_reg[262]  ( .D(creg_next[262]), .CLK(clk), .RST(rst), .I(m[262]), 
        .Q(c[262]) );
  DFF \creg_reg[263]  ( .D(creg_next[263]), .CLK(clk), .RST(rst), .I(m[263]), 
        .Q(c[263]) );
  DFF \creg_reg[264]  ( .D(creg_next[264]), .CLK(clk), .RST(rst), .I(m[264]), 
        .Q(c[264]) );
  DFF \creg_reg[265]  ( .D(creg_next[265]), .CLK(clk), .RST(rst), .I(m[265]), 
        .Q(c[265]) );
  DFF \creg_reg[266]  ( .D(creg_next[266]), .CLK(clk), .RST(rst), .I(m[266]), 
        .Q(c[266]) );
  DFF \creg_reg[267]  ( .D(creg_next[267]), .CLK(clk), .RST(rst), .I(m[267]), 
        .Q(c[267]) );
  DFF \creg_reg[268]  ( .D(creg_next[268]), .CLK(clk), .RST(rst), .I(m[268]), 
        .Q(c[268]) );
  DFF \creg_reg[269]  ( .D(creg_next[269]), .CLK(clk), .RST(rst), .I(m[269]), 
        .Q(c[269]) );
  DFF \creg_reg[270]  ( .D(creg_next[270]), .CLK(clk), .RST(rst), .I(m[270]), 
        .Q(c[270]) );
  DFF \creg_reg[271]  ( .D(creg_next[271]), .CLK(clk), .RST(rst), .I(m[271]), 
        .Q(c[271]) );
  DFF \creg_reg[272]  ( .D(creg_next[272]), .CLK(clk), .RST(rst), .I(m[272]), 
        .Q(c[272]) );
  DFF \creg_reg[273]  ( .D(creg_next[273]), .CLK(clk), .RST(rst), .I(m[273]), 
        .Q(c[273]) );
  DFF \creg_reg[274]  ( .D(creg_next[274]), .CLK(clk), .RST(rst), .I(m[274]), 
        .Q(c[274]) );
  DFF \creg_reg[275]  ( .D(creg_next[275]), .CLK(clk), .RST(rst), .I(m[275]), 
        .Q(c[275]) );
  DFF \creg_reg[276]  ( .D(creg_next[276]), .CLK(clk), .RST(rst), .I(m[276]), 
        .Q(c[276]) );
  DFF \creg_reg[277]  ( .D(creg_next[277]), .CLK(clk), .RST(rst), .I(m[277]), 
        .Q(c[277]) );
  DFF \creg_reg[278]  ( .D(creg_next[278]), .CLK(clk), .RST(rst), .I(m[278]), 
        .Q(c[278]) );
  DFF \creg_reg[279]  ( .D(creg_next[279]), .CLK(clk), .RST(rst), .I(m[279]), 
        .Q(c[279]) );
  DFF \creg_reg[280]  ( .D(creg_next[280]), .CLK(clk), .RST(rst), .I(m[280]), 
        .Q(c[280]) );
  DFF \creg_reg[281]  ( .D(creg_next[281]), .CLK(clk), .RST(rst), .I(m[281]), 
        .Q(c[281]) );
  DFF \creg_reg[282]  ( .D(creg_next[282]), .CLK(clk), .RST(rst), .I(m[282]), 
        .Q(c[282]) );
  DFF \creg_reg[283]  ( .D(creg_next[283]), .CLK(clk), .RST(rst), .I(m[283]), 
        .Q(c[283]) );
  DFF \creg_reg[284]  ( .D(creg_next[284]), .CLK(clk), .RST(rst), .I(m[284]), 
        .Q(c[284]) );
  DFF \creg_reg[285]  ( .D(creg_next[285]), .CLK(clk), .RST(rst), .I(m[285]), 
        .Q(c[285]) );
  DFF \creg_reg[286]  ( .D(creg_next[286]), .CLK(clk), .RST(rst), .I(m[286]), 
        .Q(c[286]) );
  DFF \creg_reg[287]  ( .D(creg_next[287]), .CLK(clk), .RST(rst), .I(m[287]), 
        .Q(c[287]) );
  DFF \creg_reg[288]  ( .D(creg_next[288]), .CLK(clk), .RST(rst), .I(m[288]), 
        .Q(c[288]) );
  DFF \creg_reg[289]  ( .D(creg_next[289]), .CLK(clk), .RST(rst), .I(m[289]), 
        .Q(c[289]) );
  DFF \creg_reg[290]  ( .D(creg_next[290]), .CLK(clk), .RST(rst), .I(m[290]), 
        .Q(c[290]) );
  DFF \creg_reg[291]  ( .D(creg_next[291]), .CLK(clk), .RST(rst), .I(m[291]), 
        .Q(c[291]) );
  DFF \creg_reg[292]  ( .D(creg_next[292]), .CLK(clk), .RST(rst), .I(m[292]), 
        .Q(c[292]) );
  DFF \creg_reg[293]  ( .D(creg_next[293]), .CLK(clk), .RST(rst), .I(m[293]), 
        .Q(c[293]) );
  DFF \creg_reg[294]  ( .D(creg_next[294]), .CLK(clk), .RST(rst), .I(m[294]), 
        .Q(c[294]) );
  DFF \creg_reg[295]  ( .D(creg_next[295]), .CLK(clk), .RST(rst), .I(m[295]), 
        .Q(c[295]) );
  DFF \creg_reg[296]  ( .D(creg_next[296]), .CLK(clk), .RST(rst), .I(m[296]), 
        .Q(c[296]) );
  DFF \creg_reg[297]  ( .D(creg_next[297]), .CLK(clk), .RST(rst), .I(m[297]), 
        .Q(c[297]) );
  DFF \creg_reg[298]  ( .D(creg_next[298]), .CLK(clk), .RST(rst), .I(m[298]), 
        .Q(c[298]) );
  DFF \creg_reg[299]  ( .D(creg_next[299]), .CLK(clk), .RST(rst), .I(m[299]), 
        .Q(c[299]) );
  DFF \creg_reg[300]  ( .D(creg_next[300]), .CLK(clk), .RST(rst), .I(m[300]), 
        .Q(c[300]) );
  DFF \creg_reg[301]  ( .D(creg_next[301]), .CLK(clk), .RST(rst), .I(m[301]), 
        .Q(c[301]) );
  DFF \creg_reg[302]  ( .D(creg_next[302]), .CLK(clk), .RST(rst), .I(m[302]), 
        .Q(c[302]) );
  DFF \creg_reg[303]  ( .D(creg_next[303]), .CLK(clk), .RST(rst), .I(m[303]), 
        .Q(c[303]) );
  DFF \creg_reg[304]  ( .D(creg_next[304]), .CLK(clk), .RST(rst), .I(m[304]), 
        .Q(c[304]) );
  DFF \creg_reg[305]  ( .D(creg_next[305]), .CLK(clk), .RST(rst), .I(m[305]), 
        .Q(c[305]) );
  DFF \creg_reg[306]  ( .D(creg_next[306]), .CLK(clk), .RST(rst), .I(m[306]), 
        .Q(c[306]) );
  DFF \creg_reg[307]  ( .D(creg_next[307]), .CLK(clk), .RST(rst), .I(m[307]), 
        .Q(c[307]) );
  DFF \creg_reg[308]  ( .D(creg_next[308]), .CLK(clk), .RST(rst), .I(m[308]), 
        .Q(c[308]) );
  DFF \creg_reg[309]  ( .D(creg_next[309]), .CLK(clk), .RST(rst), .I(m[309]), 
        .Q(c[309]) );
  DFF \creg_reg[310]  ( .D(creg_next[310]), .CLK(clk), .RST(rst), .I(m[310]), 
        .Q(c[310]) );
  DFF \creg_reg[311]  ( .D(creg_next[311]), .CLK(clk), .RST(rst), .I(m[311]), 
        .Q(c[311]) );
  DFF \creg_reg[312]  ( .D(creg_next[312]), .CLK(clk), .RST(rst), .I(m[312]), 
        .Q(c[312]) );
  DFF \creg_reg[313]  ( .D(creg_next[313]), .CLK(clk), .RST(rst), .I(m[313]), 
        .Q(c[313]) );
  DFF \creg_reg[314]  ( .D(creg_next[314]), .CLK(clk), .RST(rst), .I(m[314]), 
        .Q(c[314]) );
  DFF \creg_reg[315]  ( .D(creg_next[315]), .CLK(clk), .RST(rst), .I(m[315]), 
        .Q(c[315]) );
  DFF \creg_reg[316]  ( .D(creg_next[316]), .CLK(clk), .RST(rst), .I(m[316]), 
        .Q(c[316]) );
  DFF \creg_reg[317]  ( .D(creg_next[317]), .CLK(clk), .RST(rst), .I(m[317]), 
        .Q(c[317]) );
  DFF \creg_reg[318]  ( .D(creg_next[318]), .CLK(clk), .RST(rst), .I(m[318]), 
        .Q(c[318]) );
  DFF \creg_reg[319]  ( .D(creg_next[319]), .CLK(clk), .RST(rst), .I(m[319]), 
        .Q(c[319]) );
  DFF \creg_reg[320]  ( .D(creg_next[320]), .CLK(clk), .RST(rst), .I(m[320]), 
        .Q(c[320]) );
  DFF \creg_reg[321]  ( .D(creg_next[321]), .CLK(clk), .RST(rst), .I(m[321]), 
        .Q(c[321]) );
  DFF \creg_reg[322]  ( .D(creg_next[322]), .CLK(clk), .RST(rst), .I(m[322]), 
        .Q(c[322]) );
  DFF \creg_reg[323]  ( .D(creg_next[323]), .CLK(clk), .RST(rst), .I(m[323]), 
        .Q(c[323]) );
  DFF \creg_reg[324]  ( .D(creg_next[324]), .CLK(clk), .RST(rst), .I(m[324]), 
        .Q(c[324]) );
  DFF \creg_reg[325]  ( .D(creg_next[325]), .CLK(clk), .RST(rst), .I(m[325]), 
        .Q(c[325]) );
  DFF \creg_reg[326]  ( .D(creg_next[326]), .CLK(clk), .RST(rst), .I(m[326]), 
        .Q(c[326]) );
  DFF \creg_reg[327]  ( .D(creg_next[327]), .CLK(clk), .RST(rst), .I(m[327]), 
        .Q(c[327]) );
  DFF \creg_reg[328]  ( .D(creg_next[328]), .CLK(clk), .RST(rst), .I(m[328]), 
        .Q(c[328]) );
  DFF \creg_reg[329]  ( .D(creg_next[329]), .CLK(clk), .RST(rst), .I(m[329]), 
        .Q(c[329]) );
  DFF \creg_reg[330]  ( .D(creg_next[330]), .CLK(clk), .RST(rst), .I(m[330]), 
        .Q(c[330]) );
  DFF \creg_reg[331]  ( .D(creg_next[331]), .CLK(clk), .RST(rst), .I(m[331]), 
        .Q(c[331]) );
  DFF \creg_reg[332]  ( .D(creg_next[332]), .CLK(clk), .RST(rst), .I(m[332]), 
        .Q(c[332]) );
  DFF \creg_reg[333]  ( .D(creg_next[333]), .CLK(clk), .RST(rst), .I(m[333]), 
        .Q(c[333]) );
  DFF \creg_reg[334]  ( .D(creg_next[334]), .CLK(clk), .RST(rst), .I(m[334]), 
        .Q(c[334]) );
  DFF \creg_reg[335]  ( .D(creg_next[335]), .CLK(clk), .RST(rst), .I(m[335]), 
        .Q(c[335]) );
  DFF \creg_reg[336]  ( .D(creg_next[336]), .CLK(clk), .RST(rst), .I(m[336]), 
        .Q(c[336]) );
  DFF \creg_reg[337]  ( .D(creg_next[337]), .CLK(clk), .RST(rst), .I(m[337]), 
        .Q(c[337]) );
  DFF \creg_reg[338]  ( .D(creg_next[338]), .CLK(clk), .RST(rst), .I(m[338]), 
        .Q(c[338]) );
  DFF \creg_reg[339]  ( .D(creg_next[339]), .CLK(clk), .RST(rst), .I(m[339]), 
        .Q(c[339]) );
  DFF \creg_reg[340]  ( .D(creg_next[340]), .CLK(clk), .RST(rst), .I(m[340]), 
        .Q(c[340]) );
  DFF \creg_reg[341]  ( .D(creg_next[341]), .CLK(clk), .RST(rst), .I(m[341]), 
        .Q(c[341]) );
  DFF \creg_reg[342]  ( .D(creg_next[342]), .CLK(clk), .RST(rst), .I(m[342]), 
        .Q(c[342]) );
  DFF \creg_reg[343]  ( .D(creg_next[343]), .CLK(clk), .RST(rst), .I(m[343]), 
        .Q(c[343]) );
  DFF \creg_reg[344]  ( .D(creg_next[344]), .CLK(clk), .RST(rst), .I(m[344]), 
        .Q(c[344]) );
  DFF \creg_reg[345]  ( .D(creg_next[345]), .CLK(clk), .RST(rst), .I(m[345]), 
        .Q(c[345]) );
  DFF \creg_reg[346]  ( .D(creg_next[346]), .CLK(clk), .RST(rst), .I(m[346]), 
        .Q(c[346]) );
  DFF \creg_reg[347]  ( .D(creg_next[347]), .CLK(clk), .RST(rst), .I(m[347]), 
        .Q(c[347]) );
  DFF \creg_reg[348]  ( .D(creg_next[348]), .CLK(clk), .RST(rst), .I(m[348]), 
        .Q(c[348]) );
  DFF \creg_reg[349]  ( .D(creg_next[349]), .CLK(clk), .RST(rst), .I(m[349]), 
        .Q(c[349]) );
  DFF \creg_reg[350]  ( .D(creg_next[350]), .CLK(clk), .RST(rst), .I(m[350]), 
        .Q(c[350]) );
  DFF \creg_reg[351]  ( .D(creg_next[351]), .CLK(clk), .RST(rst), .I(m[351]), 
        .Q(c[351]) );
  DFF \creg_reg[352]  ( .D(creg_next[352]), .CLK(clk), .RST(rst), .I(m[352]), 
        .Q(c[352]) );
  DFF \creg_reg[353]  ( .D(creg_next[353]), .CLK(clk), .RST(rst), .I(m[353]), 
        .Q(c[353]) );
  DFF \creg_reg[354]  ( .D(creg_next[354]), .CLK(clk), .RST(rst), .I(m[354]), 
        .Q(c[354]) );
  DFF \creg_reg[355]  ( .D(creg_next[355]), .CLK(clk), .RST(rst), .I(m[355]), 
        .Q(c[355]) );
  DFF \creg_reg[356]  ( .D(creg_next[356]), .CLK(clk), .RST(rst), .I(m[356]), 
        .Q(c[356]) );
  DFF \creg_reg[357]  ( .D(creg_next[357]), .CLK(clk), .RST(rst), .I(m[357]), 
        .Q(c[357]) );
  DFF \creg_reg[358]  ( .D(creg_next[358]), .CLK(clk), .RST(rst), .I(m[358]), 
        .Q(c[358]) );
  DFF \creg_reg[359]  ( .D(creg_next[359]), .CLK(clk), .RST(rst), .I(m[359]), 
        .Q(c[359]) );
  DFF \creg_reg[360]  ( .D(creg_next[360]), .CLK(clk), .RST(rst), .I(m[360]), 
        .Q(c[360]) );
  DFF \creg_reg[361]  ( .D(creg_next[361]), .CLK(clk), .RST(rst), .I(m[361]), 
        .Q(c[361]) );
  DFF \creg_reg[362]  ( .D(creg_next[362]), .CLK(clk), .RST(rst), .I(m[362]), 
        .Q(c[362]) );
  DFF \creg_reg[363]  ( .D(creg_next[363]), .CLK(clk), .RST(rst), .I(m[363]), 
        .Q(c[363]) );
  DFF \creg_reg[364]  ( .D(creg_next[364]), .CLK(clk), .RST(rst), .I(m[364]), 
        .Q(c[364]) );
  DFF \creg_reg[365]  ( .D(creg_next[365]), .CLK(clk), .RST(rst), .I(m[365]), 
        .Q(c[365]) );
  DFF \creg_reg[366]  ( .D(creg_next[366]), .CLK(clk), .RST(rst), .I(m[366]), 
        .Q(c[366]) );
  DFF \creg_reg[367]  ( .D(creg_next[367]), .CLK(clk), .RST(rst), .I(m[367]), 
        .Q(c[367]) );
  DFF \creg_reg[368]  ( .D(creg_next[368]), .CLK(clk), .RST(rst), .I(m[368]), 
        .Q(c[368]) );
  DFF \creg_reg[369]  ( .D(creg_next[369]), .CLK(clk), .RST(rst), .I(m[369]), 
        .Q(c[369]) );
  DFF \creg_reg[370]  ( .D(creg_next[370]), .CLK(clk), .RST(rst), .I(m[370]), 
        .Q(c[370]) );
  DFF \creg_reg[371]  ( .D(creg_next[371]), .CLK(clk), .RST(rst), .I(m[371]), 
        .Q(c[371]) );
  DFF \creg_reg[372]  ( .D(creg_next[372]), .CLK(clk), .RST(rst), .I(m[372]), 
        .Q(c[372]) );
  DFF \creg_reg[373]  ( .D(creg_next[373]), .CLK(clk), .RST(rst), .I(m[373]), 
        .Q(c[373]) );
  DFF \creg_reg[374]  ( .D(creg_next[374]), .CLK(clk), .RST(rst), .I(m[374]), 
        .Q(c[374]) );
  DFF \creg_reg[375]  ( .D(creg_next[375]), .CLK(clk), .RST(rst), .I(m[375]), 
        .Q(c[375]) );
  DFF \creg_reg[376]  ( .D(creg_next[376]), .CLK(clk), .RST(rst), .I(m[376]), 
        .Q(c[376]) );
  DFF \creg_reg[377]  ( .D(creg_next[377]), .CLK(clk), .RST(rst), .I(m[377]), 
        .Q(c[377]) );
  DFF \creg_reg[378]  ( .D(creg_next[378]), .CLK(clk), .RST(rst), .I(m[378]), 
        .Q(c[378]) );
  DFF \creg_reg[379]  ( .D(creg_next[379]), .CLK(clk), .RST(rst), .I(m[379]), 
        .Q(c[379]) );
  DFF \creg_reg[380]  ( .D(creg_next[380]), .CLK(clk), .RST(rst), .I(m[380]), 
        .Q(c[380]) );
  DFF \creg_reg[381]  ( .D(creg_next[381]), .CLK(clk), .RST(rst), .I(m[381]), 
        .Q(c[381]) );
  DFF \creg_reg[382]  ( .D(creg_next[382]), .CLK(clk), .RST(rst), .I(m[382]), 
        .Q(c[382]) );
  DFF \creg_reg[383]  ( .D(creg_next[383]), .CLK(clk), .RST(rst), .I(m[383]), 
        .Q(c[383]) );
  DFF \creg_reg[384]  ( .D(creg_next[384]), .CLK(clk), .RST(rst), .I(m[384]), 
        .Q(c[384]) );
  DFF \creg_reg[385]  ( .D(creg_next[385]), .CLK(clk), .RST(rst), .I(m[385]), 
        .Q(c[385]) );
  DFF \creg_reg[386]  ( .D(creg_next[386]), .CLK(clk), .RST(rst), .I(m[386]), 
        .Q(c[386]) );
  DFF \creg_reg[387]  ( .D(creg_next[387]), .CLK(clk), .RST(rst), .I(m[387]), 
        .Q(c[387]) );
  DFF \creg_reg[388]  ( .D(creg_next[388]), .CLK(clk), .RST(rst), .I(m[388]), 
        .Q(c[388]) );
  DFF \creg_reg[389]  ( .D(creg_next[389]), .CLK(clk), .RST(rst), .I(m[389]), 
        .Q(c[389]) );
  DFF \creg_reg[390]  ( .D(creg_next[390]), .CLK(clk), .RST(rst), .I(m[390]), 
        .Q(c[390]) );
  DFF \creg_reg[391]  ( .D(creg_next[391]), .CLK(clk), .RST(rst), .I(m[391]), 
        .Q(c[391]) );
  DFF \creg_reg[392]  ( .D(creg_next[392]), .CLK(clk), .RST(rst), .I(m[392]), 
        .Q(c[392]) );
  DFF \creg_reg[393]  ( .D(creg_next[393]), .CLK(clk), .RST(rst), .I(m[393]), 
        .Q(c[393]) );
  DFF \creg_reg[394]  ( .D(creg_next[394]), .CLK(clk), .RST(rst), .I(m[394]), 
        .Q(c[394]) );
  DFF \creg_reg[395]  ( .D(creg_next[395]), .CLK(clk), .RST(rst), .I(m[395]), 
        .Q(c[395]) );
  DFF \creg_reg[396]  ( .D(creg_next[396]), .CLK(clk), .RST(rst), .I(m[396]), 
        .Q(c[396]) );
  DFF \creg_reg[397]  ( .D(creg_next[397]), .CLK(clk), .RST(rst), .I(m[397]), 
        .Q(c[397]) );
  DFF \creg_reg[398]  ( .D(creg_next[398]), .CLK(clk), .RST(rst), .I(m[398]), 
        .Q(c[398]) );
  DFF \creg_reg[399]  ( .D(creg_next[399]), .CLK(clk), .RST(rst), .I(m[399]), 
        .Q(c[399]) );
  DFF \creg_reg[400]  ( .D(creg_next[400]), .CLK(clk), .RST(rst), .I(m[400]), 
        .Q(c[400]) );
  DFF \creg_reg[401]  ( .D(creg_next[401]), .CLK(clk), .RST(rst), .I(m[401]), 
        .Q(c[401]) );
  DFF \creg_reg[402]  ( .D(creg_next[402]), .CLK(clk), .RST(rst), .I(m[402]), 
        .Q(c[402]) );
  DFF \creg_reg[403]  ( .D(creg_next[403]), .CLK(clk), .RST(rst), .I(m[403]), 
        .Q(c[403]) );
  DFF \creg_reg[404]  ( .D(creg_next[404]), .CLK(clk), .RST(rst), .I(m[404]), 
        .Q(c[404]) );
  DFF \creg_reg[405]  ( .D(creg_next[405]), .CLK(clk), .RST(rst), .I(m[405]), 
        .Q(c[405]) );
  DFF \creg_reg[406]  ( .D(creg_next[406]), .CLK(clk), .RST(rst), .I(m[406]), 
        .Q(c[406]) );
  DFF \creg_reg[407]  ( .D(creg_next[407]), .CLK(clk), .RST(rst), .I(m[407]), 
        .Q(c[407]) );
  DFF \creg_reg[408]  ( .D(creg_next[408]), .CLK(clk), .RST(rst), .I(m[408]), 
        .Q(c[408]) );
  DFF \creg_reg[409]  ( .D(creg_next[409]), .CLK(clk), .RST(rst), .I(m[409]), 
        .Q(c[409]) );
  DFF \creg_reg[410]  ( .D(creg_next[410]), .CLK(clk), .RST(rst), .I(m[410]), 
        .Q(c[410]) );
  DFF \creg_reg[411]  ( .D(creg_next[411]), .CLK(clk), .RST(rst), .I(m[411]), 
        .Q(c[411]) );
  DFF \creg_reg[412]  ( .D(creg_next[412]), .CLK(clk), .RST(rst), .I(m[412]), 
        .Q(c[412]) );
  DFF \creg_reg[413]  ( .D(creg_next[413]), .CLK(clk), .RST(rst), .I(m[413]), 
        .Q(c[413]) );
  DFF \creg_reg[414]  ( .D(creg_next[414]), .CLK(clk), .RST(rst), .I(m[414]), 
        .Q(c[414]) );
  DFF \creg_reg[415]  ( .D(creg_next[415]), .CLK(clk), .RST(rst), .I(m[415]), 
        .Q(c[415]) );
  DFF \creg_reg[416]  ( .D(creg_next[416]), .CLK(clk), .RST(rst), .I(m[416]), 
        .Q(c[416]) );
  DFF \creg_reg[417]  ( .D(creg_next[417]), .CLK(clk), .RST(rst), .I(m[417]), 
        .Q(c[417]) );
  DFF \creg_reg[418]  ( .D(creg_next[418]), .CLK(clk), .RST(rst), .I(m[418]), 
        .Q(c[418]) );
  DFF \creg_reg[419]  ( .D(creg_next[419]), .CLK(clk), .RST(rst), .I(m[419]), 
        .Q(c[419]) );
  DFF \creg_reg[420]  ( .D(creg_next[420]), .CLK(clk), .RST(rst), .I(m[420]), 
        .Q(c[420]) );
  DFF \creg_reg[421]  ( .D(creg_next[421]), .CLK(clk), .RST(rst), .I(m[421]), 
        .Q(c[421]) );
  DFF \creg_reg[422]  ( .D(creg_next[422]), .CLK(clk), .RST(rst), .I(m[422]), 
        .Q(c[422]) );
  DFF \creg_reg[423]  ( .D(creg_next[423]), .CLK(clk), .RST(rst), .I(m[423]), 
        .Q(c[423]) );
  DFF \creg_reg[424]  ( .D(creg_next[424]), .CLK(clk), .RST(rst), .I(m[424]), 
        .Q(c[424]) );
  DFF \creg_reg[425]  ( .D(creg_next[425]), .CLK(clk), .RST(rst), .I(m[425]), 
        .Q(c[425]) );
  DFF \creg_reg[426]  ( .D(creg_next[426]), .CLK(clk), .RST(rst), .I(m[426]), 
        .Q(c[426]) );
  DFF \creg_reg[427]  ( .D(creg_next[427]), .CLK(clk), .RST(rst), .I(m[427]), 
        .Q(c[427]) );
  DFF \creg_reg[428]  ( .D(creg_next[428]), .CLK(clk), .RST(rst), .I(m[428]), 
        .Q(c[428]) );
  DFF \creg_reg[429]  ( .D(creg_next[429]), .CLK(clk), .RST(rst), .I(m[429]), 
        .Q(c[429]) );
  DFF \creg_reg[430]  ( .D(creg_next[430]), .CLK(clk), .RST(rst), .I(m[430]), 
        .Q(c[430]) );
  DFF \creg_reg[431]  ( .D(creg_next[431]), .CLK(clk), .RST(rst), .I(m[431]), 
        .Q(c[431]) );
  DFF \creg_reg[432]  ( .D(creg_next[432]), .CLK(clk), .RST(rst), .I(m[432]), 
        .Q(c[432]) );
  DFF \creg_reg[433]  ( .D(creg_next[433]), .CLK(clk), .RST(rst), .I(m[433]), 
        .Q(c[433]) );
  DFF \creg_reg[434]  ( .D(creg_next[434]), .CLK(clk), .RST(rst), .I(m[434]), 
        .Q(c[434]) );
  DFF \creg_reg[435]  ( .D(creg_next[435]), .CLK(clk), .RST(rst), .I(m[435]), 
        .Q(c[435]) );
  DFF \creg_reg[436]  ( .D(creg_next[436]), .CLK(clk), .RST(rst), .I(m[436]), 
        .Q(c[436]) );
  DFF \creg_reg[437]  ( .D(creg_next[437]), .CLK(clk), .RST(rst), .I(m[437]), 
        .Q(c[437]) );
  DFF \creg_reg[438]  ( .D(creg_next[438]), .CLK(clk), .RST(rst), .I(m[438]), 
        .Q(c[438]) );
  DFF \creg_reg[439]  ( .D(creg_next[439]), .CLK(clk), .RST(rst), .I(m[439]), 
        .Q(c[439]) );
  DFF \creg_reg[440]  ( .D(creg_next[440]), .CLK(clk), .RST(rst), .I(m[440]), 
        .Q(c[440]) );
  DFF \creg_reg[441]  ( .D(creg_next[441]), .CLK(clk), .RST(rst), .I(m[441]), 
        .Q(c[441]) );
  DFF \creg_reg[442]  ( .D(creg_next[442]), .CLK(clk), .RST(rst), .I(m[442]), 
        .Q(c[442]) );
  DFF \creg_reg[443]  ( .D(creg_next[443]), .CLK(clk), .RST(rst), .I(m[443]), 
        .Q(c[443]) );
  DFF \creg_reg[444]  ( .D(creg_next[444]), .CLK(clk), .RST(rst), .I(m[444]), 
        .Q(c[444]) );
  DFF \creg_reg[445]  ( .D(creg_next[445]), .CLK(clk), .RST(rst), .I(m[445]), 
        .Q(c[445]) );
  DFF \creg_reg[446]  ( .D(creg_next[446]), .CLK(clk), .RST(rst), .I(m[446]), 
        .Q(c[446]) );
  DFF \creg_reg[447]  ( .D(creg_next[447]), .CLK(clk), .RST(rst), .I(m[447]), 
        .Q(c[447]) );
  DFF \creg_reg[448]  ( .D(creg_next[448]), .CLK(clk), .RST(rst), .I(m[448]), 
        .Q(c[448]) );
  DFF \creg_reg[449]  ( .D(creg_next[449]), .CLK(clk), .RST(rst), .I(m[449]), 
        .Q(c[449]) );
  DFF \creg_reg[450]  ( .D(creg_next[450]), .CLK(clk), .RST(rst), .I(m[450]), 
        .Q(c[450]) );
  DFF \creg_reg[451]  ( .D(creg_next[451]), .CLK(clk), .RST(rst), .I(m[451]), 
        .Q(c[451]) );
  DFF \creg_reg[452]  ( .D(creg_next[452]), .CLK(clk), .RST(rst), .I(m[452]), 
        .Q(c[452]) );
  DFF \creg_reg[453]  ( .D(creg_next[453]), .CLK(clk), .RST(rst), .I(m[453]), 
        .Q(c[453]) );
  DFF \creg_reg[454]  ( .D(creg_next[454]), .CLK(clk), .RST(rst), .I(m[454]), 
        .Q(c[454]) );
  DFF \creg_reg[455]  ( .D(creg_next[455]), .CLK(clk), .RST(rst), .I(m[455]), 
        .Q(c[455]) );
  DFF \creg_reg[456]  ( .D(creg_next[456]), .CLK(clk), .RST(rst), .I(m[456]), 
        .Q(c[456]) );
  DFF \creg_reg[457]  ( .D(creg_next[457]), .CLK(clk), .RST(rst), .I(m[457]), 
        .Q(c[457]) );
  DFF \creg_reg[458]  ( .D(creg_next[458]), .CLK(clk), .RST(rst), .I(m[458]), 
        .Q(c[458]) );
  DFF \creg_reg[459]  ( .D(creg_next[459]), .CLK(clk), .RST(rst), .I(m[459]), 
        .Q(c[459]) );
  DFF \creg_reg[460]  ( .D(creg_next[460]), .CLK(clk), .RST(rst), .I(m[460]), 
        .Q(c[460]) );
  DFF \creg_reg[461]  ( .D(creg_next[461]), .CLK(clk), .RST(rst), .I(m[461]), 
        .Q(c[461]) );
  DFF \creg_reg[462]  ( .D(creg_next[462]), .CLK(clk), .RST(rst), .I(m[462]), 
        .Q(c[462]) );
  DFF \creg_reg[463]  ( .D(creg_next[463]), .CLK(clk), .RST(rst), .I(m[463]), 
        .Q(c[463]) );
  DFF \creg_reg[464]  ( .D(creg_next[464]), .CLK(clk), .RST(rst), .I(m[464]), 
        .Q(c[464]) );
  DFF \creg_reg[465]  ( .D(creg_next[465]), .CLK(clk), .RST(rst), .I(m[465]), 
        .Q(c[465]) );
  DFF \creg_reg[466]  ( .D(creg_next[466]), .CLK(clk), .RST(rst), .I(m[466]), 
        .Q(c[466]) );
  DFF \creg_reg[467]  ( .D(creg_next[467]), .CLK(clk), .RST(rst), .I(m[467]), 
        .Q(c[467]) );
  DFF \creg_reg[468]  ( .D(creg_next[468]), .CLK(clk), .RST(rst), .I(m[468]), 
        .Q(c[468]) );
  DFF \creg_reg[469]  ( .D(creg_next[469]), .CLK(clk), .RST(rst), .I(m[469]), 
        .Q(c[469]) );
  DFF \creg_reg[470]  ( .D(creg_next[470]), .CLK(clk), .RST(rst), .I(m[470]), 
        .Q(c[470]) );
  DFF \creg_reg[471]  ( .D(creg_next[471]), .CLK(clk), .RST(rst), .I(m[471]), 
        .Q(c[471]) );
  DFF \creg_reg[472]  ( .D(creg_next[472]), .CLK(clk), .RST(rst), .I(m[472]), 
        .Q(c[472]) );
  DFF \creg_reg[473]  ( .D(creg_next[473]), .CLK(clk), .RST(rst), .I(m[473]), 
        .Q(c[473]) );
  DFF \creg_reg[474]  ( .D(creg_next[474]), .CLK(clk), .RST(rst), .I(m[474]), 
        .Q(c[474]) );
  DFF \creg_reg[475]  ( .D(creg_next[475]), .CLK(clk), .RST(rst), .I(m[475]), 
        .Q(c[475]) );
  DFF \creg_reg[476]  ( .D(creg_next[476]), .CLK(clk), .RST(rst), .I(m[476]), 
        .Q(c[476]) );
  DFF \creg_reg[477]  ( .D(creg_next[477]), .CLK(clk), .RST(rst), .I(m[477]), 
        .Q(c[477]) );
  DFF \creg_reg[478]  ( .D(creg_next[478]), .CLK(clk), .RST(rst), .I(m[478]), 
        .Q(c[478]) );
  DFF \creg_reg[479]  ( .D(creg_next[479]), .CLK(clk), .RST(rst), .I(m[479]), 
        .Q(c[479]) );
  DFF \creg_reg[480]  ( .D(creg_next[480]), .CLK(clk), .RST(rst), .I(m[480]), 
        .Q(c[480]) );
  DFF \creg_reg[481]  ( .D(creg_next[481]), .CLK(clk), .RST(rst), .I(m[481]), 
        .Q(c[481]) );
  DFF \creg_reg[482]  ( .D(creg_next[482]), .CLK(clk), .RST(rst), .I(m[482]), 
        .Q(c[482]) );
  DFF \creg_reg[483]  ( .D(creg_next[483]), .CLK(clk), .RST(rst), .I(m[483]), 
        .Q(c[483]) );
  DFF \creg_reg[484]  ( .D(creg_next[484]), .CLK(clk), .RST(rst), .I(m[484]), 
        .Q(c[484]) );
  DFF \creg_reg[485]  ( .D(creg_next[485]), .CLK(clk), .RST(rst), .I(m[485]), 
        .Q(c[485]) );
  DFF \creg_reg[486]  ( .D(creg_next[486]), .CLK(clk), .RST(rst), .I(m[486]), 
        .Q(c[486]) );
  DFF \creg_reg[487]  ( .D(creg_next[487]), .CLK(clk), .RST(rst), .I(m[487]), 
        .Q(c[487]) );
  DFF \creg_reg[488]  ( .D(creg_next[488]), .CLK(clk), .RST(rst), .I(m[488]), 
        .Q(c[488]) );
  DFF \creg_reg[489]  ( .D(creg_next[489]), .CLK(clk), .RST(rst), .I(m[489]), 
        .Q(c[489]) );
  DFF \creg_reg[490]  ( .D(creg_next[490]), .CLK(clk), .RST(rst), .I(m[490]), 
        .Q(c[490]) );
  DFF \creg_reg[491]  ( .D(creg_next[491]), .CLK(clk), .RST(rst), .I(m[491]), 
        .Q(c[491]) );
  DFF \creg_reg[492]  ( .D(creg_next[492]), .CLK(clk), .RST(rst), .I(m[492]), 
        .Q(c[492]) );
  DFF \creg_reg[493]  ( .D(creg_next[493]), .CLK(clk), .RST(rst), .I(m[493]), 
        .Q(c[493]) );
  DFF \creg_reg[494]  ( .D(creg_next[494]), .CLK(clk), .RST(rst), .I(m[494]), 
        .Q(c[494]) );
  DFF \creg_reg[495]  ( .D(creg_next[495]), .CLK(clk), .RST(rst), .I(m[495]), 
        .Q(c[495]) );
  DFF \creg_reg[496]  ( .D(creg_next[496]), .CLK(clk), .RST(rst), .I(m[496]), 
        .Q(c[496]) );
  DFF \creg_reg[497]  ( .D(creg_next[497]), .CLK(clk), .RST(rst), .I(m[497]), 
        .Q(c[497]) );
  DFF \creg_reg[498]  ( .D(creg_next[498]), .CLK(clk), .RST(rst), .I(m[498]), 
        .Q(c[498]) );
  DFF \creg_reg[499]  ( .D(creg_next[499]), .CLK(clk), .RST(rst), .I(m[499]), 
        .Q(c[499]) );
  DFF \creg_reg[500]  ( .D(creg_next[500]), .CLK(clk), .RST(rst), .I(m[500]), 
        .Q(c[500]) );
  DFF \creg_reg[501]  ( .D(creg_next[501]), .CLK(clk), .RST(rst), .I(m[501]), 
        .Q(c[501]) );
  DFF \creg_reg[502]  ( .D(creg_next[502]), .CLK(clk), .RST(rst), .I(m[502]), 
        .Q(c[502]) );
  DFF \creg_reg[503]  ( .D(creg_next[503]), .CLK(clk), .RST(rst), .I(m[503]), 
        .Q(c[503]) );
  DFF \creg_reg[504]  ( .D(creg_next[504]), .CLK(clk), .RST(rst), .I(m[504]), 
        .Q(c[504]) );
  DFF \creg_reg[505]  ( .D(creg_next[505]), .CLK(clk), .RST(rst), .I(m[505]), 
        .Q(c[505]) );
  DFF \creg_reg[506]  ( .D(creg_next[506]), .CLK(clk), .RST(rst), .I(m[506]), 
        .Q(c[506]) );
  DFF \creg_reg[507]  ( .D(creg_next[507]), .CLK(clk), .RST(rst), .I(m[507]), 
        .Q(c[507]) );
  DFF \creg_reg[508]  ( .D(creg_next[508]), .CLK(clk), .RST(rst), .I(m[508]), 
        .Q(c[508]) );
  DFF \creg_reg[509]  ( .D(creg_next[509]), .CLK(clk), .RST(rst), .I(m[509]), 
        .Q(c[509]) );
  DFF \creg_reg[510]  ( .D(creg_next[510]), .CLK(clk), .RST(rst), .I(m[510]), 
        .Q(c[510]) );
  DFF \creg_reg[511]  ( .D(creg_next[511]), .CLK(clk), .RST(rst), .I(m[511]), 
        .Q(c[511]) );
  XOR U268 ( .A(start_in[255]), .B(mul_pow), .Z(n8) );
  NANDN U269 ( .A(first_one), .B(n265), .Z(n6) );
  NAND U270 ( .A(n266), .B(ein[511]), .Z(n265) );
  AND U271 ( .A(mul_pow), .B(start_in[255]), .Z(n266) );
  NAND U272 ( .A(n267), .B(n268), .Z(_0_net_) );
  NANDN U273 ( .A(mul_pow), .B(first_one), .Z(n268) );
  NAND U274 ( .A(first_one), .B(ein[511]), .Z(n267) );
endmodule

